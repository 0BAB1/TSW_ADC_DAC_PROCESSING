`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
bB3w6vpa/Oso6U8HvvOuFoW9KR4zPzMkDxboJLfdKo5jAH1AZ0zKKvQ3VQpOR23ZZ3//ML4IYA/e
iRQnL1oU4w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gJvN6jU7WgZGTYPlWORWL2sCJeVqFotmkzzhpTanGs2ES8S0SC2sX4wznXq6/j0Qu+yoyLNeeDX3
DqG3m6VtpMqV+9fYbcZMp0r6eIh94dNTRSCnz7WfNcGURoEdC9zvU7vIRiul/4b1prSWnSmvAzpv
PQp+pq93tv0xbqFysvQ=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Bpd5n0lMjLHvqOGB8VcXAkbpSPNzWcGIuvH6kY7bnRaDG1nLwL4PrOu1KBU+/VM4sapEDDS2mv66
TUxUntOlvXEWt/RPH7J1Y+/KXtITPT2eKPT+jUU2HZyklXgn0DeFga9bKsgiQGV+55mH+KUB88C+
43jSisdvSTvdOU26pIY=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nimNs+xhbKAwhxaKoqPCURIiRH8F3C5qRC+6UsGsRobOzQHJlj596hfppbIJnvkKiaTfiqL/XRrV
ZJ2hLHV80vEog+9wor9KyCCVD/uiTt+RdNSYGmkFpN1LshEvCV8K4lIYs8Q5vSFx3oiKsOI+li+D
uBSjoC5i5sRBKoBtF+G0awtRPj4i2FlYp1O7aXvaCCwFeGI6aB//ToqRIss3ZGa1mtX+ZXE+hvJu
RRn83Kjh16LPsPDWVuRnNxeTqCIh2a5MlAZIVcZDPHLXFqOtRgpmKF/GFDHu8rbl4JuOn6Y/rtWR
yUwmOQXoYEE50HOU9WFwe+m+i98HaKOehcV1TQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
H/lhjU+VaTiz7yess64ckTbyFEL3FRoOorAWGleulrpp8+z3h7QdkU6sOo+yH55kF8FfgjySYssB
vCS4NJXHa3pmMJKsLzN1cXaNNx2NNjZF0+PXTUQgwkLhCJtEcvXdUdUS3nEyzvoVKd+ZYFvfsjOx
LhEXmRztJLSjq1Wst3Ab2u55aq2PB7x1rZRAs/UqeOhbne9dY561VGuKDsfwM1pXDD72GgjuaLyk
6it5I9AedeYxO42QXJJ0lhHY4cp5nBEY3RQs7WtpKxxfhbsqLD5OZLOUKn6bViCxnNEvoFyrM5vo
5ItgMv5CoJQzvin4OMCy5icBHqTLErUa1s+i9Q==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
xDaVGO3uvvE1L0LfXZu+8FfEfII+DPN+hcPsii9gS6vMUdQmBhSpnm0d1A7sSZtx0Ugdo1afWGc+
1RQwqroFGiP/aNX5aosV/BV0xu/c6+44bwSNUJTJnFiDgLJtHWxTsV1tGIu2WqLgBvAALxIrTQbP
vCwvjf3pEpWXpNjftlaCgYVMShwndLyqc3sH1varFNFyfdyLGItJI2vSVn4m0TbXfkVO21jOyEHH
HqwUvQmgo9Mfi/2spyRPUiXsy9iRgSEm4xQwjpYKYyIvIyAakJFjwgJqKfZjev4esMtfP4d/Xm3U
P5cbE+C7X1DMr+mUF4q+ctZ3kzhCJyQbnEnjUg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1798864)
`protect data_block
g/KvXozXI7fclKNmZqdsRFRMfrZ8i9hUjq/QhRBJVSXBvYw2fBcTj5qEnQqE+rYMmML5L3lJhIGk
QWXfeX4GBz4Aez2yqeTXqj0q9i71eUv9cNC8QTKPxKD+hp5mwqneFtQV/yHx1RZF5noERFamyXUo
jIOiiYmD1ZUFuXb1nLysmRkeMDOOWOufxjvXw4yMQuwMi9sqS4i21voS4fwhIosIluYExbs5Ra3g
HNZezV7EGXBKaCnB30h7Vk53GYRVs1yE9p9+amDi6uwqR9h4xGwj662c8n3f/pnzmUflVGQav5nf
BAt1D6bbGRSBT23B6wfHVrORSwRi560t5zY6JWvwmhbTVw8kA0ucA2y8xk9MjySDNEhmW6I8nqs+
/bXu8AbtOSCWVriLWFLqSoMx5BIaJOI0xorieOOsmJis+zxaSTJfRrd9zKXd97h00QgM/Jly1CwB
iihXlXP3sAqXSdvyzIemdGhLzEa/m3oxUEftBp5CN3MQ2gb7PkXsiNvrk+YMVQJBKON3SloibgNQ
1J0Ilps5PPxE+4RQWUhBcCzuKCF+4VRz3RWISTa3JPPLozG5wmfswOV9+ujM0H5xQbSzvxkF6esx
wSWTMr9rILGT4olf63dligYYa+9Bpd4UCaPwBdKeDPVy73lCZ8ocGznVcqnOLvIYT8GM+GXcKHm6
rDOoiog8/MOCGpGY9ekGFwJvUGanMMLrgWsvUNSD5ysYd14gbPXon/9Fd8cmnryR+vGgOmZlkig5
v15q7C2bFtw7CsCMgL9U8ooZDZ+WgMZv4xoABqDi8VN05unCRJ+A4UZHmVQGxiT7fsZTNQkWuIGK
DI2ibFgLOPdqQrpirM6zltSmV9e8qtYVyX4HRbIH3ctapxUsRCmIoyqsisfoDbywKU7T5qP7QTh0
Wtrkyr0er2uBx6GSgq32vxlNwZWol7ovTql3cuQ+WN8KcpLkRKDql0PvKnZce38Y4EGc/cFsEU4s
WPNuh+QqCScOazDfM9Zrj2po3npnP0sbb+sbsRaCartxZi808zZjjebUtuiIJZibPjYSfJTpy7UW
yYzF+8mqWYm5v0k23whSCobcyI1z50ou7Afv/irRVOGp6LBsaZFieCQP0Ydx/g4oTJFoubE2W3aJ
gmnfCg896dOcJNidm2LuHHZ5O+1lIufBLbyPlFY6gTpNaffEOUVowa2uXBvxtS/Osg8SpuDlwjYJ
2U02eh3L8Y01HfJwPP3UGEZxbIxc4voAkE66V0+7n9qdBLqkFbVF4fAMCVg93/P6uKAwYY3mGbWW
4ct27l8IEm3ZW86PrtbK46EqDoKDHZo5gQV83mLwydmbMHSmswAnfmITO+UqYpW6XHl66s3cqQBF
ANYeeGv2KpVXCphGKuyQTMYgaq3BYYC1CKUhFHbF/f0+8bARCokjRAfSj1JjZs/AC4Kub5prt2US
D9sXbDBSYg7Nx+G5pJkaMNg/Nq5zn7qYw5WxwsDMlvmKHiETeCc3G9ko2uDwfUo4Lhj7ELZj52qf
DB8y2fh8b2e0zgo1Fl9MRvN6HjmTv7GNLKW+YB2c3m72M483R/B72rvxnZmkhyOyHwGFvGvEKNz2
PFEr8Ss8kM2BarCotjh5gE0bkmmSQ789TWPivy9PxjCYnJp1mWIgUu0jlS6n5Nso4kwT4lyvHfmZ
jqD2BfI4Qwt2ozOz2Dkzm9FVMk86SO82Ymj+lJ7ld7aPsk2o2AmM/YlaIWmSj40o+EAkZsixsFyd
A0PYLwC1rVHC3C79Ch2hVW8EtPfJuoSbONWj+LcZyD57V7VVd204IBkTY5DhAB3Sv0fp+UFMrzcq
4922d9/q+5XuzXj1Zbs6EOfVQ4TuhWUzI5QYgdBaIHrjiepAg+kcl0N3gE6US8zndc14d8ECz1AN
gQIqkQe7OZY2hMnLY0j2KqmSQyXvx0OBYiMBH6ekZmBqVasmNZWfo+srhJji/k0zwmVlIUzcmGec
Ziy+XPWwkLyTUwbjQkjgYKfVc7drUvz+109fThlWW9L96MgoFOrZPlYANv+wkV97qopcGaBvbsq1
jG8loLeF3QFaDKjl4L4iHRGSu8aO3hVVIZHa1YFTCHeDQWabqqwkCtNUjJD8URSU3/L9HPeNpnRC
tlTtcdPojufULM+syxJfMhSUtD+bmgTnUlf1lkfDveNEGnXKVxOnmZ5BHgxdxWGP9Hpn0IV4F6Qv
GAP3GTB8nIH3bh30fWK9hR8l/2tRbkqAeJZKxs52FmwmK0o5cuCyqtcAh02mN6LjpKMC2O0fE4sb
g6UjXcq8/cvf+dd29jWTLav3wynfZPZyjWwVOxpkpUqX53/3zgOFUSSnbRP+a5M3/FjzzUEkqHLk
uIUTLmVowuuiiLHL+kspJSAqwrVXIhXCV7Q7xMYKKocgmnCypgF8WXSyQ8SW2gWYTakeXsNPjv9P
vgh05WGGiuEudDV0b9Cm4CfTeUXh24BlTtA2f/mPyXGwfzdu5MhbmzTwBTdK1USv78BEvMeemZvN
iSvCSZhwHb6kVLe3jkraN3gjH/7taQLTmUmgILCNr43QUSR2dQJ3XmEEyZxqfHeQ7ZE0XTu79T9V
15RcLcnRotyuSLk8oVaI6qhTHOaC/eYH7j0mwSngDK7YQP5SUGU6Gp5JzAtuaqrVjS6Pf0AoKiME
jnO4a8QGrDYSqKg8nOfOamvTe8pWLCDC3L4HzCjXFlxwCjGK606il1lAAeaxEllUM/6PQdgK2jub
EhLzJ60VXDQZUh3BzS4O9Fgq8/XHK4ehIa//psWrb0EQ/8mJlqKe0yit8OC07X1d4JTAfPa9Xsw4
EXgsdHG+yEglWs6PcaiwiTLwX7WrRIKAMDAH9XTw9hIKUM73e20B1D8cOvHG6T5bMdtk1fF4bY9o
wxqLXaq0moFuj5lsZp42Xu79ZTOsO0xWRpy679pU+WqWLJk8P4jc3MDvk++7i/2FYgrJUilZfapX
T2rYJoQyRlEwlKj2TklXyv3VXu/iRTwSRXE1a6BzPlFkr6MGAVzcp8MdxzW5yeGQmPCbkQdF28m8
zR7jGK44ufYxcmNlVkClGHAy7tIe7AJfJ5XyfP24917+Qe4GNVnDsHGHW/Vu6DMa855NRTSkUZ0N
k4t2eHA192wxpQDzIidJN0Ensp7nNQJEjAVK+N41UBw2srRvpqgVGiyBXhCKmiUYWDcbyUbYGhwq
lZ0go2c9W5OsTM7GDH21vfCaA8fZgL1GZJgY7j/Zhenrk98jf1iNuJREJ0Y0fVQg7xN8v6KMPOTu
Ib27LqV8z+uTPwTAw/xvXe1cIhE019Bmv46BcFh9mPuZNijce1+17gyOQVi4xewW7z0O1f428J9r
mf9WsB+6ngt3HBw/5OIDlSZmcEDdWzezYypcjFWqahZ3dmhu4cDCnwh8waMIFAxzuu3c3URptiu5
eeURwKpcMr871ozVAuI/2ft51uw7/eNz9Xz9oZi0FpkRruTOxIocI4S76B3EJ4MXuuPvaE2LwvVq
33Y3ARI4zHz8d6Z5InnGhMCw2ctGjowSXNFi4CW6uRJDIsX6hHRqWwMRxRV3bemDVDQp9HfXUvQP
9+ctqDfH7WqeY9J2uF0kerC48VsDuyYQ7ca+fo1++S41lNNOerIiSIhP401xz6PuxTnWpBEu9nPR
uUhMcjA8XhtVA+FkKULQ7C43ablhRg0FHGMIKjVtPE5K+MKoOxmiW+d8XxchnAgGUa8cLok5Vn4D
WzkH4Htdzqq/YbHP6d8wNDHKNs8/D4UH6nwsHhdyrVgNlHlNvwmQL39CqkovBpKU4R+Y9G3S/cUl
CxMtHP7TVtwrMwbFwHaOmf2hU9Ngv3iqYL2sXj17Y+dGj9i8aD8ebJ2MSckibGKRGLws6qpaAWz2
PtV8x4JzNSq8tMH9BqFtKxmBFte7+OdNR3pCuO8QpwsHXPE73O3sdXrOqkXIL5B4fT2OJ1c5KH6k
/KUUaMeGfVufqoAgds3lyQjRVpiL66ID5jkhDl9OgBGk/jsNf/9dnB1eQLk3Z/nFmB18txPi+4UH
xFiLPfHFOjI6oLh6zXLQkGwqIZCp7sLPp5qadCUk6TNJXQrKlbv0SKYZPFMay9ZSVV+6NrddgDPC
kb+VLnqJjxWaWUs9ifQMKoFFAnscxGmqeZ3mTpQY/i4k2B09mDKtllOAHIln/q1cHMN/TngOZZp6
be7hcehg/qBQ77xB5CnoDSXcyeywBAoz60FKUshwYDq+jASQHdumJnJ4ZgDtHMuikIo6GrKAgVt9
l6tCI/Yup+9ZVW5xzs+t7BezcKDBJpfLSngmDf8G8jp+pBpcpSW5JnhbLC1Q9U6JvEBYkfjbbA27
vlg9j+mktrp3uMAHsc+B7PD1NPZTr5tBrb2WVOXxcmsGn0fmdBxXkogWRYkckg86NPO+2Zkz/w/f
H/tfGtowXJCkTqX5VCuNC9TRuQtTidn1nqDPj0lTL6dxJ95DZkcA0Pwz1h4SZH8XfsH87IAzK01T
x1eufnm6lDzXeL7I8Wkq0/97rOjmFEGsuJZU34ayAFpU8wwyEVcfxuzKvY6NtxoADwC/UVj/pmVn
nf1gGL6dB0Bg0yI6sWp5EuxndMlfheNMHzyCI5hVfWM4THDNn9XXFHyzIfDgP6hTdU9fkiyOljm7
zK9aALwxxy2vEH4I3l4bDvA0bV3yb/tT/Fu/nDyD8R/+gLUOBynQm8KUrzR+pdRu/BUJoxBQWejS
bOGDCqQf/li7pnUOGYZWuL7QVl5WzyPeibsJw1wQUAy4Mc+EFZwWhkNEZoggr24Lu257JImL4eYN
9mU5WVgJ7FCe2ehAeaZ6uJlTT+FmG3CFEU9BLIOlQaEx0D7JVXH1FIsJYSQy2pbLzHr7QtoBH508
V1En0J1xiJFAQTiWXaQ6wLpuk7mdkvlfo7oqNbyhLq3jgHuMtKNhIW0SM6Aq1xA8AL5SAJGJqwN1
jHStM6m4wnkZaRb18W0qmP+5wIkzXG5LDGAO6Hd8yvuqDhnBOfWW/Kxpo7KSMzs6QbOMgCVwtDb2
gRWqsv8EpyxrxkecpzEE5b6c1RwZegkcbvNgTmC8YnS4YoWxVEbfo37EVzhqCRCUjLH15O3ZzHpR
7s7uTAPliX0zVMdROGAubbo3zUbGrwfvPBdz4VdioDlA0CFVYHgZkrsjZ2kyvgZIU7twReyOd8yz
S/C4IrgLowjgZPy2MB8EQx0qSSaunlvoZQ6ns+fUGs1N54SJPLzeM5D7SxT+97D/HGtBuVdiZcwa
dDLSMp8avtvg2M5bKtypujMRtyhv1IuC04wPByS5tGvMAKcDBIkRBONh5hm2Eoy/zoO/eznHmMJ8
MhFEb/mDSSAAZOOk3wCcrr9JwmZQVk4MZarWBhS0FifejzfLVwtU5OL7ElUFEWpTu0rR1d6gGxOF
7WWfSwFHvAhOmSdeV6TQS6dQ/OQPndsj8v8e9WIbTYUS2BStQXnPznqXTb1CFxedJ/2kmvVh0MGa
3vdwFi9JHdPefd0rtFlzhrTdDRdlpcqYTALyNUDVzAMGGKxarOv/CdrfDuyacqej75JztwVwIqe3
p0QeQK01YdWgyGfrYjy9C6/gMMj5t+9FXR7akWSpj4w+9TWcwr6+xifYJmk45ZfPU+hP/w4deIru
rxMijXigOi+xMrL561Fn9RnYIeG/XOjMustPgWbE1SbJqjDiXsZcCE1Ra1gR6TmIR4Hmd5ZId5YT
wh01+SHD1+2prwgX8iAjCPNhths6TsuA3j1iowycpofJIh4JwogbMkmwTRnkgddhJmel3nyCPuO/
CksMGZR5IuNIHhUPUJc1CGXHFQtrhaVzukdNCupyxs6yshx/5lezzQqmusP/j9E6o00anq7gJ47b
IH5E4o1e1RWRIG1Pd6o+Z3W9IfWbL1ULuakdT6B/YkdaaFc5d8rkeX5TuxLEVyRcvzBwFEHllsCu
JWLpG8jU/J1TOa0amRpcqPN0DRxRSKhiSG13dsJyE7ZyT9xBSOUbWCMErc5809XdWHZ6kBPGuFzS
iGk4qLWW7XA2J+KmdV5B6lzGPn/VhUoR8KvbUslpARNfCKqeYm7gzXVK5UI4fDzUJ9jnjsghmJeO
aYKmOpbaZBT/IlL9+QK0Qmsxib3+GQvODkphYr+bmTKshZMQLCLFoT0PMb9hiCUWSwUinvw0St+d
rNKWPMU8tzezJ7gtQSj6hfBalWkMjdQ1DMjgcivWY6IELznbuYXuCecCnxi1VY78R8BuGW2NQzWq
QqpLBUytRMcXvF13H6Ms8Knq06vD2nh2FqwyA3vJ9kg4R9kvWIum2egqsSwmvYZvDtBtnvT1YIM6
5jbllfJsPVeg+xwiKoRPLOUgfBWC7NsiDzj6PbI64+uDxl7d1LWZEpUUMiSMqJzchCWj44TR/lQs
FabfIJu6S0TCL/S8L29WIF2k/qFdBV2K2kq0HSaLtbxTj0lBiDvqNg036MFnC4kAOzxVGzypomtx
yx4AmyU5rwRQ2t6lcvg9g+CzbowdRuLp01cXz/1P/68v3Rf/BwgbIi4mgoPOvgUYH55aX3YaiRfg
NkBT2w9c/qdaHQX75yR+HJe4vSCZXci1QrI8l9f2QAe6guUl3+Lq+USN+kuBLo1JeLo1YUpx7ZwU
JLx4DtQ1x+XcoTcnDHOFRljW6KoZVVVDvuZKaaD6MnNE3f/tkqpwQMaNMbYC5BzkQadX+/nQBG3u
8H/YG8TWB7BnKCCEue8bHEic7HX9TradFEaUGFw+6nNFjKk+pbEmQkbt4FUBmRTHfJy5ANBae9CI
z6HBKZj6iUTmEf2dm6G6RQSwj3RphZH85lsna8sL0pz1pt9yFAkHR8/hb9BoqfIWit9WYGM2q9Yq
VO4b2ErdGzXmNWb1pM1Y137aMd8Vnwr/GzI+s4gcvqJtvO9srngA/qcrso51rObg4nimSKT4WQ2J
RPeqXUBcVl3Lz/18TZa/OD/x4XGqeuOfDUcdiQaogI/3wbR82ReffBci2xEGf4Uw35afTcYdETOa
g6ClBk5nHKIE5sf9IRC50KEkM2pE1p9sRlSTL2ck2lUUQcnrjXQDm9PKltAZatLlW7HkPnbxPuNB
OqR25IgFzVjau/3VmD9dnAE+4x+17La5BbYiFAd3A44JhKediew1ZrLQMq4hdJ8CEvXsM5NqNVwr
cgl1Dv2DNYmnr+BLi8/rZJduePgaNlZc93jVNGEgNvlDKIIEuGmsTY/Fg0Zer/WnD1qTWj8CQMzx
k9NX+8EE221w76z/FypTng4rei7shuDPYjXQRxBRLYQMbMMqlepM+0xdyjM8UM/af4HaPCOBkmGZ
8MTzNNgmHtxu9HyNDTRiiWCLyJGF6ZL260gJWM530zzFFR1wKhVz3UpMOaUePvusCDQAF2OGmz/e
944EBmePNNAvodkens9xNMIm4Z4A5dqEYE8Lc7UI2B4yANC30MRIfN8SPXa8BYpbsGBaYLHFCm3J
IROSjnmTMLBoOP4rhRVvL/6N8513SSQYUp3t6Px771oek8UNKZWmHTIpLII4ksggYR8vRAkQdUiQ
4R9hIgMmSDHVUBz/xx7l2K7fH3yafFPg5rr1D2HDjYw0gPtgQgjeSp7wjQXCZdXcWDrPdmOrJ7w2
XZBTfwSOWxyXrDchjw1KUd+iXeZq5x5xozTCAkoE0FKWe2rNF7lHvkISby3lwz0tjCgtGds83G9d
pRxk6fZ4lU1m9+ZHUsCYOu3j2qenwnj/xS8tNOMzLnqaqV2TEUG3aLObMI/r9bQP3XRzW0HeMT3E
c24gZ9Jcs5Uosg9Tzy4QcTWWrbDHIc+2gU3t2OWlEAF8BuUkPDk3zRqwEQ0sXhllfexICb8rVfSJ
vRIt3hGsW0u8OKR65RwxAcl9FbjobiVjTJKuNogcl2OKmOjgdcL6sH0TFA3euvbwrcBOMrsnam1z
OBWh2j+zoAUVdZOCjjUS3vkDhFmd9yvlYYgHlpgT+Rdt7GZ2cUGPvzU2Ftr3jWtpwlQaVDAOSFla
1PfF6hUyusVJMuAQkyMPUSidNRfR0bXGflDbhfCY0MFHVaprDl53eKtZXL9PGZUDUsEc3WZvEdyX
BjMn2CgPwah4g7bihnt926qg826z5X/6IYAFjPkhrCTSo1G7ZpbzVMtKciwmwsf6HUuFYaMm8vj2
g25qZqC514RuQYh6RI7Xrzbl7/JXvtsAE4n3sZKsNORtJApTv8gJNGMAMRD0uOTVDWVIN2T3zdMw
3Fi4Ol0W0lMvY287yJ1JYirNo9Coc9soKjuAyNreWWGMiSRL0uNjy9r8vBAuaIeS3yODaOiUkfS4
/09/5CxNYTLMBHx0cFxV5s2Fb4TAdqN7kewT9BNeGAF944IyYuCAOFAGsZUIXLj68NuL5sCvGrDr
Nr2p2IDzZF8iMKAs1XlpZdsbOFxLgvFh5386yqbYUZU+D6csllN/2I6hXC5JdfKT9OMg9PvWf5zB
hgqTYwvQoQmHZK+1fHehUC3rtcvzkMcDbHwnOkdT4rNSmIcJ8kVHmBPBHXXSzm6YW01p4JtpUYUt
bKehyTJEf/AWtBjs6cwBE4buuEOku16UUQj+0LKvo4GSW18+K4N4P08C44wx9zbpHzj0Crv3+IJK
bm+gtECb3emueKKPFakr8CCmVucBWC7LwGMiftIkN828Il7/nfotP3pnCP1UxRU4A+d8qCTpywQF
xeu3bWeXhITcFw5y2/RsdHgUz/SSHe4HTHv1ubwqBVk50YYS5w4S7fkOOnSHQLi2aoNlzKsfQPRe
BtHPArQlKEQGkqLUeYxfWht5QI3CC3oMc4vX1CRlnvJQsVhALd/a3D1IfaoTnLsOaptZhtFLsel8
auRWyEBcv8f2exZgSkc9apwecFkFv5IT8zlPDoPCrcNuAFfDgo9xk0w42SAO2ixvnXUgOyRFDe6q
737QbFCBNYJfseWZqQokfLk2GkGI2RtoFt/8o59FJTvYRL1eQVCvBwe78UlcR8CdCdf6C1sFL3Lt
ZsikIiR+1wM/gLFme2ULVtsVGTsaovaix7wLMn5HPcraqm036q/UizpXuuAJjgIqk8HcW3d8DxMk
zA4w4+82iIFOhAKzMUlVMcJvh6KKEioxzKYe8epaKp/TtvvCXJY0jGtAhTxj6AZ+TotcsK+bLlzu
mSHNQHNrsfbcYeySuXoDZO2NNo9ZbeMTJEf8b02IIPpYDW7vr+rxTh23Fr+foIu34sJf6atj4AmU
7hIBGVSg8an+BeulZaTal2wygI461yR79MgLz+G2xC30ztt+sOulSc/5TEOQ1YhVGPOTMyWHknO/
2WRevZfr/bsVpr06A1Ntj0B9wmN2iNHgtVykcHL5/VhZR4oxeCzzfYC3pXKrUaQES41an15L3A10
OlD21n113DVxhCEnR5DKwousAJV72+uZl78l7NFuQRGFteOOsdgO3FDcQGBoSAepTyy1SIzbJU9F
X/tZ/fpl7FvlSs3p/qEQrNCB48f3XWXeGg7MPAYCqYE3IbiRfdxYrn4euAora+1v6w3cnuN00yrA
pHCRDQ/e9YvTV/xNnRrksk0VJVFj9txWiK7rKLZTjCOMBIcY2Xr3tL6/0eCh2IV7kWoh1gLFHy0a
G5tp+AeRriqE/cFOvTPJCHzrhtGzDloN1Wa1qBvKcodWt8eNK7mj+uizRFbXJkcLg4ZE/RBgHYOt
14sx8+wTRFut7nFFshBH/qiJ1/vHLslRxwt1IjyTjeYdBLWuz/uZhUT3zn3w4rOvIkxFT3cAlwXe
0Tdmb8Wrduy3RM6mljSh6t2q1EKpEplMHA4ngaxlXldO0s0U3hxldgZkm4lxtTBhsWAyAsWhG0K6
R9aoWtmEu8e2tYF68K5ICnsPdTlCptdmNBHXw6eUSBaFAMCgTdbBZkH2324Qw9BVM+04lAui3OrY
D8XzFlv/DRGBgOfx8sFmoRHv3iLzed/08b6l5ofy+UdmdlKH10WQK1VvOprs1Ur3FWDsmVmTmxGY
ntpKkN1LakxJcFQlCWfZVp5q6OuA/vLw4t1K9A8pMppwLIP0Yqrv71yPvVfBD4ByCYwyjcw7LUpL
ARqBpXgMjRlWQFQEkGrWBA1abGkGNmaj+hkagRj7gx6Oy+/JV6qp+0d/bJOV+gi9f1tn36D3AhJy
t2UvSrpppxuP6pj6LSOXN1BI/L6mjcVTKfRMMtU/rXQtS7UnE2aH3OC+ERPu15AD63J/dlZCbjob
ZI51Ogcl7BhdPO10hpeF569T0W7LMrsDsKM3WIeqfe+JgmohsGX7aq3wAPf8/C6SHLQOCwCFUysH
7AkVCcDmPEZcCTQ3lqMEMWov6FEqib7teHjGWwWGHTxcYK7bCbf+GyraknHQIQ3hAxlq6vCwkazn
OmkRLBXtH7+g8q2NqRKvrnEUvfChCUY7cqEiPk4abFRR9mNSr/korH0NBH8FvVFBM+VQC2w5HWld
b+4CSgAa59/d/hoAHqL+pYUgT1aKFTL4AKtFCF3CTo+ZOGP/uPNyYjIULE/sz9cfMAEtjQcXxS7H
RIPxZ6OuMswtkqIP4mME00Pm1pK997whgqzsEvM/BCfkXKC+mtYbbhQFrCYM0OZoC6cqqiQV3wbA
Nol+4RSqOUrqtUgOvfhliJEfxCGvOF216QMh4YYXEFXaHiO/uxY5IvL6KZ28nawxUrECZ58c/6OL
vFuF1msSfBAEuwxCR7bgedtmtLElg334DgLP+NfKM1OOzmjwM8lTD2qdyzfdVQ0c05J7bC2yfSSZ
GDsvgzK5YQdQLin3jBrreo+VwAaQA4qoN3CFGR+JnBttZcY8LzAZgYxSGaDotJHGW0mEHdzYn5K7
YAylKG3dwJ8+AdFIHGyMNPzQtwaHflcWk2Zx7Ti8tIT2kn/3SmQ0BmN9GWkoqgaPHahA41DEd5xN
kwqsIgvZo/XvukbQzUs+Cv8r0RBeV2MSY/OnsZxXnzQu9FCYb+ANoEQgE3joVe532IEJgAh14brO
3m0STfiWNwkT4BLedLS7GV3qkcKiA2P/kgsdL0nFBFXXziEMGAZJ6AuiklxW3BwMBaCykycU4tji
FaRUAXWh+RPnG4mkpdP7CtG6MY30kp/X2iIPE+4npCr48PBRwWSv6j8qvi5xMJDSjhqM6hAawdoM
2pm6q7cgm1RX/kMEcCWpPr1ubbjmAgKZPhdpe8z12z+SjwwhYG+s0A3sIeqVW1ja82hk3qobu/86
6+c8MRL7woc+iKpM2Y1c00dA7qJWRNnU7WWR+12rOJaYt7Ex/3WJw5iPpbOumo8/RQRt/jdTNUWN
4PMShb8Ob0urnO+96P4QN6yP2Jg07aMS6gdG5NEjsbFcqZW54MQUB0XGEMD4TAxOe8Sf81sLEEhw
wn2mI58b4u0Yvog4ffXTM78X4mbPbrZ+mL7VAHWL6nii2gstba7rha6KMt+jFAM+G/ETCY9khVcF
xDOOOgr9SmZh0W5R7av1XOAbSzdj6VsYuwiDhWcHFMIiZaX/wKMaVWi+OvbgLXkwRUeRrzYtzK+/
0wOpjI77FbngQlExYj/ZG0PE8tNSD5laGrK7ed1HyjlpXm0G5zaKWhADOMvHxfSEbAstrAKSVmT5
zMWUNDeucz9T9W7Nm9PMaWBF17Offvb2WmrQazdz6sk7bv9d2LjR/7MnSrPedywU5+i1EvjKBLXR
YN6UFQJZUXAfgdLsaA2fdfdg+mkSsk67tND3fGPQmIS+hm9Dbjo7UO5zjH7fFFVs3rr0R2p9SU1W
gEf79bVev0a4QvuQlU/3MfS0VnvrVb2/EliCge6RkEm74jJ5gyR8ukMfMJTUhC5XkW8J/kIGVN1y
l2YYSagZaG9bRzV3mE0CSxKYdtLKA6JrdMffKOlZ9u9WfwQTjSBlZO5JNIGFt8ln1pYiAV6ONLkN
55ba93IsneNRnub2gETRw5ppe1YAzIoCbf5yuffeWf4+4MyEhZi10FYyOzvLrxraiZQr6HL5fwFt
SpDBluo5so3Ovl9flNVF6T5vyYUfQSnO/zpRvrAF61XTolBxLKE6Mu1XYZpJopJuhS2jSLBmpD02
3Ik+LkFVCh3MXY0cjMFRFbhR5OcyVBtThu1yS5+AUUd31rBk4R9fbJZS0Ou3+4gmZBKqgTzERnxC
Wm7kUyWcDSox0J394ozisjVMQkgQYQdluXuORcm16QJ2CEaT3448QXdjOTtJA3nJ0Qeyrpc6e7sk
z6nzPwVKcwkuwVmqo0B39yFDXkuJRLdnOBhidMK6sMKfEBI5FsnYUxRBNg/vlcAAmooLOEOxURby
9DH9HfJPnWJvKo/AeepH9MJcfFfGp0jNk3CHBksnyZSbh75FlGTCXiBR9SSUIT6cRe+XE3s7gKLV
Kh0GZDNlITpySu0cThmvDFNJt0T2xrB/3AO2YAnG68esyBecj3STx9BhntRt00H6WSzeGII5rJoc
ySqH5Mj9YSgZsfQtVq2ijPb16h9eRVSGcxbjXCrYras8B6k2cDUsUW7F1iOi+tmhkpBKlo2q+W3r
bMMnXSMTbfW8GcKsmkC86eXWqC54K3n19gP+pIPlXFoHLlbnhOwQ6UYdnpJJS0LRPH6Y1f1seus8
LtjeGhcVs60CkYg1HVzVlLmvDVdO7CZxAiAPu+EXPgZjOaBOIGy/jWmAiHq6yj9DzAyOwHzWI+wV
9sZINmc9q0f1twHyhc4j6MxsdY0Vmeqys3c4txveU5L4Z5kQcWB9APECP5bhO7hdM6lnCww+x5Dr
COs2BqFKym/LseghpBFp2HKZ56cwJz6o3+EZ5h0s1adFGtbgrzHwtQ6M0w0doaEGi4ui0B360xQE
M1BKdHMt6Lxc8AXIieWzY/YATzpyhclKTFLUgW8A2qKHKGQQgbaDQ9P3WQF7oCQ3CwvRZHTb8q8A
Llb82kIdnlKOM/KUUqx31Ff6pKTLmTrQ6PGMFsNmGU2GECAa1WwOYIc7HQCJuftCNTiJPkB4QuMV
jgKtyVtgWJwkLYjS+ESWBukQ94XSpR4eX2cHi79XkukaOF6jzVbMOjuF5ltSCQmsQinylf9ndFzl
j9INDOzw++uibeCyfSY/4+Hile1a+a3Mh6DMKyiITr75q6KSr4vQFYJ4imy3O5GiJizg85dNo8+z
4m/91ARoPMa86RaCD69GrfgHBQ8Z98gmvUj2TWZy6ODDv0NMksuMqsaS7wRrWM7UdFw1yjPgWqnA
6kxbBuei7TJdznVgN5Db7PEnv8nOT0qZlrcZt028m/rsfHqfzujVCKGFiJw6d+oYFVMT0bKRULHr
Y+aPa9iqruEmnkN3yNa1C/Ef9O2Xh5kKI7nfa1h4DR3qxb9lqdFcwNPsMSIVOp038zoqjMOsV2ie
tWVtq5quO4RrDElJoWN0fogugLg+G8I6yrxZWjlFNCD6zT1Te/vIwTsUueuiUc/VJe8cJPlE34LE
NY54gqmLDiOz6IhG5rSMhREL3etx1kYf+edKqNkuqxZMUSiiEbjyRnKpo5sMXzP78qj9u9efic8b
Nl2sQaZ9B3HRO1r5LJP799ePlK7Qlru1bCorZ7dxkQWgKw5FfQot+JI37ezCRyUA9YsxV0cXlEvO
FBMlWIfw64yw1xtYiFJy6AyLPj4kL5XTA16NMwNz7GvRC8U50BTQNB7Mh9WoTaGn+xPr/nzzuEQ0
tTgLKlHR+G3MtLgifrqAVtMS6N7YXdGRxWunfXHxIdNi7AOm1AKNghyVcVkWFeQKK2QxehvR8rRM
OxMyDQS9i6ZeTFDk5gaJfbcgOqWqvCa/UzgbiVY1tJIpWGZrnvk7xRAlQsVArdef4sHO2MshlvEr
uD29ULMMqmLpz/uCrcHrAVOk70hp5fzS4nzzAIrqzPuJtthznqbFq0+IhFreVS1KgqTYkhZmVigc
rE04mDR29fOthv7dwHlihFi4n+PbKgtz8kzH1dhDBgdnuHhUrQ0jbq+Ke/9d+dF1a6k80hLpBubM
pS5qFbr0sh5L2f2iK29Vs9DyAQyLIEkfePV40fuvv6cq14f+qbgb1ZckLxja42FqNUoOCi+QKd16
h62FQWregMgKowrJbjmkoNp2PgNCpfHAC+4FIhJXvj9VqBBaq7Q2p0xUjRZsNTsRJfHmqpq3fFM2
di5TnN3WiavmE4vPaLfxtQpurQhEutRR+9SlebxMKZXBrOJDLRWuuY5hAy4jCoVciRzgxZlx14XG
L632HRwkww76qbxHIGqSg1bATBOwfxOUqCrIunF2ie7Jl1MZdXL+Tw1X0cEz08oi5oUu1xrOXM2c
eKDTj0KVujvQkzQGqsMmZOIGmD+zvKfPcXtwIHqPpKqOgaKtsi+4yahFuxTUPw+Jxf32/3NRG878
R4leY/L1gXzfrrOqvfTErsCGyWjJLcyyuhPn42NUzKbnQkjif++8G37HRofw5NdgGMmXKeoz1GbO
EwFNaBF1qibCB2ZIR9jhPSbEeE4h7rTCZ184OK/8XqRNjiNx81aV3uYMeAaeQ0CTX/mkOAYY5U+T
ArN/6DTk8lWlXdUuTkOM6Hcjc1Rgl5lzePOtIHB4Gn8rPJ6CQPMB6xg1A6eQVc5WkZtJw4lip91r
fDAA2Ab2+CIPTglva78jlhgFaMHeh/i5ptCc2wv1v83tjRXXfdy91E8HeO92RNvPAtSXgwQtbYK5
Rsy9tXoBP2TCzlf+GOxsCX2TsGmm94H1GXILp2aSK6qgetKSHI3zdi1Y5sSqVFVWyhR2UwTd5niD
4kAfkQ2kG32JxrIM1juwaCLmr0tkfKgTeL6jhWiqH7IOIr79bCe8qEe1qR85s8WHw36S8EopGV5D
K40a891EiCZX/3zjZ6pyqFqpJj+gbrrX0UGuuS3iQEIOvlP6cvLhvDGCr6xaFY49mlM61ZL+MgTi
Kfi07SKC5jfzbAT0pyxpODRkme2f0ygRELdsi+TzbqShbHLv1QaQg40Kg3MENwLC1V1EMh8gWn5F
8DeWe0Yj4qaLONtk8dpGXxF8X+33iUDzMkMQO72Zmz45Ff6cCaL9dUw0mEd4Dz16uOn6ngWdPQse
3ZwLTVMhYC60J1u/5WFdFcMAKoYaWHVd549mtvT6+1k2MYhrXYR9s/FiFe3urKZtZse6zpBIZUAU
fWfw4N9lKH/Sa57Z4+qB0+IlJjGPjMCln5eSpK6mwNRchh12zn4PcPt2wWGp7QjahCTU1XXe1+rB
9r8wKplTA7uRqNLIyBmRh48D6CrP8y3DoT9B7dk9Ig6MQZG9wSwOINAzoUKVayensu7oKBJumLHg
yKVtxHa+8ewWB7ZK9nLAYhoJI5hfp65n6V5HY9BAlJmMcRg5UCsQgEfA5DVhj/VBNdkDq/LT9+se
MkrPMXoPuLAFw+gGo6DZTymMobyhQMJLTezjIi2iboSXGoCsFQ8eAI4nggpRawFsT1mckYEYS9I1
rzIK777z4zE2DFUarE46lIGpj1DS26WYAMLhLtaco1iwSOZer24eg/itgAzblxrzt5Wghwolf/ru
hFzfMR3C72PR9U8roBxRf6ZvrsMsJFVmco1AjHwuLe0r6SD9vJo4998q3j1tOE8SzQpSj/rZlFeB
uUCgUF0ONMhsHo2Q79OrmoTzNRNicWxVg+9rdUYtkmmOezoLx2T1qP8orX992huj4YZUmsntUQMh
4+6VkugM3avZ4XyNeeBLXFBGz15J28/Xz9fIsVeCix6XXFEsPPXq6hmQX1bCf7ZA9jBCT48szerU
bkl38ALFrBRgXnQBGKCaE/TANgaNpcaSNtbWNOVxk0zPTcIdyqzibM9hpc9sGte0KTFKoDTnQG1Y
fRGFIk/05sF8XJo/BajRPbARuQxCOBKgzeHDpOg4FcjFlwyWf1h63YIMCwO4TvfxiZCfkjb9MXjP
0B70GqmeBSxGOdMFoVONS1OdjHgzO6eFhk60OGb6FLoqMZLh/iL3fYiQiG7UjUqtpWHaZHVq0Rda
tfxemeCUYl3OkfPS15G9LrsnxqneT44YX+bxbeqwvMKGl+OQFxb+OkQc1RnHO1b2tsDJ5hhR+OY0
KfYbcbIhc18XcCWj0ClnVWDodk65Pv+rgSXbYbscTluz6sIlwCmphBEqkAsPE4+vxerufZTaZzbf
tL3/gbtPSXJ9uqz1Foqg3AzlrC5NRfUCfSUlQ7XuNMgbKZYA7o3A4veZgmRSwmGDXLsWC0Hn+XIp
NoJqYMnNMxEu/3d0Sj8+ydYc60j71Am6u2wi16CXZzinKJ6NP/xVlOqGFb+zWhBDGwJ8iGZUBb8i
3n/trM9XvJkLuWGX0soD+TqbUtLRYNeD2RjiJGMeJcmKHRAZTYe93BsxY3M67Nhyoz9BRkRzwcPg
38bo8ZLkMa0SASArpjAy/7pCU6A+hd+boUg9yIfCSgBiWz67V8lCH6h11tfvHXQ5cVTgRKxqNAYt
wSAB6RgiaHGuI11+uaPyBXy1a1FvR2BAhyJ8iGCgsK+BofTqq2Iax210bRrmxRFSVMJxkjM2TF57
9fW+sQISkwrzXA8jQFrOnsmQMpaNbD06rQGcVU4jElQDmWeXKTQ12tan7bDWM6EN6VUu371JZ4r5
1siZhYmma1T4DifA1/3pfUSMK2OM8abPqKUnuDvfOj6g7ju5FGxq53jv8/3EEeSeJretBKvCYVZi
tkez4G9B2UICIZq1fO+VcD/cYIr5EW4FsaOaaY/lTl0wveE8otwTcqzlnzag5aVl/J2oNXKswHVW
XYdwBrMIGVj5abH279EsYBfCiNGTVueMMa+EjxMXVOK4HeTBBzVc28ZttoFOTaO2/qoYcx7nJdO1
Fdndte0KMy4R8t2oAu1Tp3Mfz8nBoAQloSIB2HrpNRTGVhBBgFYnU8rwA2OcDqpezwbGKcGYI7o+
gfihTI24Y/yM4hHSJZRRu67ZZg19oUf4edMxBAadkD3dzWRR5qdNXuCmv55StM3G0eDVIDQQE/cw
kBvZHxcHo/Duz2WspzVXtJ2ymMhLJBJDMT6IeeYamAf7CTekR/BPh3+CBinUlyBEZ9A2AVJzRMlq
YU2b3Aka9pSEBCsvN/AEjvmn6XnxqwySJ2437u6UFhWn1bxsny3Sv8IbG3LbjSOtZGoLTEcU3u2z
HDzy3t7yzUHe7e2nTlrk+wlKTMagPEydvoLp0BRIpmsHEKadfduY/6u0j6mTmxj7/D4D3wsD2VmL
wnLBAROuLrnr3tg1nX278HxOd526Uuzn3AkEuNlHp/jSmVl62sRmYxwdetZ0VX1FsVNnZ98k6CS6
GumPBd1qQ+netjv56F6CN2+VHxr/ZGzlm2ejHSoOJFJ1nO0OogukwI92SnlyIe+h4jHkk1OBSVli
gDz1syuMW9useh4rDoTb8NuNhbwWlOgG9SnWtWM19OVTh0WJe+laRo8oxhWXesLQCR/u/gKEve/d
wIsrk09QI6f0QVWnTTSXKnoOoCtN51jQDdMkpE6lJtCp7FMxoDkKfqdPbSFNWJL+K4fEix8YxZdI
M3X5vuJ9k9PnQKD8je82KkhsRhX2WqZqwBmvc8ebIDBfbfeTNuHqxJlYDFgC9TOXPvKz97dsYSY5
7NNqWyP8EmHI2B5zDBjjetAqpTRhZQw5z/SJloLAR5Xbsg7HG7AWk4KQYAK/ZPvbkxxYPg0kDnnl
LbaSYkzD1xQ4G2pk2IuSpS0N0bDTU9YXEHEOzylo07uVEjYmA8ecv6ICjJ5wWOSlGb+hgeOj5ftX
1yad5J/FOK8ih027uAxX9upynIL8UucPzAKgHHN8GmTl/86qN2179Hyr519F6i4kGcU+AV/XZhAA
duELPPgog44UOlWrsTF9sy/B4GKeRDfHYydnZhVd5ErGsW5q3mu8MzLZuzDbyLNVdqISaMw3jFSd
SM+2i1kv/5Rjxc/tJvMo9tTrCCywc0p4fGUPzKIAYKL5z9KWC75q43luGNhn85A7MyL392RrjKF1
TeMYJK0vb5JjHV+VTrCkkXpYgDKw8sJkOj4xeYzIiz8ft/PtkInVAL5okkRPQYDc4iJeqK3rw99+
/qC4uh77au0bTXE3dePcq+m4+EGxXdZKAEMA7Z3Gjw9LyzarOada97qzsSijBq43BhvR7mEsRJ7C
CRVPXjB5b5fvto/GopMJu2e2+pwX1gIX2ErUp2oKC4iutEnJEg+2Wxd10Ntxo5dHGni+vJqKD0wE
mqhsjXHVVn7/Jt5HCT7r/Mm6DTcZW0NmWiAnSLqnN65XrDzZpw3ZfFFqXF+o5Qq02zsGbFaBgbNz
ymr387aTaBb4/y5vOETP3Kt0cILi34et29miqrJN8/vvEbQpy7zwZk8nmPMKJ7/QS0IM3weDLc1C
aVyqLjBoUCitIBniVA6rpBZOboJFg3iVYMtsjQH0MGY+LDQXHH3IbA+SfzHxmU3ceDVR/ztTHBZ1
vDWhKBaR9h/K+v2l9S+9gcNu2alUaqQRYSANxGBShzvgvcH5RyzLKZUFmerYyKTbM4DtNsGvHeBK
3tZGketjT+CWjKhdJiZtNazMWBJSE+FKwY/pA/foWk/5LyqX+X0Zjzoj7OvJUSok2L7dK//k5z21
avTcJhg+06lK01kOnCrDPKVSmTaimGNoqktFWfMJUP5wtTOnbwRudE4u39MTQYvPV4kc1CrN5oKy
YDAM+xaWahJ8L7T4m0K7mt5/WhZ3NAlW2Nlzzfb+w18TnX/kVpnpYnlEzM8rSBi31wklD8tPjUUQ
bZn2mYFsodFy+R53KcWWU4hyydjY6b+u1Nh62uQUMjJLdj3zOrqQuog+YS0g0kBmkP8Lp0v+sof3
kjPy8aWJdo/rHeF9HoaAgjUw+u+pB3CAQch+zPVx6ci91qy0WSgK9FQJQDfd8euPkHxS8gZwhXx1
mflddyhQY5CsNSTRHo3BUBhHf6A3OHqnCf9SYUKOp5iEPovOiedw4YmtIIdLonV1vMBti6oGzK09
ZCNHjPHz3ha/XeU7X0Dgz4lS7Jvpw3/PFOY40XWUBI+/TknlEJy1X//JtilU96hSP/flJRSOPToR
1bog0DgdzzK0stI3xVF5XV0Kj6mZnTxm7P+MT7wgyFHJkhAxPRvtohaQJIXFHIPCJ4GJQgG04SUu
eAwN2PyvJZK48DI3VPwSg+xO8+5qIzQTR4eIuj8Jo5yOHIhiXzS77EGylRvf+2qy4iS2u1HN6UWR
fDzSg7nERvD+KVpUUpz4nQUnBqdsANZ2nmwlMAj5pktZOrJn8yKMSIxkZHRkfu/7H9t7WFCzbtSj
G3lcIU7PXOj1yFNAKJRTMHtz2MWyojbY05sCMJM81nuAtO4mqVNTX3h40lUGojmPdiOCR5fhBVS3
g4NJRBJyKKf8kPMENTPhXe1TiJCx/AJbD3+53vtGDV+xPpgQ/ChU14P0zkaGSXEzgPbF+Bk0hjOz
L7C0z1rp8cwpBlOR1hPhXlexrZKKOaugRWDj85wUmk7mlCd2k3/Xj29LKwm+uzxu78f+SmidyWtO
KpyTFETl+anXNVRV653mI8xHjnamkKuguF5Lz2cRbHVB6s42iJaXKmz9vlS7F9KZ5+3WkpqLc/Z/
/UlZ0LP2vI29Qa7y5hgk0Kw7IkSccgCswhZRTOpLd9Ud2aX3js87nftH8dIdeaV9J7MP8GiEw8NF
QfPr9Dn7KiDKuJRW5COdrreA8spKznl9QnHB83FR7YRrkQ2JgIq49IkomLTbAiT3CWKPb9VefGOp
LrP2IWnp81KilRjod+yi8nAj/BXtYvZurVZtLx/AxCQZ5HWWzbRc0FZURZP4EVusnFMGmmY0geVH
5OIcySGdA9+AMgXo42iYBcZWXHcv1lV/ReWyVdpJ6/XtlzLB6W6CYUsdJi9BEo6W/fW6KarsuCWP
lSLwN6mOSCDjjO1rG+0lhZxxiAfsuqlMkh9TlTdkfTV6MXChVKjyl8ubeXG8SceEEOerRfqaAUwi
RkZr6tEFv3X8rYOuh57A6AmLUwF8Trg9ob9OI8P2bamFAbknz1MruCAnAbQ181XDEeeKAt3zso5Z
u9W3TGY//3ZyX1U0TH5ohsLWRgMBlazh3bZxebEp3s9M8KDup2245Acat0vWGj8FoHpqSnKe1QlO
LNXPeD6CWgK22/TaUF/K0uDc/Q72WJUf31Yg1pZ2egmnO8HFt3IJfrQZ+Vknc16GZBn7YaRMBqNC
w1OzEwOeT8Ns6UPZJZf6oY6AFWLXB0VQjDlhP1+lVp6PQMIFLOLEBUxjDmiDNPRQxXli8QyIRqir
wK6jJPZbk8vcZDYvznI+Or+qUOuqH3JQ7Ddv4czZ4N+ksr/7pZRQJRfR4hZetRYyiCqAhaQOEHqV
/Ng9G14wW+tWUdpHrENLe83aT4+H87Ei3HFhn6wYRu/cwasaXohY/fY/jg7tchJeIGKYrI+T0uCr
RMRzN529a8dQRTjc75cK9BQpFgpGsWuNs6uB7g1ApHvKKwLgl5Kj9H5i2131HZSKyhGv5cEwRsjP
WS2P/YiuD3Qe0XenychHCCYAOCrx/vL6bfoehAEKkAUgcZ9cpxcYohuWuAyemRryno+HS1vIuHK/
EVXbjBFi/uSesM3uIFB9p7Qqa1jIF9JTFe9sT5k8BgTI9oS+sCYmGcq3ftBNC3d0yDEYUBE1Hfin
TSREGVevc1zVT6S0qOZlh9WdzWR0hnZHLnodQ/6mixhsjFFZr026vbJWEIE0HqJAVEvw8B3K+AGp
p1RWbEKkgUzhESTXqNwFfIn393CF8kkBlG3DVsUGh47LedG45XFiasFMUI+Ok7qiuE1A3o6wLoFG
qq/7xEsq6PWAjRM5BoLv9nBYbR+evt0XAWOtVHlijX5nZLMP59TfdF4sLrV24DcwfGCiHGy/faLD
g//V9kTGeBvwAkjiLcuGoruLt1p4ZMpx9j3ckkfQ2Iw6bElLSF6V29ie4eCX3whZaTG6QgT2lIR2
SG30gtivbBHKkb5XGr4Iv+3Ht5KbCeMzTJzuq3wNVPWxbj6msOfvyKsJQVwJlNN0nHdiFMkAtw3w
Maxq8icmhTTnzvkHYnnRd+BTJvqC8zZw5GuDQw+0e1U4adxQpDKmTsP/IdlvBZ1GkVvDXENc9o+T
+8gt2p/hcLFVNNHDjWFgMSQBrfjm2K1Em33ODRSQuDzjVUA/cPH1Z44aWg9YGDBO31yqfVVrKSQb
1l9RIakmUdrBGfWb6usEQg1ENVZqJoCAUIheBYxew+DTl+P6XEkE8VJTfPtn6H31T6R2OKTba2ay
0cMgTOsPdLzrWfayP0w4NoyD7ayZjftJV5ToAn0oFmOb/5g6Aw5ekvtVXnKftZBqh0xgQguaIVWx
l7lY4riybQMwQPndvFAd+9OTcIZrPE90vo22ROIqDc3WuYMWyNxDv4AK9LZ/u6I9apzQWhQg5RWS
gWDkjGlLzJ2g91jBJy/UFJ4u/Qc/sMUNzECqhYHnorNVJ7ElYOypizYTuV9QmttbGznMdNm7nFX3
sZ432HuC98qjAUv8Pmp5lsffQH2gsYd9pQxl7HieyVbtGGv81sPkqB+FZKVM6rFja3OLfu5p3kA2
HjBQNZhqlmB9itonsdhQulNtS2+MNn6JcCO5zc/I05Ch6KYIPFghgTO3Dzyqn6iF2XCYFRpndrTS
0OoGAEW7PlZLDrXmeg1NP0pvc/8GmRiZmMlxZ4kz1ZWvif7667b9G/Qu1VpBSuN79X8jyo/zmr1W
Mys8ZU2MxShq14aYpRTUCg94YmluNJ1YmOsLMC9eKBQtxpdqeEtV3eeF/xFyW4lfpwSCt+W3IAH/
LX8BYmQqYlPiWpHYGsGV3NmZmbVs41cCUqd/9HxYHkVInBZh+KleBwZyLhyjM6H9YIrYfCH7CG9m
Jebv7rFnPqeKzJt7CJIM5pJ0+gGgDiP5Adv9tiCIZqGxoJCklrp6V/IJ+uWQcN54MskBpa0IChss
T5d8I9L4FMGBdL4kgSUjl5NUoVRTnXrg/kOFcSrZwaBAmPovuuvIRnEreRFxDg1e+IhoNPIxZ0sH
t3Xv1h2I4o0uZFFiMamEbdsZH0HV+PEsNATEr5pl8UdBe24q8xUfPtYXIzWBfDpw19PcL91Y9bnV
W8IM3+WGPNEUABcd3p0ZCISE5RwEF1MXMfZjOx4H7ACqv8/ToNPRQjGbPlwICoyXlKweAk9vjNfS
ViVJpm8A01PcVroYXtv4+bnpOymC2O5Ty0IZtB5iz023mzSecRYX/i0EQBVk55z4hJme0KDXgTRU
x7K+RnZpoObWyk0XMENycMt5inbl33wDvQGm0lDWSYcHwqb9wJDQEYCCKvhjW2uPaIlpRcu3x/AJ
JP0ap1mg0/M4J3TKB+KAgMVIbeQkJt2Yn5apWULJlDuzkLEZtyXTOXgRPl40EoYuWepR7IXZc/g+
PHFZN/PbJoUGoL8FvQptkSChp+aM+ofx8s8MI6zMZTwdQjj3is09+9CMQsagyN95xL0IgmO1FwUl
Y57NqGZnPOqGYGrT+CFvhknyIU5WuEMUZ2SV066iseaEd/jLBXKMDJv9hHlt15agKT40RcNdOSXv
izqOhVesZDwPpxnOqkJzmxZJlz4s3i7N53ZVnNqlqI77WTvn2WImiobWi77j4ps1Q7B2PjRiskhD
qexF+hp+9mA1qRyF00AZH1amNWIOr/iL2CUsfJ8m0vzPkYSmTzULJpHo5YZ9+0JjTMNdjszHqnao
Fcr4+SJRLAANpRbgP6/bWdbEtFf+brlr207EtuWfT5w/e/qHaLqB3oHRv384qBhelJQbBv7+CYru
dIorqTjSi6AodOwTkdgNpCa5gFEH89cEWaOXLy8kEA2GcMoA2U+xWfzsjdQdV2bNnj+OSO7cId0c
T6/Wasv7/DfgoDgzIpVbG/b0BruZx+vBHGVLwuakzeFnXBLlN9xqVY4wtS/Yl/bmzl1QiIn0le2T
0AR2opQNdO+d/3Efmn66x0jTmXEzwcYIOJIIpPbDYU8c1hLLInUarR1lv8X2tjFlYRNBAz+BPQuf
mWTMh0YS+8A8+gVDvM2tXMLWowm07ogzEAfjRrEJ8druHJfQRDRTaAuCFtdhF7jqKzMqc+lvEM23
7fDdJO31E5VI4BdzycGy/NRiVvu6S7fztWEzUL1eigZ8OeMas+5rdz4ir7ahMvyXaMf0k+h7U+QC
5zICGYqY5bpT7Buq/7QzIHVzSCn72fw440Tynt+hOnwuEwZ1t8myKsUriHucruCs9ZnvtJ5+eklQ
CI6HQbO8yCMPXaEdWkb6y0QUcpCnBMBncM/a6rfZYWPOF/8bUYr5LU1pYigRZncJ3thfZmnNXktc
+P18BlgVLpJ4MOFrxQqBkAFJ9sOSDsKkymDnhuJSytTPdLrYi4F+mhAbL43XfurxSbIth+J/u1OR
wHdahzr9Rp+t0c6xVGilKbO/JQ1J9HhrIyRENHnimf8hiPdwZZCJHcv7U2fk56NJWjHMa0CTOETa
CWaqlF8UaP0UK6OhqjTO3ID4vTVZKCQ4ngG4kcokNYJWb6moPctcC7HNg8ivyRnJob1pyi+w2Ppb
6utaCvV7JSA747yNJualvaAPF7f0ZeukPH/WZxGpzvhnsjX0osM97x7AgQEkvTySWhjpQBWiUczK
FPhuhgSwGmSh804/eq85TXplZayn/aKPadQAk0q6CuUatpqrnjUZ+rRIsfZ2BEIOxvAJsboQ7UVB
f4hDOrf3M+pfR7XsHiHkt7PdbASuy2lISpVSMa3aFoO7vHnR6rxGDjJv0/g1sk1OMdAqndBHyQSw
DyDYUuI5t/RgXwOmde7Ux8O1577AsFB+4+eVjlZp7sIlGk4IjHwG5vTvJdz8j4v4Yp/XmGtFtxhK
uAkfrsToRqIxt21mbmKQV7V9wS/UWyJ+8+UMh2oHLXv7rDUjeDaUk9xL4CyUJj2nk3F4vQRphp5K
VrZSvvs/nagT3sDVSaMEwmbu9LCBHVecYOWWaGVvNKNnKQk/C+wzFSM8poWa18hAcYoCFIuk8esA
3u9b/ZP+6F4W3K9uC+SX5DaWylLAG2aNKd+7tjPMq+PWPCyjUZGyOQ933qVUibq8ZARyUpiNzSUe
WvTQ3oocS2QbY+Gi1/dchm0rCGBng8QU3fJKWAw0JlVvoMq5JpayoBH8hZHoGiQzqOx/z+6sGekL
j+9jUSrnS2kp/37z5tDcKU3L0ROtxizk3S6EiwQEp6Lq0wO45vLKBBhA8aARFqQqaPwhx13NyptL
Vt8PfAajHXRH/abHaAphyIcP1tlVu+dMn7c5dHa692g5BZhF3x8DlPV7CNYkyUTFg3oSjc/DbSkS
cdUf8dE3LXhv2Xd/h42sVlqxtKhaVP/ZHMehySrEvSB9gsY0IDGs+2PCAMUTzALx3lipROxKuOVm
E3u0/YpLOhsC3H45Gv7xsbRms7aAM+gPY19MgU0cwGjo0XkCdV+8vFIoyLMk3kgjijz7GhSzldc6
gISSFJHzCigAP6E9QHWEL/LlntALAtMcLp+b22U4bHu+HgjgoRd/hAH4o+Jx/DIPsS4i/LnZlYg4
e5aS21pzBh/CQ6xvXPoj7CWvwjgQb5h1ZUn9nyNyZv6ujXUPFS+pod5/WpBZ9JV19zFBEotj1l7j
N/mj96JrE4VI4zknLnGbpY9TUJcaMl9b5BIHFe4IRUr+sd0xrw+nLF0FtMKfHvbLYGs8BaU61Ybu
YUQpJpw+SJEvD67Buh2TIfdRTn7y1LvSD+3YxGWtP81QFwRFHioSgXRtgkrXo5gCl2OL7edquReU
ZkqROhhZprZ0zObj56xH/Tgi32XVTRoK0FSrlUEDkLbDMOxmkNrTu6GQSmu1nkrRftgWbCQLl3PP
w1DBtHcFMDW7u2LLNiDGLVosMTuzxCUElXCpdRRhHxiV6J4WGH+2uR0VCicrCGoJ8LkmSihTta+o
6Dx+WRR0er48fon5g4jAAmFWOzUWLg/Y9uXFikdQol6aBq75O3xWniO+W+Q8MeA2BqcZrvtRv9Qx
mNU5JA8iSEjlO/q0FAJgQf7nqtHUdPnwEr1wy1WL57gqWQFfMzIsX0/7w5tVyz0S5JiaqR1H9aSV
pPI36vaj4vRAP/zyN/fkigjNE5yJ/yvZtHnDeC9xgjpvL55OW+dGFY4GDSA5tk3xEU7cRZXWbAi9
LuFX74R060Qot5g2K2a9EoPYZj+iwaCE2DWVzSYAEe99XZhNxzMn9JtEB9AmElA9Ysz+P1VCZD47
pMBsEUlp+6CfMm32/JVTxYE2PwqoZUGZvw3JTryqGRRM9WEWJiuPbUjF3bdI97zUe1ghZS3YEC58
WKb4dSOuqR4styLBVR1QEfagTzzLSF7hZvA3nMvYa7x6zmiQ5/s8jH2aM8crou32qig6mq6xEiTj
Fd++YZti6AIR5uLxmBwbNP8g0ZcPun/E4Zymvl2voChF0dGPdqwewPHuVAeXRkcuA8pmN8KB6TAq
n2o5IzsRMdHnKRO6E8hsVDKKuI1Hsoh3rTc9Itry0v34BfuO7awoI7kVK4Us24tEfPzcjf2h/W/e
WOUgulHvDX6YSY8GBEKZoQdjsY8WIaX+qNQavr9fGSpqedSbVNMcaAlkrZcLi22mkSO2bCY4fPfN
x79fChFhlnJZm/+OgEkESxmA0KRAekffK7/QKctqutEzqYcyN7iHWLYyhdT/pYDtAdwM1xme1tXo
6JZqHRC75mY/R9yyWfnZIyyI5on/juodMVgavxaKbw1MEJIR5Xeg+5F3rX8ovZ4Pqf5P8AOvtne+
d79jWS8OUD6RLqwJc7lYhC+4k1452ZpBZU3PBdlP/1D1TSAEOnkZjB/KPFM+9yPtY9eC+25gqbcN
u2y6EWbSpgf05bZx7xGiQ8+mqKNcL6h+MU8yZ/2S7MYUCHb4BQJpuE55TA3wq211BUQG6ak+FqaO
RqmDQf7E9sXU57IrfTKYnCNmT86qKn4lZecm06mkqAQAraKKnteM3n4RkBVAMTRYPanouRlf41wW
5C4Fi5jzprrhdRSmHRTs88nR+NArUN41KmSiwcSRuwwX7ru52iQp36ESyZ8173GCkE1oW0sSbNgU
RwRJ8A0gBs9/ccg350sDU+8rm4MAmB0wDhI/LG0GxE2wVwDtMahmRYD7MHjL4KHa8ZVUGVrFLg3G
ufM6FwZYkkoEf9Bnns7WT6HcHIBu8gpzQpkCw3+xghdVRNidXUWcdZE5lADz6luIsvSVLdDjw4Fs
E7DsybuJgJeyfHtkSAPBaeq+6gp2JXbKSzNo83i/Pa5nuwKqclzXN6lXhLory3gqvDTSPjWONQw+
x44XsEL93kaBU8H5mAaQpL7swZiI+hOMUPJzuGBimQnBTEJe77aeLfZBVPvJcfMyb8FbuXZozfCf
8QtTyESMNeSeSYOQSyRV9PT182cGoxsqN/WlxKHZdETkTqTmjIkA5btGqP55JQiC+Rz6ekXP8vkG
Hx1qe/fXM7O/LtCtrpsDl1wOjoCQreTfEIRoBYOMip3Lm2P2jX3PUdy7jeMdEVF//+BXVFOHlOad
igjbR67ipSwty6nC7zkYT9qskA8WuW3n1EOhKF6vta3PwdaXaUQn+klAnjQgzOJbm+Ti3HHTLtTs
mCZv5gEoh1RKp05Agejc1KCluT0Dhk4xpOvqTj71HeB1QRWmjOl78cjy8FKaStMssTuCdN62HmwB
lx6iw7lrvxq2qI7DrHaN7t+KhN4gS4TvbH/9sTaSPYPngd4pguN+XO2E0gNSEKCO2HDU4xTSltyE
n5pY/VExH+/tMAyDWXL1fkdhhf9q66LL38BO9aUX4pVEJ8FK6S/EMWWcqjAHMlxkZ5uATJsYxHC3
s6pndw4lg5pLsIoobJdXOc0fB/7h4mCuo3/zj0vE+vcCqpnOmErOOaJC2ktYdUegz73Hh5ftwaMi
DIFV7Ku5jV6Ya4+e6t/ZsClEZ5Hp3t4d1IpWtiVm7A8i9BBTZq7cYmkssBkVtEbrEBrliK9Ni00e
DYW7gTtdlskUNTwxEzwk3qb0ud/QKVUDbrghcMHfjexkBBaySrS6cayRitCfijvQxAumH2eqXajc
h6AiJomtJKk4qg1aIc0e04So0tg4Go1DQv+vOM4CG+6pQ+HsBrimynyeLfOpApFivjc9/LsjeR3Y
4l50mHRoIHCUPM+VPx+oBaWh/fMpuEFCzdIurKkWUneHBdJGfvPIH+oviu5Un4oiaI2aVobHhB31
N4T0qFkz7pEtujq0/6gsRG4xqTjPGCCEe1U0mDFswFDnDJLzC3jctOS4MJX+IbWqaYsFrKHP3i6K
Nb9lo+uIthEDAvCdbFMTbzfe+GQZkpvydBX06MqZUB3OtEZP3Xv/HDU9e1fLcoxsZAGpGfqflWIq
v5kvzXoFPswQ15v2eRwyV7HSw55YJTxVyGy5WyG5Xj+csuH9/pXF6Q/kt3iwnn08ireDCLHiYK69
ozBrZCoopRqVKXLx1rA535IVeH3n1fMllq5Dp7UCYv5+HA2pHPg3D3MM1XqWvhIPcZb1IGvzbDmD
HO+C4Y03qa+SgyleavKw8NA2f6cfkb1xI+m3eIiplSBXDzP8axlxlM5hlxdr6ADGPb20aGJoG5yT
QJ1imz95QR7X9gUF9X+45PsASKok/H3gCq80i3gEifSqZBAgpS3DV2CQNSEzdGjbdnrTcnxWhJpO
M5H9rR4iioXqdFYn+NV4kR25cNAP+/47Vs+oyZOLQH7nnSePITMD3nyyf+777GWVrZFwt2WDX5JZ
8PxTctOd8OrCbb+brd1P9YBIoQunCRpziiGt4rUcXcKlPZ/lP6s7aZxi+fezf9a/5Ij22M5C0YEn
uIasbK+avjU7FRWQL8RtHsGCwpdQiwsq1YNE1djpvlyiD9fUJCQecZjDG7oqqCWynsSI9MH3810t
2PiAy3h019vpFtRnqL4zkTq3nCo+G3YCeiyjDlLQ8MO+REkQZkTSQudusHahqufiU4V+j60WKznM
xAs2+9Dm4CwkIp7oQFvxZg8eCKS4ZrtHSqnccNhv88je1I3ufIBBAGoOhT7HePokQf02JnOqZ1CT
dmn8MuY9aQAC0NT6x6lzt5UpM68yCb7y7OstBZeikXycu+ciPj+P12y4tPYotQ5uiBcmQd4W+8Ns
aoATLsUKDXNOgXZ1NxX1U8xeziuYlu/wml48XtOEed/8Po/iJzrLDSSVKGmJhEmX3ui0AvEYRoXT
MxRix5r8iN//YSmxsRxduO0VL8lvBLtWcv900l9qz71KZ8r0gqKiH7ycYXFojxKaMLuWtGzz5aTq
Cc0jkDdOGW/VTolauhaIVfYN3JCFmGz8HzEYGagpy3C7OVUnmIgCCs5oWd/rYKvhy68xewNbJcKJ
ZqXBtIsnaIfNLX0OxX9fgcDWMi3lnU0UQj6Jo0f+wyWZoOZ8u9S3p0MqjO8hBWt99r02LvG+4GQ3
IZC/c6zJr03rlMby1RcDYnRJMoIkN2eOteaBuT4xb6TRNSl2VXEGaE58k2l+lfmwB7sqJtK9IvWO
syoii3YT6bxG7ktn/Kn8kUT3UDc3rOQo0It7O96bsaH3tSP7IxDawKZ+MK4dHaUuEqMPNjvq9BfG
9P1iJK5dhRpFtyNBZHtB0NJFiBddMwezPh8ngjyqAGQ9sUMRLIc4+gzOv8wXzv18T1ZKnVP6DF0U
ENOjoea5kxuaHolfSssl1yYPQv61iB7AVUDE+ljuwOcgQO2yq44tFD6B9Nj/zPuUZmZAcB8nBOGe
PX+MH8F+/34BccX0CFISX1KHwRGj3AcOR6ADKUkw/YisffYywd3wBArpirLvu5Q/LLX/rXrYOLUM
nw/MtRWwg8jMnWUwQl7vVmMiD8zEREiAD7q1Z1/eWINtdam1PtK0qbBihnn/Q8MVqIZffa7Mv6Uo
vvMkMrDdY8OR6PRGzfMb4E0VYs6Rs6Bsq6Ep9zRlwQ2dxuc7BpjZz/bN9FMPCirZAn38QCqGid3+
+invileBgMKbGN+Gk10J6Kbe5wJxxDPhbUlPmXanwqEI83+bQ3OF+Dpmp/hdAY0oAbVsjexzRwiR
9/jJNmc8QuV/quicd6gUdrXSKzsj8QcF2Q7dBTIqPQlvwCWqGpnXPMwKlUe+UifR4wHxkXZ0/up8
45pIeyIU/9cFluByc20r7wn7yPCI6UzvGA74mTYBuAylW5/+9QXBhfS2PYg/GPyR9BAvpNwvn3rB
OjYq9cYvD53ALGgGpBzMbPB1ZPWfdgYQG0nlef+T0BxNLgXDo1K2hN5I52YqU55Kg6l5agxLrUOu
wHapc4cERvl7StncW9Js4t1hNSVEt1ep6sNFYdpt8iUZ0JJeKV/Yx6GKgHQ2Fdva18FpEv1H/v5/
qe6FJsv1oY5JdkWWFAi1S5KhfRifT7GLFnLA5uje38gkC/8P4aM9MhsUdxUPU+9mQno1GEwmu8sn
XgV+01yiRJcUiIJ7civiazmLX05PrvRCqa8qJ/Ue11juAPueTFKN9HtbJNjscs0ZGJQUD3mchET4
hmyaPpTGEPEwLqjwAbOjJqqKFsuYw+7V6OsfitlLwHUC+glnXhVu2LUt8/Q37UsuHCki43hrEp56
pX3V7Vg6Q+UsaCP3qajlOd5DbeW4kIVWGkRyevHjtmdGdvcPPw4+7onMZ6d7ykzG3ao4lz4sTwvR
6WMYkQ3+2lUh2u+q98BIb9qAjR9jlkk6fYRBjZHXeudeYpGjsrVWYWWV0yJwJ2XU9KYXGzz2zB7R
lteUTx7/cBoPrg/mgtTxVL6flqLjycgdI3jHRWCVz0WHHH5YRYuka9nJf2QqtYb7w6POEf3sYlw8
uWYPs0oLpRlRkSzAvqrvrlyxww7+DkUxov1gMaq6PgFm8hliSAbt+qhsO9wQQMQb8Dq+5PdqvHR6
uH9E7uBt+ld3SfQss+Z0Fjwt4EIdzEsliuIiFzos/v58iKZA15q3fnEvbb9gmAy/z3WfRcbzpB8L
FOj4/z+W4JiUo0vFdeNdteS3CR8Iwmo4MFwq2EPbN2v9e+NphD4JQaUCEM9eNW0uk8ZRRFinjVFb
3s+I8an2vQMPDFIUMF0W3inqY1c/D41OkTOB3WLgM4kG27TVZjATPkKFntQQQ2N7isizy8u9yOhw
UTc1MQ1f72g3/X9swh+NIjHWPsJITtxJblixTDFlEdhhrw5jv05WkkOaDZKpxOUs/x3agFhhICxH
AdEmXdRJaPVr/Fp5MWx/G+NbCbhfsH6Ij/5UB0IVlrGHfBDhTgs86+AcAUDZAwuEnZILXo9rGV1T
fuNJA++AnHCmeGeTzsvJbfVeM5P1ngLLOhsAyaGW3be0I1C/vuSuMCcYtDvb1GsW4Sq86FNxS1DW
NgSTXQV+4JhPsG9akN7kXK6N3E4AZ4ZU3WIMwBieCrM8PBVYrXuDkUivt0Iu+BDWHT48sq5zsLXt
I5GzEIhodatLNdR4eKU0VsxHv14uieFNGfp9omxSe4xYsbV+GEB0iXi5ONXzh9ZtmJulJABFJGWR
Dv8mvW9xnf5T85d0AXfOuG/L4g+zIHBFyGHxCJH/Mv/aOJKPAwtV0a9Obxt3gt92Sjep+ARTNOvg
aFKh6WogF6s3RX1g6RhH6RPChCCuKM13sMciK4hiooLeSQ1r2jQtMlIbz+h+MeqvfpdUMY95u3C2
vjGFcpB/46Qv+Jg88H+HSLAxlP0b9UrVzC6pFEMGPa63RvxTIhWHYX5Fow/4dJq8UPvBzvMvuqWl
/A7jOJed+TRBHkvX44h8IwG8PL4LoipOnxNAqNxcO/IwNnNMDCGhwrnJlTzCGFFcyt/BkE92mGdy
sRDvvtaERmfVMcyYjI7kDkeP8I6B1tIiwj9+L86qC4fv6NPTlFk4gvcQXhsaAPb6z6Kwp4t69leL
QQj82jggHoefN1D1ik9Oczu5weaC3d7a0FE/G++uIzsSsYVEVp9alghybY0MfbbzyTzQlZ6X22As
0c94ySIXlBkpiZyNedHH3905NaDg3ZOjzqkqN5ZUTKzRfIxBWrOCTr6+0MUxOdh9oQ/66PUTaPra
WxC1JW1XYX7HvFvo0mUZjr+BRvappPBCbgv7pOnNnQ5WCJvgKwJE2t1G96QPs5TBdF3thfCYi4Kv
v3t7D9bIxnXVHf7ZyKFL7y8nzDinUsG/uJ9LBpL9Lsh+byy+niA4CB5ff4A+NqLt3GeuwV7irjZ0
fBjqiKdC0LcqG/UAwl3UXrxKSkWNHdyxJm7+uoPbAFLGVS61uVRo1OadOTkAy1H9l5QWv71uP8iD
Citf47kEKdEIINBgIzSdM36mbESV2W8K8T+e6F06HKgG24T7WpcBd2hOBnW6KR41/np7oFJY8BaE
QtfPo6ANTlOybHsigf160QNYvESbiCIzLC5oEuvtcEnuQCeXoTPBrSHpfkoTlfm31N7q6We+wWuE
9LhqvGvCjEn3OGKPT7Xa3gSU6La3ftEUEVg+/becXoRdXTOzXVJTByhkRbZ8OILIWMbPdUCoH8wO
lDA6OorrXEk+CYwMN7JFgUHsfqobrPDxn7vJs6SmLqrUjXdnhU/RjxDiiu1AneIojp7NmwvA6FDt
1Puu9AQen0Jy+crl5nBlEOEpZ7OdGf+729yg/2VCh41tZW4cuci3BwHXpm00LsD9qBU4+bZSzGTx
ztJDD+DAmVOsJhfBRYOVUK96h/JDDdlX7k/MPbOVSMubw4dQm/23MKTDMsUx/b53T2TuKIKe7gun
HdQivsSmR+/0qT+Xx6Rvp3lfUC9pQStx+njyskp/Gz8ibe8XoymbGf4SXt7Ubf1jfeTbJlYMpAex
7IZrqo9vglnfD+I0bHeCrOwaBvgSln9myZ5F5GNq1One51Rr1BEURxqZpkYstVrs1eGIDEyMcALY
PIy1FrnjOCs76D1tN53ojPnPbLS7j6zm620vYHqY1B6czT2mudaCt3oCIGntcsK2t3jGHr9zTrKO
jW/G3lS4uPdJCoYnGBNQ+o1F8wzFmLvKCkSJdeVFl1AA0K7O+rSBDVI556D7z9PrhrfSlHialRAK
DR180jo0mNjydA/X+R3lPOfXnMpWq29fxsLLshWEfSqO0K3z4dd/7y//LONbDwkdWuLA27E643aZ
Tk2SnHpkBgY3K4vxVocCjqd3lEszQjDRy1+DReIsDbmZjQadatHdWLpNwxNdwDFtjCArNAi9EeHP
56f7XQGEWixFpNQyViGY8G8ks+bRwsJeo0iiH3Q1QvM6iMYj1sjyJO0KLnu0jCZQie3/a7TI5Zr7
WElIDCSMEfSeZM8gx1ilI7DcqqV6ekyK/ACiwyRSL0HDzbY5cvQGABii7NLgnkiBKr+taRK3qdg1
5GEWbrb2Mekn6o9HzLLKhdpgGP/OfP8g9yVnWWIu/50Feqy7tbbqzh7E3aeNemoKHfmJqrY4hzns
NNOhDBw37H996YUwpcN/S1R5/9EQq6Rsq7/Vx6he7DYkYiQvD+ojZhVpDgIBh0Cfl4E/S5fsWxM1
Rd5nMtIb3Lv85ppXlbSI2aISqkrZV6SvDX/t8Sp2zOlXzl9Y5kmgKQFYJRYJ4g7TbTwCXWlCvnnc
nELNebN7DQs548RI4q3LqTuQpymWHlgo+l8WIJ1IOeFtNhR+xIAHaEApGw0Ew/dMaepKZFxdCOIk
2I652RwnK2rmtLU0VnpTmpoQ5HhDVcnkPn4XGO/iJfZZcIT/XvS4Z1MznGUI9tl7Sqw27XEyTcVP
jpbM73xo+8RN9pTbAoytOXa1o7ZQQms0jtm+YO8rtmGEBWMRFlYoid/dnnXBinr/4zIbAFQ3GmQW
th+BMoBmD1sm+Ks+vkwTI7/7o1UA4ACaqPcBZsZv0MV/c7/KojZvVBt5/KEVN5efj0uaCud2qGOg
NXFdkI/3l5oQCYacwpYVHNQMOreV0yBWGQA6f7X+IKeuxgIwgRYJ6X8vdp6s44zN/mrYnJHGzbLg
0wfG0p3yY3Jl+PccnYS1AWQtQqw1p+sWEOm40lQ800v/GOpBY5q6NOnFwc0mYZLBcS2p6Y762RBb
hYk3FzDMpmaofwGHDeyCBJEtegN8julraV1+yls3kcR2FLB2Q4OTSeigBBgz6v52dz7YRdzdfOc6
trFVU6RkC6e91gksEIdxhuvCx8jmmGCoab0kMOv7FzM4w+SIJtnoV169nXW6EoFdrVASSHuEuOoi
PbIuManumvPiCB1WeD1CkZ9B1O4lpxajPlKMQPQWZD+HX3DjfQrlMVVHr4/Gt/pX4I4i56nOQ413
hcFNzmVmQJcF+prO1r3DI8b82sIRHa9FRDginrwcdwVyfIdzg+h1uFXyWOAEzFRRkBswwvFEh7rB
AnlE1Gix+262dnY+Rtrzbc8pwuwXmDvvGvWjFZvQmYgyYqpWvTVXDvLE8dVxY99Ly5kcFc7OQ/JL
j4RxWMA3IJyewgYRzFOcUmYStHQSRZcSy/TrKbHMP0h1CVgJxvbyksA59opXmjBW/p4MBdgv74Z2
pFuKJD+wcpguT3EviPmMyX7Rn4HvfEVL/zKlzp2pX5J2ooTPXcSPds//+Uq928/v0TGZa7kI0jCx
FcueaJQuFnVIVSWHzigE/b1002/9e0BMNy1nRrdA8ar9IWISaG42XzEOB/jJOFq/4YFcMuFJWyfD
OZW95OCwqqH8N3vJ2P0o2r3pVVA+Qmzxg0yVsp82PYd5pC03cTXk+Hj6ZWgXg7EFbZkY0nmaAWew
zSL+ELen8c+7pYhIXFl3yKkrD4VhNcTxuF35VcysmSR8wPvCNivv9+sjdtmcDnM/EJb/zITagR4Q
Ow7ibSkePvj3qld5k8qsnIdfsAOh5kI5TNTwKZ+k/w4+7ADUAzNn0oNygJhPaj7iLLgc39jjTKUA
ethyY3qLv8y0hqBUvSbhQvSBd5bkUBelhoUcscG3kSYqIJHEckCOoWZrrVE4z3KGLt3HH0Dxaz9C
t4YMhoDnfzK1npy0hQROvuVHsAk3jeZKVeLZy4kHBKn6seS0d2zFyq4PlZUvOvnNRK/QfTZlRIPd
ed9Of3/mtFWhIeJIdF597QzZFxr9hw2eiuKUl1dH1SDoQm+ai8+qAUBbvWgCnq3vW5m/JTCVkNpI
BQRATY6cyeMBoXrf0cdsH5fbxxA1CNIPk2X7qUWptyiWu9DGr5xLHP6MXAXWsccLsD8GvKUrQwSk
/MKE+oWjT7jgFEQW9OCD4xO4lQdusOjs+QcHZKp03WROznd+7E8GGGjmqNQDNqVCzWnY2x1b+qhV
audUbLVtxjgpHMwdcMSkQeXVqmlt+7SteWnIcksuwN7IbYcTg5Zs33s+RWzT3mWfNGjTZyRL/Y/P
uhfB1R9/Oh1anonoSgBXYJiq57jskDPBlf2k4h465b83LS7+FsHOaLLTY+FBv2I8O8ZKPCUlkbOa
ovF2P/iVwiRSvOsCOi8ogFVkr25lX7DvrVRw3Wxre9LrQGmzHZsJy+vHdBXpWYaC+amtebJEiCke
zTTwG3mV07Fat5MrefK0mpcK0+TacYPIgLPV7lFR+sONPm5F58r7FXkdVisGiwIJsRifQerJ7vfz
A4WTBlu45xB77LeNo7qVcZCIRChU6e3wLdhjqsJ3auzcJ0/wxdK1eb0ckFO5rdE7U9HmQpd0hnz9
gNm9Sakux36bXH2NdLbXBukCZVzQlHr852ypbeCvDiT/KrBtFV5uLhkQYrI/Ng2qtECXw7Cs+tnm
YfgzAkaaJLPQ8T/QMAxo0vT9pw4HU4xBZ4oUGM/TIuKps90WkxIwwTcJKo0YxYdNXIQoe9wRHiKa
AgPC3fT4woH8NL0s1Bwt79xKi0Keo/XDi11V99+GEDj9hJFnoqQbFNP3OrelBrVF18aLbhbFcSJR
Psu2qB/kXIvTrqob7x3BqVY35fSvNWj0GO8EF9doErhSCjFcn01o+utiVffVfGbwtOH3oDr+akWb
nMUEZKTErZJfU/RpkISvjbDsRirP9S8SQrlt8u/Ka/PnzHHAj+2r2SrqnCrxeFBFiZGxKq6mdDXO
ul0i+a3QoFj0eegX9mYZMR7uaAQgSCESJIvy23yEPFt/6oIrQIvgMli20KmWRA36t6N2d6lkKvFc
0QriLGJOF9CnQRjWP0/KFtCmCLymEjEFXcCWkL8vc+cmKf3buzhqz0hH+ExIsQANrq7vWGTKCDQh
CBDajyK3frwJLRvBduOLZVtlzB6LHQ6JshwgC3zq5+BiB98TjYZE16ZLQWVWRQbB61Dz65Lwq90M
Og3eccgb7zKcfFOwTcsBrYnjrNbhTdi5W/jFcbVUoI1CEB2Jpp0qCvyEvnD4IdzTzXiD2giUMEuL
EiNbtKtjZKeyBLegwUQlWMdyq9anhbDpNUcJhMCWudPRyXtRa27/sii6cew7FALW2weRWbrMiXMG
4L5WHQzmPW8mmwHNMm69w9IctsWv8UeNv5X7qlccTkC+pLN9263P04U25Z1jfjsPegnKvoDa/x+S
YROZYJedfDjaHMn844br/7SYknDdt6/RdwrabbGQeN+F0drlESJjCEA86Aqxz0vd+QGx9SBd9vdk
5NaAf/zWqs9ZncJFamtn0szgF3PR9Ix2vsFwyt02JilA9fYpw8yFMCZ2b7QFf8y7aBZjdc3XgLO/
UvWImbp0BK1b4eLwXlKubJHwxYfU3cRBGlXBI7Xr6TtTVlEP7CuDm2qbC9ya2uaz/b9/toabs0yb
PDeFJlAk2xZPE3+2hU+1V1dTIsncIDk0dNOf+kRqdkjNEsbVhP8BXjHHMlPzyf2Ie7XdotM95urd
ZSCIH8Kw1hMfUcMdOBNkpVUfjA8Yn+dU0S4rGjws9CdTt8dYAqC4cmyGj0xH4GxSJomjzbpQdD+u
oUrT+QkbxoDq4hIAiyHaP6fs5Ne/ZsWGezy4o77//ELLqUsXXEBfhaXqLBmHPD/U3PnCbJgcB6EL
O+0+DIheqM2m5S4Gypz7XHMTDhYAw6KFCApAINnFBbaRtCcD5D8WbP00onNm/w/uaMY07SbbGHPQ
PNp5JsxTiuZsL69ylDme3vsyjR4HwgEyeTgK54DIaSkQbWBSt7hoMtlvsfde2SFR512NJ80l0W2x
3ZVKYzCB9LrqhUrALQ2F1eUChy6PVoCZS29EgsEE7SaP4CkI11O57Jnftte0dT009VqOajgXgQ3d
wFPfXM9CXkXzbKJVzLgU9doI3NYUiJq/AC49r4GElra1bE6+o8wTc3gkxJUA54Z1Jgu4vHsqoQiF
foP09zhXxR7XrRO7K7+eAFO2k1UUMnU7SjwF6jWAKvkIjlYOxjx016DXgebQitAXBmu/EzZxRvtL
zf1u8rVrQdnOd1CAKXUl7V9BhBAQBQh5PPFjCLX2v0wa2nM90x1qsXztrJHCcl6PxTnwShKnTQgf
DBCEPwjA+/Mzk7/UH4YdUpyLUBNLRlkJVCCcczCwhwU/H43ghpJLXvcuqP+Nde+LANzsL7VlmkRj
ehfdVWpVBz5lVNzsk/LxaGEgCBSzoZbp+K5flbzrTYXd7LnXc7itYKtt8YK3t93GWafnyzlrCMo+
20or67+bC/+DXugrYAqFQTJVa8qOApMYQY6xYMrnCfYqxFwKtylqntDoR8eo4ya38bu46DE6i0LK
3OdsW7EITeg5CnOvbRpHZTbcm1E3PdFB1nynpt04PQEgE5e6VB90RAyS0ZWVQMHvn15dY+P5RPB7
bBbcxKI33NWXPCJKkPPr/MoJxjZ5Dgq2NZJRtiGqHu4x1HEINV5aGNg/wHuDlE4OqCactD90vsHV
+Vgp+kke/45Mcr6liMpHWC+BHsVbQ0OmdCKLKkTBBCQJ/P/PVhrY1r/0LtuVjYWKwK4FlPsN+Xw0
gagpJkzGEGzLLmZq38trScyofDrDIsXVF9YVPxmWwH3NMCTYYNpILpZBQC6HsCFN7kCKssIzaqQ1
z6Quw6aJrACTS3k7NPB/7yFs8dGNUBQ4IUIkETSTcqXHqKekFyzdKDu/7XTeistUAgRlhqztwHPb
jsvz+NRNYpcLHQv/PLgW0PrJCEayg5Dug4/hOu/7+Ti5XDODw3D7RFVPg4f5FD0fKQ+1uOEKozM7
+IWhhjaM+NNsNkeqyXIhMd13RqnDtKSojKcv5RmsLu/c0ZHoycNePaqYkUortanSPTGkSYn72Wkq
lWvOWMfyakKNy+OfF49u8X3L8IRpnagRGLb95aXfyjLEZTr8k1lBCOOyWRz59w5P5q9NAvbtxC+e
NDkcf5JO6N9yPkqBRT0mhijy6KZTpT5l6ytpeDZYAK5xEmnPGf12X9UE6Ru/RdjuU5Z2Q4JQt3XO
oa+4Do7+1UFKJFPwGxq0TLwg0FjndP+JQp8AIYfc5MTZrUHd8NAkF7JF+W9IhmPsmD2HhRGRu4hd
a/biGMVNwcrUNioTa6QvwdBJRekvtniFkcCw05ak0Tf9NTbMIcKiBjWOrKDh9d6e5ZKmVhpdpw2A
wJbpc9n/5kWFq65R5ouxYzhYbkjgpqUcNUim6R9mV6sGd8D5N5ELlywgk/m9S28bRlgEb8ObT5wu
NiAm9TDTREdYeFJT8TjjeLXDdlT1r2IUdEQjjs00wSRCMSEwDRKp+iDVEazQ5JHEQqZwZSeSiZ+y
837IZ4AfyKJwoML5NpqUh5mPlQGh01Rr5jsgjzERnHeMMDIQY0vIZLBsaq2x/dm17VI/f4yhIB+e
pABnLqX6BHUaz9w0YF5NDZtMVdQz4Hwkv5uRE3DEFkHPCNXOiJRviNH5yYt8KeQYkaG0gHccPxh8
s1bY3tY6MNULVCbyauioPO16MvxMHgJpYtOo0A5/rCaT0KdpHQhQ/5lByCsRNOfyvBr57U77OATN
+cUD967hFl9ttzmwWiJl3pDeFcULbWefVLnr1yPD4JNC6+M61p0cnSmjm76BshaNtj3anQPMs4ku
uUSrtTU1+a6cLnN+HgHnX8ayJFbj+44qpNZ82xgQfr0Zn9OM3kGx5Ni/pdXxVCeIWQXPn1jJLVNe
NNQ73JVwHYXu2pNxqLPTyih/Yr5j7BQXAK3aEfDoHhdzWOsd5j3QYLoFEOPnbwm+SUkp2ssGNRZD
nGpdH3+6k1boqq+wYgzRfGDHBB/7/J3FXBaKE279Aubw9Sa83u2crEzqcRgb2ITbgqFXkB7rqK1E
USvGU1yo+JWs/rKjWq1kqNS8rWAdgL9YaFrJqD1Ns0LRJRoqqSrEzbrmi8UmHe+1NsjXV9d4C0TF
cnLoWN3+UkNNEYNwgr7AnOlGuuzs5LHAoUmZcJDGIpxL7cuo5k2U0grfyFQNKj755fhefShLX8EB
UjhhJZBG6Ip780MijLRCi8fX9S13uLeRudFQkaUXEerGGbk4m2RAntFqU4DVl75O54ZiMSB9jalW
YDGJLSQBWZE5vglSoFxKTatR4mf84Bic+p2rBRMQxY1RfP1xI6rFv3bk1X768SM4eGeBp9XsHaYa
MfaBYtshS7hkMmvq7S0Ej5WrhDU58e5YeSNL0qBOB+6KEQeYac0rTPOCGBLTSfvG0CGb3Mna6zeu
exeLlDdl6vO3jSTJ8siOipUBk4VDvXmoR3ZiGEixYfM7QNap/Hs5ZM7drECiIil+fIfetofBLWJc
OshcPbP/Kc8dqyfd2mQDCMkriNRmoVIlQiT3qp4kDBYQkDeBq/N/dfRurCa42uUmBBEoy6iwDLZM
8Nc48qYJdtaZRVa3ErEXBhTnqjPh5p8bm+kkfmC2UFaJQm1xF51ZizGYpxMX9prWV0oqopKQ+Ja/
V17FKAcYJDIVhzXmZocXC5r2Om5XTTGUbSAa8qsCdY+5epKst7Ucs0Dm3dcV+UsGBlR39Jh8BySo
kqHhYw6ahSLFGkSiwE8Dd+Er+62ZpVaPYy4YMKrAeAvPOclu+QLyQg4LQuoxMxlkyklRDSNSunGf
4Wpd7pqF7OmfcxfAKAHOd4NgGU03Byp0gfqZQCPVASt5L+dK6xjS5Qra41OWrWUdatO79/7ASvcs
jtIMvSNpVN224dAseYWjMTkPutgrQFfSUpepuJzUQmX5Ll7aGpLPeu+Bl3QZTTVOi5E2c2+XuBpm
YQ37OMJKZk0EvzpFk2wHOGiAlX6o8357xXf41L7Wy7VZqB+ch+5We3vluEnINxPquo+xrob5V5Xg
CdJppaj7yNE8zB890PVxOh0VoomgTEdQFE5LlWLItW3TSZHnzfmUtYbMxswknplrVBWyBblphKOA
BW/YgfaK8ekRujoU6JBxHHIYg6aMpP4fdiS4CKK+pqLJSS72Y5Nwqe20AvIkSy4SRK0JQdGOG8Wx
doHY5JAgpQ9bbszSIn4Q8ta7DaJe1G1s/V8aQbLVrkDFw8tZNJZihDL5x4nuCp0edi5VLUvMDfmO
TkjyAR0f8HyCxFzrY7xMmNjKn0U/3AIajk3SrtMvzj98Qh4uculypARlhk3R3UqTvFuNQe/AFb2T
ouAhQC9PhcRJg1H49LZT/9yikB/XeI5Lb3vHI/0qE+pg6UeuXR0AY2l3zo2vWTWSpAtLyeWUpyrE
8S8cNpsdgEwAnNgjc0iIpS5aVcZFjVzXDfWyU7fcMutOaLbZGl++J+yNCsaAMJZwbjNfGGoj2ICw
g9ctrFtmqOJftiZxR8tNQl/i3a4L5a1+4NHoFDK6J/0j4mLIQeGM014TtXQ/3mZFRknKCkYkJZht
xNfQZTDzdrKuaq3rO+S1r6jt9oCfAvPvLbXZmfZWdSnAJM0SSosa/8g1dBNCRprCmTKXeadbxUn1
TMYilwMvBrqrGRXr5lqDitGs1fv1MnOZo05jRLyiZHQyHA41eVJ+OGNqbAqm3yEwBiYjtNairEs1
dfcLzwSKH0Kp8rmgIB5LJhw6xqBLvNO78gJuFLzWq0NJ8w4/4lzxvi7iQ/LACOf7o5xyrUWsu7IP
Yr39mS/rmPF1ZBckZmsQBkn9mYZWRMEE1jCZiw+R95AwF9fl6Ltfv3saR0W+kTZd7MHnXWgL0+2K
edF+uvZ4mBcuPkT0GkHvFfsxFhyIHW8g4q+0pWIP5mwyT+/RxNzBPGbnFFV7WEyW6FBaWBAKT0qB
gz70xUSfof+qXVducEoQU5xEygeA08e+Ot4KC1GMxIt9/TXxYdNfsoxMvu2DSSZqtJDCvlbHcJlX
mEi/gMAUNCRSA2kO6GfrUIXKOooBfjNWmHrpkajxLThqKb5gxvM4zuqZm841bM5RY2ae2T1VGjGa
5zSB7689l8VXi+x7ZCSImOfnz3Fa42sHQZSJItrghnB9Ia1mGtdRvPkHpgIRxgHpmojtSHRfz3Hn
tngJGofZUSjHED8FoO+21tK7Iz2s3MHhQCnjdNMp4aZDQeFMSllV1Z9+ptu6k6iBLqvSB5934KLk
Cex4OfUoyjxyuqXZehH2fH/m8pr3N/B3GmWVjtSXR2PeLGJExR12wZUuFNZ5JixZIdCPX1t/oE+k
Ex6pcxY94tRvealNvGGON/zzZFthuGnadrR2ay1VumxyAlUlJi3AaFiWQSKNWPISb5PAh2PGYe9S
uVCYbTO4jBtfSF1vLgPYMRcFDX7GS1lglStOkUVbUogNK6jIOSiV1t7ECXQX2JbP278ywBgfLTZm
Lz62lTk5AwUK/ZUgrc2b2+Tb1nmMmKsD7VqsSJ08wxGClw4PDjcsmV14uLMKMRYKb2DS8LMgnEmD
yBVZVEU3xBLU7G5MiuxQv2A+lrDj4Ec7JGoR21xhKqajQLyO19oPNI52UDL8f2kxjO1DXEj+BHXo
XAw869oqTgsC6hFf+Jr190tCUbiPhVFYlh7vX9vPIFX6eWDQTdxzLFqendE1niNYDiRul6QFkbsd
wXxvatyBE5CfsnBQ/uPCkWqkUH/YB20Do3aGoPf3hSui/KiuEjmWQFeCIYHxE5HjXQ/5rS7v5/b1
SmHMU1STEGHio0M8gUK5tcF86B+5QtUnlDz1wbxpNkXt5PhmfTdsYC9Eu/ZaQ4w5NOdiAAo4dueU
Rs1jeUHYOw6aCYxnq1f7Wtx1xGAErwUtBCcjb8DjrvsE++t5KMIBvKas1YAGsfDO5I8UjqmfNxYY
K96T3D01b1d/Uq80W6j3eRqPl5boZMzBFReGAtM5pHeIGDJF/CIvK2/F34H2qnwvcNFf7U59WxL8
61d9Gsti6TCc5mnzgXLXqqoNlv0eXjwLiR2tc/GxJiYbuqNYyBOFm5ko9UFZ8KVgF5VbIIX6CA7/
85Klk4HOoVrvZI83aLw4HE2z8F2nqOSzehw2MgWBxAc8Qp3hUbpcFyIupgd1JyxVIfMZu3eautu4
XZb0lQ5XcbP0GwayRws6frtNJQjhfg+eOjFRJd2CHsISXscg/2c96Tm6zd3wMLV/bJWMO+meQO6h
kWlHoXG8MfF0/3IeVBe9zrTvuxcrAcUPupF8TtMHhfBF/YtYIia8j86AltccXPyYwGeqbBwOb500
TMT+sFfNXoTSvm6F7HwrhHYzOnu6UxGK4tp17VKf81Pt4Q/K5hgd5K0v8Mpbmsc+Cn/cdBFq8rDy
hSSK1HxswOcsblnqD51ynu2gf+6l7gAopBhoIQ+ayD2cg4ximSQZVy8eXy4UBCWSVERoLGEHxwqo
6JfhsUHBlwyfVSL7xNCB5iGrNZM7X3P4jwsUgSW0dj4Kb5p9+c/FvEcx8dHIM+bYbdabAYLtGymC
df+XEphiFTuP6uUEuzUlm4jCnrvHd7UXhBP3J8K2gQojUVm2CElbOnUR8w4SYcs+3SLwKzgIIoVj
bmXOxpeRAtaS0YBjSiER/NuYrFq9V5Ahtt3u1dk0+YDZz+as8WesSYkTcdD+mKmIFB5t6cjCS2W9
gCzpyLkd+Y7IiiTvYEsXfKv19BwUJZ1jkeRb5IWWr3rOxw27iTwOqibGB67lXSfhBfbkFbq134Qg
oXiCOD0NfA/29WbOpdVtlqjaXyak7XLX6/E7oV2DgM5VGlahSW6z0xQmt2mFXTJ3a0Bw0Wuh8Qm/
/ri0UI0zQY30nQfVOZgYCtwZV3RwRE14GYkNFX4NVxpCRG6kXQmBnReQRZVq+ACke8PUjLtifv/U
eVn/1nvH/zXBsuj6mszkSqmmYuyB0tgOkfexjosJ5FvA/LdiFDbgYFDPWNEt5odLfPtWxG/MP/Oz
QbReJ/OUNpIH2JgTPtcqMjdLO36wACYgG++SkbMXjtdLYNTgBJGpALSFxE06jt13kGifOdr+ZYzg
sxu66zpScdLfIHmdCGSC8kh/xNNH2U6fnL0CGYGSNJdyk8hIRG7BVwhIOAlGEfz9XAl6MKLb4vhr
nZQl4GcyZ+jhSe3qX5E2kt5LoLfDg1vfi4i2GBSNNWvRCrEdPmBIL866HCUDDhXbzPXP98DL9sd+
S+x2zHDBL8WiKVeUe9sXqKiCe7mPmCZ+6hFtcZ6cBCaZVshBrTsRWD6CUlqi1yL600iTPSUz/Fh1
lCyf0kj0Qomf1JYBj9vlQjTijcp1BDON6BE8uPu7YhS7XY1x6cJCBXP/U2rC/UmhvQWNMouGt2FS
KF4GPUvs9Xsu0BO5eOwVDAGSddpy+W9l8YM06NVmdDbhr4sYlWIBOoLyrkjWyNg79Wvi2MDUQ9Zd
JL4Pst6N/NRrSQsM4iHF0nVcIW/YcMh37rT21wv2l+XX+00ccIhqzFXH+CcTlQeANYy0Z4q/UjWe
5JtNPBQv+ki7bakY40itgeyEiDCjX8erVjfZQf2zq3pUv8GA0j/JNsmZ1xM4+jX/iF5uBqlcVvS5
br30oLsJ7gbBXROt4X5y7RUGrZvhzRE5cgXwlBzMTJvRW8hQKGmRuAjVanFJ7+yfT/M3pKJ/oVah
dmcjvk5bURm1AoerRo3pDcjFlepsyhXVDaGDN7XCQNYNBmWO/oBpGGonjg3VTkCTGxvliympqm0D
fN1gcn+BajovpzAcDff0d8kwekpZMBlP55CP8DVwtIO5DHAIyISrfMDykP6XI2J+aY5feRJbFdkI
u+yLfr9XmLEJrQNqUgLk1pGQ9F/6DWtZUGOfrPI6ORLcMf3KO/7rOrQuDuipNUqePQJcIhYxgE14
G2YigWsandKf8yz3mEh4Xt8nRFBjRES+u8jqwWAuhI/gBT+SmCIgcXco1OwQ2PK4BNX2miYmQzmF
78jqIqxXLkH/8YfvK/0RBsS/yiWujvDwwgu3R+gsgmw0kRMSyYCO9Dc/z64U08BmNMZKIGcfw66o
amarfDkg8pGTjcpt2wsmmb5MmP1r9Ld7qbsxRTDKclmcc9qJPVBLEF5SzBs4BR14XE/6CsaDMfdJ
95Avx6Q7eJ3ZzfKa7a/F5XXJ5rXLDBBRx8Rp49BBZaXlCLcwa5iCakTg5OiBc3b3loncgBBPvHuU
Gl7OHtiGJA8LDZ6wKJW2BrtZl9TVLiC2XvN/2sGhAvtIZDoKrrCwztSZwvubYlGbD4RORHitPKDG
tlsMmhtJlbcXecszYbCR3SqRA79ICwCLZIDij6uh/Iq6PkFMAfedB7afcqR3gPtam4JB6c5GkVN9
q0Q3C/w8XZ8cg5qSQN0nBrWr27JzxiHSWGHJFLYh7MW+Lae0Yhhm/g0W9UBRuN4w2Y8SNUPPawDf
NKzl7s795LuW1jv2Q4FewNPdZ0dMOQ24+Reofh8/v/t+AiLhgteda2h9zWJtsUVCOor4ZUTSZsVj
AgrBCp95DNFFCSXwiLy5s89MghLv51R3Fd0mS06c7dOYQzwyyE9ju4F/eWdcSv0rsiWXo//AEJTE
1KsEuEdfAYr2HxjrI1pKR6owNUxJjJzTcyPGdo+1SlpUB5REXadbaIBG8jFZd1b5aepPmtRhiNiJ
AvtlzYbygDacMH2dMW02E2H4PGrRDfkZ0ZULC2roMRVtjw/3aP6QR0z/ofHGuBCPpWn/k4suYlij
j6NDbnjjjNttMz2c9EFlcKiQAIKAWNv7dYLcFYku/vJtdfNNw1BWSNDUDG16bnZvWUajJXgdsQak
N1asUfOJm97pOEgcPHCBj2OU0JukiDz8YcG2C7UDY6v+I5tpu0eb3U7F8EgAal4te8AIV5zVzJnC
APGhh+gKiEpwbwR75i+sv6xPcD8K82ngy2stp7xVPW5XCtWbYA66iPzZrcq8HHmHrpz6IhZNb0oL
agMjTZOzs2hJk/naPdgOT7TLJn0R18QXl10OZBe43DCRM47TlWbY/97G8JkTi3zOn9aCuzA9ARQc
vXLRwMXfcIAZ3+AZ/FLqV93MfxUHaivqnRwAcoy14jfcCFR9AYlgF50Qt1sO1aV2Ga3JSzcA736v
qLWZWq28hJCpfLqpShTH+gL4pN7ZT7no4wP12gpg3/7BVAhGUAJyk7kK3oXDiVF+PiKLIEtLjJmU
tqYqDPJoEhfIAkfHG3JsR2LGN98byemKTbUli8HyrCh6b5qJ27rNoqmbhwGj5XnpoEpH0YmcDZLG
GfVSwwPQ3sf4EiL0EPx85ITq7J0cqMglK7n6mKsUaR6AeEF86CkhkBhL5LBZGTgfWCzz7DB68f2p
jdzfj3uQ8W0w1Aws8xBCJMU8HA88xOkoQBKrP8f4AasNbO9M9QVrIhWOhEfdvl5Zwkjy98oRuYXT
ZReTpjTkv4BE+j5Bjw7cDcQ1ZPM+C6pwD9EL7PW59qBr2Yjy/JjxgcbCOH2iq/DGpVSJ2p+CdU38
KTm85NtUe7Iz2gqKe274qsYLylMAQNvaGUGX7pyzaRbEcaNlqXFZ9wZkR0I6x4qM/dADw8u6rYX0
3DEyUxAwKOSaaqRcil3iuKDEtF8rEXvDuLsCcKQ/LSQWmJPN3yZNSnsGwWTx41ZVMS0xrxERjBUW
nkKPUimk0iAW2rXT1vlb4Yp1FrkjZlvVr7Xs7vy9zkWpsjr5sFd8qo9leBzK96Jp7HTeor3qpPsj
r7mWQsq659uzUveVsPSoeJ1TK6Z3GPs0Q4aWjhZrEb+oMUN44NOINisDt4bLEUf6nTnmc0yjWJ/X
jYhS1Mnwy5RTjQDORt99PCNH+JLMomANKXOFDbCyJhK3X/zWZDBYRtnIpy429zODFAwWJQe13wy/
deuERxCcxJwQXtN/WgwJsw+EaVaIEIpduqstyEpvKH7UXoxPeGx3P8znKXixoCpOdO2+6FVjmg0L
hbhZwKxqp79GePDciag9qNloilZS79YO8qPLRob5qlD1dRLNy+40ZsSFClHZOu82+QEwgJj9uxgX
BAiHcdU/kO8aeQgaJeBB7uu3Geyl2Xv083kvXSbtgSmT2Bx7Xpxwuy46pCk0saXjT1xzpYTnPAzU
Br0noZymzi0KpiVIwwjeoB2oPtXJwUdPXHw+n5mkSOasNL4W9LT5HAU15HYFqxXJqzUBI8gwj9OO
3QINdvoozesr0ezPi/w7sRZ+qAaGan2m/JlbZU4JMyz0G/AOw38CWiOvv2AUC0ayujmJVFNij5UP
pELFHv2Cn0YCBIguNw53NvGRX77mwyjb7RtgjDG5yp4p/jqAVpnmjJERadfGQdIxVgc3VCNsTDiA
+iOkYv+UbWoLGE+xglqiKwsVwdNtChDEBU8fu760MOq6NxIgpV8fTIp0VZDOvl3ViMLFDefRPWRb
u4QagdEwmJstuBdbgvcxyKZAX5XJZeXJ0JA7pT393Vldh5L3wZs3bmXnsl35EP+U5YOzD9R2+4j8
b8ZYX5gpUvWXYRPFZu7G7/7V9KemA7calKZPABl/RwbpNUnEkBVTk7pDlIWQSVxEkJgI7h87eORQ
eex4jnPulF5XaZwdcxgRQyufAuFeoBjwMMsFZ/W1NZeRAJ/BUc+MQBz2z3ROSLZIG3jiF1IqkORH
Iy5waMn7Tj/Jcn3sLlkkcoIYvtw/Qkw23ICHNaAhUayV8AP+hYemXT9UMl5DunD/isL8XS1BdL6n
dRwZYbvqfrXcZ7uvSv/SgPrXuEnCG1FGKv7JW/hRCz0j8wlcrmPpzDUdEHGh9qBP7kPiKh805sBZ
KYEJEn0ViN0CZNL+j0x1Nq7JFzjk7CsLSvFV5JTfowiz0FBdWJh0Vv1NuGvVJYPZmnpg2a7AqlCO
sL3krV79m0wiM6z86MNKgKzvkRqeMRiJKIDf/qJc2CHqpCqMPQogTuX9pFObazTkzwbj91eGit5x
mbR+/tMJVh+1CMheXn/g4D3P7ZkKqmMdOjs7w8SXhmPwXPsCwKSQM2okv5Fl9HCgKWpJJiV4YDQF
yF6pa4U3JoNSC5YvdBk8yIC971MbJM0ROcIFpvFIVeGmB907i8WP/ATyKylf0BgPQf3hcs7T1LyS
ELZCuuW1hhLt5NoRrDBkru4r9yKV0IRmGtGdxy3xBDU4hw6boIi2HXWFIg/jDFgJR5zaW7ZBrBaS
3iQbYNbOQQxwKjJsAI2lP2PEKHnpw4ErmoTG8mDel5iouWP7L5XdRGlGwmvd0GyXTVk5DTUUlbqf
x+irfRtnZ1DjKyPIXtHVBkyVxKWAHo0lhVIXPyHwtdfW2cwjaHa/13tlXNPs38dNla6SC9e1QPAV
W3qC/mn3ziyJ6fOALcZZCGd0jcjUDjdJkZ+Gnf9JjtDd8YT0Yz4x4zO/i/6Jb/YQwNTTDW0lY4KJ
Zzo23d50aqtfC8M1xlVWDyNaCC1vAyD2NwnW8U1VPQg5zie5UA4uoS/rPsgJ8DDNfIKUv9llGnXF
mYttNRp00aDc617szIYUWVuhSjDABgtTpC1HbHZHK3Ba3Lt0UZEVen20LD2/e/rMX8a3rn00mDc7
M8cQLWL+c+s0kzKQQtCgoizJZkwpcG9Hm2hlCoa1NL0UAMB7lfUa/oJ4b8/jchuqLyI0O3rW5aAF
6yRJ3v2DcHkSm1Ia/Uu1+oV04ybHIwfMPPAgow5PhH2KSl3fBU991JnT6GsetAWBDfG/pT+Zo1tF
ct3sLczyRNBnQns6rbo2OD8IqfrD51XgPn72/QxjYTuNMn/MN3rghOeZsl8lhENSvrPCwEwhBKtn
UAuCwIGl8VF4sdCxg9kNPkqR3daiO0DKuqeYb1WC9uVUDvm3Nls2ogEd/iwO+bqFTeP5kboP3Zck
GOFD+qN1gZvE+i2IbsrWrV4L0d2RCc3JSfsmsA8o67W0dq2b/IeFENqo+qWPrOaIhROuW671JRmV
nxI8Vi+1/t7TY3L3TkvZMFgGFJfn9A59uw8QNK2Dl3V6VUtsMMb27ScTr2EzTpOTv6hbbME4MUkf
G9q15C7tB3SQuVQ5jQljV7wgNP5FBqXtPoHnv3/bgvIP2TtUaYKrmKlqTRkZr5ofhBIxBd6o4DB4
6/fI8M1s/PIzMyDlS2s8hbTDyKABo1Cr8zKbdY6t+jlU1dvRceniUwDtjxhKsopbfa0RVoO33nd3
wbfIji6n0QhjRI2tCZcVXuWix4kuJMU81twWD8ytJA5yP9ePt6m06LRqJY7yzu0nCCwnvaIY7WNI
vermTwBtSwwa6uJ2IGkEpjNivClyuq1sof0Cyq1NgFq8KIsxmwXXB6JEP2KrAMLKXByLSKqsefEI
ScJ7OaRXRdWo6IlA4uSG96MFBX4FMVdyutZQPt8FARLsKaQSjkmE1P1huX0tQTML5wI1LwvCHyJL
cN4M5qUhVY+EnqXQ24utR1WR7nAn4w6Rw8+Rh1TGnfC/mcqCyGK6qS5m60hsdIF3x3jB1ccq/r+v
MpK2eTv/rHRR6Q0a9u8BFiFnD16EWHfm0PcoSPZlxGqhUGYyH13YnFXMAowMMl5Myigr5bAHJfdp
A6kSvDWvsJA6EEgUEvNCho3ZQyF/OpLwAhqgUhvXK6Sls5+ODheAjDF2uJBgfjTO4tL+i5BQZdDJ
LvavfY8zFffSnekcDjwPCaCuI/prHL9WAVz2oR3eiUNKHSZMUCDXWs5cBY9TAQN+xFWgamcwbGRk
VQIvjYhal7/iyvEqbaHW/yQUUILsCgzDcnvRrEGyf+7MXO06luXfs3Q9nj+bf0ojeXja3xpoQfQP
LlTACqeeyRJNoOzyOCJ9A9/p8mh+6N9yov4qMwrDwH6sjGFiYe8uga6h2nWhEKIj78N2T23imd4u
A2Bi9CkKHDD3igUkoQyWQVMJltmgyooJbMFbGYoZEoL4uDtwzOF0Qamjgmyh71vx6txPAsck26IT
IVswYCe4Yd/+uEr132MH16kVnPJ77ezc7jC4gRSaj2MXvuRD0uZUJPuq6FrfjstNfZNo/W+QmTVG
R6xUmB49O2OisqkHzPKqlw39u4XQmi12pjSp5U6EXTAcVhkdyrNbn+OniTEoFjqnUJdi4Dv81QEL
5dYwGLKl8T1it3PX0xvt8gwN1NZk65OlmV3/vmLq0gQaiC6HHkZ9tDbziT8oXbVnr1zI6nNVlrsM
LOnaB0yvkedE6Ue1I+DDSQjh7t25JlyJH/xarEra/9My33Hktr3l2kK0uqIc5W0tXOK4j6LjGMsV
g6Ru/zbE2MDrRIYYjgQ3T32xonocTdXt+AURcOqHUBIEI3B9t/oafbIy8U50VUJHXIUbtWXOzRZZ
ZEmqy2KXq/VQJPa0a3JyPocLXunOKAc8ZHcXCDn6cpuRyYjfrju2hM3ZIimh8nZdL23jsBvRc0YU
7Dz/YRZhKsm2EhnNZUcsVSuRoNKkgHzQRh3tzzvOwpl5SBUEP71P3wJIqH0Te+VnVfkk+qXlKThm
EFt77faIzcW4SnpqsHYGGf5JFuNXcBw3oC+HG4Hu1H0qJoSJgRYwisZz2NJPIlN+Gv59DyHH4UbE
3uRgdllsxLSh3CH2e102NfjS2U8+RPOMvuuvPDIvqae3z0UFZSaYquwXpGe6SRFp3IsmNIsuRazf
8bv5bNQlGwGevxAeN8C+2MMGYR80LMFGe60rjJwb/houWnApNj2v/vCb7jUCa6WFpG6lRE/b55pI
QiejzQoSxHuIKdFEqVFEH+23ufoQVYbb4OdCwJtWhh1QTyX+m+Wz1a/eVUlh/L285wwor2V/fpvE
AXfXrBdSyiknd8cuUn1izDF3rumXY/a3UhnWDe06QUFtyyglUz1fcgnTLvB2PE4zyfR3MSjvQZb2
pt6osH10MW/+PRn3zN2fEWIM1/WFgwsxWnZQ/Y1V9psYD5giDVS1CKW10eqEeUh5mc20olfWIFzW
mibzv3sJrygmM2Pqx7kx1aabQzw95LziP+wSVz7FSPkl1ulVZbF9vtZ8l/DAiXYtpSNrqkvUU2FZ
mormkcudiw5oKVFQtr3PyO+tpGKpccmhDI0rM8psUHrYESx5P+wVo1RJgRTSnQp7U9Bb/5xwsOVg
py5Ri84pz3Rsxm91LSYDfDRuiKVjo7uIsdm+yzIzKQcKgGltF8F4wYZerbexJTx5TKdftRDdcgxB
NgB93BOefQxQ1MwKp8HaVUmz7pjjdAoXsr0tH0YvOT+XLmoJgWGRa1Qr+1xqdH1xc3u4paiBo+tP
JoropJgu4ot7IOg2vrE4Vm7KtqrPNvQesPMCZKmMgoIB73KfWWLSgvjDvwEs47gPipT2fvxgHdJT
lPvMr1Yac3+8z+l/JvLekDUSgaJUjaunQuSaXbPEIIQaZMmvRLE114IX/64yfyYKAfirphEvCP93
NHowHlWGvj7hV7X8/T76NrTSeuvVc1uX/zgfLC5PGwOHsWUpn7d/zhXO0+GatemfMFCdGsbq7XcQ
5SNJ0KWEKrzpiSu4xEJBrFwq/HxgCqnZLMUQ7hDsMES0cTiKOt7KYdPsClOVrbRF965dFod6giXO
ONg1ndwK43Q5zL+VQ9AlDk0BY5a7YR8tQ1lwXMNiKgCtJwiCi36W7XHwuYfch85L724u8mVY0x20
oPTE7Jy4kMVJNpYDhmDMNt+aGAHBRQoJbbViEPUk5LnGhaKNVb9jfrOrbSX6EIbIgMGP8E57a3JB
0cg32Go/rRUcRxIotB5pb3zBC5E4YDT1p9EbnOVRztqRqSgykLV7XdM+6TrVJ97BPYFB+UZVRmlf
xLSuSiS+ofiAujghdRhqCuOO8YG+L3xYVu86sNP/FA9Iu9totRzgma9bRrcVF1e2si2SOUmhliPo
8OGtFJD+n/9cL2+aOSAXwqwUeahTy7D4HK9Xm4DGv4dgALLm7IUVJeTz6omNBaqu8dojVXombUi5
nEFq8PRG1aqwnqNBAZq0yFD/lmioBQ6KGMw5iWjX2ND4LJDg+svZS9fzTG+TM2judW2mrimf5j/I
lSMi0cuxXzS/r7sHxXVrieykqOWkNxrVIozfecaZSOCfqiOId13UmQbAWaTQbMJjfUm27pwxSCjE
NDElijKgg5Q9rAS0ZSd6WujzEPA5H7xoKIPluOSn6airCM8Ii6TnMQ+wQok8dMlAbOTglOtrAcfG
3xDGowvgVyRoIHpuHAu2gJEUYro2ttTCoEi1/xVUpXFVPOGxXRPkCf/Xy5KNcRmqMSsPqgZXi9BB
DdZkR6Qxy04qR6wRRVfojsUbXTqbYthNAws2vkd9tT0RuhXFieqNVXoYo6y2Gvb/DHHKx9IAEqIx
4Oh7JM+tOvhY0jU10hzRluPZk0uOZS11R+lzsMlZ5kcijJA6uaeXbD8vfrEoDCNbgwWVqCpjiIEN
YRsFy4nVRpCR/D+JMmPwq6UtvBXUjK0VzixmcW0Ug1MqmJjsGf5cFjxLBRZj7//dsGy91NRddDk7
htxN+V5wydY8ESEKvYQoq7LuOOc/6X3+ZumCZgf1oA2vM0V5xyfTecFiyp80Ri6SCgli9WPnktze
hRl/dgdwJoxd/fC9lJle00fcqBAmCHeddarWQqwzVZ8F2mdTGYWYwLWVR1rb8A7CJ2yKi/QnGJUW
zaaQM6GXav9gkm9UsbOSofm6kFA8BlaTltQgM9zdYR3eMw/q0GvoWBugI4uO29tz1IvGZzi2KE6q
UiMHbCSRCzxW6XP21p5yNDKObm96aekk2SF6lGb3ffsD4yQACyGh77ALZUUKS3y71bdENeqE0WLJ
L9VUathJTxl5FsbfsdH/3APOTmYcfSeDR9QGFP6vWYzXISm3aneuZ8Gy1HSL/0w+5o1Sq6XiE2bI
JFBqVzlfHRi0r3pZUG5VrOZtSh5ecjm2ZHKJdJWrkbAECZFIXXIfTHngewX2pScGxhyIxjbf218Q
cwSrFuRhQrtZChmR7z1/13ua0IObEcTmcaC/218mKYwSolKNt54ubFion9RdgdWcZgxHoWs+SXHD
EIQKM4wCOdspqDrCMDcCYlOKETKuFNm03oAO4GQIqPRZpkoDHFAE6A/53lfVEUIsAk00gE0Po9x1
1bMcMISci15ZeM0lVprxl6L1jP7NHmAC/kSU/3cVNnGbaYZJePAggsLK1KC1Jlj44a/hfjeu9u3h
JH/aIsM54Tdpz9bc9cS8I5bCS1AjbUA/gB7fTjZ4Hj+Ib021fJjm+W7M2YOmVEGMKpPqte+E/3s6
6I2Xn9jlkKaWv8+dPmpTT488g0sJs+Fkk3xI+Dq7tJPoRbA3YPcb59zgfubH4uYMjOWXH/MOClDA
jAcNhSjo7Viyd2BHVckCYqSANaI0JcEAf/OqUy8beraajq1Whp3DWTT7hAtvcavfBr2TfOjQQufA
mAPAP+Fi/9h2xDwmiTxYLga+YcuhnLbbVWFu3KU709eyP3E1Y3w8+VpCiQn0Hl8YfBykAZQBEDyp
Ro8eRJS1iuZBcrJch5Shmg4W2k/ZEJa/HSWOwff0FNJRDTtApvbSEUg8129vBZv+S97F3S/KySku
spm7s5836V3D44mdYukg0TCfOPrtOXiyKH2bhWYQ+RRco9ZtA5CEZRn7cWvh5RYiUqRRUvnUhlt3
qijn536jLAPO1djApTQjMT2A+zmjsx/wTiqycnUaVT1lOeAeyAtTd7xaZtQK0r7Su4FhKQbMZo+S
C1rAMH4ZiPPM9lYCetQAdM8URj4W4m1GnTWGBcRfZEas8Nh2AxNq+TaZR8jtLrvK5myvqReOOA6/
kwMSbCRtItLe3O6+Aj595WuEjvZsFeXLa38a0bZ3nHRFi+0gotRqmXTfHVgtWg5TQzUHA7nxRMwD
1w5mnYI5TFkCGbwJbr8oqG+3krUwyene5pbCzuFYKTSbhUPIBD/M6FPPmIC2FOMWCWy/PpmA/Bhx
MUHQAP5oRA5obmTWRZAODgTlUwRoRc0x10+m2J01qwKkZRbUOXB8CSmGLsq7ubNZoePMrUpJW109
T0TS+zyabq1eyjIcs47Xa7MKthj01Wadeu2pAhtOr6g9NX4vZUMQEia1YB0o7Fqqq9HkBpDGJH1T
aHS8p61q0bvtYHqqmrKICHY0dyJFNMuvK2P8yWHeqVGfykxA4904yeyOuza7upgFQj9+JXrECs9N
UiozNb8KchqPzRtW+U7Y+ZG2i9Ux1anDHfXpn9U7zqtLL94KZ9PSx2MqDPygXLJk8obTN4BF/13a
stz+t4MkUTkdpIQ5uzDXirgoGhayIu5M0X7n2dSiLjBZo/zqGxebKrk0HcrcO8sk4LSGwGSulgfV
TI283CZta7yVdBUle+1uDxfDh+cXSeHl42EXNMStAZOFxbkN9RUvS0+K7qVEblUgHYlxa1PUdE61
FwQe+cslPYLQZSN0+NrFPP4iAXRVBBTEYDDSfSLgPze4khZg3rsXXCFheLsWAyCxWCHrq9+rP+HL
HT1Ntj11Zv/jiU2Q3SuClSuN569V4o+vAGBDhX1eRG2cGkH2CfBgRbn6CTVB05hSesyY9hT0P/Gk
uEouuN08U2BJ7UB8xt0tglyesrlUZIHuuIK2oezZCDsuaIxRHvGAdMB6ntXOLRS1064Q1CHMCHZC
M3QlSUZNTeqXXZ1zPj01Xk4GTmfMYBxJiJdmfziusR/a0KNwLYt4BYo9XCYmF8ERhRLcO9/bf9Mj
rXguHeCr8K1mwiPrJ/4q3iUHqS5jRK3D7JTI2N5yCQ/NSENuW1rllVxk3Z0Ag101jrVXfMrmY7ae
Ii+vknd2DPjhC62Gb+9NUNosgRZSmj9bkQCkxTInKJzza9WOKy0Tqqhr3D9B+bJGwLPYh390oOra
UrRoQDJlYChCMTYdIvc73sTBXTLhNDWPFLebZHE2Hjs0BHBZU+L5auVlb9bh1ezmeNGmoYP5MS5C
/0JTOIXsyF/lk/Pz8hra9vOb2k/gpCWd6dxKO9HbqhXS+i5q53sBPWOwX0krnee2iiOcgTWZPvUt
4SB4YrKzPA6sBCeNnGsySarzelJ9Blf63UXfpDdfzl+3CEEv30mKEZ5l8qg3CEdnY12EWdTAZ38J
LAQvl3Iq9m02CWu0aqO6q4FUeJTiSlGA+37HJQctjk1g0hI7tItS/zTPsfD4dq8PQLck9ZmUkuV/
l+Zl3Pm37Zqbc7E4tOo5xxWCYI0iYqEgp2SpjeHfOZTQxTkzr8FyQrCbcKOtmWdA5JYocpsbOPk3
jh4Xr0vD1S8aB9o2DYMvOPl8+Q4vjZLJce6kE4C1MF9GddKa0I4YNfA3aPUy/HOV6kt/5Cv1oSwD
SmA/0ZsRjo6qN/3m/whuap9x5uXi/P1x2S/ra5P3J/TFvE68ec6H2Kn3M7gDNfEGSLNobUiAysGE
A1KS0Rl0lCvrHbMqLwItVlGI3HZJn1YYy2zU3rL/2oSkeGDn+ld+csZ/euriHTCpRA4GPFmVmZdi
d/qTufzrNvq0P9igLyZjy7tDc5Ct6egdD3JB2TlC70QdevRCo+AHGQnPPn0R/Z3If/YhXPBBjmH6
dHP2/Q6nxZAltXj+QyIkRfa8Zry8E0Ru4q0MfpKTTm0z6+HhCJnoim3erI0ue2kQ0S5SIF5L2Ymb
bldcsgaP4ybOYLSjZ46owNCK9+r0fRMBJUAHFVr5V6YxJHLLqwyDkdsaKMv22vELJSKzH1GWnU8A
t/HwaBOL4MyjLbDdLZkkVtBASiExdUxwtr2STRKOlxO6jP66YXLnChiQ4Wjx+SiPChMTCH2BHNq5
u0JREB7BgPXG4kjDo957t/jS3s9WB2DtM+j3t5nTBFcx2qjtBwRvWJbXWIbi0ExFD1F/qZQt+MyJ
/faRY4pxEhPBFLqDN51WDZEVXodkHMCo9W3Cf5rEtLzK7F/H1SjtRljSw7B0bxg1Z1vROB1sXhPD
bUx0h1KgeHkrUTEEUhvq2lDGBj/kIjY6YWNwGJFAJ9KV89HN6YMQdfZe9jHrGNc7eTFyJeO9eams
9FHk5H/tojKBh3pa2NEG/V7B2RgR6Tbk0ALORBKJ345V+zEiSQQ/b0g7If9+jU/1wjmzjOw34cf+
i5Rh/OxWgoLUzSg+ML0Gllgov4DTYeQ/TmfmirgZfmhOIDU0Y+YP/7Mb+qwQrl/3138OoLzahO72
w6Ton+1U6/HkD43qPe446kJsoUttzYwCG0au4bWuLF9IB4OJqx57dGVCtiWj+pYHLNLAYK+j2Qk4
HVgVukIOob6yoby8v3dE3O//FOA4nlx8MBarmOuaMc+lUPtEbuwS3kfAKAVxJESUCJNKAP3Mk66X
qcPmWI7/QHXoS4hgjrxUVmq4wmPEAwMbdpfY8o/HicyTLnxXGQK6eNSRHOzFAMPOPsx8k2IgrLsF
tT2u2YHm8VVdjkulpzJiiriMRNc+T8wdXn7B6I52O/3/OK/OCVcyTuL1NhG0v8XjZfRYgP2fPKuy
450viN/0GAKkVRbdor4q2rSIyf0lx0EJe2kcsFY6HxEhxj3WRf1NDDzo/cDAaoluHLmFnyHg/G3v
GPU/PRX67ndSp8Tok1ct5u+AiOQ4WyoFYXnBh+pdc9ZyhJwBSEGP/C8lZLaXDNcAybzXK9s4f5dI
Ut4tBVyoIYoZ26EwDjP6ZJ7zoqLltZK6xDgFvpDw6iufzghDwdLDJshtXKvp6IQUbKlwOQcjEIRr
T87SD5EWnvoFbhRaL+n0F6hZjzYTWXbxnV7eC2X5TYv2IoC1daWaxT0qxOjFpvXOuzAGedEoKp19
W4t/TDlGGNsq16v0QJ3tqhaFgthLND2QlySdsb+LhUu1HVO6INyFU5oiF9LdM2TPuvy92djt0aIA
RA6e4az4EuPuJjtigdzMjW1bSrgyWvJjkdevld3Us2z/Qad6nN/q6g/nOFmI6C+V15U16S7moUD1
8ygGecWeL6tabYm7Emj5Y10wGxBCUL5JPuEy/mjdD6UZG9poyNyehGli4gsgvb0yt4WJJyVnkhMC
MwsDCpYsTsA58jEVuiFHdFN2jRXCFysuPKTYIhRPBl/QYGd45mJLQ/kOYPFicKE+pUAlFKOjtXyt
Yp8MkbjhTwjCjaXPJwqrIlyH86zqo3VmCNhRtJdM2EoOXsosYyonD7mOaUul1ejTi6+d80RCYMBn
TXdtmXisyPE8AMVpftUGEIKhEH/QwAAE4T2sq9BW2CfpcBensoO2P+2/QVbMBpX6uZ3kWh/gkPvn
eqJMR6PuMTExWLPhRzT+49y715NRTxDAsGsKxBA2CVDmyXdmPspCuzXGab0ftOVmCUbfElFNb/Oq
5YKSlmH2wXZ0zR151DBld2XYeRF68vZ+eYjNklXq7CvCARzfUlJulnxZWt6C8MB7YQA+34U3+fGp
cgscp+R+rbWZADqTtJfc0+nB48vKVu7uVRWd6EvYNodCepNWrphV/vWA4iYhJQ8a0wDBYHY3FsLm
4hgoMl2fwwo03/rip4oJSfzXAx0Ngys3q1aVdVTdMstad0s8Azr01dC6yCOa39fDjvOljOOBRqfT
4N912UvLUV++9SZtZD5zv9K4ZhLcmMN/m1M4BvaljCqHT4S4g8mKeUgMpcj9SU/s/sOzN9gVTrRn
uE35ZNmE2IHUhLpg4L/6lH1OZjlj832s9UKq5pmr+S4Z3KWPsibgS9k/1D3sLFg7INTUj5uoDy5/
fj5Twl1F3SLtF7gvh6Xn/vNDDhsgtLpFHN8bcrRPGb3+SHLuDoRDNIZnhUU6Ij2/g/AoLES47zCK
eXmCoVO03q5ohSOt+Cpuf9eFmwYqh76drDUhcDQH59yetXn1b+QeTFFF+WhTUfwOL+Diq9G4Jvbh
Ihb120W4HVaFx9b/92oZg8fCTy6407pjrq1i4YfEdVlFB78VXKdirnGgXpcseUOU6YjJijWaVRO5
LD7NF7bmFBDjNVW5hm+/yn6usfWbVknppwrJOJowqWq5vRkrE39TvObeKTJsBg9SLRn0M+yhK0kN
LJ6tjz8VZMQKRFYNdOm6mh7evG1DillCvUB0wev+tY8d9ZJlyxialOZAjj0H5JEpUSkgFsGvZxID
dDtvcxT2HvbH7L/RfQf+n89Es5VW6lfjEOpaOHHT+JMFseTWT0yHb+MHZE572R+MBT+anJbGBB46
K4z+4JdM8bCdPx9AKGiFCVFgWLFQuo2agPlcBJUeikjebsXPS7TBalI6qPYeiq14i+quSy+q6f6d
wIMZvsRBck5IEdhu5bAnelvsiT76jGFF7ahNf+0U0qY7s+oHBQPNVqMVXb33ujzryHVwPgFpV/Cd
IsDJvmN8f62VWYFxlW8K8kabxSgkQXXHSu++7Z9RpHMV+nKnVBfbl7lhKzqWwtKRuKZ6RH3OwTby
Ezdpps+YgPMLjNoX2saU4Q9Gr33/nh/1BH13ySzEaAfoa19OdAcJaPWKgpQsBtwy/MNGs5EgwoJE
01fDUov1Z2NPX2JqlvAtRVwRRe+4YldYT4rIjJRx+UvOkIbO0GcEY0qoWbFXW78O+ys81rv14Y/X
fkci6ujknbW16F/111iKLh5Xto4z3u0gtC70rwMIwCL3ec76QcQA8uxuZSV1Q63tmE8zMCq6UMZF
Td243FzD5C7WBnd/na0wEiJnM7OrymXHgVFruVB0MalVJU7QMIls5stMXw8Q8dVMX1phaZATRTNH
gBiCJeI1pG1txBBeXlDI7p70CPEi6a8oTBsCrMzubjI1KCAGuwCVScaVI6SyLzsjmAFkMEQOCxAE
X/8yAsG5795RhmB/jztysrZUEemPWInplyVhEi+4ESShKHT9n2yvlEXbmqgucfB96BGn72e51h2+
/yW1NCVELbRx4fi/6xyuTM4v8CfzdkKOo7489Sw1KrEOGzH+YCxeplmjb9VHWUjGHTXdFi9b+tY4
iqPFZFhBvYVDGJoCu1JDZT5PUswkDUPo6cmdEaU90itMnjLipXBj24608xaDWMh0x+6tDfmximch
Qyk6bc1bUiM4V7o9UjqFnNVMMsUoAgIPOq9rFYwQY9wZubyi+BF4hkFOUBNpynQNg0wOjLqz8p5h
1i1xIaewoz0oz4J665vX/b+cgwWtw7wJoAQJO9DRcL0GK1a+KvOotguLE95rSkzAoucCuQG8ZkJZ
Nu3XPTh0icAILqTCHXE2LygrRMs3cpmjv54wLJXP8ok/DkH8El4/J8Du6tM4STKYLyoJc4s2EeV3
igviG5VC/nnlrAwXtjZsIFtK7trXpW3ut6e64U1xiabqpICz2dr+y+Rf1YxUptvSVxONfwvZoMJN
Ul+ITOMai2D46X4/uCZ3rOVwtJy9KmTwsHzNl3hOyn+/JzcQ2k10q/Ov2cgK3zbG3cjbVjEo+av2
LWfBN3w0ySdHFlPKkb1y7Vy39gJG8s7REQ1w2shFPC2pjNZ7U6ptvKthncU7NBr5XWO0fbP9BEjl
1oI9BwD6dHljYHIRyzRcernnWpSQvHROeTXMTsO68YENRVqL1LTHt4NttL78JTnK8DSPBPuC9ycJ
/HNcfdIM8eCuVzyJH4aIzI5PVrXwUqioq87alYMJ7UtX1o/qy0KJl6YBzxhgv7qTXb5/RNxlt59d
sqPeJCGG0dJm2u1hXsKVBi8GjjeGewu1Li8VGpp5ouM45pMwayMVTncUVvU2w41Hi4h35NNSRRqe
0p9D7JG1LdgOxTm/ojk9ThgEkGXfRd/KQf0ru4kIo6BF/0Bt5bggguRkreaBpoBjjxyXVaYGDt45
XXw6etQFxihUuuvWTbn61+9YvihhzVew49I3cv9xqyXYmzrVltisqxyfBD4oghnhe2TesmxbWbTF
x7zfqj5HRilx17vIn88JLW/RbMIA3vn6W77IAGMONiulPqqStm4ub91jJUaj54JSEd8MJh9/bzSN
hQejVFnqKI1xOQGvmx+MGyfUjIFPyUMSx3xU32PJ4y4ebEFihgmqiSDLNxjeRLeVtoJf9RmM1XjR
oSD1g2plwIe60SX3lgzH84kN0ScvKvTQHSD+MRSnbSCGsgOW3soWSbsHfJOqxRs3qV/5u545ub2u
gytRtIWF7n5YjLLZ0wzxfr40fGA7oK03hjXac7uHHym+6qK9tNBmqA4NXG0VcSiwZINrG4mAhPIV
XmC1JHTfct102v4wJSyDXU4M5SeDtZOLqfu8OLEPULHgB9kOFIBA8USMdGSoUwjRrybhAbAmYmq4
PlaPI9YjuJGFDzeaSbPUCNCJLw9UuWyO58yxNXsVb9vv/0SiwJQuQvF90MH3ASAIxGXhss/pwAHQ
YmuyltPDlfElj5f3I1Sw/ZmZw1CoTqhO3vmmqb3FtemimeZc129uSYkN44cGLFUJ0DVcD1IvBpEt
buqGGbs79MtbkxwePcD65qV3tQl10JJzFkq0aGFH1L/m+eRhp75yhFZxWEIHAAGGetE1kxJQRlUm
WqOR1i8rEi4bpACIEeKm9TBPqokuxyEjwgJtczTE0xttBZpr87oBrEf6gio6a6VJ/LF2KnED3LKV
to18HpVf5q2SVTC1GqM6VG5sLVXXwisvoR7QoRKQDU0oAVL7OgQTnJSPuGlJVxU+vgJH7YJ7dT1h
kz/y6jFj3b0aWhGT9P+p66ZmV0kwtWXBH7b2Dde2+f6Zuj4yfvKZXvvPTjyC34NBctlSwubTcaCn
zhPtl9uPqrPdmeTcVIfl7zwQjkS1vionuwSiatvagw5c+EM5Xu/dy3AOw9xY6xPMQEhPJTqQAZhg
BTnm2QNGYbNg5ih0ftGMsVH68hGXUlx7MgdEbcluhTQ7jlnDRibXPeW0gNVH9AZ8gJeou+BSkbcV
AXAJp35OuOOEhrjd3jfWji+XPxlncwjbo4XeiXvoLzegeRFgxniKuGO5JVs/S+4NiKV36FDt4AZT
oQiuhc98RWZNHfQOMIUdLW3VjLZ+3LWk1pH8uQtLCp458bnl8x24IZ/AGJHFsHZl+SzElBnngirr
oUAFj/MT1M4YyJ+ISE3UG73Pjjg0Z7EYBk+BK1vH/LcmcK9gZvFCtE3eNbF/LMy6sAWmmD+tV0Xt
7+Y+VKhM2gwCI+2pGruM87T0PQ7+4q9ZGovjreG5H4uNY5Ly3CgcaOmuZaU5Z2nDeQZWcrNL0zce
SaCAZNSZzNOascvz/0jUzF6RQNCE5Mq1nHZDp3BDPjuWvx2rrlrWeAZ0Gn7OLEW9KUbdZmswqBFH
Wl/siHzeiU1Z1w1BnUw0iP6op0KJdGWcGfb7DJhENWHag76SXUq0G2gAGjTgX3ivnt3xYYKvIkzP
sc+/r662GoWYaUJB/6D9P7TMgKTkUxFCbawmTjDpC1Gh1dFVHZV+SK7957uEHlGOPcaPSS+uk37S
aMk+ZdQnXqf+dU6Q+z376xjMmcem4ualfYLrpe7vq/MqYcb7cNeNT7Bc9jy6qmSWfTmBo6ptw+im
v25Dlu3ka/Xzb7mYocnGRBVrsXa/HglHEPjCFtEY6F2HEj4F2qRvcnp4/oUTLyp8BUqZhz24QZ48
OrF+wVOdYpOVzkGVEUKfwQ7oFnajjR5QubeqdCSCBljHLc0x3TctIk7o3GPuVwXqd0YXeH2sMeLI
i9UV9+uL08clnDEstAeV+2bDxTgPcKoydILjYmq+xaxawiau1se9WXbFJ9bJrqJbYMa/JOIqJbpX
UgXswfzk9rtqpx+yKleVK0XoaKRB2DDQ6pK6DBa+jcNqcgVOKcdlZbB2baBZZqWNfTv37kNRIrBU
WCrPgbn4cRNpP5X2Vy2JjqsEYyctCaMRkLBBnDRHgPmsYknVNfoWt0DP1AdHyYid4ocR7TkaSX6f
L0g9BhnmyBNM6DktplF/FVocUH2FJsx98lFBNrf9kqRyXUFlJBHySnYAOXIcipQIbEKjNB0jpIUd
FyBsTmjpwaFPMyeRW5XShwfKiuzOhqRevFxz1yC9JDOacbDR9+bsXZTMi0vRDdee1WdDXVRwl9CV
VNiuKfdaB287VcqYJXpgz2UJKj8axOn50sLn0YAFOk/nA1Y/PHiV7YDyiFShjlzhHbuQnM6N9tAq
hmWoA+EigysSABChUJqhKCp0yYJzH3ZeBzs+Bj2ueI1+a4XSCips8JT3YGjGloeOzOFcHPD0hhNM
/BpDoJt7lbj8ZrYNiO72fNqlZiU1ELahrQYWQgsYhfs3bCJjyF8dWovrblH5Hb3fRm0WZ4Uu/NWE
nh1OKrUsvqHjIGSt3Fgxz5/KD+31bnf2HlV1Q3PLE0wIbi1VOZ5q6MbtiTmA2hrFDwQD3zRJ3WUA
Gvnoa21bFRFVMoRpT3Sj2RmuKscIe8H3S42ObA1qlbZ1z9AL/tgQFWRf0/FMF6zmY9oYEnF7dcvQ
XRIF2FuBT/9G1bx+mUIKS1ejvIzHnZtVGq6hUVj1FFwqUhCjriidgs53W+xzIthYK9ChjQQYo3Yt
l4lAas+PqyZWUV99dBz0IpkGQbKcKbhmOzs+bW569lwOVqdtx9Au69RRaLz0CJaA79aq0ThjgWdc
JN1bnZdtV6/3f3mLCqv4D5qzLasbXL7KjC6LyN5en9GFfjumX1EE+4kzVuR9wm8JRGItvaI3yAAx
vzS86GwdnKoV7ke9iOM/vpyOkAVTj/EJuDlwHUn6lavSVzvAcZVBN3FHR1Nqr/rus/4ixe5hhEsO
SC5AdDL//2EI1sl8t/d2J64XbxM4RVxEfrTHkrKddMS/DuT3+t53tLpHd9iOylc66Us9CECIJ53z
Oic8kTo7BvBUke7EJGZp3KX4/mCASjIrPvHUgDecd/Fsqcm2rsnQpAGEZQwMuWvhAYoVWYwjwZPw
+cEyWTt8F8vExtJDfSWiwaONQxsWOno+qiaqGk3nZWfDKuqz6ee54P5HNHvRBl9qACbC06EOo9/3
pc5oCKn7uTkEGFLXsesoIca3D/fNNlgUJFkhaNDqqQH5UeqXwboawOoChPeO5RXv+HUdIvlH9IDN
kV3MkAWrfRv65ySHLVis1CUYUYjfN50gwYCoAVFLJ67LyWfr07//y1ml4c9xrKjeLHKSHu2F/k+3
UW6WG8Kfm0N35TMeChtKTDLqQ15ySU0Tyw5n7nh9hOBnhLYCaoG6cia1CEj7J+VsZTXq47yG/18s
qB1XmrtGVWVHex1JDN9fEegTdSFOMqu0lJ8V5NIgTQImhnlaALTPXJxzuWTq5u0LFgfb1OQ0Zx4Z
y42/lp+b34d/DAy0ez8fL2Bgm8jK2UxJ/D87cEH6tanPHVmRWTfzyZ7LB9J8lci6plw2w+SLq5KH
rMAfqgXVJgB1gFsDYdeHOQv68TpfmA2vlo9Lqhy57fRA5xY/i8SDLfppVczRuqkEwqApmIJbxp/+
MhI/UIsfFhOLeBeh4cguCHcyA9ZmiU7M0SzIfP0vF5j67bCLcOhBVvdLz3kwOKLlk2j/BsxTbZHT
bXqTgfa8awYDsJpT6e8GzOfmm/T2fVmrSr3ZT0OFhF7sg7jzhKwHdhntxF2uYOpORZNwek5knl/V
JQIb9WKH/NGIPJkoVLlzMgGqnBMC4PQaGVWxLyqhkIiWysGzxxXcEDNystyf0Im3vE4Jp0zxQdHh
J2/RX75LpuR/QNNqP6VocSfgy9ctWoLU0zMMrIixqDyn8MyBamleqqc5t0Jl6amaCiqxToYC0+SA
MMow/Vz+qSUtyvdEYnsLyuD5pUsUaHm+dD5yFcNuXwXeAZqWaTcAEkvbtJqOYd4hVnbcp86uy2LX
59VRgIJQiC7hV925QC53qgV+aLc7o+26q9dWx/RumV/4fu/p3odDB/QlN8aw6iBKOkJcjPHRGl3c
UlfsS7r8/ONcwJ2lyzzutpLZyvo0r5xl1qOkkbZJ/+qE3YsgUFRXSdJi6bnr1wj+rNelhwppVDCg
SHZ2Iw/wn/ccr4iTHNjx/XLYAph5OO7jojBFFvLiwbkshifDO+vl9QvcoGRS+QLuk+cSdnnDiiqE
sSOYWdZrx1Rtpui62eJPy6HT89bw5vEryMSeIqHLveMaRTOq5K3K1LODWrpMouapAuXr5fi5JiQd
bU25z73BbIJ4mC+S6QlW+iXmg4SmwS+A7M3XIvnqqLarVFvB6tYlWFRUIvRrhMg+12X8syONOZpU
8xaJN/sjOPNSxbVtrgxbiCFDiGAJ8Bi5vTC8rAEX8CfWBstGYr7CfSbZw3dxps0SbT1jo5LsT55K
n/IC6lTLLfSW0fFQJYTER6xO+LAecJKYgTrPwPanxxk+IZQh38dy5swwdRPWATrCmO6obnV+ToKD
hye6XMwA/AixQAxICOaEyDSPb+o3lZ41hUXlZuDeWCAl1mC40tFtqMEUCflEYWWVm/0s+3uzIf5V
yqvO6I9z+yonZyr04Dh4EvAlpoKX5OLD9X5BeS9N5x1C8oMIPvY892VF35Y6YcN23J9Rjn/yCfrP
GxIyA8IBLaT8VU9XnW0wVVZFTPztKbduKX73PMaShHQIzfvip9QKbuP+nHwbh2ZM79OS1g7sCR9k
/9iX/duIkmVFgNd1GG2y7U3r4Eo9V1e1G9Y9x0mgwHyxt+4Zf3fUvBkuKA/QnFy1f711NJC4vsGI
YlSYH410tlHH69fBjiwf7cwYyZ7hRDr17s+orGN6EX8ECeuzI3apn56qmPyCAu1SIUkb22a1fcpD
EtxAQTM7SxgzBUF4y3vr43eVsWFQgmAlVWF6ALx8F9v7cVhlCxXHMYMXgkNSdkEw9AHJT3swxnPF
mqiSvRbb7X8VH+0ML7M5pOW9LLY7rXGVXepBtYI2L0sIFcbsa3XvYVz5CUI9XLlci8fZMU75l12D
WAhhwjSI9Js6BOdkiWA8aKsIsj+YmRwC3pFY9pHlx8C4e2C38z9+Xa+5LbLbF2mm500qQ2vchQ93
9Js3bQ0KkvWMTgPa83fk49923FrhZqCzwFy5yXv/EcGvro+1hFq9xJJmDShjl5x0pppcMVJvu32k
FaQPhyhfZzUZ9iITp6ZPzUjJSS2mnbzajwIWlJpywsmdfE/uSGiQ/VQHNbDs51exF9HJCXOyvHXr
diEXBbX/Hwwv1xe92CUxRjaNPhCtnO5ebw+ahUKA4YlE01sIDPzzSK6LebnZLadES5XVI2KE/f7+
1TmcXIA2zVJmrIzx+lvAK8FgwYA6BJBO5JpkaT95hmssmBy1BBnO2DZJEK3dzAwMK9R+GcgwLilo
VsEICCfsqeaOIvvPWgP4FoCltcYak1s4aVZRzPZCJjJ5TrspEg9VjQayT+KQpgubbbQVmMVv4Hv8
i0gETUDB7p/cndmyukR0DcbF9vj/w/umTsoqTjAg3TAMrbXUxW77hBgtP6ERgq4UBggy5xuZH692
7wy13lC+iXYZJ3CCuIJQ+aytQ+xTOCN1WIUBIigW8eGeKEt/3izXnpycPnrqHOGjQ8W9xVxFy+4M
Nx8Z9F94M94pBPX8ucdIQh7GCzHa9mw2A1M//9WDP5TCL1xFxxL6Rx/81qgsH4oNdY+qQ7YJ4M89
pHfp2ezjAmK7QSfdZwrvOE5j01bEO4YVs0yvPLj6MMeMOde9PmDMJPwd6nwKlKDHztXHd/3o+QBK
u58sNYrRNDD1fHZTmxCYfxkGvGX1ClyH9fHQ+1K69vTEKBHRxt2Y9/6lNZSTqmUS7Dk7gKNrGUWS
FQUM/98dBhPHA9yDNIbYxcA7e4lTMTiha7xeTPRSFMO5S+HFqBNoMzeweutzLbXDPdqPN3KZarWT
g2YiVd4B+yFwCPR6V0hiSQuvh3wqm8kJ63+0YdNkss14szzffWnl1gqfCDBoOXJUp9o3QlxZv6ZW
FUf1bx67GxEfhR6VwFU3FhF4R2c44aABcktOGJME483QeHmgMQcJn+RrIYJJ0b1gB4XWtEutedhn
8Z7BEOXOYQpJ3oBKPDtjRznxZr1XVjLB4wavsLAjDhrjBjbwBmJdAwLL4S4WHqKzzGwvdF1I8W5J
aBLLq0dilrijR04zRy0R+DwgCK5pUJeLmsV2CEC0n/JeUDMbQVsFbQaNgysh3yRYCZdIqRyMJnXq
bkut+SiFsZquTZL+vHwDc0pxFoMgm7H+qLHyAsHSXG4eq4Yj6yrVAd1GZLDgEe7Ji4MvNW93tTzn
mtgN6PNWLUKgBvBFPfmnKoGSE9L0KnjCRNG4eaF6exqhY9SPfx4oX7nJrKKh53pUwVyUXEo98yI+
3ymKGHvYLulGQPXE0dqEJa/Qhvh4BFwTp9cDUIN8MiAt7xJ2uMpWv7qo0NMhMpkCwZdltszhnkjc
M02z2FpE6ZIWiMRoXwiET5f2VCZnzppkEujouUm/b3qu8YgjwHnmVyBiEgkwLEgLg/TmJW4NWEVH
uGy64p5mYSrayaMFupb2ejC0YXIrEYcHzxgRGdanFzZFSsviP7i0WnlMro+er0msNdOeXzQgdewb
rUIaCO3GMixAKnHQS4PgDGPugadjBv2vNZvXIt3CQPyfnU4J3m0kkRunGq94zkvz5EvAcm+MHI/+
38BSg5tnS2FFl0S5g3zTDzeGaEgvv6B5opZb04wKd32xZM60q+JBuaEWdf07pkRpH2inCcbXCZ+d
W0f9j9984lyu+9WBmpdymHGESsMv87GYYxBbMv/VVxiwq9aZLAO5Peouw8rTIk3+YVknCrqkfTPl
ai4yio/EYyYlfrZ5zW0ORdgMrYJbIX9BDCqAtcrxj5zInWIraJxygC1PYKYYMG7jn/grFwGSgboP
iv2jdwIirEvxm8/uI/efwvAKSpU3lspByknXmKQvf2yJGKx92QQ8OBBTkM9t7d49X0cr/dvamLhO
j/PFyypeis2fo4p7B/enrJjfKOXaoDcg6hLouZGb9DsvTalCgTRvsucRxy5lXH4r12xk//2oPm2h
WgsRLtZuFar+ptKQwTETGVW1bsv8ej5Q04tbIwPO/5lB+gUt8QXNo3hZYtn1834ydAk4P5raukNR
4l2r0yYdCoTh/DEHJtaQSLaJ5lo1xLUTmj16tLFiy7Q7KkM0xHOqU8IYHk/KlAO70+K6hFccOqAp
Brf/dtO/rvNlsQnKhqqU2K7hcR8yqscH2gMWkRN7kxEK4qreGNvkLGU1Au/BWNXHf303iE9fJq5d
Nic+8wyodVQxYqJ15yxtRpclNY0S9/zjnHeSWN9jFqP7B9s39oMit8ssIWhf0Pbsu3e5ns0lG6pR
fQMt92P5mIQ8M2oLChYtaS9kukSkvcNEeXEaZ2PYnf8ytOJTB8FJfUCsew5N/JDU0nnaie1CtUa2
nMN3ZJkpO15TjkQ7+0PECdY/DHVep83V+9MRYGHljLwQu/xIwEp9xUj+iPAhnmaGUcqyike3MkUH
9h2riAmv+hnAwskuGsc8EfJiEbNmgf4KTYzuCBldaWi0NRQRfFrecOsZwBrMvf/B173jBNtVOrsD
5EsAFJGQpLWsUdJWeWMY6m5PWTWdFIgjGNlsc3oohERRtDbUufQpaWfxOuA5uengjfObBl5rapuY
GEM9bpFAmejgtDT03Bq2Ho/wgejjU8f+XpyV2h/s+DgHfPu7Af5U2Ansp3BMMQXrMtmGZCM5l3WJ
egAlnX9wF9KZari1BUJTgDjtclV+LY10QXFvlT0jm+34mXKPHzlKOhz25YaQd2TyPYGITQt1VLDf
/EKqDmbCJwlA6VxmASJxquKF+Ngr71wFLgQ3SnlmULn7ZXRAC5EVWh7Ggn8fJQGtpkaWYpj75r5d
xAlfY+Q9u2bPbwsKJjqmPlMR3pW3e32A9jOVRHqS6iQPnDFZaVM80iPl8aL+6wsb9MSpIccJ5vd/
cpU7oS1/4PhTG5mRAKniN14dnWBlVOoFatfQZLJWGWrIKsDf42sVHf6Jf7QmCTfIxYZoFoLj1V86
8Zlb9AiQy5D0cshhXml7oUQ8c8UouQ0HLG8Ssnxi1uYUmUDgEJgKO1Rw5tEeFac0znHwxiNYEWSa
zUnpB9YxWzHNgJj0seTAFZ6+5lXspGbKbxdRMp3pJ+BguCFzYtqKHbA+gjIQDRLv6jaJJcAU8q+2
MRBwOP3y3gJJqdgjOAlVKGc8D3dYaRQAvyzeahEkKYNdiBcdDhnQHuESt8xONFjBbTOR+jTPDokC
Wij/xN29uh/9AGJti3eNAGeZRPHYQ6P6Y4zx1iBXEiM4Y6JWm/DoJ06q+7bp9D/eyaNWjsFAV+zV
l5/9l15dLCiyyA9lPW/yIJ/2aZzPb4RiTOMSZn1aFwnfa4OeT32kPsqsB8hK04BM6tK5BhUME+Ue
qVJt/Gnaf1crIpOqHkZvM7iR80AnAM46h47vpDciyCxpyzsf8qREIUKhBochAfirCDhW42on1UFG
LmgmMXlkvUYw9yvKlo9e2+TIf8vh2NCeeO3u5mM56yn5zVKNh6ERPHNKj9vNRibIoi5xyTJtc3XF
33aHc3Bi2Jzl28y2jBTvRF9wCIiO0dORm1DdVdzisXKkIJPTEjDF8CglahuaxPCVK2gVXNMYeQLJ
+avzDwtZv7kE4uWThf2+LCHLTXeir0sQsqjAOHdZt9Srnkl8Z0I15PkB8SA2acpN17XsaUqxfFW5
DoKYqAfZ71LXBSm4wFOc11p7yh2P+5YoOr1gQwMAL4/cUnrlgXUyG512vlihhYalhFOrOw9GNb8E
4A5AOGYQDoVnA4CP0/1hBf1CW3+N/ky5+zjsQba+Qnx1SZnuWtNxdqwq4ZBK67y25xzHWoNsGcSX
Wut2kTI45WKVFKTA/SE7XJ3kWIMuSTCDX8k7MM1yBtBlEGZrIdsk8Qor39vgMF5cctzg9+jtSPoj
dBZEDzqetWbEi3e1ZdMzw3hOFl2HHM+/6aJ0kLThRP3rTokawF0a7/6IKqD2KicUcScIshd3KNcV
ZKcuaYMFZaNZwV9sefvGDKg992bhclpP9Kp5dcCgNINnEsrn6IkZjGLd5J3D88FNVnJl1cAmd90p
/xEF1EVKSkQXs9ZFgzQTcxEQkH10JwcE5VDfre+CO6w8X+YgwRGsMvwdXFc79mQWIJRCSyRd1Dl4
uFSsTTywTf4EC2eNii2Hil/py6BzX1WdotKga1MdfvtExcw7kxRkP5DXBrNFqOTw60KVCDqQnQfy
edggvTRVj8v2PWz582c/UzS4ZkJMwl6cY894vQZJqnwdU7DUC9kFa1bZpcJg/SHWJnB+Vw6mZLq9
i/6Wep5/0KxDPRo3150GFSQEtdLob5MqTG0GMyr70p8h8Qz9uABiqJDak6FRG/H0jbq+5UflYQti
0GNvcDBT2oUiyxbXnYfS9Uiql53s1QSQyzDykSE94HzsixRv7y8dWFWGqmAEsiUFK9jmdRrVM0+1
+hauWx/SOoWlwBNzMixrkS4j5Dk96DMg3SlYjUCwN4X1Q9xGCEaXR1DyBIZ8HthxBpZaNDVjqQvW
ltCTAaArZ9/vCL30VIZRYLpN84HjDnQg46JFxsZF8+erR2czHY31jvobXdMmge32/LZZWbjIYXYS
GeWFOk2wjQYoEED3L9cpRBK4KkLt+DQ+qWnU1/PEzie5gZDCqLZE1ZBg1osTgFRVhtlThTZxLKRD
Vatr0r+WZE2XRc7kueN267WQuLX/La8aa3I+cGE6RmmP8YlSpNLuwzgl3BMeRkNDYHzkruH3R92z
P9DvrLmlmBi9vQITeDSzHSv0mY+7LlWZQhScChoa47ZeskdGhlnbcTZwo0r4GGlC23vd4sVXOixI
MLpWZJNPk7ZdebcjsvotVQqu9NTPFUHM1GqRKE/s76EPrbyXy7ybrsNPiM4L94e+WTQxKf+QVn6v
e9gB0DlWiGbST7z1ioZheYHWW54wnadBcGDyrOBgebOhKVHWwnGwtrCrgEXYlFbjsR2DG7IXsM7s
9gU/y02k2mQUw5fVi10AA9RGllJOGZQy/Kyornvju0RTic5ekkyTi39o9d/2SMf4Kd7IVNqSlyRd
Z28I+qB6f8IDPCrFqEu9WTlCFwRcVMUkZr2iF6X8DYZJZc+MBvEJgzP1DBypd6yDt2JeaqTzfoy0
8pCB51p/WIkqS6VSbhF46jyGFJy46orwXbNvkqHgchy46pcdiHzk0u1yAQ4N9YPH8Y6Wy0AyCaWV
ryMNl+QK0OcAoNqqRHxDL/4GmhJds7+YWKT3El0DK0oZhwHQATJzvhEBvHxsf7vaFfdirblJmvBz
dwUbqFitS3sCdkEoefTAuMIgL5+3qgbn9/spj9MLS8C1OJC+ijDv1ZaynLB6+Bf75N+7ZcOH2x8R
zXPyM4/MDxG8hCf50IYtiMJv/k0Ogse2ZH9o/Y1R/50gXpcGWsSwn1X5/mTvUlSEmrVZIbBYZ0cg
CrMzqpmwizTPPVzAtNEt8PDhKxNjKXCjkiojVuhKWNG6AcqwzRekH4KSycTNz7IuQBo3KmILzgS7
KwthAKh4K8TkuKZdJGWROR0b/KpUPsu86F06RJ+VDFPPH0gaAr7U9aT8n5e6sz5XLflCceitgG5n
ESPdYRvdhfzxjiH33uma6CjKRv3ffWPbivvMprScfkXwLbwOnrDyNhPBYPlPNsCOLx3FGKpSajaw
qN3lp3V/+mT3VAZ1ekilvLerLVSMr9t4wvUS/IrItbfaCNX77OAg99y2gp7JW2ekYlEcqzCUWlTo
wCXTeH3cJ0F2hhjCeYkKxgUrwtqt4rQ89hhyVBnnmoANNtEOvl4SIqqw5J4iiTWIZUkqooDvNn7M
VjL0Qb7GkzL5pj8GE6KzJR1ROFmKa2pege5p1vAqFvcxae1Seq95poD37A2Mjkg/QeCKXBCrPFOs
cZHDe0alyGxwWdQTyFg1IS0kBA5uYAFz0YlvpNMaBCi8YsX6nU94CJzz4xLzj2r87jk4/xoM404E
reEyfRLrmO84Sr5Tes0Oz35T5rH7zRkbAnU/qzZBJOwEd4MUQZ96woHMwThitGXPNpXwc444+mvf
xwLq4tAhAQ26VRb5BD7sXj9NJwZQS5EXGhTL2r8pYDEtGhrqLoisRONmYVJr6r7mmTsalJH3aYrI
SOhYBhT8k5D0MqEQUV5YiegqbpPRWnO56avK3lzTJS9FOmhIts7jfh8Mh32gHlSjwMBQBZuAfR+h
8Xq+6C+W0U1CQlSLzMoj6+HPv+SwA4Fhh+ES4qmeyETwd320yY/v1qrOUNhFWDJLbM0/2pMI9ay6
K0uyObknd7sXqaux486SUNxeB1HSWf5PO7tN9pTIU0Ey8durf696MHxz3KGJhNPBHI+gBX2o1sB+
p8HKKJb+sRok1hApEFiEEl6ljoPKogi/E7wIgkhIOWMgkJSv7TqHb07xUIEZAujq9uOYeGIK06jF
R+/jyJjOJAxps7PFFdeeUx2xRDg81DJxmx3NSOiPS5DcF1foQpnVETu+VRQnEb7OgKT/IwiCC4ds
LiCrr7wsvt72aNX2V74oAA56FQa75urMx2K86QOh+X/3VfkjQHz4b0RsEMfM6S4nEJ4JFtHg+UJY
SrpnjlbA+cpK7oyv0GOv5VPbRMfEvAdGk/5bj9+2qOYfnsYInkiuluyo2+V30GpzYayOofTdYmzd
xmEzhVQ73i7Mhbw3Ntcn/N3C1pmj9QvvJkffGC8xH/PNg1Fu/ujDWda3RpKn4a+aJI2x2U/taZ9r
3pJLjSClF4pOJ+TCWAdrL8qTD6XhkURZD2waaA13vYZK/i4a6RF3avWLloSmG7M4CTx/pRMRDqpx
e+CC+qawzgAewfS+40wW55/8dgF4B0QoegAIg9sbYYmoEKzgiMDEEJfKOqeFIRHaX1pzHo0Imw6o
bK6xZ7fGI/sd5B2iUkUkI3LZL6mNA9adevqhkK0TwcySrHFj1LrL+qwPi9+Q2EnUIpVgdwVqJAtH
lyun/3UlU5QJHEEC6CISRNeBGW+JjsIghcKJXC1znl8qCXFdKdQ2fNbZo9jrxJHTaiTFjcgfeFod
owNRM0rUaY94iQlOopAkQK2B+7fJCcKCuR968ZykdDtW2XDnN2fRI1nG1JlyLJdMHY3Y82uZhr34
24HyOWtMwdeSnEEmxh966KmbSr2EpKqmP6rpCgv+ODiEaZCrr5Vs2jgphmWjkBdcflFTKQoWLB45
So45fpUcWGNTvrIyW/j/aZgUXEu10jlMxzwHa8uJTyEqSf/sbHDlNQ4zfWoEhLDrM1sFfYzB65uA
Mo2mz54+55qRjuoHi4eilnhjNXXgs+y2TQ/MXPfv5SyT43i/jOyFU2cWDI9WTWNTmQQeQGJBFl2Q
MhFNlgasvkgykrgiufgvenxiqWNRtTSWrybFU277tuY7r/uqoNvKH0rIsgIZeGuj9T3Z2eX/PkGW
gIVwIrg6fUrvWBt2foc36FkgCn40K5qweiIWGthayQXKQZrOLWYhNoWqYGCMwOccYiTl7V7x80vB
2+vFxM0/mjIO9Wbq/Ci2cvVvP8CqcEvHo9YEAYPPVT7sVceRqFAVyliAzspJySCgRlLd07hxdIGm
OGS3hSYS0frA0qEGZDLTgeblR1IVGhWvckYkvTPNVgsihpbAB+u9Iktdwr2NXVNgZqXbUr/6nHxO
xG1iZsvSVEelYHrBgdq/rup3C0mFkzlXxX1HWpu7XP3oA01d6VZSkjMWBWJQF0EsQjjiujlo5mKG
1VUB+Twqgo+RhtiQVtGwkq74MtJwqD9GusIVgqCzKD3HymYRP9wJCBIwAMz89BQr6PjfO1Ltozbw
xVg78eVUbffhb9zEHV5Vs4CoCo3zTe7woRIc3xYGSuG3G5KBdMrOgpnMOGAZcMChX94O1wiipnHN
VWSxZZs9DDnE1eHl+rrmv8u9triZfZ8L+jCwD26xIsaAHYA1PKNwszqL2/9ysJ61mC0mcDlIVaBT
3/uak4sVFCKMUuM2Yj/URBWSx+4gPPLrVR4HSEFJtARgMXPtEC14r//HfKIyB5qEDLoDC1+/6mm6
saMQ8E1OZM1Il8tbVPsoTINzAbHoFQopFBlyXbr6vvDH697Fu6cPFp3+3KfsddSeBky7IyJy+H3x
YASyfrkWsfTjMSUwh6d0EVJUOfk0zN21FYN8wlz6VjpuOBmLHsGoBlexKtGppIvRdV7nFAFw64Km
0T/yqK33LpBQPN1WYtVbtplwj4yhMrX8y41SRXNmTWO9Wlrb9YPm6S9ffSM63ZF2c6oGkK7u8Fsm
Z1ycubH3GVE7cYwcmoN4X+9DhwREPDJITJVWA35HTcnIulMDwW0IOLO+dlf10V2o4zr1CP0TzQ+1
DKxrD29WDWnCIEUWKgkXPsZHROALzppLKBMQ3hxtxy33ZFElMbEf+PAqxOq2Rxg4bdNLnUlzHkxb
Ge3SDmu+Iy/+zat4XOBHr3Eoj+B/GOjxP+1jSYScWkg1WhdBoZdZPjpjUhhKf56R2hpKpu9hkapF
O6ZoCmsCqYhwL/2KQk9llx0Sca7OB1KeKvCbVf+lxmc+85J7T4Sw9k3tiviklOXnAc2w3nlo9JT4
XP3H0uXIVCBXEuZ3Ga+gSKGXJq0YWpsTwb7qdPh4XzsKykzHhGjhvKsvpetZU6AsB93MxlyVNKq0
DnNvw4CHPqP9OlaIOEuiHQQV1uJIsOqYmc/cFVCAx62Fb9xfwJVNslL8ZHxZ8KqaR1VVMtsUryDI
hdvz1rrBH3ht4jGI4rFLYLweaVO/hj5XHExP1DUWa6EGyzai+eXG8PwlTYWaZ7qk3Uu/tyC34mh4
99P1hD8VF3FE+lBLfXRkBK41iFC4caiIRBiKO6JyqgGyrayoPzduzoXixEo16ehncqTMQ5qrlByi
x8JFN1vzWavSTXeUAcZfvkOYMHdw+eoCvhC7HOWrYF5rUK8Zy7smOkVQ+ZCod+W9Bg4SIAD9yKx5
RSVJcXi4VtfiPPIyAGDzOQ6ocVWw5uUC3sz5g0lQE87vx6k70SQtaLGU3KyozNOvIY1+H/8Nm1NG
6LPs91+fxtEtdDAiRTOLqR6MZs14/bF299Wg7umjGYtlT5bT8biSMEz3AEiYxRwg1JMboj4DNAo1
vYZJxTNrTVi4Mb6WILbEtnY6Q4u31maN45t0F73TRcYrJrEzvwEf21JUNcA8z4uvVlHdj1U19wyt
++BNRsxpBms/MdIIMjgpWCE7l8kJYDPEtVoc9NdRRdg82xkJzKoDP7vc810AGpm/WdYz7a1QAcOI
nZPCSvyxt52yVFIFvbeoMXTPTWua6ctoF44r/k1+1Ka6uWLjonn+AHpiCoIm8e1y1nQllam9J/r/
DX8O/9O+J7Hd4MugiIePuHmaOzlf1QVH4opWiBrp+NiyA97pxjrLEtxrtmHolfiDcmcwECvKyzWm
Uyqv6WJ5UHo8oIeN8FL2OQr12wGchLIkclgSdbOkipv/dODYIlGeJH8MnAr2BYaHb0xg3fquUF9G
QqS/kB6Kd8Ahh4QWtVel23WjG8Z0mNbUqrj3VDYkf677TVsuWGxF8jekHOe28ZKh5fCcptxro7Sp
/4QcmqK7SX8QMlIaetdkGv2WWUU22AKBR3l2vNCqa73DP2zuiqVJbcXraIABbzSSWZbgfktA/zCH
pmpPfMnIoI1sSlkDLXNIyYmbXByZ7cHvJfGBPTQPszuurr42CqAlnwOOXt9J7qjC8qWa+uBiV44z
7FzkFm/ha6JRCnJPo4JhP0lzb2wZuD0QDRPS8wffwDC9Kv9VN4d+fOc7WCelPVnKDNrF96nUTDai
Fi4bVYExeC4SKP3FRPcY3For3et4Pha/7aktkEhS+7V/GkYX1pX0Ke6iT0uxWJTsTgr+0EQOFxKQ
NCVLuph75yuoMy0E4Y0rehSXdm3RMbL3e+l4ZkuzTRqoBbqMMwwBeGq7UJAFRhJbdMbg4Us5mGoJ
oB0p5rJtLqGdvUnmSn+wZlHqmpQghwIUONemZDHUMpTyaXbfYD7UkiSd7MNegasjJGJUVZ+5tCOS
97ESC6SgJIZyIPyXBiGYkc+izRe7goFo1kCmOWy332nCy3EKltQRU/IoWmX/Zfl5Pj2lBI4OSeT8
+zZaufL6Qw1l0Ja+0G86myBR6S9arCQQGr5mzVvtH9G908x5mKY1LXx4fSDL4FsHSINAAmP03+xt
Zy3OkCYgo0x63eZeCGXNxqnE4g2EDGbXs/CTK2FTIedsKbDzqSNt+7G0t0iWiVwevatigCfyccUf
+oDUHiPfr7bOmHHD6kaqQtZyUrdNv3BCGdwgVFPpZKz63w+W1EXVUsG4um62yjhLCv9AkRmJWYLI
mBHoswid4O9RGMqwmFDsm57dAolePdttyjcycMXxePy91PVIWMEvXfj3T0//7w5NG0yJoJnOg42l
JkF3l6VaMt1jy58uoIzZobDBNS42KmJaCTazoJIjj4szr8y28w5qyM3vgZQNkAXH2gObMXs/x1re
QchBOQVy1d59pTRY0rvWVNaLBYAOJuTtlf0Tjvp/Bm8acqalUm/Ml5Eua1TuoLjYx6wwIKhbcRLT
jpPRrP30f7ZlqZcYbtncBxLnnoMczSVhhXMrL3BzfKslrUGT7BBRy7e6vkfD4hr0PYZ2VrFm/EHM
A9rIYeqvGM/BH6X3spOkOcVelLjE75JdoSnZwmbO4QAMZj2ef66Px+WMezB9YNa2mPeak0LwcIaj
MSGzqZVPqc+Y1YnTY90rLocvjllw0iVcFBB/tJMLJFs14ke3hMZdQcKeqAkyBgcO3R7dHmhDkhux
9M5nA060QvP20HaxFgzrvdTyI5eAHSK0W8urRKJCj/1il+0d2pcFZhaYIVyKNbqlygwavlfnmDAq
j3gniB3Q5bWTaXwl5imnXKTfWqjVa4CWCBv3IgsvdFHs8o9rnbHU8bHPgBThQ6yiRw/9y0gMzX6x
Bs4uINVPV3RjJACfWUFoqdEniYgylYKUBwC+Adj85rrGrNjlNUWPij76DYH+gUYVd6N83G2vy96W
eTwmEOW/QbbeID8l30taxpHQqhtrJloX39U1zjspJAbtQGzzL/8/PRl+4BclTVEPHAgiUMOoDIc+
1XGb3SEOWT+pb+x078eLaicibn6/EUr/6pktBI7YpgTXASLht1imrvhdmSerwi58IpBbCcroALkv
1Mvgd1rWjrc8DTP/Q7gmKxSFUY7DU3fLv2rXuvNvzFH9+mmRmHd9XklC4t5may4IDK59AE8cou9Z
vjc/k/iKfRXAZEpHSYVa5k8HwUqvYKalkyFC8wBQNtjVYK4W3/eL2X2TcBp4eKgSEhcWDYRjBtGX
ZS5LFLpgd2a9uWUgjnyn1gSpMOSXg9QZddcGrpxZBjqnh49dCPAQtkRmc2w3swOeWLW7ulPO3Is5
5Bw3zhIWGiTUI/QY4FeBNVtzB6f0KKTZHpBjOKhzpgsMyWkFCr05Nv7crLXoJq/rwWuIJyC2ViD3
2lSmrv5HjQyF3qx7cmtWhZIW2ed/GMt4kpDXhr6B2m8plaqttUn3iPhqZJUmQs15txwR4fNJHqE/
TD27gy4h/ON4HzQNtUlJMhZQmaRBfBL5Mi2dcpHu/KeNaMFQNlBYIrigZmKu7Chj/jTZrr8V+icX
fP+wSL1qecDqUV3mo82yRZXsvWH7IwAwLVCaLNHrkasfYr+ZcrQujcuqoxaI2Z58i4xu6IJ05Ar9
J47w14qSUVJJXffi0iZn0rzOOoC8ujrwJ6NlhlSNQ8pkOA7zjZp5pge6TBTRZ3e/4+p0dER61ghD
F22uA2yTTHryKpjb8fJC3+gUBAtbuoZJHUtM4PNhpuFN6/Dcrt741gTUagfzN9n1vyE6MLWTcXSk
bPZ8dk8fmqmyUQYWpi6c+FBjax739awT/7LgMMyLENZiXGnbsg8D3Ld2X+NJ/44uIStUgmcn/QCn
D++Av2R+CaS7tf11KDYNVT2jW+heMbutrTAGekDrvXU8JpXkJMXFEqEM7orqz70XKeCK9+2dp0PC
YaHIxixiWFn0czpTlzlf85Oce1OG4/uigTwH2rEB50h2e722g08txdrbisZUcpANRsecoElayXGT
rQ3JpnRNL5DrVvijfDCN9KHeueTdrmTNCEg6HDCD1OK0PfDFjeFun2g1kpb9HjUrWQZpY0JHCilJ
N/Z+yqEOMaCuKcSh/Y/TuxMSkI1aqJz8mL6nbUXj05jln47zJVKkUwzHyhSkrf0PUo2Tb7SxPcwx
hmkcM6VtRp9dTqMHvFCqfbZmXNnH5u1gylKUzVorRn4caYLhbo1+wTAt2/tqpTkaNt5dYllVXodY
WEycTBd2Z6zvrwSkJMtLl/9l45Vk2qTUUVE3q1KMVHf+qT/T6MuRqYU9iMzlvGz7tINfHIEZJxwu
yn8hUdmuWMyk8wjZbzIT8clIkiZLPbfPkB5QO4AzNswO0FTDl5xvTLBCc32XZQVx/RndTYsCciki
X/yzFja7nm18sYOF01mvNTYTsRcl0BVDtktisz+aN282FsjyUTurULwcUDVsEf1usYW8YA5anXWH
noSWxs2dC8gOCp3teB+wo1zbDntFO4JPxQaVHkvSpSGa4a7NnPUJLQPSciZfAB6Xvl4BYem0al1S
SEpNg2eGSPRv5mul0PLi3zTdIyP/Xkp47Ioh7hGw1QWZ9eHdfXBFY9PRjFMJd9y6DybAB6Oi58Sj
EQqt2OjI4oG6QX3imCxGvXMP2tOJUYzWxvjoFLpd6aCFDoOE/mPbp/mzlZswhmPwMCujxbenFjqt
0iXrEwz/VrphvbW4IU/PMdIUuRGjpqY+FUYxzU5i0PXoc9weqHdyPis/jQzKLJ+tYGnkSG04DIV0
ZLU7A14Mo6h94jKDJkyK9D0HXUPhABPqE4XaCxwpYEQEejaY3MRob/++X5XmatgZQL2QiF2Cl0JG
QCQ+Hr/44FfCGikQ70HT7YcBUgg3HfMMYdpFk02Jnf4VxnBxcq305XlwMmM1A4OWkUpB1KQEKUwp
sJzjalGYzu1/DPqL7hLbmgrL6MuoXxfSnIXvTqfhHRFBMRR3rCNMyBEtEwnB9TX121GEqYlvzfW2
oytta7PJda2S7MKbLBPM3b7ImbGX5UVSOimIvp7WgWYBUtXJXqDYwiyO2yQwjYBRBMUxIxfRWUU6
pc6WTp+jzgEVtXU21MjxpCh1uKniyr5iRDQdCOuivxlfkLt43snbh29xXzd9DTqF2NmCrDqFDUL9
xE7OatAJeXhY8CzMZ3yVtUQ261G9L87xYk4V1SWAFiaf48/VXbHa2G/4kxEHzwN3yGF3ga05do2F
5xH11HtoSdb/8FMXt+DJr3KsZgvmoqhsYeX9VoZlH2Upl84FRtc59jb0ZEMybaIniPLMbO8lfFDz
DVrWKoIzh2EemElzl2ngqEQ7QSblwD8T7dKDirappMfFjskMUQE6ARw2NQDYSZBFKwW1U7BEzqRv
e9QuWBjhqEtGmoIxVtszKWgvFaD3n1x1Ho/ZXr7zrG8Qux1Ow0HRAeKQPhEAB0vF08MBzoUIRueO
kKx+RtPzJtWhwYM60TT7ep7raIFVOWzOxJGMw/KKqL94QulO2ZFESU70Qd0fLrqSTyb8cqThkXwB
Uu8iINhJZNDSqiTF2jiDUOOdlbW6UUWIg0EL1WfbiT5KYVQklFzgJV28fog1WqZziUfSYtx+7rlw
1iQIM9O0K6FRNWQ2iSkiEWSpkbSGNJVhCb/Tfoei+AT8tBBnIXcuEa2F9hC/jH3+CvIixSaF5lPc
Mmw5WxFhGvZbhxIGV70K7kLDN95EwqelPT83kprkIqJKg18iFzLXIMoeZwR0cIpYIeTrToEuxheD
MLZdff+GYxWoJq2nwyK4wYY2DzTaOntFeAgVMTEEHzxPgIQ1ECTMxd3Qo+Q1WXO8gc89AgHISIg4
455LfqIcTCczsXPz1j+cLAve+aSBv1Tx1+IzzsV08BYKJk7P2W/LCt8N+JH4QR7sFOuXVSy5oXr0
1gFkyD1LbFF4o8yv+w2XkNIOXew3H7x9Kjgv1pdpPNPiJSQJzDb2higT1rLXO3nJY+LppV7UZQAE
jpJjBsl/LIqZtXaXNGzNc+SYtxEGq4bl7yt6GnN9HWWdwKUzkwKNUdC7og/JY0+96DpTWEtfLm3V
ule/I9cvTCYIQaJ+7AEM+r9w41NrMQ/vL3et2CA5MmqZW8tuWUj8w98XVj8I0pTlFfhl0Y+DNasj
ES/k6SgTNB/DRRo91YREU1SiKJs0Y3uEWo/KqCRpO98sTNfvwiqMAWQSyoCHYv2/vB1txGk/rfe6
NRgJFtxWL/eoJSJFfrCNpVC235H9ys9csDvB3gbnD7QA6/WvEuqledpuTp3naa3UxTvvgktlNlxo
jlr1FvF9bRPh6dZh/GaiRI933LgW5z2+zvfyeXMXMUKvJ9Dbhb75ZIIO1Olm82cBykGqFWWmtmsh
OUfTkPTo2/2xJ6BdIRyHkmsnLUWibcIHs3u6sLeiMFRLpYTsr9WKYgDOL3So6gcxRNvBynTYxALu
tI5zkZEZ4IXJgRGNTw5QFbxsNaWu5qQJI6Qlfm61+UsAbIPyLlomrraME9MJqChCOrQWYAEb4JoE
C1Bi57WNkBF2ID4gAVmJ9mtAniMSwirLeS1qH0yp0gK+YxDCngd55cFNoeSvfcZqmB+uTyDesXpT
QBviJQTXsXV2Q0vssXe1y3PpZ9mlq59APVUu+AICeOLxVA/izc6yFqHrHqgWYA47zO6nirsP4vvQ
QF8cNKQ65XYxOWF8R/CXSCYRPGAXiDFaoISPvi+qFVHT/u7PuQO/U5QWx7VmBrAuZk9yrhWQ2RZb
FksjRIZqFrWxV7QSOnvaID4zfGi13xO65x60f/vB62SRC3R0rm8RUfdMkC7IdC2emiDUfizhI5R6
y9b8fq2bZ1O59X4rr3hituqcn3iODWTZo5zsPzZsY+tbM9wkmroVVgFdPCFu4AzUaV7+s+/gke4V
WDP4MnrCnM6IhARsNkPZWTA6PURvJLsdyTsE2bIYYQ8JzKIS80sHYTTtw9xKyjvgGgmkHhseRTlU
2ivBFmGCONjrbWV1y23aeN3VYwQNaNHPZI6QWq6HvpmVpy1FREcfKncSia2YkprChW0yEX9HVMQh
LKHgk8ErniybX6+9Oykotw4Vt4fD5AiKi5pDkBx83jcawbp6rkfreA2FBhM4ALCYwEv8Jz2/+2qU
+vqC3fpRNwofdJPxu38aJwLwQU+aqDTPLeuCw2xw4RvXZpHczakbV0Q8VoAnQIAkbUwm6h61AzVZ
NR635wDFcmyfS06HPZUzWdb4YznR9FMRnNtfY7sd8IlhXFrlOD0NGhZz/FACJSDy2iumFJ4LHI/Z
rlP/aM9HhH1jA9CzJbmXtCLyRm6tk6jONcK//kRA45DR3nK9atF5laHIFFWmjxHtPCHEvu6bc7cf
fks0vZ7OCv+BQbHGeo9fAoI41WZLUkCgBfc3fau3Cky7PLEpOgMi2xyrL8TmKTN5Lhp/rcBUUy2g
7HFm4UeYivluTlj1UWvIiBLIBskjim+IKP98JvnS2Em8u2+MhJonKfZPflUNF8FloPtBkdQD4dzA
K8Rccqte+KW5kkUG/WjL7bmDXCPVU1jIRSeHzkCO2nzKh39Undr6dtx523rMZ0RyNZ2jR61+FN9/
HgexneD1N+lFsnm8+eNydqRQaH5URcl8tTu8/hcNXGA/y//DNCRVkjxbxJw+jHJ2+F/VwRmiXDJj
GZIn7qcr83xJIfYp2OQtVLYk+OYxoa0coW85YJKFEKl6OxAKhXFQwSjqx8HfGrblwhWkxbxzc7be
GYVqzmILnphTyS2xSobOVL1FdbcV1LdsyTaMfsEVAyIHOQjOY0rCFG4Ub4Lx2aKO4P2Zzna9plaV
Pg2u10nYwMc1xsswWdGPUqITxBlszMa9p0tLlkBXVNf/3Q5SWw4IiEMl0Dy4IJ9HKubFo6QU/OyE
vMF90eWE9qOE3qfiR684xO5MfSOrC1qXChXaHhd3pMqpk4GQFqrLBPrjv2X1KIm8KmWpMYEZUL+5
IpijEFpFwebD01JUFV41QV7+d0y5dpT9qczisPhwbLACmUQhrZeMQJDIsRGiyNO4k6bS1fjlpdhm
PwmxpSOcu8TkPaQIQt3XAVChOdDHoG2fAh0HLhkkOiSp2nZCVNL9vbnKih+no/kMipYdl36ekCkN
iO3ywDBIisQV1OltVl9b4ORwtu+7+u1xpnIDDSIUneY9g6uhEBV8muyBLUiF0Kssl3C0t3qsGuWi
30RNyXuU6uNiO8rOXr/rIMkZlHgrIwiB5xWkKZT9Q+BXRLByaRVvYuANlvm2EONvs0c+VF2ntohq
BExqvrObRAHd1bZuz3yVDhXG0VFsI6jsUpDKSGCcjLR25mC0A6x9wB+I0Y9jVq+FJJS3TIgLCowN
gDCP6mCK7TWavn8tK8o449QC4rt2kh3vnrLg2hS4fURS5OLEA4cbLF9oiMXMrjG4qiSX3TPZfCee
fRyqtF8dyKMdXHha3IejbMZOULOKs2V7Bl0qdp3DWlUUUXPxi3xlXPs8E778NiRBn2CzqqmwxYN3
/Qnd0KwkKqYvSrpvmGsZhqHQAwGzlWsKa96fHs9aDrYveaQk3JFNh+3Z6LkMSp3pG+JISBp5dU+Y
aXy9t8URlflYY/V46a2ymTnEvZfNYHr2ZpuHpHq8meQfhvTzrf6tFeA53pvlj6hC3y7y9TYs8q5s
A2f81DOMHThqBjmfgusfNmgxxWTeOOrTcryp7EkBqMkMB1FtHi1PYNHWN/Caf6IDZ3Nsv9Mfnr6N
MC8WiULvN/VaoBn3/6vOablbL23AgWTrpwjq+pTD2kyrw0ROi2lYKi6HCj8KJo4MkV3onMlm6ODr
qBo8ReOAeAG8CCHBlEzmiSSnVG7xCxfyOdRbmrznAbT/Wh8dgwQE9lU//d8ReGp6hHoWLT9VrnLC
RhvVsOrUi57gas2H65UJTS+83fxV9UQ4+RuaB8U3xR3jxynzvxNopk+ay03K7PxOFiActkMe1TYy
YsMJFxwIhoVYfC+dlQzORjLy3NxyViPUzhcmKyCZmuwyKjwmk+xE1JQrizD40XnbjFvAyGALsMLC
K0QIHcGriFA2+aBhF12txbiiBWbqePav6xJtpDUSvJ0MC1kztvafMVmjlWiinguCX7EleucpX/dn
+A2Gh1PWaE36PTrRbOzbr2IZtdGBWawGzDTyw74I5AzCmNeFJn3OHJEKKXVtJV2PsP4/nhfIWsFL
hW0ZmkF61HEmg5vQD/6ohDdFhEezHCaJsgdscMxv2n34jEaq3RicR8yXRINi+lB4VBCL1tzBRazK
s0PSv9aCnDrctJHCrO5WJOFZ/QdyQllMWUQh9znfQ0RUlsG0CYxjK+uP+eVX1k1JcYXBJKP9fk0G
64URteLB/dI2ewVXUm3zI4mHGAOtEJFUOoU6lMsuWXBeIVsm3OUmm903BlEM43RqzjGJfVYbJBij
5hRkCqV85a4rQiExhBjEx8iJXTY78BeuSZVAgdgXYXNfjFZ5ptBVlU6zkpNMpSKIIYMjnX3jK/Ey
9zCIIj97njBuyHAB0/w2t7lSBETVWSOnIH1foze3M2dDKFjSSNaye9043WLxwbtCM/OtmaEL+6pu
s+vHWiljAaw7N7UGEO8y9s4Sw7tSTXdFNg7HcGCbogbxCTeFHYDXPrRjoJ2maXmSYv2g1CtmOkXV
n2pJs9o9ttFKW3MbC919+KeNfzh8e6VLAuStNYD27LqBVoJsaFU05m1e9GpbC1WO+m+t6QfrIOYB
POC8/F3v7wEFYTM3eUbv5dgQi2lV3zVTfOZt9BCT5OIZ31q/Vn72U5b9it4HZgABCWPK0nMHjxAE
e7E1BDymP+EmbU5j6ZL6Z+fRUINfoq8wZSYJF8A29uWdPQk+zVS98ITf/RHrv4PJXFn0lFykeX+I
Mebrif9Ose80Dj+RgA26IPySMwTnRysLnyaaiZJwKifL+WFHD/dvwaPgMRuJJyGZiKAqNCzJaY0b
FtKysaS5MUI7V7gzqycLRCFuZ05VKijCT0Wu9O1PLkLZPocuwgKcVwP8vjGF+ULFh2Rhw6Jhtgds
ipCFMhIc7iGncJymvDDpHkoTxrQCAj4e+AiU0vlIeIzE84YRWmwe+ltEOBCSsJtQ6iAvI5qm/1Yh
eXpCNPmYs/AJU0e5WFdtMrjn7oakddVKL7TxAoWXBh6q8CTBedn032EhClf27GubFcme7Fxk4jiC
4zIztt5CcmqcbidSSRx0G2xpIvKs6raugbpZlMRj0rxqZAGl/7+ZkqkI6gSdZxaN8mXWNwe/OVNT
d2BxGIyo5hNZpytkf9E4LoPWOzuFS4a8nqLDLgdnXrCVBC93NJwi6cGaZF4hACjX0K+7PFqJ3Eas
uVW+v30i1/sBC3Oj1lurDdl8n5kr8PRy4iQ6K9laBjUcNDMVjEI1Xt57rupxGqbuOuYZfREHEpI9
JBojUUMJv1g66BOlgTINzCTk0X+GgENwPkLKaH9wwkCgC8d180Vn0Q3+xoMX4/AHaoff8zKKV1X8
p/wC4LKtg68iUE+rJykfkKfBi0zo/QMXB2aRWVuyS17b1OKyiL0RxM0rchC9equVSVVLC86tRjYX
qFkKBjSNp+Zj/xX8algLJqmov7i+ji4RaII5HxSCQuWqzzr93t7Y6S+GvdrXs1FHHRug80kVL8bt
82Dlooe+xb+9/DBDWeXHnmRSqdbppa5SLCdEzDCqjDr0G/BSfUqF4aC7p6CpZj0zXIKJdWpu1ZzT
MThnZE76eLqRr2cOe71hSsh3RhEXLwSd3xgkUt8VgpDXXUlljLoax+E+15rFNMDGsUJUR9UaC8wf
XLEd4OtosgmixGX2D9OQp53680jtsFZWvyQoWhcC75Fnun7S8y/DGnd9Rtg7QJ/NaijC4eBDd1rA
GeabgoijirWZv/SNoBxn6zQnTPcQCTR6el/OD2UsG3SFEfAbe2rT9ed5ozJffhgMFrj00CWeFQCE
b/rxlghkVMMBUwl4j43kwSgkXduOLsQTRzmB69QpUZNe890JwxDt6Deq9DDRmGqXpxmk0ECbDpg8
EEImhPR1RmJDHV+stJ0e0+lTm5y5tnqs3NEnJglc7STZJZ8iyByCYm1P65EFjf8z2znIqf7VIu1/
DQ85pu/bddrUTFFqxqink6qK+mlQXdoZ9+qHp+Gl/GkGorhIPeW3iCWeXOuiT3wWk8rL2BB40zIy
qphCbjjNUniQqDBFvc8V6OusltbnydIp4bHhQADee6/I6Dq4IrzucLwJ+T00pGqFG2J+RIPlN0ba
wlYTXnGqK662ycvGqtqXjvN+eiYMeAhGC2l9wnAszKyYOK8Gr1cbTOPKWu7nxhTuHkoVoBsNcjix
aimsSS+jtWjZ1el0BXPCxmQ/1nTFqwPaRBr/z0+ztu0omhF6Lq5U6SjC6ZdXatAYtv3g0gQ3zoCL
Lpa6mnr218Q7YMpE0UEON8CBTVv8wsKKkhTqTYc86cBt3d3ZL+okShTXru+566f3ueZ2gR12QK0E
vQSYe7sQpO0ztk3Y4e4KqVdnw3woHGE7JuzfUqk44q98K+48761xHOxzkYs0pryiK8CEy8osbo1N
4fD8NH1Cnckd168yiGMZvpuXOOo0Yw9k3NSO5a8uS68s1Rh0Hx1TgCICEKg6KIv+hFyeqagkE39r
GCL+IC6WQxCG8oaDIvDdRpNRmNIMH2OVFJqY9654R9wLyHheLppJXXAhvFXIB+qjixiARSSZgQX1
PvQkeo0OKSqa73dMWMIRfJG7MMEPY7MD6iqncA6KkRAS7MtDJCMJXv6WEw5k2P+4ESfxcNh4qPL6
g2LBlyfQwGorsZY+7EI/sqrA2jr2jLww1d3gOK8KoqHNfy6ZcZ7KmQs0/y3xlu+YYwp1NUk7DtaQ
vRQS7kKpz3QlY+bEdHqp3jTNv7Fq3Luh2gxdCNEiYBexnocYruDtxx0PkRQLU1oQnJ1N3tbfCRmw
azRkcHKkAaKu3cJqAeUeyMhQydQmBo3m27LQMYmym0WlhqWifyuhG+FwITdt5ApnbvzcAGynt9CG
ukOXmSsE8HnzSsWUZ9tiftbCHGcOBUb/736ISGyBZThRn+kjZ4WHoT0xK+vLQGNSbCaiRL8WNzeV
ykKPlJe89crvjld4AmuS6ZkPB6Jj8qsm2bxPxH5wBsfKpZHaGMAogtdWq/+kwEv51JPJyeYAQwQ5
qKWkCZtppXW9yovS0lUHvVYkSnWPi4VuemMNsdNqXAqwZB+87RlZX1rJ+MmDTZTnyVnLLPQC2DFK
hqur+zMM2zaMNk72Q7wvib8B6A/ej4UuMypGvX1RAOPNvk6TIx1bB66QS/c/Xi+S2gepSss3bRNG
MwvjuGxXnuxpgdG71kyx5CojnAv2BGjBk2922Gs8+ZB7xRiqoAn2T0fCWooGDAbVwdDFXNt32KOa
iYLSoI/c7AE0Yd6vA0Whrz5Om14T5I1gjmrXHw8b5SQVewPzXXlYs/xG7yR5ZKqXLDJ9chnU9kog
E1tr2h2V6HjJSAP5kXjEa7nCSujbr1zLAtKEKmGW23a17C9sj+pikX4FcGWlMG0wSjNoj7IijBSz
veG6Y56F6zMKxwKR9HPzDw4vNuyJdxVhgUaI715zdiwKQ5qF/1cMU9l9ItCLFmeoOTeUWwzvx2iQ
QG0qgNznzKxaITJMKMC7/C5pJZfYkKaO2YT4AdW2Fr5OmPDrnjhlrVnYZ74vgdi8CiqgxkaJsfHg
2rX715FfGjKoGfync5H3Y9FgNxbVOB2QOyoX4SyHtGyxut8hXv7iYDpz3FaNv+NDSRjBHSGqOleV
HFfHbooe/eqB8zdhC5sEE/zzzEZwwa+keaOBJTC62dcq8800UqG2oQZKUke7a/lqWc9hrkCMft3a
ncH9xPR2uDWfQuKasNRd4wi5oYWQ5djadIDOvvFALCqNDyq++Lk1u0VdNww8fLgbXe/ZVJOIUe8S
R3CRLQijoRkrcAgVRQUPET3vgycJ2a909vu3MB48jRMZyoHyX+M38HPV8kpMfDbFe3jUmMHYWJcN
pMA0oe25yX5zl7s+Npy44Xc8YfizQCRRxy1bpxJnjDUIr+xua9/In7wOtn6jF24wH7sX/s7KVLzG
H/0x/N1cexCvDDhq42oBYgT+uAh/SM6/ctbTFg4N0vhO8qlxEygvFxY4xOux9IpD9VtO1C7RZEzl
WahrieImFr6tnrkJX50rybeTfJad2wD0F8ZXdHsDBw81MhhqgNe6NumAfR6qpU3EdQg+IYB7hU2c
g9BiGJSYx43YFTHDid/w8kk4w3yY9qnJDoZSNwxYag4bK7XgU0Q3wJikWUPBNtHnDCCEAwX8pdMC
CEZMcv/keEGt4IHG2E1C2+9l8kH9K42SQS4HDYER98j2m8/bigEnQWjyuDhqw3ibEwzpLIgFgyCb
zcCMxInZKTl6QXdEPMXjN9AJKNtKUsPkipH0C5que8/yLMLEfWnHVY8Eys02Q4XeymmrJXEnKyqX
SJLXTAL9F24/A2ZXzDogiTSc2dMnbZtVllDzFuMO0UnzQgeq8mdEfWaci3H7xXxMf7YOXF/9y+Ut
5NmVJ36ffAezhEh2Bi11r9jyKpnJ2Un+iEBGB7xjfh5rfvVPb8oXmqtekMdYBNFcZNH2r0NlByGH
BPZD2RcUf8qyeTCIODcgB2qnE6rydlDl/ZvIMX3VAWkEBkpr8+Y9SSlYMbPtEWNNPskUtzqhiCQ5
3nRMb5Qh2uJGLicbv6Hf4yrJFyOavpGdavbIev9EH5rkMrBMMGIcM65Ma837RHT4Q93ymTcT6A5Z
fFhw4+7IvZBcwv0Ws6+S4rAC4pRFRg37IftTs2nEXNuLz5+CrEasa7PxvHvfKhxyH6/If1ichtmu
hV/56rOULdBvrckOOodsLEJfcMu5LBp5gnBRSWyp/x+QdqBVU1wYoyyV6vc2Yo3JDvU8WyWyoIFQ
ukamwB0RRRsykXygLcDD+mzakQxWULX7qGvvt9EHzW6U6ewjUvE60Sc41QW4muGVJDzyDpDR9TdY
+mNF21E0DAn2uGrIRfTqJnilT2QqKGWW7XC+0LZlgqwo/yLbNWgwzitrx2n9p3BrSWFFVaUqsahA
2hHjfORqds1vpx9T+zMuzza4SsryOxhnvZ9cetT50B6Qveq98N2c66feTo6kxSssLoIFS86qPTF5
01Q6eRCvZlITrJwh+Pn1lwVrRXiSh/8nSQeM2aUA+f+EgWi5QSZfqGcEked2SoV5NUJPJKa+Znaz
d4vBltYi6CobwUyJgphe1koAFcCDnUiGQvgfK2bJLCMqsGeSV31AgN2K8JV1Q3HM/f9CKXaokj2r
AvQeOJTAvzsk2SaSYAyZxwnVMNhPvoj3vTlo0XMfdBcZ8mlHrMnWF2RvKc4QjOxineO5IpJ41imj
yEkF9IjnuV19xJwvThYq6LNjsgGMaOzd5vbiAAU6mk6SEJouMWpZDfMm+YIjHg5LQYjaBz22XcIZ
hwtep0LwX7rEvOaXEQxdj2rkuv5EFh+ss8DSrgVFPHolbJ4QPYWfPgEguFvlulfDEgoDshIvcaTn
/V1qHwfISap2GZE12ML28wYW5ryooQqvmLZ1pHFjs5GVMsNZLDHGv4ww9lHocZRx9TpBk2AL7Qqe
ItkLLxmT3QuuwenqSc7av1i98Onf1eOalpw6eBTcMS8/8KERZV3h9u5nF+DFm+wIMuKjnt3Nvrxc
8IRYX1RuG6dXgNqEC3CsC2b+T5byw5CJLBH92IhLGGAuw1Xv/sNwPq8x+5wF89QfnUlbOSd1aBUJ
4n8Nen+FD7UtUt/EHotOXFRbopRMnshMAklYkr+noUyApRQ6i21DzpGmJFhzTq8WoSoV5DP8Mz1L
3Dvcm9SlOqMesiihdAOWvt64wWh5ZznR8Pg+ZneQj/ZfSqk9+mSB5VjMEhuAx8YKDLqZddcYt5Wn
GTlGdfSdlvg04bJhUpBju4kLO0gmP+ROO0acDB9IOkFSmbQ0cMna20jrqoY6BJxc6p4lC7TiAiq9
6OGWZySeqifxdIEoX1rRJifjL7Reelz2nU62GoMUg9BVY71TdjCy1rgnxMqj/LFC95oGdzbmI9cK
puNsQ/pMGk6rtbhL7Kv+svwBz4J/cp/s2OxVcG8sfhap3i+tpknfEn4S0q65rW2xw1daB9huXJcm
fDBAldkHyvdKEmhlvhHmTWRUEL96jZ7lt1ns0ZyjsdMpD4syNQHnTN6gq0774PnRfUk/v65hfHPX
/3AGtWlBRwlOKRD6JbRW3XxTPSnbFzPyP8M+aonFJ+xwEZKjSMGMmBk1+4ahq7Jccukxn/AZj3i1
r9P1pOhA5NDir7lZ9xsHY4PSH0QSaoc1WiIij1v+asT62cMnaGkbFyqFTHrhKcn9/ZvxQEHzG40D
qCbrdORNDSyhds7TlS2trQts7eaflDobINexhZ7VyCjMxkW9GsSgb8F9EOy/wlByr8a/3ln8C0TQ
rhFYm6Q1abI1BseKXjm6c/9tQ+ZJsjlfKdfCYYGNHCKpMbSf+4XVRmSaSmhu7p31YKJiOPAUBW1R
NOm/8AUZ9nwpzy56CN06AAGyAMgWVOy/2eItZt/ETvxKLFBBazPhZPo4pD8BTvZGWVJtIei4fc3K
zicycdkFYBahWTyM4Tt4VkHST8Tt+Nq1i3yOZVi4O3rZtnhtYRzAPGKR7QeFdD+qF3ORisCJfWSo
63X5/MB4VN6x0jmkFp5pPxySJpp/PmHs039vLY0BNtEc1ULqQEz4m6ij2x0I3LwCgClnaJMVKe9X
uBVsYZCODDBMjItvpo7kB1n/mQFS+cEWfMvHf1rOydEP/LPAORq+enq6wYKxn7Q1Vg6/kaYrhfdx
Gm6STlwix6RVI6SAd2jBFoqftymAO3WLuaA7qpC8r17J3b9K4RIh1DMxlVgH2WPvGgyrFANTh1Fc
GOial3xgirOYe4jwXvZ+0PYzI7Fi2oxCSenMgNxRfa7g8gUU9iuchtm/Vepbc0vPEzJkwu4lDCt8
Nl15Jig5gBTFNefxq/j0WdVOnyNkH8k2j/vpruUnevcZfV4NKqLM5Lu+Lf4FXcpUHNCQJ4GUsVNo
7rHy61gQqD0QgA31nPDa1RcYSmhKrNomtptU9H7zXTk1+4pSjIVz9isgRdZtK3eux55brxNwqbng
FRO+7m4LqOmYCnwyT4VvWBRJu3lssrGZAO+9Sx/DIa/M2ufklkFnQzMudKHSpLx+KKQCPbV8WDgc
Y0ypJpeGKa6QTjZF0iZlAgJ0XIi0hCtYji+ZiQsuTgG/ERSAMMgWVrz0rvHZOSa2ktVuOLU3J4YR
oRMUMvlwQgVKhpsJgdUkju5TBVsaIZgOagdApATMBc+XsB3MwdG1uPDtfPjrxVVxP1Bc38dA8AAM
cYbNfr/iRcz43YXY7VtOtr/RN8eQFH8hXC0huaCJEG7umvxynbC0vXz+N7Qm0CGZGHuoM+i2ROvG
mabLcJKa21SSwsa/vGEsf5M46OGl6qTJUKaaDGzOW6bSEmVJMUNYDtUO2FjmTrVpQkDvuuz6HAT5
Iig57qWnxGohXqqu7L6kMoFcvCadQhFLSLZxg3AI13RPlcRbarL9kk9E7L9owjkw4LKasJ5wr107
cBQXyJImjmlhG6ZXpgP2O8Cb48gaPAPf6dLh+wFtqKB66SheN32aP7q10/ejnSwFZbZQuB48Fnpy
GkthJ2tHo1y3kUIRrEvK7SZgAaHhPE6aK4QiGRE+CVIrET9axxVCfcqvTp/SfNKSVbYduYFIJbmK
DEOVk3jbofTen5rKg9WRnq/VYKDXmQ2WaUMeoaFtOuXc7i1iRAj54FgbOq5POMZmL3SizyeWyfoy
exWArIiprStud0n3ns041dFmiIMX48RHbl8t+JMdGsLRlfcWYtzDo75pR1bYGhD5myH2PKkixYEz
IH5Bb2qOA3kcJ40+x6JdH8ji8l30nftsv+P7v5DOUE40KzS2fDFDCVcKQo4A7VdUXxwKyGt+yIsa
OnKGqDQl54Z2G2Zgo5Lqu12iKnrgP0qASk/CtiTIs0rV3owJdwWVITqRU2j9nh0G9L9fCJn2+EOO
Gf4FaV92u3o4S4qS4xHFPhVNFqTFdHj/lG8taLuDSS9Y5oCHnJprvHeG8/O98dp11SFVxvijdM4D
iUoxS4bKZNPwq365818O0l4AQieV7NPPSL14oRj3poCsPyx7JV9RGAD25LiKKdQo0euA1zmbH7CI
BPBicW65rDFzchMFuuxoY9/MnpjaTakrLojy5jAb62GBsV6ZH82XDU0+oiLdL1DEJuTUkRBGpvUR
J0+lCg+TQusPlJplejYhYVIgBSqASKOMdA+pnxrCT8iYNEwbcU4UDZgnu4y9zcTNtrTfPyZdw77u
sM6HKtxkA3mGwCGHXoHj/IzwAcUGJn9LgE8HTmEu3v9QQZzJWVspYUVLvGBJBZqxV/5wEp85wsJ3
xpvdNffzISqkMwDQSAqt4hr8pf1K7+LEKK+3G4QRi5cXsCunDrzNKtcMJfvco9ackadfqLzVSGtn
T0wj1arwcBL+H2IFKMjwZc1LN8BFbA456TyMpOeN+1J5tzcLwmuHs9ur2aIoRcy/RgFj7spyGRFS
xJ+nW1gCTw/6V4m+ZzaXXiGTqCL88sqG2UeUacJLS4mGkwosEIii3jcpLM/C3aQnSuFLS4b4cUeV
wbPAz3yc46b0QkTET96ZYUqPOQwvb8tUhkfjMGCArwZCKG120bAxTt2skZ1BpWYpbb6TGZTBxk7Q
LiT9DOjpqbVw1m/RX7Q7z9dkLtsMJqtQDF+hrFCe3XSC0kUT1JJibUhwC7anj4WdsbssqOmYprmS
G4wwHt/TbcPAKVzd1hVrjAiXr3JZupiGlGmRWNwG3VULcJqMsfi/0ad/XHoflSEZDMZDhD5tswlJ
eqvAcf5YMYci6dHcp8OnFXhl+cCadpY2Qmx9TMNsAsZF71V+d3pm6keV4r7PYK9+D7G9Lf702uju
GShV7zpfI5Rkc83bldXqnIhIcGVjF6h3kotAzzlmn7+GoGlMptw1+nd39qNOAy6Y7Za2NqI6ti3L
5EKXA3hGzqMKwmVMjlZCJkaXEYMJZycwgmFgL8Pl1SCrXoeb/Hy1UDYSYZNocE9K7+vZiC8PMg63
OYbKqMPc/nAuDEMaCZAiq02aJqwIDvj0dhNdjxvSbJnGihhJJxcGoGpBGalnLmX8PSbTT2lAsv6n
6qT60PyNLYerJARCWlSrrRknA+SLaIoG7WwJ0bLZdJkWfZnVyiLpRnsoKMIgf3K3ETXtgsIXszGP
4Z4NNN5qGPLlIQiR96mZt1nk30F3jPof9U3zzDeHa/RsTn7sjdfnDavl82OPJ3v/fDTahyzJp+nn
obqKKNoCXC5dEk8BESBNQv0qBD76GborAbTTIE2myiYV6J9j7LieqxlO/x99NRV9Onjwo07HFmYA
rFqgXWylYShsa1kqwVZjdeoJGyDeOu5jCBTDFh5HeDTsy/nbnIRXCeU8qQCqXQFEtOnFL33Hd6dW
j9eyNh/VUR8qiBWN/WQT1j8GDD5WysEe4JxsLsa2QJp0eRbnsa/DSNiszTBoNm2DwMOtuNM0DVEU
HyTBEQNiTNTdC2KaNNZfgxkJHRgKZQaRnwRJhjrnlToyuboCVOIK+pSKPSN59ZrDcM6rkcEy0rWd
+BBajY58cDtySj1WWQHixNQnaUEQ7EK8haoDBica5G1v1Q7/UNAY9mBpw+IkdABjxfWiAZ8ffo8p
hMcF4LxGyX6uSTYHnwD5c0/SuibD5AeRArz28WqnL9IQ9zgVK97eJCi901CiFO7Q0WjB3/9NJ6Xq
+zClgFy7U+qlN6EOdOICG8HMoiM3+qQUJdkq4QM7t+PHBENiHfEwJVZZmUmz3sTw0zTVr5g1QSfb
eVvODnbWB/YQgXg4H56yAtMyiM71s3E6p7VIzMDiEfn9WlB2kz9+unGU1PFVFYQK2N0sogArhaYD
VMrBHXQHi4RvctkKxvEbgN5DekoqYi287ThOj55nhYCT71ANw/Q91Bj30XjXOWO2iAxk9uLQGGx/
Optl9s9WVLJ5uyXytSbX5WWGPJq+yFU0c/76/8cNxfHT+uT95XF+I05daCfo2HlaHubbN1Xq7ZH7
iXqLDiQkq4tahhDr401HcjbqDKsnJQZfzo4dsIAly0IH7U2nFf3fdAtVdQrrMjQMvqlVPLdcdrZf
DbcTwLqivF9Jvsv/7LcQe9/X6+x/kepU9qWM8wIDM28SQC8z5Sl9q3zmnxb4PEay9BX0NZiJD2ZJ
Hg6vRxYZRik2ToJrhdnEvouhkcXINBaySkDyB5YFmesIfJuZLCXaVDALNtzpLvVHhkVzJX2WUcDs
G77SzJvVpJI1yKZOuFISDwfvWPc0yt+pKcQPE85ktSTksqOgW1Qfg1bcKsafp12XOj3etvQ+uhwM
rPRT/K2EYGqFqZN/bWTQd6HaVwclIed509bZbV1MgqITyL6UNzz2XkNCVKIyJgC+284hLx/6vXDT
f6vqSlvFjtj2cUk0w4b/levOvVpfnb3RoN759JM20drfElwSrud3le2WTYcqL5dubCkyqkgpTlUR
FS1XUtGUXy8LffXn8seGko/BDfbcys5CtanNwEMSbrGgUCch+eQoyyyf7olZODzQTTBQcT/QhkMX
PTJAHuzZwg8yC4btpJd9zv4hkcOkoAAVtLC6dniDXD3/d8UySHRtASCgQjv55vIbOH1gsnJtQw6K
7fwtJBTc4mOCLTWj76f7VE+pxcT2dN7ZvvW6oWaReUpHeV60QywmyW0TTCooazMMjXJvGHTlZgqP
ognPLUqdkyh36I0Z+y1o7KXH0uRhhupQHJj8S8rKY3TF0+l7erN1x/7KARocF1Ntf1eYQcpc5dl4
am6bzDQuj5quJ6diBbD6r94NuClSWDTmCJzcu2SmSuR6ILpl+bIauQmqgQHppdeV4iiFzzUZVHw1
in7BnEphhryFVT5NO6loXfITpTlouQIxbRNDUwf3DEOmS5r95QJ7fwBapTJxPlsuTs2cMeD6W4kI
UNHjJwGz85dBmB6ICO4AYoaTjzImefZE5PuiLQy68DpSexYLG9dCo0dFFPrh1MWoYRX3dNl1nAea
bcmLUfFPTNnmyG4Gc+JSs95PRi2mpBpoHY4rkxxdooBqBYgEDf6hARwZ/ihBMGc5Qms5EkjkDGIM
+AfJQUYhPAedR54snsaH58USzM8Sk+gVTlxZDd92ygFpLrEizUcYU1VHYP3zcBm05dZ0+hYQgkXF
UFTSvzEFm0qWfl/H10hct4ESA1GNcVYKpC8o0qqgl92JYLYPufV0VrlO+V+1dZLRgIB1xktEKMXA
0lfvpuiRaIJ/nB/Fd0FM8Op8jYRXo73sfeZ7WIut9AQK2Rc3rs6LZPrxE9Khm+vAs/OkoBcbHVln
JIYc+TE+bDVdcPWKBeF9d6he4zOHZAEXTIRbR45qOKSQWvObwkAog6j2+6BhGRhSgmom7x6gE9Hw
CQyYVU9DOyWSP2eVC+F3C7RGBC9gbE9q6x9sW7v9eG4KT177KSZ/5PtTo9/giLY1fr1wzrIvqVtW
GaybK2U8j/LCgjkjVT6871rmFXUDtj7Kgzanjiv1vkD4muLyGmvVa+F42Sd5OA2xucR7lN1fK2uT
HVoOUsiwLXtEcHb603duIWhppKlqbaXPYgRaxWf79qCcmTBy+loQDLECQaPzrXyzBfZcV8ye7KVX
EJwl+y6NJ0fIWV1En/LMFCyn1Y7ME03DLdJHYJWgCY0/mDImVPdv13TfZ84ddHHncdWQ72dOVpYz
5NeT5tHt2n7HFyLApxfXHQL9sYisNDOVtU68Ev0fpD/3FrMq4u4vQ1xWFAyKQn7CvEEuf2jJ4Jye
TBN7a72f7b9I0BGW4/AIbAQY3BJtXIAdcPf5mQXU8JSWWUeQRCkxGd4uKA//s3ow5BRmoYE0wUNo
gM/me1yrPEGQN6l3rczN2ySk/aTGm/aHX078Ib9jvEXa5KxEBpnEuboRLrPf7eh9opn7V53BFQAr
G1dk2vg6zGGOtMtGGt80zP1UzL3GPJIIWfoGXdzrubiPMLBXungyCL649gKmTGQBtFh5fzHZOs1B
rLeLE1E4n8vb++Mj6EIzdK2muZbnz7d6kvGht3WgR8qk8eimWVYegXKXOIC5895TYN6JNlRnLnJb
Ebt3fj7FopJah08vyDoegABUR1HkFGD9SGxFhN7x+OOsiXdEY6bKf8b/5q0swYJYsIMzsw4jg0gG
2cK5B1QrUW3hxjKo5NYdD1/mGi6nDycVrZJvGdkSzdRfUgsJPV6ztU+HWd4gtgw7Eu2fJ5ZJTAAM
o93KhWi7UlvX930dM6P7hLCQmJBprjzU0bSrsDv2PzDHIlcT/TudVsT4IjgbAM4JjV00EZgdewp9
UZ8ohkon1TsUvMj/+ewXPnkmSeVsimkGle8CJ47DUZfCdl1aDdPZ6CXkvC4btFM3ynu04umdb0m2
6QA6NM39xIBjcrCtuwdJiZF8UHYb7c31MsE1IuUuvmR+a2+XXjQHpy9Bo6UjIIIBrG4l9cdR01Gh
yaVfYF2SAJicJchJewN6wXFotN32Ur2uDPFnlbu1YdzVTPSPGighCaXEEfQwwa7gmbunk4KLS1sW
FX9tRciN7WGez+brlZ2JvSohTdg00Znn9n3jkkWb3l57E2QiaoVXP67bcplZj5RGgylmfdVXTOdG
CM5qfCvQanwcj1PeZJ6QeIujBQRXoOsec35stXbj5RWS7cCZdFox7wpI5962k1OHb4Tt5BmzvsSU
VSPVJ3Wox5P/Bom4Hkma6j68ZVasbSEXiZ3rM4hwM9G86aRKxEBncNl6K0G8+fN48FVH7+2645bA
6gTJeofu+68GKTJ4wZ6AMExB+VqmMfgTtv3QUzNDGUPOWD75BX/JaO4BG8DievWofpk1aOD6rMS7
lrfYlkwE+3wkzi/FOrqGgh6YCTcG0Ex7l3Gihdl9F9Hl3MMzHoIiTz9de6L9p/GDEemch67NhmD9
zfGd55fGHvv5XML/qCTSCvwG/AKSg5T9aUL5CQ+jCjoPKPiauh+KNKkhZO6z04WpwPqOsPVtXeId
TuowMvVay52Go4YKrrRCaUIB5/NL28W2cWBkdfhYDhBdygumntNZ2riwDlU0WEAxNcZhuweMGPoc
2XdhC/XuyzCFEDvb6SO2no89LJOpGcgzjtj7li0znmalh9T5cs2ZO/xUDu1fjdzm+bvXXlPGfXG6
YdM+KTxVyNvDxgYRVnQxpAJgLuAJpsJZlmU/I7nQdk5nMYmvUwvv3bQ0k374RV1/KfVH+ZArCsGm
IAN9vgCQUeyuQBwREy7CsYSCJWR3rcp2dVmQ90KnWfb/UWMJsHWEFZ+eY2iLYFV8EIEYQxEQQKbb
Q7wp2OywRvgHNUL/Gf49bHvXFEx0Dg5Uas4n29X8BC1TIhaeOcoEVOj4mHoMQgLlBx86T6xv4Cv3
9eVxH+b8pQGM06lo3MoDyiNxct938S/tOhqAPwaDnNXuqOBoLrdYRFfB2eLMlYfpnAGT3Ii1iqt7
pdDfdrAiBOycXbr+5CCpClKOfbanGb2FmFOz5EmVgizuo34Wk1+GWdeS0C1p7Q/aWw9M2At92vjL
huZn1a/m9I6gAPX8boKj3vaQpgMJM4aPJrbo5nFRnw2fkA5xWg8aRA1vMfAzLKc3ipoJCUVfciUJ
iZlGPNYlOqnwhqO1b1b8NRW761gu0GfsxNFabB+twl7MV7zub3/qa/jOJezkNCMvZMn7shzo5sm1
Ibyci4fpkwuhLM8UbjlLnM68cbZn7UPDGlN2WF+O+lpzMhFKOmc3PKA8R3Dea+zlUkEp14VBkm9o
RenTkj1sgSEctvT5gxi5zl6m5sbjK1SiC5YA9FxGQlsfFw5JXcKA1dt1+sRT0SFO966hdIQ1w5f6
tp+du6RjRw5mMRJ53OsbE1YbwLTgiFyI5bEL+IrLzqqAHYeXORMKEkbRiYmgvIeY10ho3zGC5k04
WdMBubQb8xBfI8DLBoe2hsg+EwJG2SdoBzOrG/hATc/WoN4xuuLH+Ox5op3b/9PCVbvuOfpAH+qc
xp4Z17Ad5cgGQUsEPgANyqO9hZMh0T/IyjZ+T6eMd4dhyazXTcEdGVWxTZ0XA6fchVUQUfZRiql4
fFeqtidcM/ccO/ifQAIdMMhR8HkbS/gOgHHyEvnpF1dVS1Q/b6MGU0PGK7kkZmZerazVJwxnLnQE
hep7Gg/cUh1Led4jqyfQRvPD4Uwdbuq+8Nd6QNnaopVix5vcKirioKMKdC8Nb4rOk+ZYMD1UASCZ
eeBviPXHshuG4RfKrsljQQJP4QDJzk6P1ZFzvr6Jg/D8/2+EZSybg/UyAkUqMG5mxm5bysfB4vGu
zFq7vohYQMfUSSgV3JY82sHXL+4nbP9VPSW29xgLJ6xvZ6gv2cyWQ1py3oboLM41+JjxHwE2ZWC4
3DIIsEjzewhopu7kUK/0bswOA1LJ7OsUXLGzw6O8SfCudI1rpLAIXz7YNHUcIN6YXO+/t4QryBqY
RTHsjKoqVlaK91bvCYu5lbsN7VYwsvldy9gp4+q+g8ySM52KWKip6y+o+87BB1B9WnCDAdKkIwI+
u9Y2LPMU8F5aCvh8Zet4DT6XfefVBKSEHef+6rgLFWwUuUHNMBHTpp37vsZrtpFIhwDRovQDBUUl
Rkla/KLylu8xWtr1dnJ0aSfrpb8Pbbi2OXf7oKBTm+OJdeRE7i6Ccv1aDOOUIZSBc2s3YmsglUPj
l73yx4So8Wxq4nd92DMAUOMHPUAWjnMIrjKF9sMD+8ByekpqwFB4mDo6n5szXAPt6/mCUcIbCDoM
jeara9FeGznH3i5vjCsSlGF7iB7jbUE2dXh+r4x/rE88gJSwmtL8wzg4eynHtyx/oP9ZZk4Vzian
HAFaRhaF6/vxLBKSdByxKqSNQI0d093+/Zsu3hWOTDTsXucR00XUyFu9+Ubqdpf/PKQSozuXNCsu
vy8qS+20EpGN9Ka5JAoGNPOSX3RfaAZQ6GjLyhiwHQ7HFWwXxHjjnIFv0oi2nDKHmrrN1XIXVGI/
vNJFZk7pGk8YMdDU4rCjt9Ye2frzV53ssEGgAN/TW0Q6F+Sml4zgZSn5Z6yF64YutiHcht8GvHaa
FbHZnIFytMqLf1Z4dHlpowGCugMkI54k1KNHcOBbKItybnGWIFGrRzfLbU+9xO3hS5ujc2xKpul9
+mH+a5MC1g1uWC7BWIHGaIJp1kj/tq2y4qykgBLfJ43tu5OFPsc4H66hUI6VI0XgD7lDAPzERK3E
7+71oXBeOIRdnV8toF5YBG3+5mrtpWjYCC2FwmyRqzY5JtUZEm4B62EXd9pTwtmyl9Gr/Xx/klB9
4qkAJNeRXAtTWUcN9bWzHN1OIIub/azjCKfZkE1GA5td6pd5A+xnMVyVub4iVsHJ4td4VWhWO9/E
rt1RpvceurAvC21WYm63SKkpOgwaBmz/JvwEAXmu6qlggaxTExq3Bp8EuVhURGJ1tIlLvuLARhdI
JdXT+4dEY48NeOcJECC8/E9oF11MYKF1Gxj4OAN6/UlaEMenmA97w+P/dFOVzQwaF5ac2FAKv0J+
ucYlbPs76Y3urG2oJu5SoBCw1oszegaYsMtKaS/8m31PnLrunOAnYW/YsY7KJCx9Or2gHKIa9aoe
is+RC4LppPCZeu5s8/iY0m6K8ZZJoS1+2Wsdjk8uxNvj1rHmL4qXWoLxC5By4onEcOP+lyGgZto3
F8c0eXaCDLJMxdnnDsJHDBcZz8/8+BHkv+0hUo/zNBFSml7U+tZCUlbMnmfRCfpYvc29gyftMj00
/muHPki/VedBEqm/VfD3aLUrJ26S46U8I12qkL72lwCgdJTg5bUHpdv35H40I9cluuX4SWyMqOLN
0MLuSuxNkaudEg//CdQcUgM6pGGOuyQYkWmEC8RLXU2r7/tMj4IfjEG8IcQtdoVH7TCqowqFQtQH
lWUFsEH4AXsi0sbmeMbuPHnlOkjotp/pguGazJgdPoTtY9vM0OrP9qgEMegSbzm/FV4l5BxukABH
A9OlqPnBplNog1gzYd0r6ytthC6N32/M7cmCPOePKYnY4/tF78chkGZLJ1ZKydnTXHOyoeaLlM+z
w9AYEhm44OTz8oO8n4whIy9y443i0XftgrPfUjQwOS9Z2kGNUwRT3Hlu7jubIbZ2xQwvbBU87vo6
Vx+GyvOSPKuwgKgdiPAVB9BiA09JoVgDcIYP7Z6SzMXFXLPGUBhjBjixMkGDc3Gh7HKwQpgSGCkT
dg18XGFya9U0MSwX7JKugwZqGfMgKSXFXITftzgkvYgMSqjn/9KpW+A1WHTgGFahbo78vwKprk83
qzDUNUYilqW2CAvbG64/NYwwBkPMi1ZioBdywhovtF2HhbjaUXdrgIyfKSr2coznAbLapme1RZrC
luBCuEO24LcraLG+6SIkLZpoHBAlOxaX52OcioSdPUz7ownUdhxT8KBmCqJTc3l4hRYR9jfQIzwe
4ezcCHdD7+sJCvsGcA1KMH708WADNNYDYPctdPNbfcHlveiebak3WuGa/2vw6pawhuCHJEk1PRwH
5nd4yF5+3AVNx9ncZTE+aBKej5OAYsvsNmalTCnGEN0a+/0x55uiARAT987T55CdY9qNrUOFW/FD
li+Rm439Y5fd0FLPNDa8l3uK/DAmZOc0qlMvQkD5+BDGcwRPknZML8Q1/MltTtvuOTDN5p4I6Aqy
bpf1DTHl3puiD+TonZ6xq5RpwAeCXPmbZ83KjzMCfCnk6dTtfb7rPHnVWU3VGww7AngYqHafbmea
sELMzlIIYK4tRhmAmHDzUNbZTWBVG53dmcSfvqxmer1A5xFhgMU94dm4+sXU5Tmsq6vMfWmxZtea
cJ7Zw4Pu4LzXIQJMeD4AXg7ev3IKSWWptufRsOJJrtgJWTXyEevcHv2byx4V3d3ZkPjIFAwXyRj/
WNrGJ/k7BYrW/DeIaOYDUjomyoRhYg9Ge2yH5W9TbDsKj5kfAXOFMEQ7cAUcR+mQJ8MXo7V4OuTi
d7TLjGRUqY5qU2+LarSQf9YkkKQu3mQo8QhZqwQ8NWHx90ZUXvYnekfWxhMrPAmtLh5UpfzXFzAa
zyg8c+lz6hVUrjGh54oT/tCn4uuP+Culyf1cDvMaBjnD2IH6OTXgIeBR8wvix7XgzHG7hjUGvfYU
g8lEqDkWQaFO/LawZbfJK5yMA00ooybuswGhFEQEUtVLVHbTBMBEo2HuRNG61ZjUGLU04u5KYGMr
SyLuXsO7LS0IJKM04nl10QWsU8XKhfJw57ntTnHiEUkLxYmZ8A+1ee6qDIbSMjJKzOI4mbzOZXhQ
AmxQgr+Os6KXWU2KHdczrZJuQ9+WH/Fgd4vK96q5DvUqScr87DUc72OUJ1WhwqNGQjBRun/OosOW
PKkPqDclZpu67w2UxGPid0jsl4Fg7PbHx4xwwBw/oLAr++63clQnzJ2Xa8eufIHrW2EGpyeRddKo
IuJWIKUjKDOR9QdoiGDtkruTww1ZB/iDRs3tV8sQnvJO+S2FZ14abaquUOGacj4+MqvRsZrMcB/k
emAHVrawJJNJCELyAnOXh/Jd01lPejR2+HIOVLF2UU3kCUuxxC6qYRgwos57gAPUfLyjrejvSQg2
WjIQodgaqPdDDWNxh5uOp5o8VRmDGmBy+fEtMaqJmaUg1r15jD57GChi7FcvQtw8Htpwt7h7Bv3p
MH9wgyGZL6CYyXGkfOUUfZwTRM9QmOBcWGN4YGK5CbbYWy7D0dspMq1dBQ/JXvXo8BkNDYz48XnX
hHYg1xJd4WGTs4Xt0beuuFkSxr84CGo4hyWisIhXy5E1zSK7qP0gYP/7yUB3Z0iOn/0i1NNH5mA8
C+cey0OeOrbmEsLvqnblHbMfuacwhmWv663mwC8Le5ovhTbqcu8wpifXvXfO7hZk1ri8TZHWzqps
sYx41XwU3fqCtdv5bncKGLCiLHtvhGq8cJBHRz0wU98+rRIo7sJpvOAfL8PQyBBKqwjg9zC4TIKa
1+8I1JljfPY6WqLYlHXlVRhryefgxmRtLFo0Eoy+LN6dk14XpwLb51eAg+gNFvfUaGpa8/lr6XTz
f087pas5FDTmHQv1yv5xmDo+FCvTt6yxhWVlEF8HWoU3str56TPKpjNhn/wZGR8JQM6f4kQZ98MA
BpZBPtNbV2DDIZJFraEDpb6JWN55wTpcuu1lUXPThJfxrMTGJHF04iX2yw+ZPeAIsDX9tHHDfxAg
IoyBdT7NxVoUBjsDU8DqY2QwDdXM9qecVKmFII977LJSt1dBZYFWU3X3+a8IwxJlGHpcIhBxh6RE
CoW7GDjcNb+ro30cl1uSIApiX66OCZ0sWOmArRDIEyv7+khrrJGVKkbW0apruCCCrFrc55CEPXrD
qF6tYWeNh+q89zMMNeDh6Gh3pl71QO/lNXCu3UhINcxaxXxinmN1VVz/TrKZMhLinyGMZEjo/ycf
vw7btTzl7fQq7WePkQUFKMH2yZd6ZpZZxoeiu0b99/yrCqPXT0oEFv2f3M1F6fOtGANIzKmeIIpu
vzGiBy2aFEPLoXbjTf2wtEKAapdQpqF1FK95qCkqQRLZ+VLor0izuvSIDancMrHcIyUSbr1isdR+
ycrheRfZFwhs0lzu6iV+1POYazK2KRgBgQzMS4SmaiA7MMa4habRIDQe94hQkmrJwsxsY6MZmu/v
BEo5Wcn52B53j42CLri3+Djsxat1W2CJmZIkh5yDcnYXiN6OxzBGNJzlYqWtWb3b0748ltB9pkLt
cLnxgbY+Bct5BkCY6CsyOeQkKyOZaEFs65ROmWtPHED+nR7oZIa8gik+dlD3JSHXjB6fG81h8OVt
bWdB4qpPOjpDNJuSTf7DHAw0rPy5olDCIgRYsKSnZk0qDsdhvKeDGGIpbZCEjfJgVJTkJX1FzDmA
lmVsh2IcitEIC6U+PeeNWlu8TnFqynTjA3UhS6GiIMpBzsxN0YXQdDiI7KoLycQGzuJrmI3xdTGH
5Rq/juwKSUtjFo8nlbwzoBjHQddXgnnUPlixqKgjsFmDpULs8kdhwccqt3Qi5v796URpp9KLawYi
iPId8hwelYADQD86eq0SpoK+O4LFYs5sDWCc2ZmKLSwYkizu/3sP0tV4PW0qluB5qj225jiKEzqU
/x+xkJc3SI95zYcyvW2ZSq+gl+W8FayDMQHgNzONZ64HDlVw1dqcSbkKXhbxos5fITJD5fgnOlvD
zsc+DP20Bdm0IDV0qVBkLb55fRagsTtLO3yCYxY8mOemcCO5X9Ty4+qOqART08pxINclgdH+9fEm
yvFoDYsOBiPouKsQ2BDbnO4g15d6kDw+9FkWpkxEAVnkY+CZp0HDuPk1a9idvZxW4K5s8ag7jnPd
hEQwV+pcl2+397JMrWI9GauOy6t4TCSQXJ6MoUmS4RCfhSD+tW5YlUg112k+xlkZU5zRlDIYL1gp
l8s+9YIX9sql+rrLwKIl/KI6honPJWXd41Fue3MYI26bM/r/qius391rPU9WYOD/w13I7IksyjGf
+Xp6IncLVhNPucYF9VE+Ks+a2cuvGFL79GxoJ4/ghWxD8pQro0lYaDJCRaCANgvjswZEa1ipM2Ah
Yp19bGwCEkxJspBxqEhUBJwJ1QfgLDDKZBL6n+c6b4rBCN6Kx4r5ybwtj19usSRWiZO92aWOl8Lp
grzsqITOLYe1EIn+gBWKdEkRMHuuU42neHuA2534EFjCD0mEinyQ2lyERX3henKenR5soLnPJLEd
X5ZBlJWc92jxebo03zG17mccHSp/23vXjRejMChyaaoCy9k2QNajGnfLKyl2YZzYz3gzGxEYtdgm
y3lzEdzwRA88/ZOa+6FTTMnzufUrasHod1zXpD+1MNB1CejYI3l/a3DHx1aalxm/GZi1QLvYT18Y
5Eym9CZ01OTWaa/v8cKnJSDkS5i/Vbhx2x5XQQ4Pf9HOFQmJsZALBoAsGLuKZhj1pxU9L8eMEIDM
ALHvbnxwil6istLPSYo0I5Pms0sDwzjEG28F9/yBA15qQe72a56SvYwLnRRycVvTElo53/mipkah
z2vqQKaykwPiilVfcJMgECcy4qqxUSXcvx29xsDSEy4gw7VzeE7Fu1JPRs1F8NGtMAMuRMtd8JxH
E7KtxQeCHdjtWxZEmRgw94lT0sJlARQKWmS/rN/0sPO4w2PFHOpQs09lQDXNg1TWRHhRvQ8kGkls
9ysDzRSz62DpMXxa9eOPYIH9Y8XHx0yTMh5JIpaCF/aD/82AS+2EDm8wLuW0rd/niJPnPlcnkSM6
1g8OnxZT9GMy2oMKZ40fmLQc+z0VWTTnGRkG7VaQRf1FqMZKYQceQLxiZ3GXZfLNkRKIXVkeluFM
8LS4mz4OZJttKyWYhEQQ+Iyvgt6v+usRKggxXoV4OuMDg/hGCtm8Iv53Y1NS5+R93igQ5HaUQBTz
xyJwGlgQNU++hEaj+t6f/keNlSUcTL9it7c+WFEWmjYNv6ym0Etw6ZSD/N7QxjHcJbXq5+v8wIO3
iyyGWm2Uy2hO9YNYxqdn6iFT8Sr1s8qMsQ0l4F7aVTjp69w870yLBSt9HSk+IH8rgoOzsOWDJbeO
w4D0EdHp7mtYXDR/VU8KxreQZdNjLRY+GdfIj3QdsC1hzkbPXmpKV24pjbgcX6CehsStSpbePYdy
jJ6V+bRKs54W0FSkiGrK0UwJEht6ZPQnQec3vrDguMzjyUcin1PEDsYXIVCvVY+xkp0ZoMNTsOiL
MnmHp2gpY+d27JhAu4NBXl3md7sjVwamDr2Yq82O9mtm7GmnXnHZ6JRwFzr3E9W+U9rgZP9Ep60p
rxfXBWkkf+ebP0QE0UbaJHUrVrr9qNO272c8bBqhzTIqTBgTZd/25YH+TtEq20X3JvSv+x/L53Ob
Jrs8lodmqNhF75LNp/babut3FZ71kSHe1JoavdaidwXEmfW5yEc8+g7nsG1EJbtDmPMnG3clB96j
CypRPt9pRdndU09e61IPTyGTkn33X4PKWapo5sXag7uvYi2AJlJ79Hs9Vm6WIWUZgGRqfPQbqqZV
ZDgp/uqVuFdFdl0yDODkYMQzNpXiz6UYwIFhL5aYd7Su2A83bvAUzXdTxr2H3bMsMeZ/AcOHfF0e
1SPZTOF4qgmOyyXq8A9z/6r/AUJKv9cpJGcJSX+2Oh3s7M1KitcLKOvHOvOvDDcCSgc0aQZmlbge
fHWeTggfaNz142Y5FjHz68uhrpqO6oMOadZb7BI47BSM1rleqjD7PPk+nWe5aFszuOneyvMFdgf3
cEnRnbpYOte10c3kiw/ATC4sHJPSBrYC/X3m1V6T3GGxy1DglAPdR4fIYYgrl1VhcFl4q/ZU+z+R
2e4ZEhgNbfiwWjk//Z08/JmOaIYF0VCA9m1uCGl4lgXLp63TuCpY0bIYgw1wXUcIaT8i3zHmK14h
UTUC12uFljXZ5uqfZRhm6hixfBdF758lMPFg+fXooetMS7wLEluX86jqMDYtW564ZbtS0f8N+U6J
XqfSp5/f+OggvDpTjCiDxrAw00Jor8eAXslWX8MMcEwv+pAKbAlb9+cfcgkShwTmL+TcezqTTAHQ
AbHr4WQ1Cso15p3xv6wjAfoTiROcAA21MKmO3EWAuCiHtKM+OaKSiIqT2sNaGQy4+9b1TEdoxxAT
yemzxv2kpf4kSQ/j9CB2HjcL0k4fpruOYLUkrYO8pShEp1F9sCg7I7pEmiwZqBjVVHm60iA+x12D
xq/5+DCIHh6sQjadfmxYQnRFMRsWA2fbad1XNFUIdejQjwJjzl0kh9XwNFbigN60F0Jbins1/2Eo
zn/6hnlZznFVGPPWJ3gFrid3tpGVQKdM4YxdS9O+DxNOURCWsICVaTgCs6fAtWcsdCIkbMQG52bD
hXG5HY/h2ImVI9aYnjDzXn7hSeg/qJwFmn9Q4eIp5TcASeDiUwNF844H/l7gvuWE2PYW2SiBm91x
iVMGdUe9kHXHwYzI3Pf+RYssGZLXnObgMCQaVSfiWaExF+pq/ZCUPivSC25+jFxZAbuKXkIr0Ry3
ZdDSv/OeKOZOyiqdenGPqYtfkqNTsItMPsdKVmOnKp7TxuIci1sQycCB0Ugkg1igop1DvZ6m8skS
KhblssjX7fsum5d2KYdOxGW5gxeznRcEsjTKxAPMuTL9oRWeWzm2wu97BIjq5KhwAvFIRUL5cw5Q
8SClOsjNLf9gepuA98+BkIlUMNN694aMgkx19v/MM9B1Msk46C7f43YM7XuRQspMP+hI3+cQaxFz
yzSlL98nF74T9GqAJIFScJB9/ib3TleYkJpJAfnHZR1ENRgkS3qQBxcgcvZNjYf5N67+w3BtR+1B
Y+3U4Nj3HIKnJ3mafLDac04T0+Td+IkiUL+PAlBqG/JfnViUgG5Ram3c2rlxuJo+qWwT/DNzBZnN
S3GzNAmQt02ZqnfzTIJeoMd/kGXbT8QcZJtEvYR3yAbs5OHxaMK0sKhWssvo1yoQ/SZP2qK73uev
jn1sKvY74MA0yL8UtmYBG/boB8Kf6k8YNJq6pXL1dVa21XfM7I6lcmuUkdDBzYItW04+n4upDQz/
D0ReR1kZhIZ/QT+mAwu7nPHKcgW1DWkT8FgttI5M8uVi20EnfjAnsOADwYAhvMWxwpkMuPor7fLM
VOM7hTdyh1tHaZZiCJxqooicqBPW7CZFKvMv6Te0IKspdMM4CevWVOLDPauRdXPzZgCy0qlAP7LZ
g8GOgpj3Y6IufRPHdiT1wP8xJ72q3bSQgY9mYUkKPmzkVJ9Lmidg8+NUEeG53og709Q2KIT2iwUh
jItW+gZmAqnGlhR4goytH/pm8zgP/uUyWwb2Kpr1pQRsPWOd+DdpQITHNE9QXOMIDI5OdHYdsQsh
ghxwBpCZnubeitB+bl7binKZN2dZrlL6mvRWTOd2taKhOII1c/ABoCfebObw7oXySI1mNjoHNCZg
iGEwPg07SJs+h2l2TAKYdJd+Jtkg4dCsSv5I2TcS6aQVpw10QNzs0ZFV1UsXBZm8blRTzVNo4hTr
LuYldbiYYDPL4KoUys5w5wozVgSZRX88wBdLGPzXdNEmFp2iGptlTjEo2Wu0G1XHwvenYrxTj/j1
Xepy1GwezPbh9hQ2JyXYEr7Gynw56Gkzsmml/XRC8bCK8l+FGPRKHOmwQGWCMR37xFgYtqWMgJeK
mIdIwVBvjuWH4tpMy0Akdal6LFUvvX2L33IGgEHFY1zX2/kbCuk6Pm1D1f3LXPs11pfENa00HQHT
j8vrPuKj27JhrLibXYQeNVlByHN8aiv4TBvvyq1lzcl8rwcY2b0oe+/JYKPTpIHEvDtPDWUiH1V2
8Coe0zmia9A2wm3BCduCaxZA3R3WO7vtwv6o+G9cf7cO57WkSKiUHkrCQ03XWYDIBHCxUt0+7uk8
BVMVsvtQ7WvbOLbmpUFVQ9/Ld+ExEo8j1K/FQ0xOKMmVxW4Vuz0p1iaI6Ur1eAImZh9dtEboOxLs
XYPcN4j2yy8foZG9GgmhDnuy+uy5QiEpZU8yQ7kIgVHd26g4vLGIiXZzxs7iRWUB7Jysi81g3fAw
YmJuuFXHs2nt3+xFeAsG4yC8s2vsvKSPxOnccWUAMD9bCSuwMjXu7t1Dwk5ehYV2jrd9mkj9hE62
CAPOBCk+J4+YZusLLCx9BBE32TfdrzAK6N3NdmOp3iCSir2fvoXJ+zDtY6P+ujcMTS+A9DxB+ngD
3YTuDILqcP0yiVKMmhaj2Ajv5I1xWWu1o+uXA/byGwUh8/ht/wqn0hSky2mJPKpIsip8L0mIzQEt
pdpp2hCWNQ4iwvQKKJI4mTA9Xmb96IM+zwhg760OxD/R21cO74PkbgLuv8mIqv5DAGE+uQpajUD+
dGFE8Sl3VOgJdJhgKT8L/M+3aKTEqRgKRnHcYFnA2/Axo7FaPhMSrDHhApvF22cVYWXMaAeOZCYK
xY7nsh8ie6zYZd00l6vb75eh7m10ADx+QuUOd/OI2pBLCWhM7mQYN6FnQ09bCIplzC0kyIrdyb7Q
cXJhdSCFTJbkEJNEGY+HTrkljaBFlQtBO3mIGZSiYQz8T9fQXplpW7K5NcQrad7vf86Jdh4cQZ6a
GgrjbYGfZOPMwq6FI9lj/3koCwTzljsVttDYmZYgrne5sLoOXQrWPoS8L5R++3oRhebjNzpBQc5G
c8e3Dz5DOgYUCKxxKcpk+ki+/4LBeuMffdZZOdmtLGneUe8wWBxrInbGRv+Gvbn4UI1XL1Q1xaqC
ZI/SdzjfSMYxY5pgODbOnTKx9N43muhc4tNRDOFsVS3zlwunUZQ8sScvh61YSnoRnRsEWIaKkHbT
Wc5+X3QR/NTsNmjh5ra9zGXVrXQI9N3Q35MY4RAtGVbqMkcAA5lscUh3W6DHyxTefztF8eLNnbTv
e5ItWzCpoFofWtjDanuufbuf70rpCHEsEXP2z7aOuzRWJLMEi+fRFRL0GNrsKni2gcqwLmthcwap
PXujoR78G40qIvC1gm7mHuB3RYqakkx/WtXgdfo1LjVk8xO2sijJN9oxbnLw/sFGl6XuLP6ou793
QfREDgkGC7UYbnmjA3MLk8TiBuPVPeYRs6xQVOB1vvQGjY+luLKasa5jt3nYtKRMF3n5Y1w8Qrs7
v7dF86KBWJQO+I5P9Gp8uBoadT8niR4fezlvzGUM6iQ/xmLwFpV7Vx8b/zlqM9fGfuyh4ez8PfGd
06Q8gwzbP5HrF5KW9bdDYlkZWT5dk7ChHZVs8PirjV1fLUWx8FYLPQ6hXJdCkOxg+vPvtfMpv96A
12FEGsl4ZyNI8zvhiluXYTzXVdh1uLp6iWCS9zvXGMPXH5oqxWiA1uVCVaPse9Z3OKywHIxteExr
UtXpmBVnW5i3v/435qKyrU5sTaoNpKXeG19pD5qd7V2QUxKVKzteIasU2pxzhOkb/y1INqyT/qDi
TJ7cTcKxBB7eXhAWOhXJK7cVYEoKXTKiYufIBufQAqFcCv7cpbmTrAPVzcWY0ONxVpFcKqNmnzHT
/gzOJTo6ALjhIBL3w7Scd78zmyrDQtV4CEe8ra88ITfiBsBKe5Gw1ZuPAG8X52+qY6a8kpJDDxtG
Cs6lv3bj3JjnE2UzGlirsTmZ0IB3F/Nrp/1Z61uGDeSE76AJWmH5JuQCqhSoIiybIiMGjCrt9WN0
TKrCzVVUgeKMO4ZJr+HXIsjOUbby7kRR+jHfbvruUg/IB7Si2WkBwHyh3U7dgUq91//WpH59W+ia
OBRUWt+XAdPE76rYutFkVV99hjKsJWg+7J4FZinqushIg729JYqk201NUbgZppmbd/EKz6m8AN4P
6ZD2OBfO16+h/seT1dOn0fHDoPIIA0dgqE/r4vjOsG/tc+sl0M6pZf7BY2ZpGpZeowAy4pejCrlO
yrntj0QHIypijXT0iougVS1gGf52OMOe1PmbZOmLFO2Qfsgya/hcqxERVLxkpMW4cunZPmIf9eH+
3GaWr9Y67rQhjfvxDEvmh5uDIQjyW9Xn52HVHt94V6Mq7NkO7NTFr9+WKAMdrZ4nf5A0PjaG01wi
YBM8iq01qYYEI+k/7TCWUMC4gCZSTzxvKCjio0Ft6EmX8SmKIUHGp5SmqodxTFpg5huq5/mkdCdY
NtLkFKw60DqRSZsJJ14wk/vE6taFY6VoqV9v3RgQBi92uvPWLiQ9mtI/xo9fU7zDwNpeaAWbQlks
h334yw2crvt4W0C+8A2V/JfOkzA10xX5n+fR1qQPIquRRJnUnyyjhcPyBd3sh+Gq7VbggwvTsz7Z
ouNbmsFUC7Wgw4nItKo5i9ujY0bRFewTMEA+DiVv6nl+JZj2Y2Rklmhy0B3mNu1MX1lv9gbwDf1N
9DVo8p3Zxwu/BXITInsVKl1BsCu+UP7tZu/NIJA/uI/L1fFyl7cR9rVWirsX+y1n1lIMfhpHLvTg
dECfC2NS9tRbqNv822Y2RWNbnqZ/L/hmMjkOPuBAYN0wfts9+Bx0Ex+5Enm4LuZih4l4zsQoweUq
/BrtQG+pgrNthoSEz0ZnuglsC8lRsdD2lunUWQuLqDJs2ecI2sRvLE/vmVwG4BaFcrdbGTl+KY1K
01xcMA829RJoPjq5LFWTqj7iP1N5pMe8axn1e17BXGqOHDQL1Vumu7f0kennBMOup6H3kf5tyDc+
qPTM6itCSa0WefKDSjImFviRF71J+DziMF9sJUxawC9pimcaHZB+WJaoiSRRhlkj/RLLHv9Tnsgd
ENHc5nBHWOCyZgqjrYeU8fKVbkHlMqsXJHfaBdhzrgRUKQkAGDowigIfNr4ODef9hI1+XArate4w
rQXWCbUIcUXVH1xK4ACrnWvOozs9cL5C0bpZSSuBvXJ9JQmpzkRwWMc9u3ZPHnYn0YaqllpoRHWd
IFt618Vc9b2o2h8Tb5sETXazf9oRpAKr/raTZmucLFB33r/FdfBfJPTV4Igcv87MmgSSyaA6bknH
DXld/EIMopyafc1Ky0kF3x3BYDUNiSLAmcdwXWlLeRJkuQEcO6nMwkOzMB49VUzg4AGnCFJTy3Nq
LwrbaM2NhOwtP5clQZ9UzdeCUPHUP+ypmuwfeQ5JhHYaitszwaqdcFVfZ/QYb/QBMC4cpb4DaoYS
1f/xrP8shQ1lj9zmE9rw0bA0RsJcly6ydbzSG5Lsk+wJYBTkOExAxYZCEctXhztLtPaQ1aX8DdlC
N0QqFHgg6UT6okYRTfAQEzS5lh1l3r+BDbpvDlMgboDhoZiQPstDcQK36EgxyJxITRQ2kHYor1Bg
rirPW/QzBGBPGzbplmrFEPrh3RnvIvaEur0idN72vAEDVlGQjd0e20ujCxOSz6n/zzLM1PZNi2OB
LfT4QrjJgNuBVqerwf06BQLJoyKfTadTw77ZFK/A5siGRLn+5QHXe9Fw2d781yzRabO3il8sywo8
MgwOO73kmJKhzWAPvlwc0IUMnu40+G8ptAqe7e1T+YoD4yP4ynBWVudBF+jBZIW1yKYnoAFoSKg1
8afWHckrjvslEPar70JIBMAHatAP0+qDGrp13QSUYXeymZ+MMZ2TUeZ+2ufW8DCUnJSBAUNoDHCm
gk8KJpI0VqQ07IEXgcq0O/crpqMl9IWY9WTkHZxw/ai7RaBEhCvaG0QGL7+JcsxFpp1Bib7/Q8zR
Yiroyl01LiradWnazXM2Q/fN0PBtHgCzIg0ujy/4rq5KffD2qdGUMF3S3cZJuuvIr7d6gdANKcy+
2emeRRpolY++i9H5BfwMU4JglW6RwEn3eKeW9dOFjE20TGekeRjyhPlnpFgE+SJUIlQYWAfwAWk0
DFphe42azakzIjc87yONpGJUlttaY/yOj7jwlXJFKl9z7xO4fjcChu9VaOz2sGMSFkScSLPngF0T
IUcgCsRNfiS5JQIiW4XCYB5+WW2S17jIrn6fgnodBIkhS9u4LFGBeWAp7o5LPMyHDeYl69RvnXF2
/3Kma9Pg2TFKsQpx8lrUwmLdGjvHrPxIf1VlA0hFBfyB09jhn9L2mobUUEU8empSa1wDnDY5gsch
Lf+gwyR8eskDTDA2du7vE7gLkZgbCNEsSWLO/868KQDjeqR9JFydbL1tKe98IV1MIVOF/Sktyt/s
iyVoHM28DO5y9h8yaIYEbtn6QmbIKbNR+8nn53gkJjsX2QLl/TBsvwxj43BEN6+1PuWGyi9c93DV
aYG0RZvKqEvc/XJCgRdiHpLLcEGIcYgD3bt9gwPW46cOVqXhcoeMrgtCTaDUkatsENWEGUWa6EVV
3hs3F54Wi8COwLyFteqEzV/uleFe7X3N/Ri9A4cXX+Af/gX1GlHlClKwsGiLl/uFKajzL/l3XfAC
VL/WwBz1Fdw5umXElsMxr+24TPf0nWT7EG+iLNv/PmPTxF3nhyKeSX/CciCzSp+GWteedUvi+sjE
0pdVvcBI9inWCbJFKDTCsUc1yFFVRhrxWU3JgsjF9APwIixT0ELCnCP4vgPP4i5ZQZiFNDfa8Bi6
3K3DoL7DB/Vm0NDZa0/D6/1u8wKdvzcaFahhPNXbajxarIQpijnLgmQ6sG9ZqtizldCZCR8sDeo2
zyfBY//Ljrv/JrSdoI8UlpxZJN3ecatujGhpSLGoiZcyqC2JSfLY1BkFMMhsNV/rmzIoPV+TZDr3
9zTZ0Ak+kox9f1L8vRed+9KgmmgD/v/xzu2jVFm8XPdXBWYHzAauLfK1w9YHMzecMJsnO7fFdupI
LZrJOxL6njnFbcRIy3DVzfG4SfwKzfM60uPW4o2K7NiuVHEKw3W0uhkz4hcPw+ORl65UzwvtWJ/m
6Q6wJV5YszItK6YZenwz1LNxZv3nJkrAwo8hu4gr2xKX9QKszppqXJht96SHSaVVRsXCONRUThVB
SthgYm7xzd2Ru/jgXjtKjcP46eKfE+M4DVTBEvo5nUreeSW6p6pmwtUy6GzInA4mGVe8375CqrmN
RBJRvPdHqAe9M7CiG4ubJ46RXMF+S3br1A72pEYzPgrcHJn7sJwhVKOIFx/pGxkqyN1+sZtDbpmo
3Zfo+NrqX92ZdeanFjcrdVzEjD6yVS+gZPaxTzfdVmtTEnMPrkjMeukVDYzPftHjfZeGUdKzfFOL
pDKAXv071ArXoG7VU+c/0lH4QmHu1jM5A9ljG6o8ce3sCFQ5L6r5WffuEGSfjt5gsiBe+tSi7pmD
eWHIxPaqeV6fG7/G42qHsA7l8KiLuZ4g/J+kt9XEQ/ro6WS1LdgfH6rmSGe7QvM3SIErH+31PrVj
K56Kh4CkCG/KO9MxWqhgznNo+df6O8PR1eDsWvPehZhS9UR8Y+FP+H0gZhLX1G34ICzKTusp+dxk
3DbbsCuLXBKl7wWp+6xWrNo6Z6JMM6lZeAmLt4wfwfbFBnrkSftwXxyhPzu6zqZP8F/eHgo9pZa/
DKCM5kaHa3WrsMk14/feEjprTc+QEcVx67iOTMgWjn9O4mZKdcxp1/XZqYttpPNHv/5fmNbFCmpS
eBmR5C20i20UkAlb3T2w7zQeUtiZXErS4TwEP3zna20qJ4nDAql5v06sBjh773W3xvS4tD57jbqq
CXH+K0hPRAP+4K+P3kSyPaKvAHFSziMCLp1Zgt++u0SrsJzOVfJMIGttXE2/cpjamR+LSEMNgJU0
mZr/Xj8xhRVZLargQlRyYeQ4nXUDsSkGKK3IJsr9bJcExuhlPeuDiYEcnPYbehzznebADBfpX+PA
csFFLX/TbbJLg4xwMSaFXmbWb5u5PLp0CciQK+6QeNGIltT2gT/n78YjvWiFvYaBJrH8577q4U6H
n9YmXEFxknh9TaJSjeEvJ/aLSNTbbKChR7eC5/PC5WRo22kXrg94SdmulboOhAk5PG+hxkffUnX5
srpZLwSe3aMmG/hpvov6hgzQBBdXfmkMyctgjjCLl/3SzySX5qCT5YpDuqSJrERQU+wnPtwt+WAU
BW73HnG20tDiyP6iVFhkMp3PSonY0jplb4YGPaVdH2mfqccIIZ0NscBoQuIbLOXYFNd/MZ3itd+y
mol1U0OVhIniWB4LiEa9cXQ0nrLR4OnfCbpXHzu/cHt5dPGfbPdFSEJxWYrP7aa0DdCbBCbtWK2D
gfUAodyDawV4Y3bWKmwQA3jWbYu5DAqGGgqcscsPW7r+IW0WStC5meFcezvK1ywdfqlVh+Lb9y/R
4PAfMNPqXw/47INuRgxdWglz6tg8FOeX6NGOzyJ88Ilebp/mjQAI4fPJ06NKsLJftnhYIJYHsOkv
Fx7dx/8N5pqFxzaaRyP/2mlNzBnQUDCYnvH8og+5+o2zD9J/+ytDRL8JvDVGtzF3PqVRb8sm1/4p
hIZI3K83g29OC53h4xEUKomhLE80VGqw+j91/rDk2xugdGP2A3TbYBmePruDUGS0gJcA2GuFOiym
khSKQedjO1sljjkU4hhmXUA/dot9lJsQT6cT0R70517a4hfK2tepmIeNpCV4GHVMOLOEtRhuxikk
QWdRC7V3u0+9XbAtTEZWEbfQQewFE5A5ZOd3XjZoxEXTn4xnp/3JulZFgiA23LO7uMu+XVGnNiqi
xXcglDZd68AMfKZ2lmUPqbjmystekQdMnkIgJpL/yDSLM6UA92vbIvBiRry1Q4b9S2ta7+2rWDFE
Ie9jcNhotmuCs+t57vzrU1SXVACkbWm7T/P8jYiz1Tog3b+Ggz6RCb0FwQ0u6M8RDC4EPNs9+AKs
Fba5a18RJYIN1DZdKrHx/d36Eg/98VKCs+CT62VHwarq/SrLFmepchkfogRoO4r5s11iNjIxepKY
3oPp/6nEvxw6wloKSDQQmFsLsKHWthRj32Ry/TVJcL+Yjb/ZKOHeJMrHzT5llcKXe7Ditz/t8RSK
RlcMacBjSApf5ew58jrWOHN5itv+0rj/dLFIdPbYguMCZ/LiZ5ENTt9ZiHAqBO8B9qwoDVPTOrMy
O2NU8rSFVh9VLCndiGZlakufM3u+RSoBlBGinOgSqlOyQulgWZHyiHYDHXUakr8OKkCZDqm8+zVv
XgjV6lzRA+Pkcp9vo9CoS0MWmbYSwLJZQxQNPe8V4pvPH7roC+JmtEANXOBXq01nPf9Y8lxleW8o
rNo1s/mpZ713NP71TsWYVC/gH7KvC8yEjvwmGoODhAB+5TtvU6+sgjGxeVf5Wgpoxrio5ebfKc+G
uiwxu7Chxyvn9Nrkt60KY7CMsku/iTx3wk8e5SFDKhwgqRi83Ml41HBL5DyGJ6RW4Pv8anTUlFmE
gsiO5xaWM8uANahg7P+NUhoRtbJoqe4C4PMvkqgIJ+JT9hqQ6XYo9pB8VAvnwh+pKia3IGxAovOG
d/V91IsMiEyDDJrTkF1EcXCE2Rza4QQCQ6ol+upLQGqFp1qj+LSryeQlBOthijkX/pdlShPujSt8
gFNQ5VmlS5V1TCA18ORY8XTZRd6uZnENShL436ogAyAHgu6ONADezGAt7b+4klfKzxEkXz7J2C05
3TN+8o9sW7MKJlbKzjRsO8wVqQZ1nFvMWl5ns11MSuoyPStzvKpsJp4nApKIPq2eQs3sUQstmWkZ
sDLrdkKCUyPx05yF1nihInhlfMx+NmSrLbE3tkFpUuhskaJ1EjcCOS2zkfqffVjUrOxgeoprTUbS
+jdi4I1zrVxmPnjEcM4xGSsB7QggqrHBHpu1ZYY9FDiQ6nU8rhSC+tSSPWx9zyq0br9/ZMpxd1wi
j74CRn2at1ksg0l33sDrohzMcMAbAjLR5vLdOeIK9mbFFzR9Qqfl9/cmlyNiIKJ9OtH8Hz0v1e/A
bIGh07Fg7d/Oj1gLOUoMZPy3Cyk37Qlb1Re24ADnE6TN9NqnBDznJ/NrWo99qC5Ql/9oAyX2ubME
yyG7oAPo82n0/YGPouzSwcP1HyxaZADmFKeMopSbpQrth2mSKYjVL6fU0LGQnXgwXkMF5My1l8xG
77mgRXp3kEB3JYUtRcc1T/jmTJW/OikDm3POsDdAg4/I8VUhV8OHpZjC2/L5hDOGfnbX6mWA6iOx
Eicumy9bvUTJFP7rckQhCvY6Uhf+KzuQ6SEv7UQ4QL1Ddx6Z9ZyMsHac4qFWgfg77Ladc64WH+dd
v3WfVSSZgE9og3+tMtORbKqh7WZRXeMpxskqm3prgyBP0dLtvK7VYT5WS6lAMkcXk1hwRp86C8Cz
AtYyjufWW1B/HG2CatCasrsb/L+f4C0t97/tFboOEG4ZVJH0VrDolRLa/FVgBZ5lovSCHC7YJFKN
Rsr/+U56E47M/qHgY8TWhTefGa2z90G65wc3OIXLduZnNrH7yACeziFvU6YtIRZK1wuCro3gNB6A
5w8G3X/1iBPIwIaLI5CIY/9fjz/4l7IGL2vhysA0dE0dUjl8SV4O/HxvRTLfVPFkN7gBeACi1jRE
WViI/z5QGpamYVNeiKzRr8dhJlPWbAoEAREZ0JXFXJLV+N6B8c+PJxMAdgMsX4GcNvFURz3u7/B4
P4be87md0i/Mfhs4eKw8jJkmKS9ua83K5pZOG4r9Duo/g9/P7Yi9XOYdf1Y1tgy8tylT9RaDDjoS
q/9yJ1qBcGkQ/Bd1q/cZct6j3Z1IQ1gNJCEgsdcWHYJ/LgOT8jQU1xX99984wEpt6CYsUC4sbtAa
dxfzCZNTsews9K/hB91kVUQQu9uQjTjYSbMetynujcCM5EXjdWYBAS4EFuvAA8zKeRbB7VNexkjO
7LKSO6KCNdARYHIhLErHFSZ9p2G2VcUfWWc9PiHsdzEm6sHJ5p88kFTp1BRFGWpxAR6UTIIczVDU
qgzgHwkzX/SC4sjhFTJFlFrQCE11LlBG5ZniHSOYYrbSsEIZFBr51E65sg2Tcfh2fzZHzvPWFGkI
ViJ2ud1P3zfPhIQ8DOc2qj3wIhZXQTlKoWq/Qj9bfZtOEkSLtg7vFyJq1ihnxk2HN1wXXcdF6PnB
LLtZzNX3xMAw3YKx3QXOvgUx8H/1UKVloSYXzjBFR7pm//GFCC0QMeFZie6Seq5sJ+pPllivc1RC
D8fYKDwp/UDQ5W2Do1eYJIewMyeX24P2YThz/EIj2vw0SrhnrkAj+pNXEbTuI8IkJ9eXigWug2hN
hhvd/t9qCzPbWGutnsONO5sdwDR5FIEsDBypDpRU2q2JFA2frZFja8isTxxCGdUYQobjGOOpjGKL
Kc8JNNg698m8kIgHMd8s9xiNA1CkXr/Rsk+WwYYhskOqc5++rwqv6gprQ+Sfz5VrPIFFel3Vy0a6
5bXvPKZznO5Ff5vM/iM1sffQ4/CCk3oc1PH/AeiJwVXzCczbBwfUCK4JUW0LHcfxRwj7kH7qDfth
HByYlybMYY7Llh3dgzFvTrJG0RLYyKFa/LDg5Yq5Tj05B9atlYcgU0fTqbdgo8NY9W7aARFlPl8N
nFhnXvRTwwaKJsbBPbcWo9sqVHkHrzVrVdWX0+PAE3v4R+T0o3OZ6BDzii21T88vm5oOXdljINRv
reCtPH2qBuIH+YsFCL9KnsMLK5AglkfNvpWhSXW6i0m7W5SDWEWvJP6bOj+eDfw2V2w6KodHNqh9
ZO4u15at6g5t1Y2GgQI2cix7C/UjhSpzUcQaumcqa3XfawEyjorz3w0nO2rklBeIghbmgsp5xVnP
CqL3rmVCPbPYL+ATEdGATQ0v9n8yv4fMATtBgrX1KpJWsnc7JipaW9Pw0ZoOn37Ya0BuoMDxIye/
LNb8e1cEqMAIFSP3PfQjhKFRXLeSKzg1bsfaKrOjVSbIuVbDi5nF0cWHdbG0ujfzL1sAAYs2z8ia
G/grDNbjfhvhkKLJ2X7B69Ro7NTL2FclGTFWvSXhMB7c2i7HUkT3IG2eIGCmG7CTYU0B+CIFHKl9
fem7GYEUVf0DpeviB4hv60HRpxDIb0gfxQJFFb7V3KEIC+QdUFpc+EJNOaF/kxd2Hiy5iMXdLQzZ
B7TgfHLG7+MFynwEKk3SQFjP/CgRAFFiEwadBHki30a/UUD04iVueRPXRKsHFk5uVVAigh7kgtO1
R3GRf5DlN/ZA6U9O1QvJku9JoB3fnlR3bBLW9iW4tkXDKyegOEsBPyyLCsavPdckyn9SJgywPOkx
03rfqUkli00ZvJZlE6jRy9c/Q5T0Oddmh4/kmDP44prxLAfs69T0894rfqaFFeAdiWmx8ioCLVIG
uA4ueZdCWUdJjaQ7uW6B+qaFA3QveAcRpo/TFgmoPGsgzcjXAFuiEpj8gHylgH6fMITYt/IU3Sar
6DpXCJn0Iuw79e4QBn690ZIoiMh7Lwy4loTt5463UDNc9Fa6/Cmjk12iuQ3RE5nYcezwteJ7E/J7
fyqRRQZ9kmXTy+cLSxLvhLl1cmupEi9H9v8FwT5M9rq2X5dJAayeC9ejIPp9ePq8+kgRxjHuiAce
HdA6gwcEIEp6Uww6Zhu5NiXTrfoAuu3mOEvyb+DC0t+xZBExRbTxvSvwiYp2ODsxij2s6KjBykZ2
B4Vk9XpD1vJtyUExpJEKFyhyhF2KlE99aU3pNmg6duQO2DMNUCTKRy/N9B6XO6Yt3qqNK6u5Qwo+
0iXLMVONlrzlz+TIKBTdPJ50zj7lTBsCDrlMkk5FSuaIRVzb9JtRnPVobrpDDpw5c/vpv3uQf7wF
1rOhTUoytl8C0kK+TeaWnL+ZZdO7UVdn2Byiy7x/PFlC/v3acGvqdSLrSWtok8CjD5Wk04GGinHf
6VeqWGVOXdTjyasVWClQ4wrsvIMf1NoRi/stSZaHJ5fEBeaLh1/9+K7VAwqnYPpNxfmQS0bM3cBY
8cQ6Zd49KuCW4V07Am2jbw/k662X10pIxILPrCdkCoUCLiZ+19Kkw7mjdtz3SAfZH7sVxx/VXVx7
AMl8mec0zOyQnit/qLsjrAXifSCUI7+gWDhsQn6d+yygWQitatYzqkYAeS0lewuZzhtFHTqiudZk
HjI8mtBuBuInq0/1vjX/FuEsYXOOXFcclTztjJw8gMnZ58vdp9rMEMDeF959atRbVmU36ejKmXFS
vyur9JgBpHgw4HIcXQ+8Lsze66BN1VFkKAWkPMgCp7luuo/7vXTEVx0oILu67VTcuMYy0amQ3H5t
+W0nLxkO4p9+AwcKAJbhfbE2ktKoNQ1UIgllaDbfLEphTfQUY2xbIRSpzFgH/Lhy4cRcH+nsM/k3
p+fc6olSfZVbF+5E+SS2Vac8qTexTGGoIjmXCOXXH5eh8TDnZdbuzCQUmOE2lzxbX92LAuopuvMx
C80bylHa2F7OoZ9b4+CmbfV7+I5Gz9Lm7Bmmvxb/luckB/uro9UTu/6mM+DctRGAf6TgIo5WFcG4
JN0E/jH+m1QZzEQwxAY+U5DpmGkMjkC/S7S6pGnScuvbWlBFr5leeppe8UanBxjqn/37xHzBq25E
+uopaW6SNcGsMVtOYw1zayL8IE80mJqLjQ1LO9kWSAdRLUzn0ffkGfTI01nm80AskgpGIRmDlIzA
n41jXAAVIbUTBXXLEQlrj945EwM4uPLymWB9bpwcoDOntuubD9odaDU+J/vrByFQKMDgwTUHYWNa
QotDHfRLKAM77LkwUvJs7fYUNN2faKqx8SoFrrM1IfyZf6QCggVxzETgOWkQUxE7QTy/UNZMOwx5
/WgOYoTbFazyy0qg2jqWXNx5Gin4SuyI77LeuKp5vMYpF9nB8zZJ99WKpPd4HJ5n7p9z7WIdnFx3
M8An0//ujmYmr3fc3rTnhS2Y8F81a1hPHYIK6IC4h9fV4MwBa6Ut339mDCBttMzTUKXSQ1rb+AF4
5IhPNc6TODSXcmY2SVicr20Horn76ZeHuypMD3RR8+hHrC2lODHNgCI8jDf8VgZ/fUxjc+IZyebh
7x9yoDxR/oD2MRRFeZHVxMs6+ezCzMrBxSz7iR0jaammXtHzQaUAJLEmLIusCnHAVgqe+hXJp/kv
e0aNP7qfz8qtQ/7Z1rm2WYlZAHYoqCevJ4czavZhNZThOEqg9bqDqVcN52xFXLOwQg3yMIPvcV++
vGFqa1bFMwyC1vFD4N6y5HrYx+tlskMy6bmYQnhqp59WLgf5nxGjbYpVUdJS93b04hZk3PtaadME
7HKolA3Ln2iB8m9DCzpp4IEbay51ZFfxImpxQHHyKM7KCNThjNHNetccU7ZixaaqAXnRpXgUJjN5
3XbexhVn6mgHANnv1Z58V8XmRGKiznwZ8QFiiOX6LijUPfcW/N+qio52NFH77tZjCRJdgTvFH3mS
bXfx26K3sDXIrxDdVkg6Ic4fuIKk3v8WNR/Rnr0RJzK9e304lWSlOpSzG33JBzW41Yy7HQUjVx1g
xldtmj747AUGN+aIOj2tdJgAzhnn0rLcrpIBHDcih9y3syDXOquruZ5ynJYnc3ucAvDf25EJRjY/
bIzplVf34J1cD6BMjYxnnmyRvGtihBXiFkHMM9eocsoMDEG2A/5UpJU73YbwHuqZIY+QVRB0Zqim
+PzYWnslkSSWP4PxGBIwRq3MRvuIF3RNQtQZ7VUKZPu6Fr+Nku/v18wIrId+5a/FfstIpsSgSr4L
M4z8LfB5o57PCaRQDkPFo4eiwGttuP2B6+qrZad6YWV15pIajAeepDiiCUKVKpLdePYgy2VGu5Xd
sw7peQr8UhP1ykvaLDViBTfhNKV/xCN9KEi+P/gla6/QsHZunbUQIyV136pIv1O5Xmlg2PeFlXqb
IYHEWwJRI95A6WCB7coISmw9BWn3PnN+3Dgx+cQJrOx782Qt3y/7LOMmUISo717cFjsuYbnK9NZh
A65HZtgIkcaBiBEzm0o0cXXOs7wfct09BwAkQSAoEJ+ufyAi9xW1elEdQYxMkZYTsYjnqqYZB+QX
k7yfekIrkmDLUnlJPieOjsQbEMGQmeGvArIk/04NNBktzdi7OEvOFcDQM6/S+bUQ3dcxYn8OBGQt
rIaeekYZXVrJoTvWHKnZhaFEj1AHPpo4kkCuiZ+sCEAsUksiO78XQPwZt3kCV7ZQ4Hf5I5HhiPMQ
+iR+fHCjJJWtP8Nc/x4RJJyomFLWuxHo+7PunJ2W3wNO/eJ5BPVMjZHF2Z6WBnTQ9Npjsp56R5z+
0Q2M+hkSOi0haAxSaXxBQr0MWSoYufm0MGNCrS+x/Wksq805pk45PYk5kuI6FCqSB/+NDFgYf+uh
I0A3nGmyjzkMgKvuYKfZHhAVSaoac1A5OhSIZWGCUJwMGRVg5XluJf1dRtyrwD7EXcg2+Jk84Rtr
0hHKO21xR01ZU5hrWgl0Ja8D/EnqUe1OhRLnbkZVghKmRvkq+QlBTTt3XU8eqhsOzQLft3+dvkZ2
aq0ofpadiSfmIhTC5TUtqBpDhk4IdBezPEnkuIKfe+ItH++G5I7nz7trv6EGeXcX2C92UC3qc1hL
WsvkbW2YjYPFCOsJ1QHvCSh9HQSfgUqnocO2naWjhKXA286RgYAp+8kGAmiF0o5UNfqxy7yh73L9
TXlOtp+KVYJWsTfgp5Jwc1IaWKaHoms87WBO91Li5+/6NaS7kqm4ieyiGQ63GJCax/4NFxyexwgE
z75UuZ2vRuc+NOIb2cZtcbkjnsSGROX7OPeM5a5kM+3fKNlSj1LYBPmcFlQd/nYqcUCAHR+VSyeX
9Xzvr2Jq1RMSi/rosTvp8Ku2ijXnORYf9OJXCe82+QRCFsot1Nj5R6YQirDvVrZM8r2h0NmWbIYl
XPdCFhLSmz3ANatoOPo94HKSBSUBEUuHaohM74RMv3EtGIUhvnT4UMc81fBJ1h5iIzaozk1ihyK+
PVEGDUot8odsECgBxmWyw7OQ58YXxJEjQpUyCrMcL0k1976WzlnmtfCFeWvZ0mWwQ0F4Bq6bqO+c
2GWFo2qu8hR1XiA1kKNgLd18k7JwDBDnLJ+yytmHmZHIqqvgqm6VejRoUYZWvoCOc3R4RvjBQRKE
mL+JIoFTS0K8U5MK3unItZ/A10FLL0uwXOA3//oIGoDUlxB3pj1cktulEeTotMBpbmsyhFgE5Spq
iIyAObALAM6FGUH/Q6rAxdolMM/AjaIeTWCguLqEzY0IKVBaiqGcFMAbUNaIW94qhMJkS/YGXdC0
/MTEyk1qtDNLVvLVNF8ewJ+8kEk7SYvYQEt2mHYEzO1M8aH6LUGWZkPecARm1FLaXEXVR88HCDQ2
+vkmHBX3doDxev9m8XsrRiDbU40qjT5268GWgU+u/59LNqEXz3jHRgF5qhvZeKy51rK62eJM+buU
4MMny0FoEmQHQ74X842Weqc0yXxLSHhWkZuWsQXW9BZNoAzTgjHdxfTgPDJSs4Xwchg7hObFn/KD
FFuzuBqb3u515Be1XZ6v+BIBK+kMYaOrRQ2ay0Tr01np/WXe4OYVdCcIfVkNpJQkIpQ7EBHzL1py
0jGcSRZRgGj0+C3qFQfQ58sMxKtqH9xhLotQjLX/8jqK6VD9F//87HpCtNMIz3ZeWGdCTksSt7Td
uYrwfAulUADvhN8lT5jsATmJjGiBwFvaK2trLC8wExgKo1cOXrm4zvoYI+x+Q4GpHeRDoSlWRmQz
WV9RFIu8VKdOhf8pspvt7exvamIwvZzfjIEBypSub0J0oHDNtlXCO3ahIe+YAwFfrMmKL+iGfcxr
klSR7h91g9OmBmw95Ms+fJ1s+MGqgMx7OQkJ7BUDJA0Hy2n1SuUfFxpcH4E+F1bixDh+S8s6/dJG
hcKy5UpIQziuvgylWIdOwROjkTqa9RuCXGX+Y/4wItoQ6KFoFVLK2lbaa3BHZfKymM7jS1ajyx6c
o1izZfmLWaKylZnb4HAj2AbZIHVs5DCNcwFF0k9EHEiFBvMfpwshDPtANEsK+WyHSXp3bO4pPwI3
oMoANASw5x5c/O/UtbNpMdhgBUaFBW/rxxC/pXIpCzofr9PnY4dRj2S1J4Fad1D600qCEmx4PMj2
SJxe8zd3cHdlSZmPfvCqVJdyhZKe7w3JiFtTQxsVaTNBzF/OK55BKocliOoiID4e44dblYqJ2071
hQrA/cIKY1jpgQJ6KqNDubWQ4olnKrOiTnzn7KjlBUGGQxiFsMgiRcSnUH6N1BMvE14ljwUEuj9Z
xi0pb99QLlgUHwdrzgiun5+LPs+Xd4bBcSI7B5R60Fao1hqwyO34s/j5eS7yhmoBvoK18OSPrC3u
WJXhHc0s77JPakavC86xVMYF+DEDvBi/NX7JtZUZPZJjSbuMlC9zHHNIF/MQzPVDI+rH4zGNQGpl
N4+JKw5RCryT5kaL/x0CEv9cnpvvbczXqmMsgbQy0xTeSqEguRx+cSRM0F18TWa43LeequCTOgyR
zEDSeJTQdp6Ng74vJ9DvxFyQ5CNntJmCnxAXTk5BRnmj7A5bNuE1SaMs5X8hIYMeFIzv/0U1THiG
eeGWvPpiEiH1nCYZuY0BG2TvaMyJtU3E5hW0ajrsO5TE2h53ZJhn3HsjfEOujK2Q/25esKjFgdbA
38ghLaLU7WoWcJAJjp8nWbhohUdTI6VRu3fJ6+k3qErj8j6ItlmZz9m5xRXB6RFhGVmO93H0LlpW
35SF+yC/l65uUUUASKERhUqjHD2BAYaLW3YBnZI1rU1S+LXRVHmJm2g7AfRlmWrim8p4KpFZsE5l
T1FvGnFXLXfGo7RtKOxFwxF3OG6t6tlBbv18nfFBKrWJ3019m+UqxHb37KerFAqFXLYX9nYrG9Sz
4lCnrfnDAaxu47CCr88bhJuKOFIf8b7YH9pxm92Y+nbRfAeE3hKp4GzVx46lJJ1BgFlO7hDtgxVF
UPt33U4LcvlUMO5zIZQVBNnCfJG5rzN5BAAwXxWgWGrZyyFPQ+KH3uW6sSyUcpX+153sOSdCGa2S
g0iKVTL4JeCPCoPKePtaAPlAvB9epZEkSeJ5b7bK6HxgmVUEcDyOxKZFc9ajbBj9LUgdIHqd3STJ
0BnM+uGpMHW+PJYlHR8QUTOlSD8oheDauTI2niP7SO46g7tcEjBoc/D4V2+TrSGeurrjOO7qfy5Z
WPSpT0np2TsAbKMHM2swYzNdI4rsvN2fXMF1lVSSTNr/gbMwcP43Bg2d2N4IGgfa5UMNpcrW3Lgj
KMA7UwAwL5DjltC/8dvSVZxNFHThqdSlpervy6I5PPkTP7lmUXOfhEuIJTWCN3GkKHuWgmZwnb0G
9mPJmQwp1+0CLJdhUGjQWy/taLA6GEminJHruuVyImQn4M7ibu3gbToKGFzTPFSGG5mF0wDCdr7P
jLnpt8al9YJOJOZzbKv3FhGC3Qg/946GVtIhKNQDumeXkRR0d7omvs4uEt7QCqy2V7g53DUfsWkD
NdQfxfkRFPjBmww6HM4T2nSkx8OQBp51LU/yVHphZtM2ErNaHsDDdFZaeFAc4HTa+hESatqqTHpQ
tIrGFvioud7LTiwKWPobaH9X+e/uUsfBOH79Dh/ZEZkF9wOiHQFpqoO+Juxrz1raDtE949AOuHEj
08kszlK9D0qM9bISN6Sfblauf5iaMgqY5lUnDttEj9Y2Ya5vuIaUYfhkcuh0uNZg4haGCUKLAkYK
39/ouNNQN7w0yVh+2GMNRF+loBM5GBEWyfzfzCfb3PI4Fm/j0H7xbtu14WYcMPEEIV+mdmEieOU5
4Xo7+br3Wmfy6XMYKFBvx+/SPWglSHeQxdQW4e62Gw+tqTP1PdNQhW/6WLpNsKi7qsD6tDs6EWpp
rSvzctrUBYn5bhIGtyX1NdyS64YETCsDuluo6tFJKqYS5oNZxthtvWfvQpZyhKmmGEO3eh+3Uxw6
kckQkiT9WFeAmghzgfKnabbaNO1dGVQGfsMsjkrZOgJVl+S/2pYJMyrY1bEC+JrYOaVPcg27f7XJ
3LLz0vFVrwL78eksfGp9A+VW9BYkLN7ZxnSiUFyoN6fbjHeOCXQE/DH/xfVysWgtDyqdNiesKYGS
ALiiBC/TMN/Wj74K53Y1EC+HLibzb5uTKbk2bIZlWJiM0I6qN0KXbMugmqN+7Ta835VsPetM5RD0
LIqjJUNof9o9aR2MnpUE6iHmvDYyHyrnokVxvwfxbcIrpxhKUpn7nuMx/3njKs6Esi4Mc9ycHDCI
n+QsQeKQ0+aNJjZvmJBE/GKQz2B/OXCC4EzaNGgHVBUMiHz9Z8IRl43Oj6Gh9FzYaMy2I2hIlhjY
lbn08x0FeiqTHIMQTkY/+KHhRQ9Mm7PXh0aJU588in0jUvByYqfl1PQPKfY2IhrUlrz5Yu3C9ltw
LBLde/xQMJ4tWynFR+LqR0vQViPsQybI5Ma50r3KFlS1+EvqMcwch39BhFgdhmEM40MQA2a+88fk
/F3I1nfdxECRyK5/ZBudeRnYAdq6GBnkApJ4dNbyfe0Qm5L32d03hMCg+acPi5u7k5c7YWEECmhT
2sKHop6XX/Nx/JlxFQaE8wrXCiFxIJLWc863SZL4zDQ5CnFEKVkNwoqONTydFs42T16B37+yXLHx
BlUv0Kog6VgjSLrl4MC52xCt7gW5q6uRP4zGZAiZ+lOCMpWIe3JUaBesqn+6vid1E5LviijOS8QB
w1Px5Jx9GvuYhgC3ONxCa1SBC28b1OQYCykzC8m0rb4XTjzg5aNFD8gWhQ4PLIzpxOiyVLRSoPNC
GJ2XjYyjC23J7kdY4gmbOPAVHslsTvPV3JXiJzTZ7rqnjCU07DclqU1lGVfKPBv2FJ5vjWxl7V9K
sXsqbTZzlDVb4+1hhmgAlDJQT72A3rzwe/o7HN6D4ukIp5Y+mva8tK2jSwkDEEqPRJnODzrDKn0r
V9pKYR0NzMgP7zIpo8+dQkZ0kgdVUtJSQHnTZA+VatO7n/4TWC79SrBXx9C4Y0bFcpEhJrfPyd5Q
I91rod+af8E0WOJYTAIgxp2E2lqhpV61e5Jw2+8GD4X76Lqr22/BAWleyvJAr0igXGhLjNeZK3aO
gWnrsmsIHfaF7Qlc5BqNrwAg1c1yYYFHyf/1ZS2z39FC0MD5JWPsZT2k71YR5EWPCDP6wpOvXmpJ
wY22qcyYOo6vy50+XlWGnJ0yck9ceN2WBXpL7ALB4ZQQFf/7Xi6/04zU64rFE82v52UTE6dpLrHE
7K85yzL+aM/1MoojroVSTxybcOtuKgKtSwel+fPDPmB1KwWXKm5DZklx5qb2hQa8JqwdrmMIqlm/
PIkrE4+UBbVENmKKnttWuuPuaAf/bBM0dd1W0j3W5vbI8xvgPDp8KdO+sbRje3o1InSONcMxScwd
dq99+z6kiucoCFgNQXWyiQeTW2th6FxW3ZJ+nG4lksoEln1hPXQqobd1qjFu6jWQjShec7XEQWVG
gkCsYmt7JS+aY3AwgzKktk9LpKIxzULdVkwrB5tyj8GY71ZVXzLFj82XqCx/Yd2eDo23i5GPD4fy
al3fyNi/QNOirVxPPHUr/FylPJPs1wI9Jem14giTAZYwUVDTY5XCoyTZug274G7INvsPrH/fU9E3
VCTd+z6v81YBBEtJjYFl8akkAQWh9Y+c2OCYtBp6wGAQf6dgXXEoff36+8xzhyJ9EwvJapTngH29
uLtGO3eHfPlBdpL2OxkzaG771cwo9E4TGxxdvfjxFmeuki0I2JlZYaBmNptlv3TEKWLvBem7lxbH
O8/giF14JKdV9mhOSoz57PNyeSCq0mXLT7ovmCiHjZs3s/tbb4OtEwp03JRMZQNbj6dfxsxvvUFi
Hzb6d3C4EV1m3ELRdp1LlMgzrh9yplh4wxKU0gNvMf9EY0UVxNx/4nMiKQsUgkXZO1eg0TNzwO4b
757t7anKFXJZUxvRb2r16faL22/yfUyfqAAjBZdIVLxk0pT1MzPr0GF3C0EpXRFUYcWJfbXqqxJ5
7+1WJacnKXCZgQ2WLeQmR6jwNJNr8W9uGUMO+adI/z9uo9jBRyV9aPW560ZjZQfp+2TGLAQqw0YJ
MgzjmzcreEbCuIxq3+J/j5njSIhGM+8OPOCr5tXCm+MOfrHOhIeHFXt9AJKDd6qHYRnOUS9bxYet
P5wQmArxUK+4ZC6WVvWFaAP+AU+59FoH7mkqZ8wlmnkpAv+49Alo4+TXUFYACfoAfFQfXJdX6hKP
6PFVWtRXQnwXS8INsMI3PA3EGrEoBoVtW1OApX+ZkKtYbdanh51gCtMAhU/8vIz/6Q8dhFtC4L47
EjwHb0+EJCQJvDsVTIPIVFSWAw1lf19l97ZSFGrxiD4wbNrGgOgIsBDgStU/WuDWQ5EV/k5zlj24
BdTvvgelN26azSEFfBluRu3NhkkRoW4htXrcn/qELCDo9EZZZAkvQJAFcDlZF5NoBRxDoPozw5oD
PNI73lPQ67GDRn/lWWuR3HoezPBiWPFUT5tGAqBS9mzeA0DEex7qLdbbH5r7ODE9ww8oEK8awyFx
HOQi99lpxjWcIrHTlHlECFTle/TdmwsI4pBTflaPBrJJfut5QC2bOPGR++aMZvTqElQDY13OSQVS
wDe2Yhd4xHVzyMz2jjh+UGapC+PBUvM8EHD494vDo9NtpjxdiakJUTxokAxr1qGNbVT+5bjpdhHW
fcZYO2H3uxXSsSAGYgVi4xr19s5C/SWrl12Pe5H7F3CJfLT7rqXdNH1TkIEogPKcUuyiDPReAUDi
gGKrxK5Aofg7y1t7leqEDHh18+x1W8cwnjqztai46RBAUEIfV2szfINSGjKPAtuzWdjsJPjcZSv0
LgTDqLwtE2vyt2pP6p+kAIuks8kiYOZ7HECHCZ1o8+x82+LUX403X1LzTxi9UCTTp6dWOIDc+P9N
aZLkaCU6ouiyoowpWpXw9dGS9jXC6ytL/aiiT5RGQpXKI0MumTo/P66R21+ZxB1P4EsOpgRK8H3i
P89EAeA4AP/TprilFWpLHg2q21kMzQoDTtlJQh4vOVtmlFggNGvHvvwFShL8B+/my6Df56ZrjAf3
MinhT7jbQr4UG9AzB+9UhURctq8PDuAj8mVXxLvBI/VkgyT0ix2CNPfZfTBP3fNrLwhXDpHm+Jbz
1KBBQGwiO5De1+AOZ33bztIUvVyeK3LT655b6PnbMJgh1PYXOU3QwaFGNfVKHOJkb11Enzc6QDz8
YnfyNcD9gnTU3K0I3jRrV8Tyqh5XZt7hWT/pFUjDTX1Cvk5rzOXtG3awa4Fbt739eUp3FEhpCGA2
lykzR16kX/uE5kF6QCq5BaXOlNqXeIPK+B0WJz1ARMzbinUq/m4jeKpJtVeWwxkFOPoMWOVWmEFn
hpkCSjwMTbH4M+bVIu143EDgNRFh/Bxles5MVi6hFYhmJmXg4ZUmUaqmNnx8U+NUuKm+o4SbxbLH
1DLOvRuGbZYh0elTI/192rWUPYtdb6bbIAIH7IokrGpuFNYXJ09u1uD3JqVLn7/Dn6RE7vVhMVP2
P+CpXp7nIML39wtLvl2VOB0HVdxVvElnF2qsZq+FhS99yODpKQ7+3Ks/iWlvLOB4ovs/fAkGpW1+
iWccdAmNgFnufvbb/PUWp2mEO9fPqj++P95LMYU9VbJlCLY08Kt3t0Z9Sy9pnq4B2Fd9qUDG8V6O
SBSmk9wjvKPbkss1lL9HgG1VmWev6O6G16Q84e1FDCGDxBclJhEVk004az59NLdQh5ekRByDEZkm
5WMNw6UG0CH+oVFMGhavv9jgMyH6KDEC5Fo7+bIe1+UyFfrGrOYSP4vKjerXkIRH7KmkGN6e4iwn
JFNh8wAZkEUc+EI8q42JM1JoRVqcbhednitEAyRxq5KTZRNPrgb59w9YcDXpRv2U+/J32u/vH+2G
ppTPXOK4K2VVTV7zmlu/oAcj3XI9TO/xTHPP3i8pvMCTjae8Rs+Rs7XSFLF82nWyH0gX7IuVZOsl
O22g6IthIPiWVo5fJIOjWzevDw0nv484q1WWpsXbx7U4fb8k9I97CUwjn5CjsVMmWgAvLYtVfLIh
uHzuw+qZJVRq0OvPf5qo9DLoNj5q3wNUqf3he+9IJLsgn0tYIFVwqIyNDg519BSbZGKZFBp1jmpu
HI65U9SMhuSS7NDeDnMNBOZuf6aQVRga8wroZoJbTyjj10hpmoqFaUAzOtzjAm8lit5MUPMn1Aji
GtOCkzK9wv86/8T9Dd+jhNoe01JvlNPQf8CfaKx5PSzUWKNL8JRY6wHltjjuOaSdPEXHzijeaBHb
s/+aml6gNGvLX/9vFtjzHYhbvE0bFw8IhM1Ljx+xl61rA2gVQtGfYp5P1HGGAdJoMpZghzVZLQlr
2EGn5fhMxnE3ugFSFh8hFwQeqYb+ETl204rCwQyRpZu1ROLNGp9oOT7jEJVIf1oV4WXo2Oj+1qly
kQqcH84Fb889BLhGaS+jf6mgL08MTWssAOpIXJS2xwf6c5Fn5x1EmedTLWXCFqjpqL8UqJzXIrG5
YYqSTpVKXHRzHKoRqALTeffkLqJJrFvPbx03qypB4xBG0JJlPHwbizXUskfV+ZQCMwoWjVB3u1H4
H+YYCOt0UONL/7rnK6C628kvemHLR8c9FitK66lmylMza81N913RMz6VdLyfMsVErKDLkyIuZnYx
WzBhOKuJlrutXowpy5ZzKtnAE2g87npH4vRtWCT5kD3AyYORNaSfbOTsCBW2LHGoOJ56QwbfaunE
Ec9voqBFn48OWH/I7PYiou/Ev70Pu5Y8ImTUdGY37kT/N++J485fTEtdb7RAFIbA8v9PLiS5SaSG
vMBuBVOmaBsMAxj1QERoeoSHjiS5sq4EtYHNxUqdUcdHZpkjJxZ9O2+uiwuDwBtuNM0Q8dV8xdjc
mo5NA7Zrdok73o55/NHkL6ohwvBcR4xDIaS1Y5zUzkgKmMbMR+8exSD4obezbelzhFZK1hXDndmK
nb5y4aDXGqzYdX8cKxycoIYp6Mq1saVkuqvuXVMJ354pm0gpaFYGkg0k+jwGf83Uq9IpEOVLfOu5
hP/powtlUO8dJfEHKkTo3jAuftYdQgPQBN3KWyKZutDgyqqeclY+vQ9NXvMuKAgLe5u5Qd4/K/xu
thsyRqoQiXvcrZTIkHjDPX7JbnXGvAYNelrl6S9T/zg05C/qcTp/BBuIgCdeGd+i22df1Qk+7ph4
CzlOiioz/olJfPkaJt8axxDuuk9UGY1/1wX4f7tAtwIzcf3JA5uCrAdTnx+wevtQWABJ0wQ5+0NL
s6FVkwoLu14SLvvttqrpU4U0IO7HbP48c3Cjw62iQ6nNlbpn/Lb/bZvppZKVd9doGvywJ6LGSr+0
IX8Knk8DN9KhYGim8s90BV4KT5oeWqsYlv1gmwMbYSxLihnjxg1VNdAR1qm5mkaQXFQBhwGHptal
cbRBYRwyFrNe8L65VVYD8Hl5uXHP9zImaSFddO2bMr09T+/LAPi8wUWPRhYJXhBoNqZUqBCCEIiV
M8n/DgR6mLCy6c/ihE5cTwLgMFv+KX0TY3LQzg/5cLXO9fsZvBxP6VLQKGBNKWJmhNbCPTqazIhw
K3TxZ1vhifXEYI2o7peHbxLjBpTzSs1Ew5y2GKCHt7XGMMGffOtEFm04cfNpOnKHQi/cD1230jLF
o0vxz0ek7QYluqYL/vjYGOelQ7CkX5C+r7di+Vya/vU60oLsIWfoqsOYwPtpHp1H3RxQRTDZ3UsD
Dh58pyJGCgs9GgcdnenSZiU7cndkpg7zFt7EaEYUJUhCDa6YVngkHaBqjL5DtBdQ5T8AUsNRByrQ
o3qItyEvo+8ru7hDzhFm0GUWwtoOYWbhqt63x+VeCeRBs08p10XosLB9KRxpzWt1Pt1TzFodAMoW
UQ2uuxVwOl3b4nYV0nSiEhWjz/JwvX8VrdgQ2mQwZHSXap8DizBuqiuF694lYxZsKAcm+F7yxWh7
IAQf8hgaVtysIL1BNelyQN/NLb+rIi5sqZ7D47KudPMfWmXBkZeQKY6brT1eIR921CC25UgalBuF
CrG6DNZ0vb9ClF67zRVy0Fn6W/YPL3CP6EA33nWEO7VAi/GK/2ch/7GgxoQJcp/DRML462Kqp65z
u0PQgOcfo7RnGQhav/pjQocC1K6yOFOk7qFai0gUA1UzqLmmoEk+m2++A6VxighJ5bwcxE3vewTX
nQEdgOaI4dcGfipPamImMSfHCc/6f7aaIFyyCZQV9Io85R9T8hygtBwFKpd5zG6AcOAWvJUH5Za7
j+/mua8JldzYS6630frpr8/jCLQVIDLN2eJQVykHARwYx3x9YbXaN4CGoTBLcqrtF49Pu0Hyccsw
1Yy6G1a14m+lKJ2dHANvBB4dG5Ylo8D09oD8FahRHro0C33J6SrYkd36Tp0rjSSBB31c1wWhBamw
L41nT5yBqyABIpgdTC0uZXsp7tZ1CIe0Dsllz4a3VXkw/W9iE0+1A18/jklU//5yW9gu9nWNQJyr
EOQmBJEjlP7UL6dthoR0GQfcy5kfXoSIZ0M142hV1nyzDyqckABc/lEEc7ixcbjnQDf1etGCglDc
HxoG6RZ5pp7ce54jQEZWHHkfuvnzpbdA1cwj5k3fk0HoSSG96SrLCwbZWbCc93GWHgoua/w9m9VQ
eUrpvI+HDnDOJeInke6l1fEVG78LN3N/NUjJyED1fuZXa3OkljfkcJ7UXKzBlkNs/Iej5WOSQwSI
pl6q+c3tuGhZzZuMCzk4WAODXfzxflINKL0yENvRyYO7ZBuAavu0ZB6Cjz8NgtvFZ7Hw9HuqqKO6
nbikjNrHDDslVgQqktsRZ1SIgxdoBuiSkZDCw2JU0Ydt/2LOz+AEpIAZuu7zn3Zsnm1AN1y0nPOO
oGKgBextLYoZC0JxPLnt6HqYv+bctOXL1B3u57PPvWRIcofvuXeH/a0hRq/GBc3UkQ6vtR7q0hrs
CdGBYdiEt9uRnPGyUyq2kol6gFvdyCM8DR0uCyzkePJUagOX2A4dMqkZuLxXIQSHKHq13G8QHz/W
O1E+5VPHihDRyWPCr0f1KQ7IlDmItMeAIVQphKhoVj2/7crVyD/1zQJjKxN4mokxqQqWTrUdAYp9
7NsPZ9RZXnsqimQgvb/hZyco5OGNffTeQvmg1C4gFLIxEH2oPxV5CPhwtwQTKC1/tiwcnX/ppoq6
I5wBj/w6CFuknap4RoPBR19ENFcANURYHi/TtiboGo+i49EC4ZwXjEt2TdbdK79w/DnRsC4WGjXC
CcSHPpm+KXC+SvJbRZGd86VEz2oHSKdHNpLjawkFMb1dFfegKiVBNA13DcUPuQB/8DVVTE66m0/f
I2kh7kn2c7znU6clv2dVmG/siCAxg+lUV0yBBckSC+uwHXNkwHtCSgLfNMGpHqZXWWMu5tJaNQ7S
gfkLF9FzBzgABZ8mh/tTRTHS6fEPRWvttZsC3rrWl9BjeAzTLfjPUr4HbZR/Jc2wFHob85ORx58n
jppAIrV2mHikJC5qeKM8xqB8TMKpLK7DHT9szRLpN3D3meU/0a8yHICmYILgZAk6AZVMrtauuu61
vrnpczrWiU0fhTvH1osFnpPWAxMoUTvU8gIRKbJ1Evgef8FUAznuL8rPHLEOUt8IROV+e+fvQBvV
cr4SgIlzLcE0XQWYxokMSCremuygL0roKTN27iZ7tPEKdZDcvb0VN9y/qW6ao3kNhkTeaMTNmxCp
5aUiKkzFxd64AK9ar83wkkmiVrR1NBzeMFwiwFEZNpT4K8aj6GkA7Ap41O5BaP8Jdt1SYxb9idxA
vOpv0zEV8HQmkwgwGsH5zXr+M2W0ryPUbHkoWZyOH+UDbfsOtGS6YN42x+lWcFykWSPr/4NnPyEp
1UFGuzpdOtwYZ4rrKyeNXamms+WiKdikvLJU/UVv2XBYqOTTKH8L45SFSJof3xFbJGdWJxXCtAAi
PBfLz/e+TSg+E5aP6d2CRI/1YczIDPgc394tme/bIQWrmA8qLwnt6O3+kuMbi/zT7iHpUfKFIpVS
Ll+NEV0WXA2hdePRwUpIxewyR7nWI0UejoyD7HWyuhPzuO7D/3l7jqs1ExyjoZuinFzGzSE9T293
pzaJ2vOolcNbhVZhAY0ruwpeLjw/q/9D//Gz0Q8wDtqQspxbD/mHq+FrIo/vN8SwpVGe8lXQLdmW
UgxJGpGghFFct9BTMZD4AfLxlVEUQtzAvE6nPCOJC9HPbUOEHHrWGajTev3vyOZU85y0D6sCOon0
0rSLEZWqb+owQ0nwwUgpuVa6tp993/6MK/RRXlLBQe7YwaUkgb2Ofk5rBU2TC5DH/3kr7GkSwa9L
QaMhMbj/6j3oZwTBAPes31d3t0BD+CMLJWDXg/oO14n3N4dMEJs82yazAqgNDCzMnZDWYIzKDTSk
29MIj/P5amuaKVbnf9cJ/mSuavbOLSNPfak4D4HrGpsrR1knoiK5yA88+1pzbXd9NLIuomq+sNBU
CnKcfugE4FCt2C8eePg8eoFBmH2Rcg7GajG4ibx8C9No3T4SgfZY+9y0lQPT7Yt0tBj56z/tgE/C
3AkUuBCF1c9xqURPys0J2bd/3hMpcwLKDfJ2M0LJCl3ZdpJW8pUyDAixEpcF9VTppdM0tPSvETQj
fn1GhbJartYf4+FZiUK6f+yNz8PO/pA4eKTdZ9eOEAONjnug7rBnLKNGCXhGzgNTqDzgRbgsozjJ
S5qNIKJH1AJLaX97CAZEDXfg+D4e3kelQLNUCSVy+Fgs+aMXosdmjjH4j1hJmeyqw+l4Y67tjOCE
oh3J+yHd08HWk17/3+8EQO9mKkYzPesaUldoA4WM5/kPOU0HDEmAVZ8flGmbz2nskMqJ7/peNI23
K8zkEDe7sMywxp6K94D/1kXAxKHFxULIJSe2OmehCnPFjanUekfJeoQSQhIzCNeohfqU4eTSZhEF
5xYjTBju8x7zLFbgajxp1W087pHbgNuo4rHGz8UdfWQ6hxOZK4jnrVYEqo/WEBcNyE7S0FefKuk5
6fC/VjbmnWXzeW8rrxVfjicrwK4+kKc+ZxPuSv3AiAF6a2asbPB0exxg3qt5Eftsu4Xy0Aq8KbZz
d30qO6i1LwfF/9/vOVlQMoJCrXWzFzlGJhuzLGndKJyl0rt89Aiv/2tlBP/ve3aAHjRE0f3J6mZd
DCaHX7vXsUOc+bvs89SAYD42JA6bc2gnAfFHraqCHlgDBWBX05qOupQWvxCjbyMxZULIP0WdnRei
7ww+tRVAoEobwLBFvnggZKdvSnSdFJ4rnyB0KDRg3aOdYQIg9dLSyXbfBhIsD2N2DoLXD7ZYpxcX
Wmyh6BmDYW5G4Rzvk+ppSFW/EogDhqeAtug0mzj9oX+39ft3zPhx3jpwdSjoHtHuaJ7nIQuvYSNO
XJDvaNHLlV82H2dLQUm3q32eBpX0wBu/NtXIBe8BsJv5mfMjnDBurlwnxxUtZCwy8lozEgcSRgxF
QnXsT+S5DTC594iTuIcmmif8glZrgM0yW/wyHnjYZ4TlYSL/EhvN5YnrMfge+wlhDzHdtM6W3nCB
sgg4a7aKDAT6Kp9mna45XedlTRnDiPNwCMSIGRRFoxrTrmA/o4REEqyXF4+yBRe9aLmRRlFFBCLi
fnmedYl47G7BpE8k33jPxW9LhwRhTf2SPI+0Nhov34lH/usI5p3TFgy2TOONummkXtuaJfaINXNr
uEhNUTzjty6G4EPniPPXyQZ2u3pbsyMOSAWO83wTrc7bctM2pobQrXHIZobyWmp7IWBq57kal55c
16eUpr6ER0+Db1vIRz/zfaN1FwvXVsyct4QkEwfjVDzyWAthyV0QxWYaMhXUuiHpISBbW7TFR/aa
VeNmNXAYhWjpzCRuKOmdaOX6yqZwxSj/I1lNgjhwcb7gRyDRTZFdcNIu0KxLgVwR/HbRPfqDHB1R
eZhW55mcfn7GVgDXRzi1rOmtrSiSg3IOEmr3jxXX6EaPy+LsxslVvWqEhgd5jL00mZ1vPlHV0jHB
NsEV4asOH8jFGW+URB59+ofuI0tfSdN+AurkRtyx1iGV1CRbad7bDPhox9jtDlYVr7ytAYgtW3uI
HBrU3TIu0o9U7ca1HXSV4DmNRBbgD6C+hJ/uSmUWtZ36STi6nUoNXdOInWVrri2CR8FMWMPsT6c2
VBd4pRlBOGxLTUGO8uW+74ScolABgWnCUujya5UqsJKbhRzSOhr8zzBscOG9XVRT17Am+khK+buW
jBiOA01eHRlJq9ABU3loVYVXd91bDE32+uUF0dlLGTYT9wkkbEJeD01LhvtGMM4Z1q+he5PXIQ+I
v5gufUzZiLGGbFSs5Y77Mt3eOayagxUCztP2p7e839P6TlTfI3ibEDc5KdydSGgTyDpqeR4GuWpc
WZStTqQdALNjgZ6otu99pCg03P/HCKIHhBL6BHQTuonCEU3wcIdZ31llpXOQ9EQBOM4UFg6iQDm3
POt9LHy3EpwJbOe7WP8Tu+OfApuKvnw56hcz68strbXYLpfz/NCMRCrG9NOjz92+LwIWivoi+OcB
2YDpMqv0JOuFptMHlMLgvBsDke+99WmVFfH2D2F7zfOHsMOcVWus+TglrFjeQleei9LhnKsbFsos
Qu7uetT3t/Pz6Bm4Mii3MOyP59scZGSqnusc9arcEtUvDBvXaW4707fOlShNS4tegIhEXVU8AsmB
JxbfjYeeDyJp2nOrmlPyBvlq7ePEpXs1iyo11bfM2HH56AMYQUg23Tmmq8CxkuXORa5CaAHsDpgU
1WWPFOad1DFHb0LBE42H5ZeIHTNdxrP/F7DhOQRAJ1BstjOt88b7vmR5I1ysTeN/qvkoQw0RK57y
oafoBbumAUYlXq5P/j2rw9tNhOyKSQwlmH1SLWBrVuwm7TjH2xLpNvFV36cBho8PPIiqVEjkX7OD
FLrN0wkpfnI4h2BTOImwaq8LY2xU5F4lg5ootYTossoQKNlNkk1D/i/WDkSRQsNhidRDqnHVqsyZ
+NitCys68tng62J0fjxqxE+h6I74u2eh5xIk6SZFUv2Ffv8HhPjEHZE/oW2z5C5f4UbFTQtgsONB
FNMI7txrtBjJ9Thrn/pBWSL4W1E9eJygrrVE7pNCFSYnVUzbVutFS0mYQA9R1X75P2R3ca2MDJgc
QX/wAtPweKfzjJ7yXbJGLs0S73S1+JCuCGCoxrvkdebc9qCp4XZ9rNCELGXB5nY/637XycBi2VYQ
aJtOGqke1U+oV3J1pFCea6+74EEKEPs/CIIacPnHIJ5BLbSD9O6+2DLFlj38NGu1mKLCqlQjOL5T
VkHmNA915yYBHULcY9FKU6s0eO+ivJl6VP3iSmMicyWhqFuqntUN7XAvNQHEXIn69oPbsELDxDD3
HGaaWaP0dvsx4Tt13IiG2zqkDB0vQlIZ3TZEfuugd7dDFBFdphhyuPCG0j5oaCAdveWM5ZUw4FmC
2093z6h6k4Mn32BR1F5PuoaXcTHEYgOaDeHCiG46Ckw1ELVN9KXSdAivlxLJYwpnja2IS8DYgbK2
uih+cUwxenzMsbjr44Vdg4z+oxT2bpxM+JGd6szu3i8qccsFDqLXoX8rpbG0Ysmc+OiQ6z/1cd0B
5Gy689sm2/knPQNPf5Ijn+uf7JNU7vIc+Mczr7CZfT1m8Su1LtScCM8n6mdN2qJr59cLOgXF0G4e
S6KskM+H6ZOLVC90BpU0eFJsiGRrNleDX+CrbzfWCNjIUoswRixUl3gRXFg2fr7aTcL1Jh566Tso
qOlmjx84uw4NQ9YUKed3DS9PyChY5qynmScWdX/UxuBJ1J1mx0+0L8x6uc04iVc0RE+RS+402oSA
5Y5YF2MfZx1peYFCzhbwQaBGjowD6ghzQpjCAyKD8mzGXnH1whIwXKDEhLG9WGcSel27dLOQZJdi
UFn93AkdiBAWQ9qO5ryb0hd2XmzCvy0Xx/U6fr2NVZiGYo1F8y/I5uB1EljBOFk+Ae5D84+vEQ1Q
xMwtNqBk6NKSNM9rdRuW1hhreH1hUahM/SIHE/ZqyJy7mnmBC2pcbuIm+T4sT9ZGTU8pYNZ/IPNG
5k9BP6Zx70725SAgV20nCjbPDr4tsT1jHMCYOEXCyMBJuOm2aZiy2uzKIQo0lwgONh4b2pqyPU2T
6WNBl5l4l6G76B4vXZ3Cd8/BISUd+Mx6v4ggHZWziHMAr7DVsWWXPZNLJxfvBYtVdSWKwvVzoGyi
lQKWwuhaTNNk8dOw6SG+b7kSOHRuKYcL8ZUmaFqP0E8H+1PaSziaNrxU4azIP3eY5drYjeOLhdtI
6XhmvLMSqaWwRbL0v0i1TFdS+IxP45crk385FX6FNu79Tl18V3bNj/R6TnNax3YWGhONUwNeCcEC
+AJm9T/1bbdWZTZ4ujmv/i+LD/3fse1I2hE+9Sz3PqKU9bZLSIZa3OR5pWZbZvhms82+vumP3vOS
fqgDKRUbTpsWsELnKEgiOT3Q7/jyZ2mhNclmekCFfBsG92x+IbI8dNiCMrIkJMSeoHr/dKjO6KcD
souVow/QitwnNMwrXFDfQALIEEn8Jyde8NyFSPLVP9zNZcQOcuKIeIf8sqmY8r/PirrPeCjnTheD
X6lO1KxKQGtTzIa2JYrhyQKMnY4vHQaECpSGB5KwmKmqPmfPaQFM+RnhTADE2GFO3u71RPQK3/wK
hnC5cIru3lzFeUUFbRzUqpJYrrzpqp6wyzYU9hQ3iI7iU1f2QBcD4oQzLi+N+O90hRuISjte5bli
Zn1tQUsmlf6hAjbM2KN5nDEfDyEEwvZLZievAVkEVAMV7apBtm7ZWCjgcNk3KCTX5Xy61LM2JjKj
OFezho6iGzqtDo5DPdIxOysrbFUhLaIbTiTtR+akjhUL12ix/gXJ21LAkegqImApbpyoPwKRP8+8
t+71Qk0ulm6I61scf+AQcIrHkWjiBdEkkN28B5+FAYsJ3q8Pe7eVl5snT0tLw9KHXvirJPptaI78
3ycuLAucQMMIHCsbB7IkT269y+L5Bkz7UdBi5AgCN/n+ZD7hTZK8zEwJa4IPyBk2cGVNGjp51PFx
8gUpcr8U/oejJDwOe6eY0IewQ/0Gcswhf0aH23a0UEtJYRGed7qWXOqkOuTl4S/+Ylz7H2nOJD9E
yPDZqQObh+nFyjgTG9q5yr2FPKXNqxnD78YTzptzsWzjvlz0r6KjPZmGr1ZKKkRa44v5AJly527X
6/oBCgWx13oAX5fbAnc+IfHMEq2znCOqqvUA4Y8bpKxXQ0mU3YpFbptnvH/x+EdE+zjAmZmg4sJV
7vV6B3zTzu/4gp/bW7fRldgGWhFUSYZ/tWANBS4ByVIZP95c9ovubqQRl2LoMtXcuT/8jksySmTI
TwpGtUpfjjqjSY9N65HePHsIh0f3VJNm6If4n2ET/vD2s733xutZpPSefKWjwB4xc2na5Xhv+J9o
gCkY3oiwYdvUaWLr/s19NC1ePqjw0LhnuUr2jvqoExxSqwF7zgQAROS39UcheROG+s3E9fnIfv8u
UPpT/K6QWcJZTqEFlRfiHW3XQShQE/tw/seJNJ6nnzmBHVoH3HIAhGqiXhCGplzdsrhvkhnCZAbu
70+BeeVrKnne/Xy74eWsqdjEdGrsCs7X4sJqA4roPLl7OnHRe3rKlMUs8LEhzsvJMAADsC0OGzph
EbF3/IKd4xGQCRD7M9RAoEuAqPUhvcL6uYhKrkqiW0CtHZhGkBAsP1OIcAD6vup93LQbvv2LkUc1
UuKuhtvZTBN9l1bGzL8rkBFmK1ZksDerBBtvVGtFmqmETjvu7fesVg0+bLuBbNy2nVhF1tZi0teo
4DLTy7fl1RMJiSdnNW5hYvDuRbWM2ZLTbfEK1F+xBU7sOazmJVdy+trht6DGGG5a+c1qs5j45r+U
sfP8ZKwYhTr2T6SC95oG9IGkXp0Ut7Jvi0oTf6fG6DS05Ek5kDcxcP6Ld3yTFJ9niCYi4h8p5Sr1
IZKY+06l13zXVPiD0xjY+hRgh3IqKM/8E7HKtAlcxBzAoxb/8waz7VbkSZYVepiN0IkXkcNUbj+c
5hhSurvrLzEop0lYNiFn5O4M/kehDr98z8kuk3O6/oH3Iy2sYNStXgkMEa7pZGqaXIcJ/t2KsiF9
p+H/0Z9+1DxAPXNL6dIAKpLZnNTdK2m8E7P9Hs6zpzAJIpSIxSun7yfzJVh264QC4ViXT1gXKqWs
uSUKKCQcKd0Av1PB2vBORkPOu0d6rOKEJDtjLcivDfNwKWGxWrFZb4TmCa1AbxDmbgnh4R1WEIhn
cwMh4TGax9eXgwqeRxr2t+GNsSvkKmSd7M2CB1ymbC5hYWz/DfY6bk2ZUBAdkGRqoz8pwRi9zfdy
AUoCNGGwSLkChXgrZZrsz1dEOzXi4yGMZRrhLMgk+6/d1wiBH1mOytfBtfXPW2v441gCHcbvipYe
mNEhbo89StP92XOimJMb3HyKpS3f7Dwjroxm5GVfE7wHWXL4WSRUoMeppz4FfAmC0hy/YCQGblSs
cVaG+9TkobT9BIQsv3OREHSVFOHZAjEFlA9hIHqLB71wf2cWc3zvVA4pjvhQuoW1MvV/Ic75IsiH
LpGf4+XadT30zQUIcvwsHfa3mkbKGQtQOr/QSfOA+VY1UhvY0UsJHJJuz4BpNGf0Eab6fJCIjnpH
M/F3uaNnDWPRlBUaLjzz+4s7z/pjkHhWrWxm8YTc8PSnYAZ8ZAgra20PJUNb9MZ1uQhE8/7AeFwD
tR9OBkP/ve8DoDcddO5zQ5I24wpMCxIaUULcI8lbtXN0tzsaTqzRdLA5W5Vg5I7rec0q7lvF3q87
Msb0tXPEH/vEy8Ak5Ht07Sl70rFrE5MIP9RpxqVIIeOnAD/13QvkPJuwyDIziNeQu+CEZFXnNajW
pBMgSO/FPEtPT/KKdLrx6IkbV3xeEpwp/evlrOHmyCK7B48yrIa/R9x/BECduHWlLZU9Fv3IZyQS
mnzXypwrNWRFJTjPWvmr/HVN3h1veVe9q1yoe35jO0FoLA3MLE9B+fVlOOnsFCAVEz2EPiu6Tij6
2twM1/heNeaGqXv71OKyvixTBj5X1mZiNq0SJ/84r61C6o6UEB1q4jxL78X0exdtzwFJozEVAeX5
ihfyJttDboGmVOK5J+H6JRjJC0DbQH9onQ4pldDYZErtIZyuh0hL+2gvOgruUVamUwOD7tLLPywr
iN28YuXwcnKzkQaYmEobzDBp0kCj79hlZY9L5MWP4m0IoHFi9rUu4qwh1CCMUjfMLQLd+2eHAUDe
DxNJjopnwXmvfZUDT7vYLZO+VybZPkX1oRhwUpexLmVnorLIx/smqytG0Ax7Id0FSiYrJC7l33eR
LBDYEcfOeA3DlYVNHvAOhKIFqSIjM0pE4T+sbeLNzIV1+BpeRtb5pM5ZoV33yBP3GfmJrcwS9PFi
FqwtnZZlJlG3MqkSCanhWogA7UN++ffC9+/ymxLuUsL2Ba/6ooXQnyEFDC4b0MJ035xgmYtXF3k3
4i1nbRTXfdOb5U38sSR7fDiNvftFrKRCOV+DMXcpUYcsoJuDsS9gsn2VA5u2RuDcsm8fevslqR5O
1ukuuGIqPWVYbPmNUfpqrjQiZN4KIQdB2t39sNH2eAlZ3shZLU5JlAc26tkvr4BTOm9km3UoTLdd
PsIkc1ZtdL1jpydXo4DjW13hZ+HqtqjYnHohS55npFmMgypYL4Np7Ap9v2bk1RnBfD+1Yj0LVc65
ScHWHnwPQzNIFpzS0gyqGNdE31ANILD78DF7YOFDQt+U+ZMuRkjimebRi/fwNMuQUUmLYvk08i++
48UV1ty5GDV957b47sXTkMx0hg20pcryQ4K0luVp9wONSMa3rHB6rxurxWUDLrutNgYvhoMIAamO
zLfGpZMpJHMnmBOrGG19KqEzDX+/8l01dVCHROlBXMLUtJvKRboW9wjPkdecsyqVBznw5UkEQnC4
Ot6kMGdo0I10Wws8D0MrPUtkMrNeEWfwysrxq9K27yYQl+Nd1Q3CmGvKSDhW33dif9ZfpRV2jx1r
mzfgRQNe9kHqOzKRbjiw1Nk4+rVeD656oBPm+Zne0LdGtIhjW1VpkkgJ1pM8sPeoL70MF/VrU3r3
tgb5aZl5KemOXOCdbIB1qgvoX0sRDEy7yyKrJvkprf7IqmqPpBcUt7BJOlcdacjhVEH8MB5yWrf4
LVJjWCvoTK/vPy3X7pJiSFiplZXxqmyavEsfrANxQuMLWREcCyXNoTPOhjXHpcViHyXGZ3xdqm4B
yjaIBUktdpQjO2nvKDS+m1IA2qgjd9+o4tE6mpMRwvfPbGtPAlOdbYzK5qbWQNcd0wEwb0RvHBlJ
GABBfiLqMMsq1LTVD+TumGWE0jb+a2XhoND+2+aBeMwvg6LPLXKbLcZgO41YM0N6RdJg/H88jKe9
mWro8drePrV9I2/rxya6+aSjUXkyeow/TEFk0ZlfhZCKK1t0JdIoxPTZeUY8nz05dWzIW193Ml5f
g3h/1NcuuMXWiNL0dGKLLbIpl3ZUNEMz4KdPbg9XS7EPT/ckw4OS7jqS5QVhGHLvowLvKuIps2Kh
qpNwsJZB4p6/1xtX+CnQVLu0qCCvTrWQIFAZU0jWdfSxrEYy1rrA230ZNPvGvnPJ+FDXSb/JurIh
QVSgiiKEELGL2cjCFsmh2k/uQLNE4n5itLEnboFyrlNNYdvZsOhuqdSBFV1eoZmtqElARqsLDPeV
xq6PfeCmjfQzEqQ2j9jsQoZRBt5RcSGVL5f/+usFjje4xtMc1VF4KbaeLtZ9Hgy++U3ApXXZG+4Z
M1BA9ZaF4ii7eVS+XDdnx9lICApI7RpKKrPcDh+M9qIksCrsEJuDOLnRXEWYlokVWH/IKBpCK9lh
LdfITKC727IfrbeLv0/H6K8H5ibPdvOMohrBaT+ybS+pGpdoRA5oM35/JZHeLTt9frNTW4ZA/2VE
65QMCoyfenpmpt6I/w+Fk6hR0MQpndhR7LyNn+YsFT6wXHvvjfAUADmJNZ3sC4IwDVlfc+TfmWGB
92CcEGBH+YJrQnPf2UOZ2Q+AcSH8X/TPF2pgT0aKeJDnXIHzegWuslIBTZ0nU0h05KuC/SPukMQM
U3wVD+lioHcHDDgDO/Ei5EVHkDSDV7dHL5un5wAyKqCtNIJTAdJ7lDagfPp2MiM8WOzZhAJkOvbN
j+PM60BX4uUl6YeiUTUs9aZ3IXzstgEoPTiuYfcEg8KARcrm9smcQy5ftebiPQPoR3LgdSQHM6Vz
zQg2bLYyk9lFmCg25JhKW6ZW50QFbKEErZdCRLc2pqniBvv5mJsyC5cL8FQqB6KdkQ8VS7Xqoe+n
Zeu0yYXL6kJ5LB2d07HEJQ5fOIFZGG4x/MWbUrT/eS+duQ8ESGbm2hIsqVg1637bKnGpD3lBV1lB
thh5a+EsWflPP2MdE/ZpEQ8ParOhXVR9OONf93IQXEfJ3PG3f8YTZpcspHk8vd37XFt/qJ30uFg/
eda9EhEJIyjc3d/6lH5GoF4DTsVub0XubZUDUEw5yWCdhgTONvmlsEJuyssOhN9tMyjs7F21fsIn
YdJqVGNuTkT8RRyWvKE9pUSGkpjME4yPSF04DugRNFqMBumKbesflm2bvpyK/3L7aa1WzBpHa0yG
+dY8WL5KIsweNktE8VWwh4JonxL2hYcP59Ubqph9ackjryCoRB31c6orMif7cvGuEVGebWenAMzS
xXGRiz2ClVb/uf+mqXnXs0hY9VGIxb4bN06teo02b2UuhMERe2K1/kKm2Tdw4/cR6oRjrHF6hwFB
H9taDNjb3rFwjBoOIz+tgkRLTLzazG2IZ90jOCmp1SbMKZ+OQwDDbNCyu/5UBSuZKdUe22Bsz3q1
i2EPz69q4bZMedCVnsvuxFe4nmYec8tjy06FQwTRNUla994ohpbIAjSrVcxS4Y+ABK8Jq4hqUpRy
YTrQxrATxkZIae3ajc+pd4EE+FS7hLZji0x0nh1DS6pE4h7HBV/tw75UNjrJxAmqyBxGK2G3L40N
kXS6jGQHtOW7rdC69ibvuXoA+w0/f6oQgbXGsppf7O2Rk+VsK5s/ixTZWO+9yLZjDxRX+k3L6/yl
wkBBQyrOlcXEbllzcroyhcOeLpB7BKXm62Fax7sppSF60lDYCDn2JdcB5iRYC6yNs5y6Jt7LDs6u
xW/Iy5ggfbSauGzzYAJ9dGySAkAPXayqMi2u4lXZk8BDMddhelZvMFqKhEWTCwXP56MbWYLwlpYw
43qICzP7v0Hv9MEdakihucc0bZRIi/Uxf74+4P5pjm8yOaNui8OXYMuRUx2kUdSY619baVGdh8UT
SYlOOoh2dHtzCxuMRVCAHTTqbk37+75qQJeQaUuRcMAThsmFjVVEYgvzS+dls2d77fF8ML3vEJJs
nP0QwmzYaNG4o98rjHyRmgw4ScW9zh0kO7+bP0UmiqpV6NBTEI0QiD6FtmDH32c9xL5aycHb0bML
dL2uvuFwYPjD04yPazv+k7zyGIQbl7zFkSoyKHL8oS3ILr6y6XXHqNhjVk5ddzc4eCTjPKC95Ax0
p+CYvlvmW/btou/K3tTNrU+pFn+OwoYKgaxF2xyiBAamM1IJmoOgAA28LqKOI/NYB8qYknNkUR5s
xCqq7AqkMIabVHokh0XM7iZlo5ZAOfjKS2PPA1dLVoWMjJnQGOupin+ywPTyZ5y5ERpF6mfxGMKS
cuQviLDrF3yp3HEyfW+ZU58BmwWOgZ6mYELuWOabIlJmD1DWfDYI54bOaXDsOoXSVHEaxknYIG/i
pBr69XHbuSFitLMEKA78m1HlEczCLu+g9/G4LVCtRS2som74nRq1DLk3iV+8dSH7Rxegame4eHXB
ofGGqhAZme64JdRtwlQuapNu9nLRlgmtlzYBJ1l1MXfbMVda4LNrxr5CGutzYIovCErWrJEk4M4h
nJzMRLxlXx6fuhYBH+nRcUnCcj3vkuIddZiRbngo0TlWITiZ2VkY4pB4xbPD4lzxBWxZvkboWxWK
Q8+CD5YcFo6aRzSjiQAhMOO3kDFtcp/yPkUF2Q/NtdmlNBc2IZfkt2DDYTIRnY/8jmIPI7vpwYpF
HFxpH5z6XVkhKtO2FlCEJFZE9/y43B+tj1cmv2SkBDOoOigVTGqLoiQ87hjND7ggaAyKaOOtHLNr
JViDXdIZ7eRDdXqAEDkKputchWouLfnIOeOUOwWZ2xClnPqzEkW2bAhU1RjyKBPOg1p/dPMU/jkx
iqvijyE/KSBQ3Hys1cPgpTENM717MzBmUuPVDi/mculjedI9JxDjVyBHrybx/19ne5/kTpCS3PrF
AHuzdmjMVKtdbNTLe4pGQ/xXA7eLlzRjHNzXlZwiBCOrIJkQiHwL3tHMZbI4M0Xr5RsJM+Qoqbsz
o+XhW0mY4Y8KdkALWtztYZQ2+jZM2FvIgxDILNw+5gM8XgLQJCLE4FgtbWEnUB9lwGv7k7Ghr3YG
oXr/yp2o5j+N5zOFiZAGW/X15tjNQXnpy5g1WUaCPeXyR64rx8APK3DwXt7jxurgGRk7cq3NbfRN
ZKX2hZNVirdREb8+rYuyATiIaaBH3F0j+TtYUjkPqCQqkHC8BCFXFSdL5qladYNZ7Cb4LdjnW8en
QFp9zTrzUCHoQ7SSIPf4KRbnXfXdTfp2FyVod95kgAEobpxA8dSRKCeIXnqmrFLpOsFPey8lxPhG
6N4qIwnQjqQK/VA2m/ajq9lVQBPIrAtjOyuKrLa8tVvmZAiam5BGOUam6P7aRcpS3CAkW4IXGR8d
heBAW5egPw4amZZqBxxkpj1WTENYljjYcGFb941xFPGcCvLa/HpqTHTivc9aVdIC7kdyXm3YG1/m
0JgDp66RVOilQS3GNFe5NWMuM5tJo3Un2la87UMVlEdycYVmrVOCoBXitOyuKSJ6pk7L6Q03DYEk
0rcv836tbCB3M/GU0ZEyFOPcrEu8cGSth156t2wWZwNyQczb44z5sV/joLqGgFjiYPDZVVUkG10J
OAzW79dhNBOrKW1vQkhEirQvL1IIKDZdLeRmZgssZXBvR9iK+g+qUJu4uBr0nZL6AgEy6NQ+ujCQ
eAA9/QD7JYzEBsF3/HR8TUYZqEqJzHQD3gGpL6so6+At+LwgtcdLEOEIfthKw0mEgtSva6bMif7H
kl02mv1bT4D3ZN9ZbV+nfTDgnX/64bV6FU7KzScVwTH1erGrVW9MNG/K6G4aVCx3x74rORYa77jN
qirxBTwt8+nxkQ9iVlY0sz0EnTBzoWlVhAyLMdLY7piOVvexbOguzK0wk8vOENA6T1vtqQLK/fgk
ji9KoGfbrPN+OXB2G64ruIIv1fxIgl5zzxuhpnuIE7vX6edX1dcZsu+P21vbzKuIgpFleXQgAbkC
j5R/pS/LS1dpeFTPvre/pOYgyf+5R/1+7tcBmYx1/ireCebcyqoHIrYsEwmD+Jna30ky4MmEtvH+
icaUmBqFnM7LpKK9r7htxcrnkUIz+jTROFZXaZRuHQ5cqF8yDRqwYdmhfnJv6EHQTLI7six4fBp5
g0Fla66kPW4wsuFlZ/ahuRnD26eZZic6fg3zt8i6vlPDk1fqoVZ5KBX3eXEu/SlLYnvEDAzCIXQM
mg+upPkZhpA7eVSCxhDatlNELiCwt8tkfaAuuSZ48fm0xOLtb/gLzdQusLzHQpx3IbgbQVDw60it
qXocEM6QNaWGHmMDA6DcO8mh/yCFFN3fsbKdlMIBi9xdTiSngpk8ObwyMRk77hkBfeh0WyX5wBTr
bEz4RygJdsDPhJth6n6DxTjKEehmEgsFYgyotmevQnEIVDilIzTswqsmfzCk0ozMAt3bwBu4Wayn
+nTB2HEz0B71EW6mSnf4u2fusuijXfvlyFy7sPgCuXnuFgpA5gjRHtylohgnbavX/5n2QEJWFXPA
E1DvKBtCrpM8uyEVPMLc+8NBi7nLxA+uLKYHzb7PnxX5gM0X33IVIB4wznMP38vEW4wAN2KLIOP4
+su0iArQM98E6qkdDfBe7OQXSXnb0FIHlLxr5oJDNrrZu2FXGTVVqcfB23Mr11+24lzEoDPa/3Ru
d03l+aTM8fGCl1Kn6nurszuQMYMycYJub+jooUus0JI0WIwvj/X+uCeUanGSTASUB8UsMEu3ad5r
ThjS0JzQXvZ0Yue/P3Wt3vHfAidZSv3Ayl+eFYLnbiX5BGp32bGjvJ2rdnz468Vlq8WUy3CNqVfe
6prLvAY2cLxOlep9IAAPkvm5h5+mAR42ZUhxXnmj8FSe/oOGePJ8S34YVDzNO2GGI/uXT8tPRAfs
MH7yU2RcoX20y7BI7ATwpYE2CuSI9WM5PoUvt9MSReE4DaLhs822tb0Th2tlpl6dfWklv+vT7RTk
V9gwkGD2bNIGJG4MNAbRJSVZOmMnC64GtDAyCPrMszU/1NoJ6Mrh6eIlFMP6mtSr4bG4b6zRbky8
YIu8TxYWJ23iiRMDvgWjwRzTYG52QMLfWwYLnexqT0VibPEQUDQDn7b8jh6tTevCfSQhR0sTdMbR
8k3+4Y1lUnRfQ4b7zF7vPB6fNMmkASlRdQMuba1kZe19IASO5stn2t72N5ESEHuWXpecZtec7Nb3
3ADhZ1dEpnJfkBchZqLC0+4E3UMtIM6NyB/NyvwRihRs5MdhWa51BSGZFWHYJ20iVvhci+WrIJOh
WZUyhnF8aPiNclfRtQVF8DeYxemcLExrJy/5dv0/TfTJrh7FqTMcwiWySJJChq00pnUK5tZ5rzK4
2xL8KgONY5k+wv06gjGXPaoZqZC+TuNyw9xj2dx9JFcKa9Z4O0moL9kZc9bsmhmYzSGm358SRLI2
ihgUP/BYqNxsLnWkdnoK0qEe9AyTx6hHmkGWmhIQ3jlnNCbqmuTkTkdL5jBHztEt8VHpL/QHE9Ww
VSLeZDaAO+sYaBWdVOTs/14uc34b82+kxrq91PYihXQOFHxmx2X9MxT5Jn4MhEJtFWpRWJt08H0v
n9xvo5zaD+K300EWTXSlrMudrnl2YdqFdNCGalDczwg1qzA3SzzEe34c7povq3XRfax5ALKfyIS2
alNMHOhs9ryzV7GTGuW1xhExk51BTJpQbNZF0sVvhrLVzjiBCe3Q5GVn3lOXLgsTs3wg5G++m4mC
CDlO6qLjjC3t66XiFvRSdiexKqOttiAUuKv1oo6pcLLq8p3L8XycrLe1ohDRpV1C0DyF2MGBcOgc
dEL1NP29501KtoOf/aMdWM5LWlJYVLYnTKDArLWdHKLudssoZLtM6AUbg2TEAyf2l86r9xALztEK
miaVAH9UhvzYqNQf6lz3OF+WylkZCUibn6h8Bp8IoLh6KVqMDU/vzaGRVIEMNaYe9exPZuaRmqTl
Q0TIbm5II8QnjdtoalQUmhKQ2y2T2gqmcswikFr1gBYNnAMFts5YgYNP9/D+hh/4vVAenupiJG/+
UanVbV3/0h2j/9tqx4WG38twuC+EB1twD9RZ4feTfZk49mZT2AM0qsnlynan5LHT0avK8Lx7nWZh
LG0rC5zNkzv56J4W8OyCISUUWXjI+ywdp3a8cGgwZIeEcYbwlQ/cFnWqDypBVjomGbf/8KmwBlYV
46+YyJCL5Mhz7AT7HrwGcUAx9pQ1pCLCODTbZHkfLFHJeoY/eWgMce2OQxxs2QhUCYD55Cb/yYGN
PHMInWNpRXu6duh+gHqy2ispaXr5D3VwbgDHNwBslYDjYCMY/9u4MhbTvCtJTp1DiZM8MhXoT2Ok
bh9d0pnWLOXfu9JlhmQHrW0yMyeny1tPbBgz/YgsXZftp0wnuvC/Pj3qLSRr7qxXPFWtCAJAwiMG
qXBb0xqVYlcALbeI8Msz3HKIxYIQV6bQrlnFbUqSnQaF+jsmpChC6xjmXnJELIyU0ECEuPgakFEj
XAG60bCMI1UGZUf7P9SJmqtArSQXmfTrnHg8qYvGakPKd6TboNhlCnPWLXmrtCIe4nHOSFYUYK5r
YDD25O/+Ns4zqPC4uL8rf5ZfmDU8Pwsvtxj7rj7lXFCzM+4CTATGpJTL83wXikvrH6PIi27efdD6
un231e92ScpgWAvZsD7YsokZmABWdEVEy/WbVmGIZrCm9nDdWDbLudmalX6NI5y2q1WnpxYjcMpR
N6DJmrtI75p2Ush/bgkD4f+6SktQEkAHk/r/IFajAXF0qkcokR8qLdEoOU9F0YzP1yaVLI2/LvOe
JP4XwKYY/alobbZoskaBcWY+L4StpczvRQ2hwg1yDQitYZpBh/WyL3M67y8JIPWmCT0CpK276/zE
iIzUGdGYgaUGj/pp4S6UkAYH7NjEns5koEW7m4w6fw20Ydfia0fxsRF+/nVGmOwKPobHfqw/g3GE
P9hNkqFZru6S0gSYx1avb3E4m2z6GMHhlHzjm6otOl6EnsQOWj2T7gCCd9o0PViqxBx0dwNsb1sc
2wKOVUQ74qcE/IkheTM/8ffsF9vA3aljLiFYgReyaDuxHKMyJ95CCFJO/y9IDNc4253GpHsubtPw
7Zn9dA5boT0YIM9SjJCGhd09F5wzgLqmApzVcQd8ZpjxqWcSqmy/NwHbn67VpVgiQdVEpLt7r827
y9DEAOwi5NNUttEh85JoRUmhTQBB8webbdmCcK34TVaQBRe13PJTcesYtSfZxTcZr5wo8mi9Qh3w
o/FF1XMXVoCx2j2EnvDFSjP9nmmBdGczmRIvzwfyEQNe6xoqX5p4aAaan1EqUcmCVq7o3LgpuvoL
BhV6hUpfxk29dOQ+WCFEaeujW4OUmR5zM+nZxaBzurqeJLv02AE9OwXYrQKidZbwlS9XylO4kZj8
FVqJqyfOrlXjdq1trMrX0887c54XL9L+/SvTSKxl7FR3Lq31fEyBUd7yUPcSMotEePwP0Wqr7+Iq
63jt71/StgCoDm9MHtWcrDHOMKVIGQRXh1eSCMzDxXXcaLXVDfoxpJX78A/ytbeCi9yprb1X4vVD
JPMIoS6IBAYne50sxmv8M9vU0wj2C+vdLzBI6ylOwM71KOyfqhE1FVUfx+wzsqXmy7Lwg8Hy3saC
1NM8emxFXo+3mAlS78JyThNSyoBUcNi1qt6l3kVUd+26DtehNiiUAtmnPruMqVYQSbzmDqv/zMm5
xi5zEV8ZDFWSMnYh/ZVLjRG3qQsaS22F1SVOaXvWY0WfvurXIouauFsE+XxfWGzIYzcv7LdN7gq2
Z5msftIcnyGBROhUgvoM7X1M6cExwo6UzoJzcNmOQn1g1BIxJcIVtex5TUQNmyX7vv9yyrCzA5Uv
014/03Lj5PzIdtPzGK/xsr7Ns86BvKXu0hl2m+kxq44RdrBeFITe4JebIfF0roc0nmkVieE4XKQ/
x4ZgJeMD5sr8W+7JjlZkLJ7q0io0dDvTz6s+PI6T5Rc4ajOaOEbwEy/r5ZYv0eJIeGMsQhdte0O1
oQyb94vM7EGsx10mamVIdJhG0G/oN1IJ3Gb5C1T/p1pcdQwV3/3TJVZbju8c6qfJDFjELKzO/OOt
xEaSBBlj3A98evIW3nYzToN3B6lsqhg0pE7jmLhqpbVDBvrB7uW4xfXyrnPS+ozj9yjmwaJaY1Fj
dzi7m4Gfz4hiURWYuBOIBHfFtXTBvKmWRSbdldWzsXy2GCyHkRDgr7YfcaY6u4dh5mPeOsL14o6H
x2QJ4BrOVN+2W/zAuAiZItC86Sw60JnVKo4lGSd0xrpHLfdYbrda5ugvRagzQHpox7gOtr/L824D
Xvjd5I5k5T8NulZP1GW0aJiLdMR/GUgW4xJh8QimZQ7jo/UTnrzky14P7WRBkwS64DgpLrBRh8qb
vmgXn+GOGDypx0choDod3UH+EsIvk/Sy9Tv5cTw583OAxFf7KfjxA/u+P6TdBddpTtmsLmTbfOOI
5Dcw7NiXveuJM8y4c9S7ag0W9sunLbVyh2TeWZNoGr3MFGfDHpiCQqoXqgjTZofnm4DyFKCoUtGC
xxes71IDPSqJ87Jc0eETdd6SIO3sikUq4ZE7gdMwYOp+LAg/JrNMA38jfjMEkQ5GNPunPlUpXi/T
wcdeBK8VTbQqDh+tja3vNKp6/tdAcU79zFesMjAZv51Exx+3zJzOqChk7JBlzu70pZnYLETPnxCC
w6OTYm2Fyvk7u8Kfxqnn/3zuZUfBdjgC/qHWxbUYRWpLci10Tk4zbUJ2Bz0eVqTlpCEXJNUSDKu4
4D29jdHNyN0NAevNX7YC9jtjysG3t4rbYXdStyOeCdJDBf9Q8Iu4jWf9En9hyJshqAmX5Z+52si2
wlY0c8CLv1/2492tfiqds/dAsvtCN2B2hRzpR59g6KSRUHvCQKC4vO6HBM+8Vd9CyPmxwOwShkGE
gbx7lAkCl7y6tQdBFZ+roktsTXYxx4lTRCnAIbiDvB8hDJpklqaePtMdhCPF4uG9sVlR0xir5E7p
eFifQreh7EqghrLVF6CNWbHc5s5qEoX627/7q9dVltAz448Nh6c1hcIyF3bgSCL5YSp5VRkGGBiy
ag7zTyKTD1Gp+yOa5Ymc5KaR+eVJDQytqVL/BFg3fTKgk5vcqryAvg3NwAiEgS1tsEafQ8BXUm1v
3Wan/GB0MoD8+oeU+8jG+bwCL62o6Xr8YsrqwfsDsCnjfj1RydwovpTvpI2aLGqKRDG5/33Nfuq/
McmR0DW4mld9QHUweiLE4CaCqyNr4O+Oh+rs073jxfPb2nUr4i5G2fDD3xxEX3sQ/u2jRHdItYaI
1PNSdmbBqz1seCzXF/EFa/32tri3B41TfJ6+avPvvjIYVsh+f2/7W/EOGx0n+d7s1iE/tUwZqnnW
q+DWLNAlwl5oekcjxb2HThiLVBka9wsKOwYBRCsr67LjbFKFu70DMHhEqFC+0mgFk3WhUqkafEv8
XRp4j6bJfsWhsiTjAkvXY2/2bu39U3ZPd8X551v/tyffPaG/+TbWT5jlDSB4NJrZInKt2R6vy0Rj
+Q4suQXz5Nq4YEOAVgnuTK5JDs1H5/gT1k+qx8rXkevBTWKBQIIJTCIJZZIkX9/m0KHIo3jXridM
ljxDCskvDpNTXNfBaOkuPU/l1hDK/ilkgDitppfIuvLYt/n58LFQgTfDuG8NX4FUmM5MBTam7MxM
TCpy1n2z+0cUxRPnCu+sE5J1m+KCXBrjaur9l+lZ0wMOq80z0Ve8r4SvW3LizfOi2Wcp7FiP7Oqe
7KbdtdQrbRyX96LZiwRPSIZUCZ0c3/iWFPUvxuWPXMf2CkMHGQ2H1HmjLt6u4KI2Rq0VzDkP6lzm
ITe2G1QZkFeqat2YF+LduI94EYdDzCwd52QRC1HXn//ZERFSiObIIFDY7ol9ZNHrz5813YLCaPf5
2a3n0XVYyvSXP1u14QMBpalpvNQVdJfWM+RJM3XJud3CNV5M9vqF3ifCjTpvCEiN52hNDfbgsJ8+
eg/eWdtxv6jUzcbwCfhjGTDjVmttLysQiHdkw9hcg4PwinQN+S36itLTDSv7vfKRSTvRkVs1N+/E
IBNVTtCkQLgwzlti7x1d2JTAbNlX+Mi3f0oUcylt3XRuu/oovfpaaNIXf3OhDYNRL24DDCCZtbWT
VXDs03o7Joc5ZAezKPzPNoocnmAhSYkckC5LPd3wYsG+HbjKHLLrsD3PLlTkhiAa/yXOQ3v0FDvB
ul5XIzGBFEDkfLoap+AV75uKQd/AK8+uaqlt75aq57lQ4F/Eaox1nucCq9C/JAExpJjEndZ+ha8r
sHwrcxy9JNhSulRKoTgP2VhVyL2XpkOzFC5gS8ZN7tCxrgh1M4d1aHlSip3y4/IhSm3Bduz3Y6k6
x/S9w9ZLKvfPpcCdsBqCiMvMb610z2BXM2WvHeiU+5Co6Ybhfsp0S4kmVhFxtotNM17fFOcMG569
Sdy3q70/x6M9VTOfiT50BLjmuYM4szZgi08CqUUYL/ZBHDgqow9OGJGoW4F9l1gSt6CU2O0UViHj
RdpFZtsA45fElEKZNzCvh38MsqqaT0ZRbi/hbf1JK6nfNmrccfKftivxt0eOOl4esM42y9BfU8t4
L4p/RvbJ7ixIy+TVVV+5K1jJqcDlDK++4UuX00pCRCRUaZgwdjtlpTD9oepctpZ5tpCND8o+k8+J
ALSjVG/MZWwl0gMqopSi2yMgiT1lXCHyJVk2hijh3E2kEBxzGwHAZpR2XYNi+/apGKp9GhDGlUN7
lsixU6TccoK2mhODgjuHemqJ36CfP8CPGJKjotdmuCiEHdC66ndT0jWaoyim+t/Tzu5nL/p/MBAa
MRzaLQZ09lxzeUJo6wj+ddPdpPpUQKNE/fEH3Pmfvxc/nlCfdOwuFUJDvT2uAZPxiUCAcs7NL2Gq
CZ58CTWOoiMr0q2DT7op9A1akIkz/2HzmuINxhfL1BoyJtUSPpWrtS/McyRI67XBUpf22fpgJE4E
Kr26CPoi/nlC+t319BWXqXw8t5wl0R09vnurWoemfuXQ8cJuDujGW7gzxxdMPfFcsyrG+Xa3W98P
TlPC4cl8pjR78HL6Jj+ScREPf0WlDwNJl/cGSc/NXznFRcUpnX4wa/54mkVMU/wVwxPpMy29xWni
xH6mw3eEWHsaM7TTG5eTv/wd5p9pKbqoq2X0xhVAEsnSiVTLe4vOk2e9TbISSb1WUHaBrKqUVT2X
Szv8LGP+Z8JnoOuzfa/+9NxuTBWI6ExL3LaM8d0qT7rEzi1AgvXPnh/tQmAM/QpkyXrdL+6hkIjH
DAKfQXHUo0QqPYVCVKYBk3U5iQQPZqF1VgPHnhkt1xG0h5JlmcD+Y5jMA+2s9fPKyUTQ8lTFSDoX
vfUWvNMAlmD7Bom/snrQx7XwoZrPk40BWblAU14O2F7Tuc1cEbfH3a6dvPc4VGGl/8HGWZCg7gWV
e4RGjIpOsgeq4Gj2QSGVNNbIB1QNbYeH0SWXLSUkOlk9dQnQggdHKObGRQOYGEI67qYzfMpZ2WDl
Qf7U16pFb6EALT2zeIBEVsb8cDeR1SxZDHGHg34dl9CoQvqVm8lmvCIVX3pR8iDrn289YhvEzJRO
yjSclI0NGOAIRvFAWJ57FMZScKjN/HAsVpz5xvVG2pFrRBBQUG2iaEOONoBYtem2OXiKlBCIxEEW
Yf83y6Qn0Aoi5WxldC421AdbleJf20Hth1E0XppYaVDQnm0jQXTtjeU1Kx/avdSxjpKv5ROToyih
xvxDtxbuD8aRxF+tanHnuaErYlszEBIvMZmNen8zY20CIPUkGtNAISEwXBXbfnoEkh7xlTURZ0Ok
CVReUbAKoGiaQdAtY8I4u2fwD12HXxogg7I2IukvSDod/wpvpf/wd5OjhRAmy+j8bwr+dTetEL/N
XOAtwWTLjIPNrWcPEnhI8qGnKDP7rCR77iktH/5aCf0R2Bu97+fRom+gz3NnGqsrhhlWzuXm75WM
3kB1icdQuw0YUZrV/dmsX0/xES55VvtxAqKoSueCMgIp9JlH+V4UHI1qIuH3UxHuiadAZNzSAPnS
57MdEZmiSMJCqvGFC1agxDeqdGPuvsjz2s6cHsQJcDFhToYp5mPOMa8Y5xpFVjjtGKW+3FDPQSFj
dl+A9kdXOeK3qNCb/HGI09Tgrm9rfB2jmb4Z4EsPPG01q+gIjVUTzRHlXRgnpisRZXSyeugAwWT+
I/7v3ZohXl86eG9ptY5WE8s31WksEdHj3MmUyyR+aHfP1ick/bIw3fUANYGsKhtFUy9xT5jxhrV1
+LHf6nHw8dD7W7oYKSsBaX9XL9fCzagTG1aAOyId5+w5BxNFGTKW1D1SkWpvVYVrb6c4+n3cIxkC
0WCwbUyvuoQHbGJ2pv/WDBak7yt5+PRwpcbi/K932p5Yc+OMGJZ6D045G6xM4LIK9y23RHRQu54x
PeCNg7onamCZMnMGse7ikfhNsmro33/Fg4e5rnMmofwaND0ic8V30Eu1mPFcohKqmHnB6OAfeTVW
q2oQZmDT35HWOaVIshNdLcqZDsbOEWue/twXbX3XcRWBrFWZAXFwrCfeYgBKrbtRaCQqAqFRWnnt
K3EKkXPfLzFUIKHGT8QQShHkGkqH3iRXYOX2HXNYwkKTRMH2Rf3Ug9FXMNxYPrjQB0Gww2yAfGxV
UUBVLL2f0LtgySl8E2KqHjVnL0tzGl05LyW45gG9rSnp4KTFxCodv5gyfwjxAzdvN+3c87CW/DYB
BqQToMzorFMmbvYM6zCBeiPnKC9u+ZEe29+ksFEtq8eRAa5KBL5YsyhDktTiLCMaPtemeypeByN+
mIXJB5cAvlwjXvdy9u9AeK0iHmjDYEbd5WlWSRECGW9zM4tRl/oWCSWYiba/s+SnRBpEBOqMIYzv
2OnN5JO6UNRfYjQWmepJH48T7OXbtNjkS5QGFGoqPjc2zIaI3QV7IbhWoJf8C1QbWbcOzTbwzxDf
NWN3u0IB3TFb8+DBspA7JbeErUq3aXt3G4+s8ChkHc87HKS22W9OHtfvMIK8GrhUFpIe6G1xoTVD
UQoAnVFUtMg2wg33M1O4DaHdRoWp1jxrlIJoNifm4Fv3cvwRVrlCCuKfidSwqBe0ZwDQkJ4Kz/ut
GKNahcr3L+TZCimvCcOnDCDCs+suwHhW7FbHwfMpcphx1LJMVnWuH6tUFwmieZGxxX0YvvzzF1Tz
wMTZyF7Oa0OOYhcf5lLgS6VoOek12VJCPTlIznWN/tuaBEWWZHxpMugpB7S6iHk50F1uwucz6DcR
hifa2+6JXbh5QEYLFkUmghtR8sXZ3x5OJe3X0jExYlnaMEtORz+Xa8BUgBKtR2ogClt1vrYm1egH
8btoKsnbiy+WbnDXPmeh/71jx11JOuOgzL2t1L8A5nZgD6bzy9DvvU91XYgJr2EaO43lm526Uj2V
tlk0yHYCvpniYlucfhcbCTmUAIZ+8/1rpsgzYQ9l+LcyENUvJa6kzKiAJAIVpWZwou+nDa+ZfMkN
ql9MyhH/U3EM77Io9+IZQgjmYjPgjjC8amhsNRZLC9FX9XrNuH+Z37Rw31n/KZYVejdL4ASx2xvb
mKhAdoJ3C8HjmxgqOBKsMaJaitgU7V1kZwt+grbg/pZ4RJaaUE3v472qGobl129EdwwBmYqye7Mc
AFg9ITnGusmc/HqaFvB6I15BK1y8IQLpZkjokfUhMKQAbeuA0e1llzZyAvWFpslN1qWYvQMXgRm+
WPFCuxdRYub0/6oKUU7QhIldVm/k5+h0PnePQnM48Jrc6QKSYPOSw5m0fLSd/yTlBxK+1ROkd3+M
523SYib+MgyJ2nUS4abifaGxwiCs/a6gQpdRXwZDqsUXX/qGL36mRn4phoY3ufOi8tAiDTf3D6XY
n7qAH+cCRKmru31PbAdb1MJAJdcP5Bzt5uTfXbqvjUm/6K7Ro3uHoxF4vMN5CVH3ZSUGI/8ssaBP
umUOqFnHhaSyO5SEZCeH7VIu8Q2cX49e4JsoZemZjnA3Z0AypeRS6xypmACq22KjjaiFHF31Jbm2
ZNpVVtovD0cYAMnI5LggTkv2ZrC1W6G8MBSLVRnrc64gNO5td5X9kobWWhHUF1vxxOzzPYIjMNRM
aQ1FPN8Yj9X7lQ1OBmUsjhHn2ez8a12yoi8BfAKs2rNz7o7tb3m8r+lmYNuiW1COKuCkS/ikmE70
dbj0psoWw6cEeFbDtIJdxFDzs4H0sqKev8GjyYAg4aN6lY0CDq0X1nsyNtYk4o4v0EhfIi0QfV3A
UBJV6UY8jJwlDMlp+wF2Bd9fELbo3G+G0/W+WkmEWF4IbZdEUvXAtadNANPoy2BB6x6e2EzELuYX
e+ZTKfE9cEa96gh01u9hsR1S3T5gGFrhJadmZLCPS+xgH26iUy0tOg+s4OK+YDEc4CPXwotC/Tsp
qL8TO04aQ5P1xpFwbx5GyX+L5Jm6wSMIcXGCdB436hQ5ZPI07PprtC1pMTJXeKMOOoIadcIqeu0g
m7PhATZauZIdEkx8Gv1omkbtTFhVX0XP1hoaYOxIDE6EcOxpystVZoTwhACcaHsnSrJVPgWxPsZw
9vYZ0hp5lTBeUdLXWZWMc4iCPSDGb1Y3Ar9+iVlMQIrqW9SnaG6HWvrl5uXd0O9uhZzlL9T5Sr3I
IpBT8457vxvf5L+egSWV4fLjUSuR2aVp/LWfHavoswbdyufb5XMUzZ3zdZBnfgkTK4eI3gLQCCLI
19VSqXQiyAj4GMEMzEMqvyLSICgMYnvTEGi+6EKI/qo8aD8aU+WzdX2C13gItIBG3FvXbBSFSg7h
W+4nmuPqLlBV8omy4N23E3ffWLFHexSK1qwyzYruGStrCcTT+RgiDUmcH53U+c2cWjnk9hkbYg6P
ZlS94G53pLdeXvsxbY67//Iq9ZghjOEujvK9DQ49pas8KAWT0nijsB2DpOuQetS78fLIJMT3N5wW
gCoTbNuxoeTmGCSAF/UyybGfcufnxfoMKt4MRYL1PCjbcf4DUdvYEw/B4wflhf9658qNciSn1OVK
XuctdLHj5WOAY5m0YDnYiBuYv29k1U/wB31MjwOOCkdY2NKNZ9tI7ECNS6l+4RCk/FrD2jWv7pRi
sZuJBT6CpWxoCGCe5DO0e+oREJ4mXvPdtp0EciNQLZhAFOhy1yqJvLgCEf9sF7p19zinETd9c4rB
1Nk+ve6wT26NlXwr/0sNmcRC99o3nrgkkGsamXOtPgjhAijN+QiNv7npR4i7fCDW1G1j1r16/F7K
dsMTmxhRNrm/R9CA5qNEgKdBEtXRtYq/O8es1gWqLP+4GRHKcsKxn/7ARKFddIZwm9xiVHuiYUIZ
EQnQQoUWU573RaTh3FpAgwUoVpItFaYtkLH5y8Ys+tbrtF63UkriyYR+pSymTJPM49a6VjSXazGI
JW2yeRl5NJtm3XN4qMnDiHLAPNKpXNjG6rK0+vxFHR+bcMEqdVafdul97vsLJdYaG4TqmXxW4Rh3
MshaBhmXI+cWxrG2uL9r1j56LOqs9bUxR0957aqDCy5+xNqenvWw2qBvAUC+jd0AiQsVGIurAAUd
n4wHAYbrwkvT1ixtaZKpmnrycfB+74RCfytdOzK6sHyHoUHbTt+hkei645ldrslIdjWv9CK7KKkc
XYQ25WYZro7X0F8iobfsVwW/TC+m7lA2ZjdkyZVHsvrKJRXOgE/yBatThXsGXdgPWJGmjnWuj6bO
JWZQ/U7raexmyY1+v8Y0AxLoi07rkNPkV1NTBu7H+gJnOfhP+AJUu8089rdI0WqNtI1RKMGcZ84w
A89mqsYMBiqrXyosePtcLZ0nl6MApuWtBCeszvJMrRX7whHoaozh8HwAa7OriI1rc37ezQIsCUlr
9sO1QC0CKZuRUYNPD1pJtfzFMzGRi3oi1eH1nk5RYfmnxww4yHWmP0fhj2zEtFUoybE+2VroiA3j
3fLhnWUDVRqeLwBBVTjdHrcy+p5jeNSMKAeFqj8cSnqI86v38MFS+9g9bYev0MOp3bi508Xl/Nza
TigoaW9b32Wy+Ca9q9qeCXir72cBeUbN6/Ts1Ogep0qtUd/ztIViIHkE5XfOzs0fd9Mf7evW1ByT
9H0UJvFBWORBlrXBiKvEZ2ix+DxY/SLhTna40br0fHOhaqLwFidZxztuucRVUcgOm0yL+5ddr+f2
a1RlnmVDTIl1SQQfOmgTBw8lhoGrXbcj7Cd2qpUvNAFRg0CMTA1tZxNaOEeqbjScDkdrk2BO40Lh
282GXqaabAysUL3SbyniUcOs4+N1E21Gh0RD66Yc1h5yDZQmgK2rwBgCSE9jT9MV6njXd3AkWz6t
pawq/96ZRxBRZgIF2yX1k4WLP68pfrDadK+goYKywLntM8hr21aJhFM6hdFSwbPncww1VwntP6mm
Tu5BvQ5BbRbx6LbUaTdJIVMXB6+kQEhJAu6/JqwlWVCe0m/bEa2hn3x8pMQ4X9NxuEbJ17W5cehm
mx2+dkCdgW3901G9qbywk81I4kjnMK5FACUOwDPsoJAvHtfp69R/fuFmbDKzPMNDqnTC5WfEMIns
PZHZOV48t25BZraMKQiO1SnH2MrP9r9SwkoAIKKpm9EONQQBfos/KJAyX/hxknxWA+jvN3hXVtmv
9AywsHDWMXsJ33r84nhIvqU6BSOGIAhEHWLviD5/Ng5w/heCDxHFl9e1Ek8/pudHoqo2gqbFs9/V
CW4TYkF/0hoQq9o2LDVW1hnqHRxtppBOWyM6Fgd/07KESX6gE563IKtyIX8jLdhioNym+NydLY3C
P6yqioxbFT9Rm4kt886njnccO9T5T1SoBC+8hzabuVsHPKRsWdFX1bA26FhlJ84uLM+wnS8wPSx5
k6V/dtTdX9E6ueXjzt9L1dqOY/BEIOKmqFUymrSjxY7caNRrIKsZsuUZ5bt76qd8wCrCWsB/b5Jn
X7uTutRiUV8zfDq3W6VU3ty0QJMh221zAR3hCyIxLzrJLZHE3Eo4VaqDQlgnAPCH10VRXIQa7Csf
bZsrQY5JPAtC7/CrG3xDsXsLerNY7Vf7ildI6PNjY5Z8/ohHVBEd7cB0LSqoBzz1sQIRBnoe00Ri
0bYZmGW+6fj0deDi82mLczxX1YRgrMhd1Oz2kLMtziySEXJTjrsmOBbHEiQ6jKaWarr8fmjldQNI
btPoMNF4CZ/7TIBX9NU8CLAwgdoFYca11hVUtuhxO+ZTwE28IzcebMZ5WaFO+BdhE40FkG7qTgLF
M+kllDLOJApgufXcnlz5n8WFpvZ6dD9+ICw83X+NikYQfR06Lk4LGEXsabob6syyaN8FIensY1uW
EdOksRM/ZB4+ijQa43CguYDEtw6cG2f+J+WEOnu17f+gqjV37PFmkIYCRJ7FG++OkdlJ21/TRyo+
rDmrqm8DbbcAJApN0WDgtFjA/Nc9Jx4DNI/DDcwCI0zsX9dkC15Go4ewB2d3gw4EqgEXGmXDGvzj
zGLBksO6uQVpLS10/EORo7HdyfHEXK8yMYIc8wwC88RVyUjRyvE4O3ju8pQoXIFp3nmdq1gacmRv
optNX71T3H1WOAzzpNEuAVVLhYRj235WKr2Hm2CRP3yRRbqtBOyTW6WvVkFpSrLTKbWa9aqnjCGp
0zNGxkIeVztS7PYA/qOfiVdw0LMTMsCE64P5nZT1t2CUpEyoCftQ+xw4nfjWOXEXBzh+lEM2z3yV
HwLrwB8hzxvoxbwMM4Tg1PjPOleX+u+50nCpBQrIixP/+97RgYobGAQGZpSP+yYCtm6b1KmwVCz6
+eq0pqmfrROc8Xze6W6EUhSjmxoofQErUPsXU+Df7KN7Qe6tlknQCdhEJpy5TkYU/PBenntes/hY
zofvD0Gw5Dn3Ms7682pBXhqfvmEYB3pLwrV+/pmGAPJB40tlCVWB7eFkzYx/Jt5C8TV8rMcrp5eU
tXVT6R0x7TgzFRheV68PRggS2yNLWoKf1MdZFI1BnitHFCk0l9Xx1FlojOzjHK3aaSkjx9vmRETH
cXY8hUZEYANifpJMAyLBCqbsRDhgVE9Ygb9WA38VfWk+Xxp8IjNNZPVohJMwwRvSe8J/RLjZcWth
y7NZkHAXKrVhW9H9+W3dStCmW6QlJCNkAFoZc3T+4aOZ9sNYxPypFN5qnFlESsTQIBSZt45mFtGN
Lp2t/fjQ1JbfEoxifjANg4g1nbXdpITj+DSCqGVlNRD01WErGW51RyWi4aINdLrkJ5cJ6Kh8HJS0
nYPv/+f0Pr1eF4Nrwg7bgRZeg2PHrmIoGgbQSIpDCnBOeeWi98iAnmK0rHYQ7KM8Ggx3KX7cAYKi
2PJYbDknxh0uf7p+ZJ9Mi1pebk88nuP0LE0O7PKFqBZqUnxYx870OiQEMIF/P/xGLpSyiRs1Zujl
6zzuE8RiL+hUKWQictD/OydsKDLHbEZm59iCO5BvfZW3LmN3zRpO0lOFtDjwuaLME4B7fonzBivt
3hs975Gea6pV9rL73j/zHYJriUA6D/ZCS9OkeESuDgyHBHAi7MaZZ2mEir6isWxKAeKz9PSOcgpy
vnJYyzyD7nuvqrUAwnvCt/QfH36j9OicDrlph8orUa9ak1jzWUzDYJqblzjG5ixgn06nAkiHn83Q
JKL41HPw8UOJ47LNvIvIMHcO3iERDzrdJs0JfqmsGpy8dCI7GGuw3+Af6Zwmde+gf4MvujtZtilI
h76jPYMfE2rBpby7LxcOGqajI7gPl8blaAGpWpaFiiUSNkWck+rePgViRyMv4obgJrKAdmjkXnWb
B2cpcIN2tXTwR+xwf9cY9QS5K2NZ9XgPKNfXamAtMsrHbcvQmKpxkk7GRq9bDVqEuBC03fziwLGF
0NmkbW9YmHl/OlYvSEt5kjfUnRml+rsC81GzFtifvzQY//6/I/KmY/b0R+bKS6FlaFXWogoalENl
EPLGQOkeTclBHGV+/qYp7r5+aHwDXdywrv6uCETSgp0vPNzrmXX+HKXhANMAwQeTjwtrKEfxROXb
AycLTAQfQ7R2obXoVyVei2xoxW9kYlJ4Qjanh9AJvIhoZM2TmWQ9TnZ63dB5MAzl8+LBufxAdbs4
pJUKAJHfZbliF2JUvKbWox8AT7ctMn/0JFsGxTGkRAQC3HmxCNTRb4Z64HSMRa+9zGTj3eGqYkWk
fvfjoGeuquK2ButtknWUx1cRIvbZ8eeDCLjTXByf77V1DegdsFtB/hgRa3TTAuEPZaDczKYp3y71
jE0mJTu5lbCy+nnSEns2Kvi47lOhkFtmA5mjhWFBk2HscZ87FclycSoKUUtmg0jmoCvAMoq5b+j4
UX6Kd3mHc+7ffXI6cpPFhZVynBeEndavRJJ7NfgCkeRXtMu8FV0je0hQzLhmBjwi/zGq0NpPscFp
VRenM00aR1sksBFQrhxeuFGrhXDuatC2dZTgQsnW2tWpsah1UTwLYtL/SIMUnnO7/AZVHFQXt115
0JdfzSLDZb3EN0v+aoptFwIPn13/O1iu9rnBxbbo1uZ5erNJtOUqNDlGUFzAqUqvP672Pm4xTxh5
QpSEATBezuoBFhD9ZYd0Z/N17zPK5qYvB9/Xy5c56bSlMcf9SwT1upgE253RXCSKUm4fppYSEduc
XjMuDh/KphpI1EbQNDzTV+/nhDspxSHtsZWRIybUoS2UkA+FGbitRCJxqSl2dcgJnSZ2PGM/zu2B
aq3Sg2FlXgjQX6MHvVy8AgSFvXHIQjapblZd0cS993fl8Wc1SFh/hxdtIeC0fbFPwsTFPhkZYulq
GZXEKSHXBCrHgnXv8527j3Y43TQoJen/O1FH+NyAzBuX0X9FuDwHBw/ZYB/FW4hs6Mta3/LzvCZU
bduCVHf1/TNB4e+g3quzzhWXQMrRBxSZ01/CEih1EKNdYp4W3yuJuQeVqxQpenuy7WJz/L/0g02o
SZuEJCccygaAx/ANH8uoexRJAAwzpqtBWUO7Xrwb9xnB4INLhRR+Lavum7syylFK9nTqJVXHMdjc
UeT1zKUbwFOruJ6M70R8dQFurw8BnaEGauWnZB3DqactDFu2pQVd0KcLkkRA09FjVRm/QXObIoUP
OI5TfG/SEJtNA9rg8NeSNiFQnohYgd+opuS408c6fExqK4Jj20GehdtLik15sVprx6yXpIp2lJac
Mw6WStGSvJGTys1e8XecQ9YJ0thz15Jlh3Rffdx3daKF8LAlqUhRDb2r57ovPxaHz4kJWmq3bh+h
WLWhB6QkM2Ny3zzGFFJ09FitthJlc4x/HRHBGdII/PRkctBrN/u2PydBm8ske7s5O4kXwd8GPIIf
a/YlWynJ7hXWYzOsDLDn85F5kjvB97WerkBuX5RBiqLcRDMAm2h/e7b2z7gxUm/o+TsLcOBr/VU+
iDt/MS35Wi3U7oq9ZYmZ1msJzVK34M6sZGUiefk26GE2YPWDJLLVxWbkaKOMiNNwZXXlYBCDpAbm
zpXtaf2UJckzca1y2cQ3hY/Va+oaT4mgH3rbOc+eFLd+HPyB/SStae09tUR/AtpryzF9CNZkVFZK
DQr2ZkoG0dGwPjROQJ/96cT0S8R3EmAkHILXzoNLHcYAnrxdqSwP0BVzm8ppSf2MqQ8etW5Wc1jM
y0HMWRpQP/cME75ISPrZlRSSrBipK2d4ao4RGWc0DeHgNzZ0w5K/EqxG+vd3g3RQY2n0PbiwEXfT
GHk0lmxMz1TWkJkS5bh/eOOuh+1iUIsd/zMgNa8ArtifrbkFW477gE+eiRWbKCHkIYcfZxXkUqOq
A/kBHJmYFjroYHPblHMrPT8yb5esQVai/yMwpTbEGrQuYNPfTj02Oc7fFdhn/Y6GZNkXHw35E1j9
LUfMOMTSpFujwF8HPOs2Pvhg7gJsEGkNvdSKYQfUx25MbMzsHRCsN3z3BcEy0X8bzY5zFl/ojyg9
ltitjtmaZ0FFmYxpyxpZh+tmal+xrzhkKYMnqDD0ioCLXXjJ8H3Qextnkfvdmhme7bKQ1Q4wd/6B
hZSDtCp4IXegXcwtn/cfw/i8eV7iVJ462/RkqXNd02sdSO0i5rpxLtsv2UjU6pMyMWxkU+Vxx7yw
/vMv0cpvaBmCQJF3OdkkZUCPq6HqyX/qwRl5FStCg+J2u5LIxHz057j4Fo5mULdYzuin1VqhG1C0
UyfUPJlqCe3WUtiG3D8e7Le66/hPfhPwPJuCeLkJACWcmFPyKQaoid3TacRNE46RtxVlbzsAelmg
x+TVkVpd5O4C4KMbGVq9sM3F3foiv5ivDXeAX06B8NNfJ4ERsUnbQM46K3L/TcOxDHbbb6sfDy5q
hCcQIQQ0G4NZQgWPZ8sPKSzxt9unq8kebM32y1r3zv/34lM648NQAwlvlt2bXfmBDVaVqAM7yEuK
AZiWF/pECg5Rrq6+OY4WmV4YgCYteQkiuephNK9AzZ+C8eAM2QYDUYxKxRFzUZpV2xW/hFpVEs6x
R1SX0GCwI7MkBNIAzT08/rzJV9RA75bLoIlIKmtrTpybU3AIWY4gjcLa3o7DenJ8kcPCN1FjQOSz
E1h59BUbhITD0sbZLV1HhaOLS9Jwbwm0ya+w6ohi+zj/vsCcPOiwYxEIRuoLhujap60JA7kGSmLi
EuOMxAzU8tcdz+PYmXvFj6nUJLdB+tIW2mmjVJTNiG252b4GFOYYfLIcbqCk/uRNfhgauFvG6Ljw
TDxJgkrsqokdIdknorxWnyENH+pYsOtkbHhnY4ENC+WP8NuwkTCKEANbhSduhz5x1h8XXIlE5QaS
H3DdKdG+pKCIvxiBx4PBVjbxayEZr7AmA+b8TgUu++XRhj3SdfMAKjM3BXszhl9R9VhPWOD3BTQL
YwMMdi2zujk1ILMzlGFlTTPA9l43kY4ww2Jilxz3O3KaIKRM1NvySxDTsQN0bQTGHpeNxqG/M3X6
khHXEdvm7IHFplBXsNacv7ege8bONkRB+InDj0/Kgov5W3SP23G7X4KeVdehviLnRBm7walsdKVD
B7Px/oSMoUH3d9hwqtuNBAB3iuBX0iWFJSgX+qgVGJ0bF7adX4w6sEE5rl2VLcSPEd9LwAdCdGzs
49S16gyAmVgeRfl5fqzuUzp53JtEIYIUcfz+ory5IwOpnbgEA9D+/gbKBCgjpvqc/lhF2R8noDXr
jHvHcRIcb+LxHGcxuYV9VhvKJWHrS45AJv7+YTPvgaZ460EmG2ccZjB127i5t7gKqjRf3lvqNUx8
IbR685N1hUjhP9qkQK2BMF3ca+WMmYhCIZmzvMIu3UsthNEA7ZCfK0MF/830jaugFI/vCIk0RLoW
XDUCQUdNEr2TtQx5aIHoRlNsdAq23z+hALvlqcCQHmBR0m7OmgPP8Zem9zVWw+hPwA8xdmSrZ8sN
cCfySM4WmVxgaynq6uGAZb1Lvo0Xwe9nZHTSQi4bMMO6X42R9GL7xnQdkew9qt+4oie68iac87vX
XQANlbzcL2Zed09yAFxVim251TsV71eet3QwRe6cSlx1rdo1Gc8Jp2A+Q8h+6jvn+dy9qqpjgv+q
8oxhsoHhEmrMbwWqJQ2iOeiP2QPi6hcodYabGENGhLbSuQNYfSMFKtI94vncmzgQfRJFCMwNDGWD
hLKeKQD2FsSlE7MkvuQHFSH0TN3Bh2wmWedDCUIC3eREreC3Jx7Drrqf4k2lY39XKsJA8iK/Fet6
Tdm1gIoDelOHb9S5EvkHVNl3Y3euMUb7w5K2BZRW9ytwxROQww/j4ppbJ96VUVdZYzY9ZDW+aywI
s6aXv/QURwQZUZqWaRdgB+B2n4Nx6ETL73YY+Qme8H9c/ORKqAvDtifE6PLQ2Ww+rTQLazb9tuzN
V20jFueIlPq69p7UposQESeyQvby5ncAEXH7phBSIKoTfTh79fnnhjbw1tqUFB2nKBam5VPavpdU
CtmyBJphb+7gKe5NBwZqpt+TZfVKpUuyFkWnvk/WquQ/PZuZLSF0dmxiJAIDzDSog+IEpjIwgUNY
KcOtsZJ/fZGL3gCOcea/CDxM3t41rjV/SArYrM88Xv0k8shsNZ+GTYEDKynlVxf8bli6xGKQED4m
Oa+nzyuNmSxmt0TWBBzC21h7oFTPh9tg433D4GuHFhsHyR4Y1C/zbakQ9X4y14RyOimVFzYiaJ3S
VxddbII/ZLj2Y2c/pQqY9wqRek0bA6TZdgJlRBt98xxZaf+cgpPJBwD9hQz6OlxyLcIr/+Y5Aq5G
a3PBhwunnF4Q2tn1A4Lcj8CaqCulS8ER/9NosOvJ45mivMUfc2oo10eokMLbnKiP0/rneo+KMD2J
klUV55dp/mJaTITWOcGUsS+PQW1ZzdCMUfR0Eek5FVuf0pLtX1ibH/mHQp20+z/FVXlLG5LXRlj4
1sCxBX0U/f8QACu40+eYhQSE8g6iS84ko+JV8TL+z6o2Lh8hguDiNgWTjICmGZ15XCrs/LTgnQWU
z+YZ72qcVTRln5zwQZVhECFLmR2ZpPVMoRp3JVk+EWD32LNCFKJ7XnMUo7lcyEK3Vzqmp22LWKK5
aoqm1dXWFG8lxyW4Z2rAz9PrWnbO/7EN2i1qJHYYvemyKalgiLkz2XYsaNK8+zE+zMANl/r7+9mR
K0it7PJSaIsldRiTTfMSIHIJxQ2zVWViGSjPGaJ6HNl8ofxorDbaQKO+7bWBIrbdZzd6yGX/qN9N
nXEDXAglP96iIwcpMBZiT6cSzZbTJe3Wcbgz8UPYwBqht9p/KNLEXdqOxIHpcsVAoiUEwuq50prM
eLgY3vROd26gNexL1A34PUh+bqF+j9ee0LiUxJpVgqY1q7szka6b2Jc2UfRL9YQhXYxVOYMChPHH
/XqNT+EqHXsgSLEXsuNf222fDAdYGYUDnhfNsYNKZHzECckNjBJyS2B10KY2hqRNyTbscXJEGArQ
sIgJ+jtPoKkNT896EULLae2jMaJCqxcWd6BhSQFGW0/lXubSTWG0+3yLAq4HzsrKGVygqCQGQMIf
v3eAqoeL0mlnayZihAkXn206xElrQOo+f/kSJYuKih/9B2prOAQDPz+bc6ElPMi5fBgU09t8D64x
a3wfhWoQHuNshiWrXRaiLsMDJv7P5SDVcL9G/4h0Xs9OD+wTfAdhZ32OZRfOKawqg5FWjbFeY4cp
WLYs+8qWslSwwzCL8unV7WP5lqTkilg6ZWaDgrskyb7R31lXDTpzGYuhYUPtAqkH+u8wwU+e7ugk
xFji6LOTsR8leaFuKFcswfGDrqzekJ8f9AWT0Ixg4PLzM683zkW8BGp0yySMX+hdiFgzBpKJvDSz
lQxW3fvOfHqHP3glYBjpWjnWZ9zkz8BhTbpT2P9cA/x7CMugGSV10id5BrrzvlwvFVI0cQto4EGS
VRPDTt5+a1rmBugrzjwfoemiRRFlvXdIs4EkQXwnnXmlX8eG4nWN9ZDxA3rs+v87t6up1/K3TtJD
Rf4TBuTmyVdr6EQJVb3/C4wWTgEMB4kaZXnOp6PgdvhPjn6rOM0jy314ERJuF5czlgEJWKeXl9KS
MqUN7RoHpPNBCBm78WPcUT8e4KhJk8yRn+wIZoPSFoTMBUOmbpEmFCJ+DkXtaM7vqa+OQwbg3bMc
HNx/OwTaynmyiPPaxV6o696ZrMs7uk7uI9VfqpcnRJYUUGJw4CI33wciEiJL0wwpEpn75xGtZEUA
jfRtsXOBzlLd3OFZogKzInBXYeRDmE+NsiE6KSIVzp9kkfeUAAloNZyD9HvEP08vmE3bpBJy2a/l
l4SzYdi8JkWeAkWlg/lVc/9Ejt156VjK4bxkCcQUJQBE9wjrStcJTU8KcujnHEYJO1ZZf51EpqcY
kESTZHeN/yPskqzsMGuIcMRyU7Tmo73vmdqALR3a8yJrDpOiRkFRnrk6nu5WHINIhsa6yg/iyrRJ
bnzggRBC5aR/PpSvx6iV7g2Q2xc+j+2muWkHcvgVdJA9evEtjM3SEkRFyQ0Wykt0NC2h5AsVilWq
Omj8d+MZhSZLt5mI00r66GnPie9g1K4wClK7QOdCowIsMwNuuq3SCMizJ4WuUKSdXHwgQJ3Jn9rL
0qtaeUmnjBo+v5yKCS4Lgl82GG+bBn/LGjiyRUt82knlhwRAcfGB7b1i6WZmcGNgx0y+fIzh0/nY
RcTBsMluKg9LynLllfCeVwxYx9foedpkHYYbmNDvz9L2ZHwNidMEPcdhNtzYfwg7q8R8b76H+j8N
zBBxXnif38cvEFbvJf8+x02c9uMxm4XlDEJPJvD7XaEUYrG+6PyjD6wbYmSv64AEbJXGdqpa/drn
/LD2IzLeuW35vt1kJaDKw26y8rDQ+TvzOjn9Sawc2KNsCFo+dpobOQr1VXL3GZ6SDZRCLyVGCBqK
ZU3R2Y7TveZiSUCdiyOF6nPO7Ri328X5VYu34rSQLZ7A2RfzuH7mewy2i1f/IJ+C4rH4Tu6TxaDD
2AkJg9bXrGfldoxnz0cyM1n4M3ftZBnmlnXDqXUVv3AX1cQQSAHP9fcT51AlrOZcleS7Wx6QMw3j
0ud+ysF7ICBujgEbai8s8H/ZgOvnaFjnSlJXqDccgwcv/oSQaJ3uPlQju3yqyO6q/5obmrKCGXuk
2Y/6dviSqiMCbMiPB7aorDVglaX2lx6ciAJJnzTf4DnLpjX5OTJfrISPqQT4QS6r4NkxtIyIDcNH
v+f54K4GBuUYQdanrEda3bymdneRN1o4OQawrt0Ogw8QclGnJvcI3J9Qhf21UuPiBWiRDYmxzc7W
d139thFq+aQq6yRtqf5PbfHKuBTOS8gYz3eJ3sKWGKsqQeRB4Mf68du2DDxUqeTgiwo9G/TJOJ1A
cu4sqiw/U0xFuc+HDmEshs0H0EYeB4S/MyxlqSCQs2KxsTwEzhS5RF/gUK1+zx3nNLoF03G7wnhe
uRJ3+0BM+K+1IHx0qbnCNdqNaKdMC3OEXPcuzqON5Q5juDTFFG8A5y7Nl6zspNYh3RcIo61r/ZYk
PGxtYSJENhqSOXm54yd5eC+/hZRRWweDlkTQGllD8+FC4DOgvWXRPmPs+Q7c3Xn3K4XXdPhdpOjy
kr8UuBJnl0+8eHuMyGjICwA9L78yc8IUFVnu48tDXpjGtDBY39DEjoAQuj+0faj87d9eCfXrw8tI
Issh5x1PehZh+wfXLuhHVLsh7AmnEHYFcNf+rk+ofMaIiiwe7Sso8mHrh043TAG2KSZX7h2YMsHe
dBqDIg3j/9p00t9/7LEkxHeWi1hXaxWjMPherM41K3vzcF7Dn97oFnNcK0U31P4dUt/dyGo5O4RD
WCgJCyhtR74+k8OhdvvJ2avBBWLNzHdho9SVS3hGqXGuoQ+rWfYWK90fmqEWE+vu/lWDoqt3FC76
QMTU9otyve6oJ7ZCcasFML5xPX/snL+CYqnVESI6r3dBKXbcVVLLh5MU7FmufE2LQL7iurlQDOqy
SwEuttlNgBnkTuzTsp6H1oqxj2omnfGQRReboo7SxrVUZKN0tcuSPsoGe3gDQ4RpM4PjYHr7sUcx
x2tTXTT4nrfgqpeg2Z70GbdijGOJiDaLnBKh/1RMgKRjb1DtyEk1UWZNl1/Yx5Vy+4l1AmrDB8RJ
+eIJ2RzMPTtkJjZSTt2mPQs7YUM7gy1ezNR4l014cqEFLnMydlbSJBxGjvUy4nBQMubF20ZmF/wz
svgwkfEviIzXi9Jns3u+hK6rKsF9cre+f5L/j1ACwrgaxkmEHXam6HRi9GmRvrbKLbi6RQlfZodz
1M3nWLwYHHTUG1QjZM0wCulaoCjW9j7jsS+6U5jGA8pZGgHllOl+Xqlpk7d7N+4KnypYhGdH5zwo
z6t48y7cNfoQS3s10Rc2b+HM+9XXDttl8b7KM3niIUIte3/1ISP+5Qpf/q8QX+ugN53iK8FcaZ3t
MO4JHYO1YGF8ylJ6b3olL5B6cQkwWFM+eQT02mLoE7TvrLiHL7eUekabRQdoCyNjsC5OMcMR57KZ
rg+LyLCwzB+9ic8ikuGh7mW2z3GCqjv8AFDoReGYz+NR/soUvSPsrREhIJmcmOWZm/NyPBt/HtUy
IXKsy1LfbtgeIk6Y0mwPH4jHKG0E7UUTiMy61fiwN6LibYpi8hTZsji/JePvv/DoX3+aLLkA7cKQ
ZDvFxcQCDWBcU3v5R7GgC3oGN+cr9TYFeQJQArfkqwrYwo4AC+Mwle6EGzkRnyseo0iai3prlU36
1WBJCqG+1moLjGtQ3tT5tibywT8cztHKb5I+jtv+ECVhaxWnf2lYWJHRteSQH+EDzTxJUniZo25v
iSaWMMEi5L8O7oGMdlQuLnVu7AAlmX9Buiimptet0rXVLrcCvDlKqOYfqe7JrbkS98YuF+iyvwpv
zszaPpxCiD2hm0qAnM9HBV9b/TYL0HJHV9CtWTMwgR/JFroDuhk2x3+nodEWWvhuJnVVkE1p8BqZ
3FYj5Mg1Oji0Whx1E1l4HkR4jcotGXng60ANhUhCXATBg7sGglKnzETyZGbrqA0wcXw/EHXUAAtu
IgLwlLlTA2J7QChECQ+BfERyrB+B7kf85LGtPIa+n65RBz26cp+hExVPaXsPMKImDWiKb5kYpi7J
I7U/iRjeYkMyOU0SeZSmNF5AcQz286SBHebR81p8cw6V/JgI4jJQ3l+QXg1zOYEQjj2bLUgKb72T
MXFwn947F18rrx1jqc/L6jFLjZTK7egMKQf/TfyUmAJaaSVCZUwTczulOhR5ySsoKWnGTT/mIAeE
JDGaD9TYOXX5PEUE3wK2M+zw+Z/JoJHdTQTJwfj6ybGMSzL3EsbyMC/15tVOF/7sN/uWNELB50Pb
eKb1JnhDO0Rhi3tK+96B7duMl7LlyvUvnpSBjXPiyjzwOKfVJWXvGk/TIQYLKNzpoXfc7GR6vPx/
qwYLt+1O9gLHYpvL2UIcbDl8xMjDgdUiwoN1BUBpH87GpplknQs+TNFrlCClqLKP+ReGHTZzADqF
QPood4wa5nRaNFZVgAOnTyHwpwduxHXmxwtP6TbMysSko7p//GjkeQxrX7l/BxyEReT5Hnk1at1B
OZZ35HBCLHLWTEBS/iuBhs/NH9mtiszB6+q3aZi5YVIGPgB3W2E0g4Ui2VR2LCVTc8UbN+hZIw1Q
uzIAIWjErdTGwRAQC0M9ojCgDTc99TD4PtJfyHIlMTeJoj5UjGIhNi5NVwUYR5WJmeL70Lx8w7WK
Nm+owJP0GnI41vlSoz4YIpfC8K3+TmqLLdxED/7qsvFoXdJREJtR4KkrG5Yji08FjfSyRFRl0Qb9
ncWNf2lRxolfrj0v80yucIfJcve2ipE7QHEiu6uDkkfAtCwbPaXrmIdap7miv329j91Az/MQlSS9
ECOg8Xm3OWXYpCYBrVOSzpY+2R7HYqgbK8ZumC8ii/vspNkPiymcdO7/k3sT9S0CnAmmvdiRyU5n
9Pg5vvbmatt5JkB2hRd9I+I428UGtBGqrMnJhcQr8wxVZrZPIE/X7ZNkt1d9T05Xz5hKhFdjX9nh
M070YX6yElk74lAfFLTJkZc0ap4jUK3ZHDOkqGtEJ+n+V5fJl/xwIjrKlgekalxVlLWRVbPqytVj
AKtx74RD4tnSkSyRPhUP6E95M7QOE262yj3f+mcMiOmWqED4d3Klv6453XXTkcfQSsQUv/PSVHEb
LB5C56P2AohC8+oztYWLlC1r0hbcQf3xcJDyRSZpDZFdPkZt8bzO/Zltk8GZmAY/VF1XPHOPJ64i
wyb3daH9owAY5WkDBZiEuBq55+N1ykWATV5DBX2LGZM2uo0JK1z92EDwQcyc9qOcW588n4I+cx/L
wYrZe4PMOVF4P564heNOyh47eqCWHroFZKfBcXffLA8CFLofKi8XqhlLJGWgF7EzUxtUnj2peapz
ns5tNo71C7eV3nOb5JnMZqBgn/pYNwuEa5X7tKAbkEU2YynFANSmFzohGI8qmB1IYlLFpSDnNVQQ
8AJyzohTyEbGjfAaEGC33nWAjeszV8YibJ52TblWR/cGL7hiSZOZ6wxIGjdS7ef+8s0J9pPoMcru
EyQvoRpi2oSJnstl4nxmbAonPJhXhZ9QgBTGUMKGsDw5YOB1BFPpm83xkHAUCPDZZSRmG2jxzwGA
Xysc8HKtmhfTQCs/E15pmbErtS95meumHqf2GIhBAZT5sYMndx+ysxo2TdzpbImOZBBGS0s8lOHh
Z224+yXwnIf+oPcS3zRY+pYa5QJrxEIhU1L25OVi9lXVnOowOc6UbsvRQ/61HMWSVPuW1MrFIJeb
Feoco+Qc/saceMBsn8mjFkK+ghF2Is9dsleMGommv+RKHZkDrT+zIiS762wNxIfwwoERzhapQi2h
/QMB9NnJKxlZc6hL0HNj3JU4Bm5d6VYX3fyb3SCECgULMAWCAYevuPeaQEGOv3+Bs7rOnvHPfkEK
f05G12UvJambTv2Fo1jtXoEFb3LV6/CfCvnYsCABf5JG6+PC7vjscO6yef8vN+jnIBRRdApDyo/b
otD0WOvIrL5H0EQhlx4F86gpd0DNcUlj1YEC+Cv7JcA+xlZIDfw81hWdyk+SXEZneAyZJ1WHPHw7
+tqFLk3rIid346R8kTBsSItGxZ/ZzSAEY2icsmtvakc/34hK7cS6BNVW9kjKhhq6RTz/QNqrXV4U
y1lgobGtVlcq3oFFaCfR0gZn1cgjvz1Gml/Ee8aSE4qfJ6c/tKWdnuzEWAMWlcPtnctJJsO6kNlj
3ZMj5I7x38She062Smh4Qra9SEzi95TLYsG+nu0OL2395ur/E1dTMy/t1pMkgkSXPINWQkF/8cAy
/QH4OoBmRlGHW+ki6rViWKpH+9f4MuXIYPbY29/IqYWdarE3gzJKidiJYDFGgQFNIqShmgDIzqaJ
IHQtwljd0O9afRTJdQtGVR/kBtlArvpyrv5CbZjyVdK4RSFNSp0wPs/GjNqzfLGNX3291bDvpzmM
PGzI7zLXI8cPY70k28mYR6TdReqdK44vL2rvK7MpjXAoduq98JhpNgt/Qt8WpF4uVNWSIEUmZX2I
qUZO8niqIkoSBUDfQA9GYyE4ac9SQvme+RQj11/+vlvmBZdrrm16C4EAMgs/OGk/mhC5IBoiAUUp
PgSSjUMTEXNvddHzcSNPc9Sabta+haHsiZ6Xj6u7kNuQGQJ7jtIO1u1YBebFKuAf/2OiO0lVjUan
1hNco4kq3CyzM12dHZFH8Jk5jvSuWCekaOO11ld2ha9v6+vpXWrYBNRR1JFXD5jXuhv3tcWoEjYJ
bwCTBamkErjuGq4UMyO/02mZSJUvMPO19RoMdhI2+nxtdSkZ9G/TGeKSCGuZ+awq9FGHRa3CIv3C
TtvvTGPhiwkjM51Vcq2XUZhy78LIIksvhhGNwha43pv6zbfqG/8JQiytFIA47tFBE1WtmVbIinSJ
urUbWmt8jYQuwVtYye1QS6FnXoMMHE/LRTmNVOKCwFeCQH98LZvMkv8FyMTyS4x4d2AJtb5O/2Pr
Xst6B2lyat7ZGzTSPDh0Wfu27JCkkk1v+Zmh5iFl975c/iuA6XvOXnM7rkIO4sGlGEdGUsx0RYf/
mzFtkYxH2XXUukwfh0jlAgzDzNGnXiu/WSGOjJpGdPMfzq8BtmoksZQe3LTbNrQ79eWEKqZd3gzE
Y7wguNANyPtThZwNkY8zAE8w3JnQZRqZ1X6JZQoP5NY+ZN3ZLi6YHAki1inItzKDGAQv+ot400AK
0EP8rg25VTxgvqDdMthPbOTtr2k36BekRHnqpb0w0fJPwoo5cH3Wfm9VvPofFOKVzpJvCdppGGV+
8Y0dR97mYaUgsU+DYcLq4A/kfPW66UmQuODXt9PtEcVut48FGWxuXh4QKIl5A6ALHt81/ngsWFwH
9lXGr8lSphJ+2m12Xj5UR1hquOj4pI1WyMPPDud5VoufNRTUeFxKX27/4ztzDVh8H9JPAuyEAP4z
s/uvvly1UjMG+/d2RkXlWef6hUTbFw3cwrrnbwfDsmQhAorzJaC4xNChYzz0ScVKR0b+pJtArczB
h9pJk4Du4A2UU2fFfTwHONqH3U603eBSxiAL/kHGkeWGs/YWr8klaIlv8CUrN2jwC1nKze5qgqoB
IhOyDZQ7B/a6lkXi/LkxsNyQbC8ZhtqWIIucmHYEfOcm+TnDRj3r7Cc+Kr1LeanY4rUiHeoXRBkj
kDi39R2QUcsQff9zmi39JZd2Dgx3ad4qAJ3C6VIqrqNi/srT4olbArjBn3eR59efFJ/EaPPwSrpT
/YXDTm0dz5dNxqpif4p2uicjK2OQLxnudJ41OGYUEggQ4khc6K7w0LJg4Jd4MJ3ekyzu8gfZOG8K
YW8//KI6Vhns1z0Ire1jecSD+4bq0TWkqdaewFML5lecxb1rh6/sapLRoiJkuSTxeSkRLb2f1CO5
UM6ERx80fgC591Iaz21dgboDWDIusi6l5BycrJTfEzBajFsfPvYqR6NNoHkWnodOK8EYa3rMsimy
n2ZZaO0jevznshkO8yMhxXZhDVb6JPWKPz+sAkPkFMWqxYNzV6h5ApRVfbCB3c3xju2/aI8zNP0I
khm7dRu4FP+ZPh78+SbI3gn1pDbihbrSRHCNUC1wQQ3l0tiQHyWrXgknNKMFHEOglcD4Ol6UT65b
atRAxDHYUH3f6anmXXOlR/jk7tEV56T6oQVxYr4DXH3C8V9uRkb6tWirYhfx42rg4CxRbknfjU7B
tTn6kskz3Ewx/cF4FrriYdaoFCaSQZ3vKWM9mZPY7gpZgE6VmFSNM1zvkEu3Gyte9It+0FWK1guo
OaDA+KCzJIHEyZJCj1UFKC7tygf1KsrTBfQ6KEdZhkTKJw/xKqvW44HPIo1ak7bNwqNTi+UuzXLw
ypU3QzuBaAZ7IWeoUazfzmnzObPlUttuX/+Ut9aoHpzD/uAdbQJWhI3KpdkWqZdmv2mNQS4r29NP
J8ya3v/9XTxnSA5+pN96YW8UXBv92cxFg+JiekS6y162pkfjGIOBg6litZhMrzJwxvuioWq6/pNV
kCDexCDxL9LTFEQCQRQV6NfH95t21tNIov4H85IVZsJTTmTMsxqYkQZ64SPZoQzEgPGTWxzI2OAh
im8iRqoUhugb4qA3eT9ilzaS0F8NzGdOElV3acDNyuLr13cdg0Yg69GLCeX3056i953gHcY+sc/m
EnG5WWMhEPOgqHIxnvGWWQLMdGqKk7SpBTQXk8hev4c1+jv0+zGly1a4AX4yKurq7rbQIW2Vbt9e
pz7iOi2aWhyy40F8aQ5+HxjIpWTKP0aJq0FTu9+AxBzjCdTaudUUTVRh++EW8U0ZX/OacIaMpGks
G5RqHHvMV45d/XDbfRsdi187S3Gj714llC/SABhZa89i7jgnYbN2COPrm7qnfaNr8f4BdaZ1ytU6
y1RUU7jQmwOjFDuYxlcCk9KZzVR2QTPtayXNaS0RzROXBnUsmby1oPfOhCckh7a2qTUXCYVGHIPa
NdPDfnX+ytilBv/G4t+iVKZBVt64MUBzXugPMZX5elcgtfaurWhYs3NnPNhO+mjbeIpCm+IMmCrK
L5rOv3ILfWT7F+WdW+UV7ArowuQ9THfVmQIwQkAoFI5K2tBC1c/LFBGVi88/vQ+OsIxGSgfcKwOw
Zo31fcPU3rs/yN9UThOEKEqqpmd5Kb3nw6dc1cs3uPtuYL3xyR7e0JqRaataXpedtDJ1tjNh5+3J
MwdFdLuzuXt9K+DW0dCTr1Csk+9BG+OB5RwgpnkXi+iPgTTl6oq5nFveHHMnqY53zbJ7HkTF3LQX
1WgkaUKMs6gyBO6Ceg+vBfmensTflQUOfVeM9ApRbpet//WPuNyd2H0EhKKZEWi5mhfLq8Ptm6mf
eCDb6aTROnGlcdbsFGnx2tVAFUUhkxrhhKtZFyMGGisADDoUiDgysS+V8svKDoAxYlpMOobkr001
FkS2ZMkWkhdCn8fAKTErr432B+IxRSuqnrtvqAE8Hnkt/qZizLBCngTldF2vVAqM/2ZpxMJpBE9I
JhozhRPhW0s/Copzdex94Vn4/0QaZhD36SK+NlHXgAZGZIGi5QLtdJSdj9pgnzCm0r/lAm+vcGHk
GskGv5Ow6NFHELjdvEnIURjMb3tjFcYOvlFhrhvJmx3DNTI85ZXrJHiopCcp5Y7ejWGe+Ggpzg6l
jgl9mjYwW/m653WV+gbujeRaD7FjW+gz1M4rMkPJHK24jxmO9si2kZRwaz45emlge7wnJnrBWmK7
vIqjS+hYAxcfVINv2tNeR02iZRAB2KaMvAi5GC7tk+UgWdHfu7OAC/O+FyCWwTcy/J/e4COof2st
6ESFCyDOh0bUXbVFnC8VsXnweqd/TRToXZnzFMKnR2qRZ4Ra4kQ5GXgYeCK2emGmSSEhcpSizpl8
k2skQzu25zyJ7Ydh+9oyQl3/r/CWxirJefdTWMOZ9POzGyHZkh6ETy1uAaxf5X9TOJZK/a4ilJaG
YW635W3tSrIp+7nt6F9jT+KU2yAmJTLZnZ8oN4Q1+I9U+Xd09LEiPOA4GeG25A1T2vNLgLE1La2m
+uAaZnB1fvn1u5FH6Rk8kMfYTOu8jFDZc4iM6Gd84VawGGSiwHq1twG1FfJs7udV0mTAJtdH/wc5
iq8eMPjfPHjv4v7pFVsvhyi5vWNq94hlgxTIPncFllQZRvh6l4jF9zkT3sip31wqTTMP+0o8OWeY
IaSP+L8xsZUq0ltAv8OnYCSPa/nmzAE4SzevJriNSOt5pMIM7RDurZko9GuhIpZ0RWQ7B8G0IOBk
mM+VpirvRpmXvJ4xatRA1snkMB5+xLVuYeboDNcfQceQk3FE6GHMsTD75pJV8SuWTWWrUGKy/wLn
5ZI4Tr89ET4PaPglKlEhCob4V/khfEWsAc4BuaT5Cu9ekcU1qqxmMw2Vltl9wyJAxcCwaXvx+ATX
32e/Ypq4gqcwZoOJgpGEGkHH9WND9i7vDoOD6MqqBz9Ew+O30vd5NMccUxiRAV5SlwYG1AYHZws3
kfvE+Rp6mNRNK7mw9QpEdtyvSkgXkOWBOgCx3GfmM3osds51heMfA0aUUxvRy7XOBPt9sLklJSAA
tjL9m9fYBXJC5jmlg26tRX0wykS2he6Q60UhwdqNTqXsYdAs9YgaDvbWRBJ8sUrFXa93mSAsuPKQ
zQcv9olAxPb8Zl/hG1L16zM0arpEB2clZdKlIvlCgnMBhwgxC7G/5F/CAzGazlyujWbqpX3Nv5MG
JK7c078RylTSSf+PJ32qOy6oj7SeEuJbYjqTCjFcoSMMmR+AQt0TDNw132FN7a2PmqJzQ7b/eZ9W
3xgHRK48V/0EEYlMVBC5MPozaenvsT7drk6IXEAfJTWnHcgExZvwo3DgZzhmA08hTqrCg18sC76M
GAchZAS+3UmtWABTXX9HzuvZ49x6CNJeUMVHWMc7cTqnHx5vLMlmud03i2dPRBQ48dKvFaZOe5RV
PWyUsbk/DtupBDIUaALFAcFQGbeTfmIkIL2/wZLQRo11ZFQw5jGr4VKqpy01pomNuObyyHaKbgTb
o1QaPsLLTwe+0QFWQoPGsbM7ZYbQQCH4PTHSBLtEscCL1vXjjPgbfBsqxMltvUJ7Pa+rmb2mARHa
dmVfrrMswaIuDEWF2jk29nwy6bKveit1uExaZal+MognHrOpUEuc+zNbJNhrA1AQFerj+1gpfBXg
v629jL+RIf6KEN8phg1ORjwhXT0jbZVs5isFxhwGEzx8xE0MGB4xjfm9um6UWHv5KNhpN6xg2lrX
1MAwIM/UnEP/t+y7dWhwgM6uNCrxYA9aE3UtN+RJqKkdc1ve4x5IGX14aEVNRKJRc7fTXe/30Pc8
OUD5MTmRTwoPmE3qYzl6GzpcK/rbzHAhFG3j1Hgt2G26AgmYlCSnyaDSnvhez9gSkRAn7mYTv8Pf
yBKIdvZxz8H1v+Yk/QBfyy0q4h0RC1ELqUQZBoAZQlwmDO3+yMwm/ksOQn2SWO8scAiQqOrTAnYC
xQmJ0ovKD5jlYHj3wPExk3Q3FMZDhgYy8kBtSyPjbI+4/e1EFI3wZBfs7dcIqCRB05V6v8yidcq7
hQEA5wDnwN4tYXgwAogSn1mkLD4rmVuERlRea0IIX0NQssrI7OxU7h6qV+Tjtl4epuKlX2oWkJfb
frj1I36uD8oxRPcOxGe5pDRiXT7lCYTrOydTXXZXutOvhpEoji5CpvpcI8nHSRDCsYm+vs9gx25+
OVCmMNmbCDo9n87j1EUzMNd/uCZyUM3Jf0ffRicBTWUDXKkT0jPSZfpsLGdxvQxAmin9Z0kVQyHe
U1M42DIYofJ0CvhwyXHHOssyooxwwPiG3I8wSYmkeaZWxTKYMqNi2p4Djgg1OCF8+usmRGIfBgK4
48I1oMxE5xeOJ5Y0so/jAz8eUPWf7Wl2UT7czowZlxMfEkytYGX9TMxTntS9TkUzCdR7H8eZLp5j
3q9JN4IotA5XEkBEZvI6ABvIRk7CFDmf0NGa8PVqQgndLyZW9XpbeukYCnEiJ4NIERMz61tDv3uJ
lyby+IvpRoP359S5i+53l9R2wm78AZloyupnEN22Oi6BTBD2dig8a6G59JpaRgHgrJ1k1yTyCxWb
5xeN5g4ZfPEKZO41sJidW6+/Ib5hD7o4Um7bD351bH3KhCwt2vBNrGKDMqr58L/jcoWOKOFVExQG
VuRRklzkizpYHiSIY3oYRxfOvXlxneI4IXt7yupfq2jV6Cis/LDxe/cDYhpjeCq/QVxpgJ7x/B4o
07T8FBUvFvuxExAywQhYtAsTi/U0uM8t+4ZSMLbAkcY4UNCLMheZGC8BrzU41at9gGHjq0g91VwX
0Oze91rR0shY5TEDSlRkmQFtRWga5Tx3wcnyTfSRbkn/0BL0/qfoSgk2zjWsL/mI+cmNbi0cjlBa
Xji5YqKcub0P1p92mKqLaW5Z+SQMnD5JIdPrNdHyI9U+UsdAXuJadA4VlLWmA0ZoZaD80ujyQ1oa
UeTMd32KBlFvXuoa1rM1awu8ZV0SZsipyI8sJtHpKHG379mdnockkTINwi4PIi1m7GofuFXT5Gun
3PWKBw2mummxcKCwRxsopuXi8FKIuGKvKCuD+T4hkuTxszzAG95p4M/L64J0vKb3XmV8nT8zf3wJ
goPCzV+XdtRgrWHrbgZ6MheYptRGDIDv4yqxnddlFMoDVN9pqaQxbB88Uqjz23+kdG25FXN4U/+o
uotwqnD1AnWxWymFR35Gflc7ikfy0aVS9hpwag1cmdcAfPhxkYK6l5tXLdPS7g11kg7WBS6hI7I4
2YK6CJG4s7xlCRPJPHVfuRopFd2ihth2C1hv19l0zU0cFUpszKUMyFJl0eghYoGPig4vCsZmpmla
TauProG+rQ8hwd/x4OLYNQfcxwaD/4SD5ep6ucPqCroBTxm0iLxqW6AXJy+vO4qcIimxpvkBC9ex
klANjXBQfw/OHvq+AC+SLlauEQm2+RP12NNkmsbNF7h8bVyVxeDbFZmzCSUe+rIPMjeAS/1FMZ1M
XwYP9gu7f+bsjtETA1SUOZlwIGQ+ammpzPsjByL/3K/x8WHQmrtq2WIU5rb4ODNZmWEz637e1xkr
JxYbwAOfBXxD0aT1/Hus5gARayHwF6dJvA8uk/J54J/LNJFeqspd/DsCwJVFhzZI2IVJ2OKLOOsu
FkhRMQo8kNKPOlzeI60ICsoobLozD/oxs6/QAd7gM1OmvxY/x3X3WO9+u22UukVu1cChrsUfke7h
T95+XVxQY+XH8g7wmVSXeNWOzmlPt/S59grNlLas3xr8UtNpLiZUEG4LPk5lpgg0g6R124kvX0H+
1BdejhCwvs91lPpqScXixzRB2UEt75GAVTZMsstlbmVzi9kTi76E6d8Zv5RSuG7jtxGYh1D5yVie
x45u56aMjfWrP6VgQITGQ6nABnARUIstDtSlFN5FJqpVCHUTXtXzZVdOWpetO0JAJpWBZ+oR7yae
Bwv0/Ua/EzXphB+DGNOcJFwxZxnDdlTfaUf+kElQUQV1mXeh1xouMVrmpx7n2VzKqWAe8esAbPot
2pTYyL38aVydAQCh3TvUxWSImESMCJyxbrvRA8X611g27BN9q0BvoNwPirQCZJCvmKXMA0pT/JpS
PpR4PH2lBoQSbPWjxtlCyABHKQaKOPGlYSB4MW+jmFt+nStSauh/8Ao9cU3QMq+LHh8BhN2Eq77M
1ePl894HgcuGLzrmYHsgG3EsKUrYdpYaEZo0rHb4KI921yd0ijSFUO07T7KU0l4rxOyPeQWjVF7d
3YIq4PvGgrFVhYZvBAzsQx1RhXeVDASo8zbATyOZb62UD5UNBeJd+qVr2eSmYDR0qdhd7O3znq3X
1JxLX47lxU+flSvBfE4yl8JJLu1icHAw208l1hNkZIMaskvLq7/8pYCD8Gkx3lygMv8lZYVDQG20
dieupY7n2fctrCk6xsfyE63yBAQt08w/HDNKOfVg//6i27YRQaTxw1LFKgwpOCwWPLYNafbUFlFz
i5n/rHuo0Ij/YL414tu4vv6YoFluLBrgZS0Vp9ivHBI1jQi1MCnRrDHvPgHIFCX0u6b7wQ1HvElo
An+5y01XsOGRBSQDo0rPEjNzvb9uqenvRbo65QLHidJ/u/ZK0p9cLLse/TWipYZkxi30sfec9bT9
79AaY8pVrv6NDVoE+TH4z1iQmM8WNdDgJyRFIbVpb0FP5z7bEtwdcoouaBYroq0+dVRooFMpI4Rp
BmuKFMG9uvI9bFcLcw98JnW2yr01eK0cRhUG5ReXEUdqcRw6Se9xjbJZiqBdKGZmsYiJ6mLUq/jA
QijAZBvdAkyTvUMlgoIe6a+uFi9+IxSXyvCURW1MdpI6n58GaakkoKBxeFZsKvRGGAwS6y22yIkJ
nETsPea8XZFj/EZHtukPhzkFl/1yeEIKfiFfz5Ii9L5MvdcnoMY5dT1kT5RT/63QaZch9Hy2NVrt
4R2gXIOcEHC0Bo5ixe0Oftqsi4fOFZ+8NQuF0yWNsqNlRuuL0snvToGGu/Xlz+PsK6s1quKgaLE2
ndeUj9lVyLL0NzflKCC35rfNI1QYbfdSWAnFcnHQhcXy9fYgV1bl7Nxw74WzVjI19WdksOMsfmwp
HdWMNuHA6Pcf9vFGoMm7fCAu8yXSw5oAEVYs5o3hJ3UFnS0DmXCuy1r5NO9tHPIu1MAnUMqXxBw7
4e+6saTaaPJs7NcCNisRb2qp+HA0dOSpxkepSThcUnKlc+cYYxVLbIgTEsEdOtMDyYP+4BP4RboJ
DQy69ciaMq0XLhO/I9dq9iS4YOLoo2ECb0pzj8eBthNz/sU9TFK/tJx/5hqWA85Ph1O7M60i6Ruc
Y6arib9KHNUaWdGdXDCftbSSYfFRJ4PxJCE/ySWt0uY78Ocg0F6Tb0TvVX5hRXMkIkzzCcdmbyVp
nmm3sCu9ZHcfUNOFYoS8laFt0TWc90L6j9Tzt7jSZGV3a2Be0HdsoXRS3ym3zW5cxs6wEH4QBLQY
LiLz27FbZiJFTJsxNGcsyLexnIXWVPuyxb5UmQwqIMtgL2QlvJgzNDVq6uSR8Apd0FlLMECQAF5L
LuLVOt5fhH5MI74KeTfrpuxW/2bPk+kjyjJq5J4JujTGUtbZtaXJiBWZSBiUutO5GHW0kr5BRUbT
hU1NeFL1FYHLEHw6fBzmQYN01CyQyCtX8Ikz26uHlTCyEAEhenzoxwKjAhAKxXNEt1zZcJlux9mi
T9AkfCLSpbyQPbZRdkxzRanQTpdaQMacI+NzeGb3EeFHa849k9kCtpL5Dbhyz3Be1zvbtGmqw9Te
xX5bTpRIXwurJ91mK/NoQwZpRmTczQAPt1lPmkQ8q0WzIiHpH7lZT6WtXz/iLMUNfPTQeOb6BY5l
JqQDrjr9nKoe4emf5xfOVMBllMEeTvYZzI7oJpDACVA/L/lzX4sIarnINf5RHmWwzicS1aepFAOr
OrTNmZ0b1b9OKp0AJFemFt6xdULHlmtdp7G1q3ovlHyfPoXVVBqegTPIZr5RWeDbxSj8pQZuoH85
0xmS+jWHOCuZwAV/dpo/i+kf8xBb6B7lmAscY6Df3In/ccLoGOyMccSaukHVw0C8BIjYgEvx1bV3
AoAkxvhEY2U9GhI0TKZZP1VSujtxpZiibc0To7nZT8ZdCgpkLBOOf3ypN7ZHgJgBuDK738DEI/PX
pWfeHIn26kPvGnsyylfj8x7vbUZnU37IW+aFeLSIW3RiqQzUr7gXdWl/0+y4e3maBU9H0wfK6qdo
SKy/nKN2U3Ct7otY4vZr65Z0BJqvVV4KmgMasrj0iU5m1xG6AZIBkdQ/v8328qoKAC9bRgQ3BCyB
l2G30po7G4OnBFubXHbcwedVA5xwuxQlVCWYG1mD7mwHo6ykHkt0Fw4PySVvSDCWQPbzHBfT2bvB
S5FPhMCajntymkY99+p4i/6v/xorQl6AFmPzEkLvsiDWlTglRyr2wHKz61eE24TBQwvTo5rXQOol
IJM2EETFXI4oJEp3zM33JcG13s6YrTdgosh61cFz5YMCQg5BvdbfrcoEjtE25nnNRjv335DaPfnQ
j3M3FvkfyXO0hm8thbAhhniPPaM8YAOUpundkyfG5fdXu4pTwUsNMNqWAiQfUIvQvOr3dK6lTidI
1hub/iSPair1rOWl0ZLZfZOSPbiUq9mdjSOTOZeFaLiNXuEKEY/ZCmcInq+PdhsBU7aciWBGHGyL
MvAIl9mF3NcegdhMBgnUGCJ9S55pP3yeqjTh02YfN2rWKcuG/XnM+kckCLzWw9PeDJO02k5PhhmF
SV9Yfvv+kT38Ypuc3PA85YflS+3OgxjBhUvZYeJdkwTpERqTaUiatf6dMd8+CTMMLvlclKLiNZno
L3EAAAPm9QKVqQ+OszftueVjc0NbGO6fG/bHMrA3Sh+2/SzNwJhkQ4EoDKPM7NNiYfUoNJtUuSIC
Y4l/m77mQ+pIkLQz3qhEEIwkJnvA9XAIxGzW3IlHV3vZeIS3XIt74Iu+HZaRcTnKY0zHkKeWkQ+V
+9dUDeZ8yoCN/3YDw/8K7erGDkfV520LbLK10QU9dubVZmU8bddpj6rfNa2Y4ABFU2mRxrCX2yO4
Amh/GmaMWQpTGRhFTVZWgrJk7J9P9074hMdgSsGpAL8rbFDpGI49i/5HE1YVR/BwxzRfufBv7bRD
q5kEYn/j6gRR33r0w7omQfnwXs/dypsQrEx1dNNzz5xm/PcN5UoXiKoWSOfGV+N5Pdk/dVwZJC1o
eHN1Smg1aF5gCOBUH192mF9jN43jmZKLhOhnJZgGKZ7woLj04Qk7h439rKJiwysszdpnL6nU0Zi/
ZX2WSbE5OF8FWV3UUO3blwpC0Vjtcn9RJnU2d9kqGiOny1BbCLiSe5N8YECrGMXAROwubo7SLh6a
Q0bvlUEXMq4YWj/D++O5colAzqBNULzptgEOZOqk/k03vGaxjE6KY3YtkxjCMhO/gRfmJ8NStoWQ
zRgqJbrXF0RbEnmu4kM4vCNt42p+s4/6UIrnyUJ+9PavQG154iwtz2kXzmtBD3gyJsJt6jL4FLOZ
2sHhqcZ8suQMr9XPyelS++ODSuaSqmh1wJCv/DsFm0Lq7B+yTvh9jiXPRKcxvpQAKN0HL1gCjpRn
b2NtQ+MR7WFUYzRL8mPk38pyY2hOr7qCGRZNq5ANwzceyCOQ+VaKc0bzti3UIyB0Z5S5LVjeDHBH
dIjaedjx0/4s8OI2tUYKuvQPEVUmDwHdhO+pXEYWxsNeqxlsngeUtlmWqbyGFq4gDAJljZ0CPEfZ
kqabGULcchaf5ebZVb3V1lkR/kz4/LqvAr6bcapkVwZ7A3WCabGnB9hM90jm6FOAbfo4AtnJJ5Fn
YBAa7nfKJcTlL8GtjlSGEfFu05f3bc3sTubjdQx1G/YWHxhHhQ0Z6IVVs/xlTvcHx05bsxq0CUoz
7HRnzJHj2StOd51p6Iy8S/MLI+iKF656xnmhE1Z3wxXKwYFxON2m2wfr7eAnSRxEBRoC1WJ+xX/V
gTHXuHlFGgfrmIP3JNsafXETn83i3/eEMQx1WfsuJrQsY6C/nKLSgJw8HArN9FHQ6/+hBsbbuaSA
jxW6SSjkyb9+v2LUdQr6CbUhLly1QXuXPFKA33aV+O4GI+i/cV5F3qai9YHrLioehq0Z5qJ/zjI7
8kPZcVAnpkx3DtVhxTcgToCu1MuOKzjJ0dvBwsDSZnMVShQwl5MYVZvQApd+3IHymd3cBmpDdhqc
6YYvyxjdKEhGqk0kLa8mU4xyUqql5qYWt+w1lwPxmo3oyfCd+hJrJjeX1EynIBsChu2Pgtstzmi0
lyzvveLZBoF9WVGGPe3S4iIkhOnwD1C2a/JEbRNesB7JI9WsYE34PlqBlkg2RPDfWudlVkXO+KoV
Ovww0uz2V/tAle2P4nbknyXzwEeBO/xt6s46sgd+gN/6UYO3FkALgdH+heoLcwyzqAd0pfUmfivG
57Vq9bBvT8C4rcOMJwpfA7jLl56sITaYLR5DIQyRi7EamhA2AWbN3XnjgVYj+YjGgQjqYFu3vGFc
a53EqinAaLFDDGhOJRmbVEdshDqUcYqEd5OtpchdZF8KyZT0YIZ2D9j7ALD7qvz5yojEAIAJiieo
lXC/XMI00t3f+hgqJQejQhiUsVntR3cqsrejfmKqiLhv5GPP0pNewlawvusIJ+VTpruAogHJbS2B
XHhx/EvfGOG3RNhUzDf1N23oDuXV3S+f7O8rWd5RnNb9NYtCyycjjtjRPJVW2VaVqVEq7JPUxy11
se+u/Lh1F5Lzc5wMmpIeNJZFRWDasSPxmNyXqpg/UpLeiOfVlpPV5GQNxl7he8mP2VcYh7ECDG9Z
U3XX13R7Rq2Er90T7/MQz3qU1aTA4CatX50Y6ui9gvY/KCdN5CLSb7hTdIIVSlvVU3AD5kaAnoh+
bRMupqjexJ2+Tc91FSTwvmcjj53hMBcTap5S2v41/xv5V2bbVFuDJjn+Av76/HUF0DROysCUMfg9
Cah7UccsR/P784Q6FIcjFATawrH6N66X0wEzfBWqS/rvTB0Y6YE3pF45NUMehat8UpspBWBPJIeH
mvXSB0Pe5noVoDH+Xw/z+6t1REu1NJwi338UCDNqB7Siy4usG/zTdQc/7mI1TrILjM6mB0hH+Ig1
WQJwhpB6I2djfuHhJYMuFs1WIY59gC5mSC3ugjaBV9HA2OmoWMWsRWur0PzgHlDryQn7onoopXau
n8YM0mhkgHTkODqZ8HR0CUL6LrGD1e0Ztk8IO2ngtQEAQUrcB/e7C//lqmO8+Dkb6ejfcwkMiMDf
ZgOduSAinJ3SZ8sHKFNIeDIGbUpe//C+Q8fQww4hCDZF2ChUvPknRwKSqqNgyzjPXr1uqWZo6d8y
ObBrC5KIzRPIejQR4FYqEJpHAzatfBg56BxPu1WXlu//hV/KA455wxW+Ji1CWVUcWpFRzUMfqcLJ
mOeyoPQ2v3/iYDAyWVr7H+0mysRdpS2paOQggwWUJpYI/Vj1xGSdh2D0wTmufYMcuWaelw6jIC39
ht9wHVErwwiIpebf2XsoG8ruWFyAPG8b8HRYpyVDUq64GXka6Cy8OF93Q3jRkbm9FqHyaXk5bkiS
zqa3FgSSKvM+Kk6ykpyGAvI5BgKRVeANbM+jE2L+XT/YYkxgRpGiPdDfryK4MwXM70oXcJ3XEf8O
j/B82Rw8unPTA5GwjDV6H1gKma3jPCjcGangWYsesayzYkleFVqooim4MtFgu/AcWTRfv/Zi0wKd
NbhJZp57CMvxUVrNiRal4xH+fcvzBU3BQT32TtEwJt3uSNNIuIQWkdCn+ivVuN0Z6orw53uLUw0/
GT1xJM0hh034tuPARyocXuW7dEF+PVEp2BQCX39X94yEQ+0a63/qc46K2qLhUi8AmWK5Vq7oAwdg
1GvDf7hZFXE14pl7CdtxyWiyHTLKIF7O/f30ufSSNW56E5Ml7QhbIH0We1R06Wg4uuK6ER84ECzW
yVr0LzKv4hWEv7mv8n4jrWyz+l0/5jpcS45FLZB2Zfxovk93rS/o6fldPShqlzIUsrMum6UQ2WrM
rwwB4kkJwdcJAfd02iyx/2gS+dcfe7OUPgwR0bpnZ36kdwzVR4pCOLZPL1cLQyUhZtN/B/oVt7Ut
1PH5skqaGcvwgNjEAOUCS3sapoJGek9HrlqYPxpWbVW0UKiWvHVSlBOagxy2yDpNjbSR3ychI/7R
HecfNkfd99B1Hrd4Y8d+MH3SsejfZH+vfsnmwl/eq37xjAXFITl2Liz/wixRoon2pVv7pL5fgi2D
QWT9AlsAax3aeGkO4zccqDpm0TZknJQ+hmlm49YJuBzZLWXhXapBT6t0sS1OkyzhCFplR0RMul0U
8vTrCoFoajsj88IxWuKxOzRUtNW/OuQQ1vCSpBRezuHnGvXk2NGrIcoC0JE/xkC9MMrniDP3sYwJ
kMT81Sjdxov9H1O0byKgaU5Yk8Hz4WtRl+AAJ0qGwN6ZhyrF4ONuY7+JoYvmC2vdn6rJjn+sMr9z
8BpzB5iuDt8LDElHsKqOlFpiyzoOF02UXiDyvq/0VkKKSVibjeqTyoZthtFHBkeLyOBqCQTDLeBA
nXS9LMXPd1A6ntB78tF24KK6Esyq8Pcmsn36hZi2FMGXj0Ha0AooXePHuOfBrJI8aE0G0vgrlMZX
r7402dvHMXdigNEZk+HlTu+ERNEXUxi3nu2LviHylDA/dPWpGVQcK8b+J16MDznAIkOKiPfVw6ij
UqA63oF+Cdp+hv6pZ1zkHTyC8QxxdNg+oWKzsYNJvrQ5IIQTZMVIMBneV+uh1yyuGtt7S8bkaSkf
AYiUbE7UmL65DYJFl/Vf8pziECorjOXHn3nCCh6TaFKYhW56LwSD5TrykYzF5XGWCGOwxtsDel8Y
+AbDDLVLaRb/ifzRC75UlY7gURMUur922hIdE+kG5VEsssU1apuUuhBRNomHAPcYGSDhjGbgnMZ3
7ceVZed+H/vnRjPKURaDDkDIA8YuKayZuLGyyMbWilFZ9AL85o0kuW8CB5TD2yNVYWk2D/6PpSv9
JOc7VLqKsFJ+jSwsr4m0Q9iUNQDVZcnoElf8Z+UtkbadJorXKjKOVUdId2zZWQCbZhUc0pOmub90
m4Dx8kOKcJ04jlxsprwL4MgvAonwZ3cMoA01n+WPlieNTp9hzFVjKUCRXqFLTyoIAMB4taQwFTMD
YSwhHRr6IQsGjtI5tyvQoifokwXm9r9+YZAk9G4PbC3bYkEbomGIrvRWKCy+fk6B/ZXGUvj4o4yh
tieJikdf0o2It/XgJHyaKXBvrfXqMqUWSPai1sknzgrvBs0bJSpHcJdU5XHOpEo/2jltLGTH7xfj
UQhMr1jVg2HCX1rueOkaXhHk19UIqnkyQW2QmgWG/YpQt2wW7anrE0XkGQFctI8gOkv2IkNe9otA
NrVTCoPFLIu3lJ/AGrNJrGaw7ymM65zGeYI4AAVaihLfekR5zhVXp7TwiI/jLRKpC1OpxFDlDKlP
VxfKkaFvOLQ7PENicIeAdvfbM7DHM4jqm4XM5NqhJoayD41Md4w0mm6DuBeSr6DHj+T/gg4uW886
LHDtwiflmiuyNZVOW/eLi0BD6tBkJhkQVjRBh00oiJK9mL1JIbvvn/im4gy9RnrSFleD/RvkSom4
GfTK6jzO5PLFVh4CL9xndYcrVDDUkW2vyNAlz9IJQrwcX3jIReOMRBM7QDJ+C2YgzgJckbjmLd7Y
nVpCh4nfeilD7Ys7M7W01NTfP2A1BObiEHVJeEiOCNKILueD2Et0Red7rPtYf9tA/cFy1vkLIcy+
T0nfnCVaA7Y/7aCy6Q9trbmZob4GRxTbxKhCbk1DpiV5mXxpdo0Sbn/Fo8z0p0r6dKLWVJYd2gQd
GjKps1YKw+mEpC4K+VCZvTucKDO1/0ks0T+mGR6DNY/Jz+wndUyEVH7S5hoxH7lAsklHi+NCsnvO
+K/B+JqaLVmvVWLswWGoxwVEHQkY/waRIq6WFQBXsi5cIvsrmQS2sJ/WJf3BZ8iHZLvTIfIxJgT2
58IkpwPv33UgMbJPhSSIcJahNZRcp31Fr/JgloIClFlW5vqBLvLhk47WA3dLkVQLek1LUto8j2sR
hoW888KOjHOyiGPzQ067bCvN0tCfKMJzpeub9dBWZja1ZioiTYyYkD5bi6SsE9TXjoibIJij3jHB
9Dd6myXXKST/GR1YVTx5PMGb0r5oYusw4b74NApCIf8ju7S/ShfiMRuMvlTkAt70aPmurfvecUtq
+OFFFkPlJKxCTdevAUm8p1aB8Ze2MnfA71swLRqaWkMxh99LUHeSGbpqFW380CyUoOva7w734row
fvO5MQprDREvSPDOdVAQStYSlNigwR3+HlCQTmSbqR1TzFIl1h8k0F3rdXUL5i63iIYYZu8suGqL
czX23Dq67duT12HGXQWn7cze9BFcBYizX6l7VKcz69QWBFB4bnaaN0Jg7OJWeVUGxpejhTpIOktg
ZnwGC1rHrb4qRTln+sYRcJ52/sJPAAz/aXc870tPQY+UQZC9adYgI8lUAbLGvEWu2x4QPIxhnXvZ
9zLjqK+md2yWAYDs0+2J44gP8I2lqj4NTrdvbD25sI+ERefDcA2kxP6fFbr3e5NbIxSzLo7PZAVy
PF1niecraYthBKZ3YIYQdvbJx5ZCiSD8+2lBH5q6wiInfTWfYpJ5t12vEv9pERwxMOWFBnsW//W7
atF68OhperoHY+Go+2BZ3qjhBfZ4NxAFb9nHCEymfl/D3G0UCcGIG8d4aFDpTmc/mBiP2AdQ9/UT
nM7zcwDnGEd4C7V3fIqT9klYhKojFSa/r7t1vcHViF+Pe+hAAApkg9SIdWGPTojQ6gc8YewxT/NE
LDeOBonXr8We3rTAKa5US7FFiwjE0Q+xIZs3DIJRVXaKbWGJDb+OEsdHrcDV8usSnoe4V7QDLF3a
fIBWBUWTT4K34RcAPc+PXOn7RagRn4NrNkMYsekk9+7Bu+qKFTmQSVgAiBelhuIJ0ymM8hEwIrnX
dDo11ffU3DBcKq4/EEWFMWVmtj8oz7b3feIocRaN1bSOvmgn5WNXmYsfcPyVjCzVL0cT1FYD9HhT
Ca68s3UkFvPxCvVDnH6TGNw2kA39JWP9MSTmDn7zsMWbPb07qDkGiVLetxP+J6W1uXsU7WOWxeeF
f6XrkGms+yuOB4YEgXK9U1GMUgPAo/ZvHnoAybm4VCL7ygVQO+TnDcVXcKErI2pRDDnb95/3FWIW
m5qxR1qghEyqb97KjRz7QSBXf0+Kx+lbEICwmhdZ2lnuzb42wBwUK85wGPWd+2xbDOfw6+eDKtA6
BZrYpqAAzCZohEgJwwqCHduJgzqXPedsy/mOKD0RATI/sn5rdv8Nv6QiatBGSrERS5UiOtrXxFrL
F72f+XhGK3zH9ktxbK7GtAqHazzeThF0UL56ZTdYRmV8PJwJ+TJOPVs8OySGkFIqjbaZD8SxvJTV
zft2ibLdk7OzXFGeRjI/9RoRMawrIG4g/+qk6Dv0AHv6uuNhs598qYS5hRSfthvbCxbQo/yd2eff
qHjnCkkSZJGnqGq/hh7h1TkuLPf/fi0qUHCw1exslWIYA2OdgGAYqSdNut3JfFTliSfQJRYWMVPp
TldtRo3SqZA0ScT/Phyc6N8zBigpTCcGxSTO07Wo01udKu/QfH6wLkReB/3SOndORpUw4GGcP2G+
ohvki8ztsKy7VYVOiL6zmwWxzsCAlm7W0Zwl/ngqgXkwamk5wZrO3lmwIrF+xNRlzp9stXp/6sTE
/Ubte0QsJAc1+9cNbpL99FMXY2PfgwxZD6rjOjiNgTjbZWM+XQqSeH22641AABekP/GHCZgdnJoA
v372guKUiBA0y7eze+/VPGTQjKUzp33fxXfcqU13qeWmIhqdGv3A+xcNYhNirMrLocPzs0PT9+fD
zB3H22NkGmXhcKByOWVL1UPXtg6hnqKn6p2Spd6VdbykIcTA1MpxlJt2Y6wSmiMgDorLCJar9LCg
wQAyk9IFp5y6/Ue5XjTBdTTEAphy4QqBQI5nKPY98H5lWVap2wVPgKH2TzdOhG7UB7/VbR7PF/87
5W2m/tKw9XRH7s1kN4EogNpIewwy7DaKkiORcMImRTcC0Fih5O4NEPHrTF2stecEujqQcG1YBDy8
HZBKiIqxejJd4LCM6xTsPOH9qdL1M8LgSZSZEpjQD3OeEJjIN8P89WrnRmtSO6yA8S3KG0xp/HEB
4CVA4FSgnqkHBXJJKZyCSZVrzM4vq7PQVYSG8lYUjxNzeGSj71L6r3/m8x0eiHvyzZNyxOOZVAgt
uU4RYGbHeRoC2lBzIugaQbRxrrv6RI+5Tf/FjFaTsp2lKshCeXYuV0BGyRbzVfL2IRr5u7B7gddN
8tpAaB5yfXIt5mL9rvYUGACdny9pnOWbtQqIT0aqs5T5tblLqP8xu8jAnd9VqItjVmmgeawhnM7t
CRHJrLue8WFY/g6asqj6UwfgV+Lk2CKKoPQ3E+ID70EBYrpPT/AbvpdpkY7vvJ6NllHxAExXWWo0
zFDrOmGOMFbcfC5Re3wdeUh2qWMByjxFLqHJacvD8vZOMZ1qY1A1gAsu5Sm6dEHwXcuKgwH3LbJw
O366ItPuOb/OyWnajzUXjy/bzhBRpft7DFK0kaYWkcTY8w/1RtQNpEYQDprXDVd+syaXJoonVZj1
gwO5ojuHETeWFBJibQLjmFE/rzfXWKCtVf7YXY5/ak+34LN2D9aWp8wQ+78TNBMC7+XuHkt5aI3o
7V0xNBi0FsSiVEFzlNvj3W39TCgFxHylK/jpdbFTucbQnJ6b4sK40vBa/EKM6wyD/+VSwXI4hAeL
UruU50ZqbysCHDLTmq32YnKg6A9mHmpEJQb2BYsStC/omLJBdbQXSCJ2XCkgoo2sTwtEMFwaipdS
TwtCv/4MOSm63qEgd+nVkhaHtzQuRRJ5KdUzS/ZQFFw8Of406KpDj3YDgp7JSkgAxesLiqeLz0QG
3wOE12OpHzBkw/Fahly3WxS8oFREyh0elkZyGgDIUzurfaYp8IKbMOhymz3r/aSX0m8sMWDR2hdD
Lts9Vci0lwyHstQz0Csjf0o7BRVAhPihrxyIeySFeiZXojhAQKvMOlsqq8cuZe80Jexdh9KEq77l
GHL3robVMS0FXlOROLi24bqEybN3p7pb/+ZGG3AVQCicWE+JypN5+UFVRNG8jsCA5ns/D6pb6BbK
olXhPNGFYGc7kDvis+0xH+r0l0axAvE13u9rvTNgrTTVoD8WgfppJO6NHPuMsqJ44lnZ4mwd2jIQ
AP07HwjG2LfnRNAU09GPWFkkPVPs+NB7POdxTq/DP1+/rCtN2lxBE+mTf+w3+/q5X9YNxVN2iz6+
zjoCEjVc6foCFi4ToVBoYrtK24UGExTqujCjGSUYa2bFETasgF+PBuXwBYPs7cmzt6OqJp4eLKg+
xbCIZFPR05KykqiborzZdcs28zTvuRs+e1zEdpdTkbfnopqimCtfDT2Bdlz31CS1q3OrR084uSRK
54OWxyvgHxOLpEduhQ3yNwDaYQhxe7Xixe7Eb4/AoVaDUwW+sriiw111rpIUUNctuqB+3uuzkDHj
U7eMTtL4mVYfaEQYh5+KdCErRD/NRYgX+0gU9zt6/WAkr6102x7S4EbyajVgljLQdq+D42rR4TXu
4vkJ997V1RW1FM+S8/xhco7LjcB7Tk78kvBngzkS2Q1UpuRymhN43R/13Mh0b8LFTfRUUjZBqZzA
/D/WKDv1FxCFLacDKTjMDmDJAnRhdtilM4Aukm41Yeaswcvm1j61apdhgc7KpnxSZKOFjMpprDe6
k1p6uLubilE356yEHg1P2oOBLEeieZ8BrV2Fg/NmayJA6WBB9UmIRp+DPkGDaTgBCC9QBsjdFu/0
4mKO8mKwkMGjZ1K0hSb2njnL+hbtmsh7yTsf/AdFPD1oNTq3lEL2bnyrR+f2bKQUHXAbEmhoiNiP
UxrSMTIVXsyQiwZngmIugrHypU4ANREenkq1KQN0vKA3SkQDhRrdz3j4FVuzeGtDgzkZJ51IGxJj
uHUcdWvqz8xkpIq0jiK06tK13IY81bQKRGodMLYLtYMDU6Xr3l8UKOjnyFX9LO4ly4VnCl1kDzJx
BPEOeUSnYu1xl/9G+0NL+QivK3K+zPjVn5XwNNan4/KxpG9rVijk/UbxxHgeq5hSSNjke80wqeYh
hq0OhAkx3S22JyHPg1tKJl6buTaLRExxWZmuEQgZ5DhhOINJ/P6sM4wa3eBvVYImkiznAaRLZ6LW
V3iLkMzCx/dNtqS9MUPmm3mIZ+N/SNmud5y/IJGD1fBTOAFSaYlv63EAc34lt3YYHKPNLynO8QmI
k+LpaTfieZVi8NKFChnd5bctyvN+Nq9LberSjLpk6TGviEw1zD9ZHPIys4Sy1dfctS/i7PS+MdyF
igh/qLdiyNkS54p1Flsb1IvLhMWyV1SJu4Jp9GN9ZdFNCbA8nisljVG5+wykTt4MnnWdG7xv2pCZ
pLL0klmbjXjr2RalhqIOYr0cHkwZILwQhaXjclIexJ7X1i20cjmxIBqkTM2LOghCG38PRKIwnTx+
FBdcLW56/in6OizMPZN9N8FzmbvkaGmUMM2pLwv7+GMXwj0CFpXUmkFDjrIBYW6C4nOVj5eN2oG1
grOFVdIr+OYc2EpU8STKiP4DuUHRHZSfMWozdLrXPt7mWf70Jw+LygGxe9EupL8hD2f0nR/L7K5A
6sm7IrRXxExkzrduZyfY0DALCF9XwBLDEql67VV0D3tpfLeK8OUd+GIGzKuS+2pJudSUxGAzoLsL
x2t0ZN2mG6DBn0PxKqmRgHpNdOeNAWWbKLjIIEErY8yjriSNxf+Kbl2DUlSf2FdQicOMkmIXswHa
c4grheIUFlpjlsUjSCa9ut8tR+gxVZiTbjXOFOYyikKpEYMBdx7NeyTYjrPVacxZTrdLIxnMaXeD
aec3BG9WaXqBDty/bDw42D9dgqA+wlp+v/xmsxzn9Zp9YXdG32JIbKHg2I5MTV/lHyJn1ZrWfvh+
cnwkipzhZ01qBSXJX3GR63M/Zkae1YsX7nSqc+ucGmqq1rRsrcvFdEmYvMYlIV4J1AHLHCQp7+6l
u+VrwEkJEqOig/ZXs7xw3siNgyPjS0j/MEQNAzt6YksqgwztPvSG9vNfy7htx3LVUt/wS9xWHDdO
2oL1oJYeb95tUCtsC2MpxKBNSmlVm20fBPe6UUfM1yZc4NCchFQ5ggFH9psjkhVrSOkRQpT7ypEI
9A4H6BOq13gmCe4HxPnKJ0TmDFfdqOXQ2XtLCt9s/+zRuiyipwM4y5EzvaoUM0kir/3XdpKEngBb
upDh8lSAGLDt1+Xt4hJStrvW5oQiONsD+EKVp/5Dwmu467C29e5GlDoU+UC5M7CsBMbYOgbwiD5h
qnnmfAI6LdY/B9HxZtbnFoY8fyb2qkJWBtHr2Ma0EyCgf+iLYlfyv+omGpt98djVXkBvmkX08yIQ
2yYQrnGaiN5x58CWq0wZ+J7bXTufT6NLqi6Lc3CndmTsj49UDM919Wi3qJekMuZa3dq0SgMmLyWj
AVsmlkMVUi18azsw6UUVbwY2jRlSezpdyS2gX7XyhCGbKRW46C7i0umphoEEDQzWwXfTuMYODYFj
WaMWUs+rs/PQzi3MU4R2t01HxCh5gPFG5HOdwAH+zDzZLkZpo0W6n8GcEZdi09oSaEqq4Tw2nDmx
CKvhE4VSDz44UWsCZ9/X9r75pOrLlxjM8rA0aiplGuE4KZ+jPGxPxaGPNzunAsPgRFEeBLe9TnC1
/ZGgKbZ/fbvwq7V8idqZworZ5/EUObCYAmvI9WTOwPpgU8kkDC8yeFhcH2VRBBVF0sUX0GNNFPGg
tuPJvT5O0cpUZRJ7VrjLZkcCRWyYXrtKKE0G/0dtn+oxagmK2Efz+1mKT6L97nJHapimS7w29eRe
YqroNHH/HRTjIsyM4ihEIKprq9iXCi7zOJAFrgyeKU0PNjdgdpyoOiR+Ft1CuriNdMSSflBdbTVO
f62zZv3ivyHQsv4drC4tLpsV+m/VmImYcFzJnxaNS9MQ0tSu8/GzcTb/KvM0gv3VBIoeJA3i/gFD
RbC/Dj7mCkrpz4JMBUd4LYqk6ZshMxQJRmja+xitNZ+gQuAXWDE8uTxVNKZSlGndSOeEZ/29aA6P
l2sa/D1WOJWHvgRbUTueUiDkHAv4YcBjBxhNZNNI/gVf13xb3+Hro5tWeVz3pA9mHIgubBdNNH30
U64+oYpEsBHpn7LOBbuLgR5+uUhwhkqhLGQYQhCr7SMnbxRQSTQx9ww9nEHs2BVcbjzV5V9bWoIP
MSuQApnromz7yswOm/vPSIiqWuGyBdUAIke0u4nvV/ttD/UFdOXMOuJfEG7hlsEBrtyTlptqVn8C
JMfd8FoLmEjnOpHcEgkhZMQsgwiFRtVYQ0FDa2H+No/eZrUJxFvAREz/q/fEZIkexinOp7dJQ1Bh
atTeVN4AQZJh8zW7vF+mb9ODoo76473RCuVn0wczjv1PHDZPWbIHw0yz/U20sLIq/S3AtmSoC0S1
Q2Pl0EHtn8bccSnNhJ962ubSv6gjjPdWZ9cU3Nvhq9x/DSfb83XYV+9JhyAi/jenTcPFAjV7VIxQ
JUKvzNHqfJ9WCKagIt1rc1pNiScjTAhtbqbChMayR4/4QO5FI9v4maA1MrMpHHToifypS+oCyEvJ
bhDS2FaP5ESo5zPLgLTgZSOswjPHdVrtbHmnmNvme+JObf8Je4aE/JzL4nBBiUdLO5vGMzxgxT/p
9T/huwCSSSp75asXAS+IpT3UUtGQVslJ4oiyw1pq9COmhf2yIKLmieaYJtt7kgwZFlog+VrejXhP
NtRj8QxHaW05P7PHVaRoguoZPPmX40xQAoCRIOHuQJpQH2XByM0Sgh3SKhKLl28Z9No8lmm+3+sy
lW6I2WYWT6NBn1aXG6UKyp/11zYVbhFt9LL335pHH9x9Ohcsnq0/3/pHZxhmcVIT4WObsvJstLvn
FRvYO1xRc4UEBhscbIFXmxTZ7JBIZge6CslsHjP4Q1VnrWKBB16VxY3R655rL2SuOeegFdIm3Aij
uwGAsfDTg2Ro1yr3frG/3JVhLo+bSqUumlbKs5wFBUDr7TIyFOySiBfae5ip9ivG2eR0PfU+vNED
oWM8h8NwAvvfE/8XTcjdD3AboH7jDou76KXFEQdQNtOmfKq3+AgV/F92AdRJeMpSCbcOy+nSkAeD
QDwbzSAmQtwtjGHqQkqgmhVXe4OevQbBkUAdAeaFUtJk0e+vsRtz9j4JqE6UhtfZcT7uvj/SKTOG
PUOUVhhizTZUMCr7mqSd4sjl/qSSrn/pJJ7WvBYs51/vlnwC3PG3oP7FP8stNj9G4Cixt6rwP7wf
rKfR85qAtoldFIvkVukDaX8liIe9IhDFRpn75/jbbFA1F8GvGl7GmSlaii2AxnyU/uZdSlVRoPaI
ZUECUheEiyG6Dft1N0zilwry1NKhgKVzTjrDYB6H1L5qYFgwvWP/MSXyphwdizlYXDtZqgH9vY39
DKYvAAbnDCR1xckGGAVtrgLM6Uj9iD0Fri+kPaNzUSdGLrxQT9xYLV5dqEGbs8p06qUSZFieqRv1
waTRR/aXPnMORCguOp67Uwkz5IBTrMM88hMzwOiu8EI0sC93KWaapHqnAXdhYU2NmLcGouOU3LBv
S7mVHqpjejKKnEAeXhYJZpeR68fT+sKQhgkyoJNvcOkip51rn4gCExVO488PokR2dCoqzUYB0qPH
56JyDpMaD+Bir7NhiawLOtcbLZVScw3k1TS8RPBWAh3pAvg3UoGwzEHsSvG9BrgwY2RtN4w35nwg
4pR2xNpMi5jMLXT6WVni+pKSDX7EZRzornmEWx6gGIj0ggGb6Kdj4EB0UA10FDZC5mqKsk2ZPwUZ
CfdmY3KjIEbeWhhzH8q/FIGfMvK7GqHEXZ30FrbRG2/pLrC5wdu43/nS04i/VdyLAYttxBxDs/yp
Czfph8w1HZ3OUwMnh5DB7fujHhyY3X07lySeITmdk4ve26VN8nBLii6qr9obj0GGE8tFf0/xG1+0
PgtOjvrgTU2rESVOtZG1Jgv688p9r/m7wEEiPpSt21if3vETO+XFcKIfHl6xGpIvkGhBOoy1xUln
sBvSW+g1AB60V9kUB2GiMS14HyjMy9VKLTn8ymn+mdTXqvC16Lc9/7nMpJoAZyHlzjYr0YZa57Vh
yn/TcMVtlQYTBEf90rACTzbcl2h+j3KRcmWcX000zgrSQOuwUAJnvq0qmD03sRtxWzqdiqCw5a5W
X8Bjt3+E9UzLWrH9apKmzq+DGXuhlIJplm7fEQszRPgC8asqvLKpsYXD2aTk5E2AHqWSK5Dj0eNJ
QMJcoI6qxhKdMYm++t2LgWVFOx+9AC8aTFTAoPdeal4LqDZJIoGxM97oPJIDw0qpDi/qQPZmsSts
I7VH9XVZkn4K82AYOkbmmPRgyNSZiT0/9bssIt2wjVw01ONm0HEaXbsbf6PnD1VCNijzxeF6oMWF
RSl+maJIRKvrChRZz8fTnW3AHHEtECvjUZaU9UCww0BdesF+XT2SAp53lf7hDTinCl3OUAVXytSY
Kekww1+7ZLxjh1bFLhqDlT3kz91nynVX1/8NEURyKFsaf4WcnAl5TirGeH5qAClUrtrxkA5ZSwFk
3RdwAHFTNX8v937331IeiNH0ss6l4CKuKJ6uZv0yB/F7Kj72KGri1VBuqu8KTv7MOG/gcx5tZgj4
VeHbitDv+bBkED4sREHabIqLMaLpnHwm6E+6kNGSpqiEJaRoBhuLFuhTQHjqoDRHF3cbwsKxD3ip
HNjNkTyU+TJdxyKGESYZeY7MlgoQfreAiKNw+h/RIN6+WeZ3wvxp1snL8ZHA7aITHE0j8xkK32El
TAfcEw3cGVBnbQ2Khli2Gqm2EFExQWUlnw3oetepQzaHVFBOfY35kK8LEdArSspTtj1SzSj5wajD
GoCRV1p9eYF8FK4jgsS/yfueaOdrr8UKOcbXA5kEUmfwdH2r0hG9y7ARkjUA/AqE3mpFHRho58W1
g9gcYjEFoPtM0vMcGYcsXTnkEjvBfLERiJRaGAWUJpvO5r2If2U2iDnpgzym2Tu346qV70M9PJTk
NHLxKMKQsBrO0AaOv6qrTDZBghOgqoc1WBkxdaeYR+See1VyHhRL4V+QRF/JAf5updNJ/dd/h2Q4
8WTmvntLFhWFWRYxc+Ti8eOUeouZpXjn2pu8sNxGYh+XBla0bGB0DeSBb16gjOWcxbzOljGNPWFN
xzVu+NTz6R8CFCkTEgu4oDVoVExZ40YTS6Jim6fpMCesXUMIj7pOdEsAxpFIpD3qiNAOTDUgs0Zx
oGIHpuisO7YYoiUY7pbHePKylMhHYQBfv2chQNZDWGKyE/OQ4ycfZSgvMUQ92abBEoG8nf2JmUd5
mKcCXrq0zexlVlGv+9pE2/xm0fD88tPdoozV8WdGUQ+5G51r2ebse3U2zTb2+wJLAxyetJa3nqnv
tEiwjqtRCvwxLsbzpPxFDr15cokiy0DEJgQYS4tWPGyq/GnazZXKuEuxcAnAXskzXQvl+ONT++od
5OR/+Op4imp9PQ2yaB7GU3xAFh4IOpMGgYH7PqZM4ZtSmC2osWR+4QbcnfCP+LpvDJAFOjus0uWB
9ob67aq+KSJp5kNgHhcE8FvK4c9cyzdIBGPcU/1n7t0vG2OjRoWe1Mf32rF2EcxTqmksExGMaF2q
T1Jatk3voJFXu/lxQuHYStBCEbDOzALJ3xR+NbvgNQ9YJsrsfJProcomosepzOYs9nBJ09uEbogQ
5Jzie7tjcdQWZpAa088hSm0l5217NrtILbC4QKr2PIx9bW9OYMZ/5OiQty+//7fCiKPhIDbSSFnJ
SQjixag7Nv09ilHN7jXNTf+//uk0LY2ytRfwkKeI2Hqi7VtxpQKMxcvCUhqsfOQG2NF7iI5GlqqC
JBZZIcS1uyXAmeTWKr9vRSNRJBIRWB6Odd0LardxyHs1OXwNI6JSWZrA9sf6FqtVb/VBHiFkoSWI
y2n0dJ8fruXcEEvHY/nr51/yQyTJT55JqZqnPefgNGpGYHHszYOOjFCwCwevNyrQoWgOvbyVrzzR
z9rXo8e4Ggm7oMZRcBfPC+8o7BcAhMehKomGOwuoum21GEasdTP7VlLuFFiY8lcGBRM41Cuw5xxW
POAKKl6suXWw07yZfikxh0DyPNwihuB3XLRWUS4LM0zl5SYq8zsnW/I1tTUxaR+kBBithTIIfPt4
fIhz4+aDjWmH2wjcXaFS6WK8t/ksSGO94Z1IxRPUj6ymMXfQ62UqTkwjdLy7M8rOE85VzcD+Vp2L
CNbRO6u6yavrez3R3QMtkxtTc0G9YCSUeO2ZHybxhqU/U4Ggs9MJKIWywEJ+p3irpFv/C03Z+E+S
2olR/Rzyng4oSIjMvJeEDcV9Ag5M1Y7mnbsNv2GeJRQZkje/cK0pOsseJLvmMiP9psSq06kQwKza
EDN9aQqPmEhVw/1Jb4d9lRkQ8+J+859Dpe29eJ2zvL53eRy11UYOry8qOvzp6akHFr1/j1SAwzfC
xGzu+6x5o0IKGxsGiDFXT1YBPbRSPJLtwqW4UMRwmLcGVrjM3w2/BxtmqgLo4a8NylqhvpxtnDW3
IXIAIoPevlyQsa+Se2LzT4odtJmk/fyjlzHenfgQY6ilJSL49e9x1Te8ZYNR+HwpIOS4s+hk2ert
l/D8E1AENbor/Wf5wsGEwpHm/pW9FBIraTGB9CoKLr/+50Lukk73BybAdDlW/zYwlAVl34v4u4cr
7MK/SK73t9f92bU/8COrFoe4ut+m3u3llyYcMFJGRk51E2c0fnFA8otUzxTZL048DVPN69DNTemF
+ME9lLpD2RMiYvEjm05KlLR3ij2Bck1A0V3qjeud2jMX9J4xhaleQzSX87FgPG5f33iCzOEddpae
5QnlIPLX0vfwqIX2ENynB4i08tVq8VpiE5tVAbpixNFUl7+vqC9qSpv5dqSn5WwCXBwAgYrRt+nf
MAY95MGM21W+3PPryuzLr4k+FsOB0uunSySSqLmC4s4FHINl1cBMCPUgNdpFQNp38UcldeT5OHHi
vb+HMSlXHXEwmOAbzilCrBzLnr6nkJfOMIpNFur2wZObCLILTGa8P9/pyUX5/iixwB8L0Asnu+Fg
VQqGJOYtHMd8eSO7/OmY1sCv2qSt5KKcCiLZiqd90xbe84OcK007yKy88ipWLBXmPqIP+u/+bDZ3
mIHjGLZ19IYJ70/VGjHu593ILS7RNl0/ADrDkplLkNhE4N6aydTTga/DulUlfXCd2wFup/JXs5jf
Fp0uXqHzY3WeyckebV8LRs35zR92slqllKi3mV/+rvtB5TYvQhK4DaF6hkZAStikkWfCNeMakUSo
t872oxvnd5+UXIi0eqC9BMPnUSS+9jXA4sBHVxYYw8gToL+3tJuMZKBuc2DbWW+Xu4XfP9a1N4Vd
lFkNCoVSN96XZzReOa++/VvDEat5tzEMfLyZxCOJT6AHV5qhEwJEucm/EjFXDkUtAYeIoZeUpqdP
Asd1TKZJ5/jE2v/bf7q64H7lsby8yEmXFZ3KLzvPy2kGtv2oOFBBivwQxmoK4Z+ppR0BeKcgSyp+
G/wWmAQfMYYhyrpfcbygF0isVG0bT12VLpKxOpMvb78KGk+pS69e2ubDAjpYmPTfRhAQMEoo8k0f
ja4H0e1QdBxDx3dhMdF2eXRg3UkopzSjUB+IggzMNF+K+7ocDQsM6I3QKAj5rU5uo2xGXitF85w/
VWctSQELV57l3X/8pLPzHVcKIIS/eUL5q7kuiiQtNy7pdFV2GtQw/QwmmiFrxM1BUo8OHYtzeK0B
olicWLgfqVPsdeL1Q7gZ5V/rFxuP4JKchi8lvr87dstBqJHsjrD26x/wHVutUsgAEDmo/0T8n5dU
JWXuyAGTyPjYCVVFu3jZAfVOguZVWS8Jj9SKS9Ckqwhoq+XpWce1wFahXqSS5Wc9sx6c3ScborF4
OWEwueswqVqoG5fK5nNNtCxqmpPJWpDqrwpFr04Tj2juTZS9aWobFW8kQyh8isZT/ic/2i1gwl8b
qeXQchCn/bTwFcPSMxWo4P22IURTSnI4frXyQNYblrgwGye3rvnwIsrl4bB7UJhm3Zlh2HbdCLhK
Gzul0e6FSqt/OD/7cU/5yhpG/5ag3a9KasFu2AM++/qLKsQXj6lpTbuWf7ycgTDsVAF0eaPUdWiw
/VTQATes744ydHPO8e+b9PCWbzAbL+WOQkjsKb9Iigp7TYTz7ty2lj/Lc65QSjz9tyOL6n7jccSL
/Gip72xJCG7sx2g8kHpddh1E+gSqNWy8Zyehi9oysvVr7lMomXmpQyhOR6NEcaj9NBEZsBIIDHAF
M3EcGI9RDVKMNb53qXAm2MqB1zoyg/U58COMW7sUskfdV7Vb2g67IUkElZhESBTLEsiFN0ugfiq+
JmIktkou3Gbw9mIoBoxqyo6GFebm4ZMvX5gPm6ZXteClMuWuDYIA+ylTKqRBc3j8uX+N0fK/3R+Z
YoLwIoGYRGar9hp8vJXIDQ4+2OFrnPX81CiXX6ueiyktM5kZYeSu6EzR9Iv0qsDwMjm5umXKX3/V
Zm/2/LpUCX/AvLhMrh07u0qUyOSrjsSkcsO5w+13FOx/a1ertAt2lGdbMM+comlz84ZEKV/2ZmDB
AMBQzXqES0Ye0rVf21jn4Pw62Yeq2Yi19r9O1qYdaKCV2q9JhwWl35r40b97wmacWV8aPIlU2srd
qXaEltJsaugvxDlGn/QMkgGHSz4ZXLrQ8jPIAzhowLmsccfaJlHSbR9Mn9b8/ueORIzoM0/lRC4q
tYPAcNZKCOiPR36EX33OIZYPbCVWsKPqLqYz3UuQhxhWd6jRyhRzbCpQKlhjiRP3u+gCF2hwjr3f
ASRQHznw22HIy2TliLwtQf+himevYlWeDiGDUFqva8IEBgNdvC4ZUsCxgy2pw7MC7QUawH2Y7DhT
0Waj48G3yCBt3OgkaQzRa49aX4qgeIHjTiceoOdLxJlzaYMh8F3pLGe4vNtwO3h7n5tHrphmyGG3
AhgG4UcPLvETMY5U3rlipkB1MJ1v36fgTPt3lTQOnJjBIS47sKSi6Eq3r4CG89CXc5JwkbEp/C89
Qo65uB5b6i7Art66dyGNmZDYeCkwtF2QXfT4aARD4H0+rpxltsoG5XC8+yZ0Vk20dfe03XtRB3BV
sPNBQ5p2uNTRe8J1JVlFw17PF80hB5Z9UHYscGm3nJL3Lh02JSqmJPEla+dIpdqWQarSvMwQHoYS
523kWOr6ZMSY5Y//0ENrP/iCyp0NNTa69voYZvRFMe4wSbKelm9qfWGP6vRCi4oZ2CIzO1Q9D914
03SNspSBG6qJM1CAmnFXT1OrcjBdywVQL2ZLqYfieU6YfPb19dpcQ6/GSK2MSCsEPm+pjJXEMYUY
wg2RxigMvWHeP+rxvowSct5PeZmaEhAYA9T1BDxknqeZ/1LxLu0pzjRK5bupZDWwDGG1Gszp+O+W
j3OXNYw4keVezYxaXlSHwsB2qA7ApcIu3cH2jLY/Q9ygLv7lAn1pzdu74FpA1LqYr9TUsJJaGxBu
RfJ8WhQl7eM7OyjLMVNJDlTPLiL/w+8jPIWGJ1ja94u+clynnMjVrAgurctVoOCbkUTMsB/0cB2v
71quuBOlIitTFCYWiDTioJTTZqViXANLiOF56Bc+Zr3PyKtwYSgIh/B/bZa69pPvHviWOkqZIH9C
3Vl47n9pYa3PW9tfcH0jtm5vNZsWOEl/fFDHH+aCS7kx2MAdund3yUQkLnuNK+3DsEcqKwdDFwim
QVkRSUl+ycF1bN30HPLBsGwIaZw6U74IewvRdhvGGSkCWJpO87GfojnLRHNiODnWxQ3SNeUzRlFw
/YtWswiNSgz6AvJT8v/+htjIdM1Cbvs8EfKhu5wGOebHfWmK+EmeHraf8y8HvzIi9kpWGOolKZIp
bulTWAHqsUZmeEE9AGVRad1O91JrS9QBoBDsiKdJlYCF0ts/o8PA4/WHLAf6hc+a5by/rH7Ewrd1
UNhLQbhwE7W8CBrlLZ9jNHg0aaAfM4ADeXZvaGD/EW7P/jWoxnPn04PWIDygIqzRwnwZ4oMT74tl
/hzTdCC/07Ebl0kxboN+dC2ofQrQhcqNGFunFlyPCKqcf5w3N9+nAhdGaitSxsKhkdxgvU2Tkvwn
Ru94/ROIBK2iP8LCb2dmpFaYwYleV8Gzh85cOlP2FgLGvQMPMnrtoca1zcpkX4n9hUK4uQReMHK/
lNlr+CE2DIMtuZbF2Rt24KjcegnzRZXtAOe3FhQFf3qcihSMbwkxPFaiZcmP8j8BTR5XnVv4mkff
Rsp3as08OaZGRiK+HuhTPI6iHAmWwUE/Gd/RnUJtbBxZEXYhgphNwif+ou+zH9ju7thunLQCWDI1
bl0poitzzxxZqkkTrl4SMZHWk6pCCqcvQwwVtfiASEa8YyvrREZf6Li/K8eFLlqnTdj466yzd+Uk
QWnY/i+Yu3FyXv4vZ2JqJ8Ss/Q/Qsyl6LuGwxR7DGGfQ4uKI6ZVApZOJ6z7EYZUb3xiGDugAp+ZL
TCBzEBIoCZKiLnY4nNpT7mUE7TDrs0CWbf9uYPX3f9gpKCVHnkpJCwLyN7sk+8gtxFOeb2L0y/sD
LJaNYsZGxqjyLlJIOeRbn7DDdphyo3FwGzyKO4RapY3SvAc0TZhdnQmJWN1ImNsAwiFePpAaCn7g
9pDf70pguSkmnb7qxW4h1o49TXSHlxL+8k3STDQhuFp4F5sgWyH5u2YZHGXgh3WR+vVQveKRK/fo
lbVOL78wc3hfd1mPAPzh9qIzspJIoDyMcihO2Ta6c+Lwidqc7lgskm/NIdmrCXwPSF0hcsi9Q3r4
iitAdaPdi0/+/9lrh4dZud8sauzF6inqGpzhJvjdE0mq1J3Q/B7eJSXLrLvMCsBumY5KHLie8BrX
BrKKjxN1ab6clgAa4PXGoic5220ZeInV7WRSx7SXD1wx6so9OINZOg6gKr0eIhiUM5WW/NL7I1q2
PunbhTZycvOiv1wRcVPFd7KOTwjrmt4KqjJcM7cltL0B8BGWg+o3ROC8zQuQKnRz8xmdGOpOK3z2
RS5+c5yT4PFxXZWc0VqXbV9tjv0NXrYea+wqCy2WVMd8bDd6PkPEs/bBCtzRnIhSm9qoePWyoTVN
5ZDx3Q2oQSR8GmS4E8HPxjAdud8tt3Mn0k5fpFtf10B3cmD6TjZbRIgS2zDEKL6bEv+aodGclrel
8IS8rK9mK1QkkWpaeduOSEMioCV2h0DX1yu1KW31i2N5PvSE8tIOuKngqMDdv7qTfNkihIMsABTU
b9PM5uFd5WD1Wk+KmQi6D8qHz6SPW8vTv1UfLXAZbcF/AfLlcQK+cJoVN7MpLBS9U+LVoKq+Xnp5
5OjpPPckQZyJFN6hPWZuLHmHEAkt61b8qW4RaHzdOS6FfQb3KE5FC8qwVKNfDHEp3D6W7a5H2Kn0
PG5mKd8o5+fFEu/pGut6a/Tyx9JUF476w3l7RdtqEQmLlXeOgcmoyAsnCMdM1RH81JqmA6AUb7Os
taKk2M8RMCtRVERFPxmDoZmVnAR4mCb4LeHwPrM9Y/EmCLQ8wnNNMIZuflHt1GjNPzp539INyFVZ
LPsRorZDVSzt/2XiVqmsF7EPZnjqm8rRAgJkTesTwF+3uLzvS5oYP8/odBSn/GsSZcpMLYfYOpL+
gusr8bJPHkSYYahIi9QskZA+Id4+ExJjyXZDxYFhkZn9PwRKHWICo8hcq2ESlsaGQkXVPnJOLh2G
LPACZH/oPR3LW93LhlXs+oWNxginLbN3xM0xUe7JOqZxzwYj1MYZ0aDfx49k4UF4lyksnBvkB/V0
oWfgmHVoPjuxxpIAASlni46WmfjoxTgEkHWvU9btiXgDYdRC3SmgVKxfGgKh60EqnUzwaNR6ftoi
U/XN2Ga3+CYobJwZ9WAdHundvGof944SXvG69WEuJ4Q88ZRkkPQwzKdSJJfs5TgdpNv89cQOJWgR
QaP6JD4Bfcjp35/wMWwmAE+CZRtIeMqi4O6lZR0+w/kbNhWGfBG5b4ty83ZhURSgNnlaxQ/gFmGK
DJaRNewc9GZlUTaEt4OoHTV+Z7L8yprdzN+sUOBgSXEpj+4ShM0fUwshuhFfmPBRYEErzEXTF1eO
bCYoCpSdbc0IZKbmh465nxnJueXedcZBgaGikB3BUuEmzqnuuCzOlnLlCE7ix7pFfd8a+W7xDJ+k
85wTOGRiVGmBySFY6ig01ML/bQuBnxOv4fLomgBLXrhQyN0mlNCQzpIg0FsCnyMJZzuwtWWw1xv+
PZwnROgMeoVoj1dpM6rxIu9aor+8Sr7yJqc1UX1HHcXlsfJiOS6wPy6G02mu5VSYifbpbOQIX1cO
Fq9jXmcXheeJeGada32u+DVVq8Ke0XrGXqkJNTQc5ZckEh+kESZMI/hVJDD7tUmltgcdIlo1bFsw
pAj/QUFuA4YzabnDmP15ewLj/zpN/K66KAkABufXoVOYy8pkTwexDioHP0bL4J3eHMEA9x57xeb1
b4PlxJuaeSaMYa9WxdD5Efv4PaGFWB/A0gCMhmLHpcVbnrBPhO4VDAh9LpGZd1KB53EYW4yIGvLA
m7pWY1pMqUox2K98wiirHd4yx5NLoWpNodeXsG32H/G4dO9lcrmSy0740tjJhEClfY7uXlXVaASe
LXB4tKVFs5VLNNRNIaYVUUq1q/8x01ztMDi6a/Ifbzr1ksQIMJ3vUFy333uepAb3EyjX2B9as+1b
RGD4YitxOoPZJyg4DNyUeib87sF7R17j1I5KqF7JStEgeVomD5jxXUQYo5rf2akFLxPSygtIa7gD
X0/yY77s+M3ZBNicHYMi9ibDDREUGQ9rvRsyYH4Sg/QcDlPQLyTXW3wc9O2FpsgtgXnIwQRXxyrC
pz9XbiA5mVRbbbhGWNM5Kcv8SgFD4Fg4+g7qcQ9/msGPubkTqOM5FiGh19/hS3/hKzDhuU6/LC5i
MUZW4Hu0X7q4dxub524je5SR6SL1q7hNE3ysmi7NibWhK5ogERusG013L+j1gkoUoACydsdAfX1A
133TT+yr/7DdrZDiHtSJ5PY9mF8GqsfsoCpzC/Ck8mYGguva78T/jVlRFwb4j0H5bd6DP+hZXHtU
/Wy7ImHaoqmnvVsVsWDKofaKi/dewxfRBWDTe4Ly3jgnid99gJ9nnCiCuNO2p/XZURDtoO4glph8
I7KU59VGG5Co7mn+FMpHKzKAq+oChDCbyr4krkMU44NhVjy+YIA0CW09bN5Dgk2WRrKSal4ZTbKT
8Vy3RN7dBBHqXSgvrO9GlA8OQHtcDvD1SGfrA+HjB2mCAe5k/KT3vHal3lPjJeVmaook1r9/ZMnb
m9pE1G6S3SCPFkr25dCPPA8Ap1HVOL8EDyAXZKpMRNo0TfWf0tMc6gW1IOJLUqd6hm/MqhEpJ7DK
nF7A8Lw0/dkNztdLEgPw64jUzpscylcRlBfxVAx1YlD2+N0j3NptSrNZy2hDanw1HFlhXUAWMWZS
wEYeqzxRXu2jyMKTuhTO7HCRWIMa4PLQbb/pP79CQ8qGQ24xPmC/JyBtCLXAiyipmhocEbbD0UcH
1/Xl2ekJpVMQEZF4aFFwouROm5S1UK5p9s7Dzi//aahBlRaBS1rT3Znq5jory8ifdT58CBoIAAVI
iHrB+x8Ue33ehF/FnQcBTbLk14xlUbXInwSgp/RGnRCG7zMoKi1owlz62j4nirHprfjwEOypK1dz
RuPrIpyGDWTvbEYdV4r59SSMo0zL/oVYfrXqiCVVV5/jTQiq6dQO+adF3auURdQaHTjj0R+sxKvM
eG3coFRYvhT3eU8gYYX4es/kFOPz5buZhmK3CMK/4a7S5H9HQF6B8Bd4eut60rkuAjlcz+H0dhdv
XNxpOktznL/BgizE6mqrm+GWuqjumYKJUgl7ZLPgvkfihVoPr0cAqBb3jfxmEq+2LBJufzLoXA0k
cQWkGyYz/AR0B859U3N44wWdcPhcT0wOuO/oAdLLviQfalLpTAk88Z7XXpFGlSh6PsqIM9RMNtEk
6BkOafD56929yg1gL/243RAW8uWuKS8LJpojwNVnBDZAcWQY8bIYtI1WRU3uFYI5P1bvn1OyfYHb
niiw51vw1dsT5m6Us6LLeUSOtWTabQiQzrfnHQqdhtDzF3eevhRTVIY6sfMEKUI3PfkcfjKcMVXl
4Zh+RWAshGPj5iG07Oj1b2Xz1emPzJoG65oWTYyMvmux4LbX2iuVNpRHnfcKn9S+0RBy4Tl5CHtJ
uHsp8d2p3rJhHClRFX3QeajS1ObqhF32lxh70SVDySPj3zeuA3qIcPyDhqwIqEJotzuTm/CkHQFS
VMB9qbA37mwSIjHoDpa4MKn4jH8Xwi8v9IdSvHOUTdzb7y4V9R7lUTWfYfHIvPO5FxW4W6BdPACq
c0V1h9VzQXDl6S+dNuKYqiXSeHXnegbRi9S7jRGHdr/EMWoWw24F95vk3kjtCWOOB6RU0A03Gtf/
X/zgF3psPlRaFYvxhstyZ+1c9pTTGHcCTzrT5QRY4CSAsJnDv9xo9aue3IzYkrBwrXJsnDw+9HAm
SBdYdc3Fe8vYTRviurMborNO43OfjhZq1lJZOIQOt1yqXUVr5twkyrqRfWm1vQ7NsDhMlx3IJ6cq
EOdaeg6HFRJNzTfBsPx8AUjcdvyWFGFGaFN3dBic55bScKEzL/lJ7hJI9v3VE1uWbqo3wO1PCKO9
DNNiZKu9bgNRtvqc6c60K9RyrLWKeSN6zzWjpazPOXX0ZxB9cwEozXCTql98qoXiazdIuxSc+F0B
jZ2ilYxDu9f5uqmC5CfrRb/VRP97qUSBatEe+vta3+VY4YeZemKzp5n3uZyVNYXve569FJxM+Whl
OlHfDFkMoWfdUyIxidPu+CFNAEE6Ra+Y7P4ERnT+5JSFhiiTLLFoPTAHxM3tHw3HI8U35MNkHWxj
J/tetk1wj1FLa2T7yETlZ/dNhvWGBs6w6gkmfvjvqSsV83mSROLt2l7+IKk6LEsCT6NI/iOaqdh5
3UlBhYBTd0HcfJGrm57g0h4aSNR+oUn7f8QDILfYuHG4qsTMV8OH6xVwa4eIBo3LWpDWBmiACm1G
xcFK1IzE3WwphZs/SQD4DieZOnzR7Hif/Fpz3YLAZ/XzU20skFFkFywyP8WX0ZKFRQVvQDn6L+9k
7fRM+wHcxqiZ6tacn1ElgDt9NqBnJFmxZNLky22Z5MwPpVggtHU0evd84qVHjmBVGqfLqwofdc9I
FC3NBn/UyvN+w4c1OGuTGsuO7khD8cwfOvexjTIiQ6wS7+yr0rBor8JURD+8wUVbf1VkEG1tHBom
hkXJ7nB1Jl4wEHi2NkxLHSMaZbI71iR1VpFT4zJglIIPkvgzbSL2GCNkZWgW1t5GR+yJf40V6Bdi
FZe3NeYKel0Lp4F+/kR0OfYbqdRjVySdxIT6zFTjN5IwkSTGtj/cQZmUfyNTNLJ2om0bLhIMfNE1
WHedl8q0aW6dI549jciDaE9s7rJxiCRMZ5HOPrweD3BKZjDIPeqZWvDLE8+3SLaAYENiqDx2o92W
p5aKDsH9L+xZof6PjhPSDiQNGeMpKHO+yibKyPkqzcqM/5JPAszrcAeRTMb/w5dIk6chm3Fnvoer
LBx35FjmX+YJcy5gnpF6sbiqkD/S/KOTqrb+YcPpXVyvJy79XedNjOtlGN4IlG0kRCXAR84Y3/E1
MJW0vdRJApskqAhLlIDqVU379wh/tgr+duTV61mBiTFHCsRSaSD3A/1xn1WmgznpRhi1zq5ea9At
/krMUTICH4Q5TJNAStB/quUiWX8SQLm+wnLPkgP8PJ7pi4YVQMM4/tm0ZadQfY4vngLhfZXsK511
i2pYszkP5Pgt38m2Gon5WRym0hyeZ7bElFCRNvdko4Fc90XcHVyMXgOrw2GKgyWDa+I5Y4zRV0gB
2DzFzgKKG2GGE7enKoULQmbGG4CHstq9c3A8vDeBS/H9v09VMKB0JElac2JhDiL6ofVVflJ5Mmct
ZZl3khW56CY8bFtu8NzSonjq+Gncg5lt4yrOh/KcLoObE9IKDDAUxhKr69BX2YrBLh//2Rjm6mKk
8W0jepc9oHP4MwodkuqbBGg528Rhh/xLffU0BkMnthoh2ZjKPdh4nPxuqYidxzOdDRrAgIZ/E2Is
zy68XuVTMQ9Q1k424sYqvBaYXPsgtYCowB7LQnwsFr1g+9B60nDByWL3TeY+EiP35iGynmWqYaDd
gJvo7K6v/o3xtBt9Wie3tiuS7WgSvq57tOn3TR00ScgNSzm9FFAkgVLAkARTa53go8swO94DsrgG
J9kzl7u5ISwHk0Ktrrlls6U7jmHlCc5qxtQPP8Fto97CS6oN2iVtiO8pV6Lma7Sbhc+1oa91UUXq
BP/KW0YpqxUGrLakoferlN+VTF5SiBSBrZ6PRrml2ENoQAg+GRcyyYB5EuwMxOCTLEaB+Hpsm0n/
RjrU8OYQ3K1SYqSq1RIzPT4+/h0XXSADPna43BySpf5RT9sGtyF60DAbZzejjo6FbwNqhTQU1LtS
jsEj4/DV41DqdMHo793cckRd9mleyITkMXXGsVFM3KAGBtbWw6o6n2hCFL0U9PuYmGQkGjZDEbX9
mIB2DQpfpSppTUi5E/55F4vJlW8dsaFwskcJu5jy48NSyGENrZmkYrcaflC+pvrn0oG/YzMdXIJG
T/83mzuvrfIlmlZ4392bs0UWl8CYMCn/FukJfRgDt1Qdjqhbpd0WzgSiHU0aYSCxxwiwHPywSkPf
EENFpV7ROXjwksEpKoShg7/rsjkDd6yLlPh1KsHPx88DVMK7xUGHgPu4oWCH/qUsAIqZI+py6CNp
s8Fwbx11RATTU3qpa02wwPZWgsZKgfk/B1q9GN3Wvtnaug7fWmCG5zRhpGtL17/dadnyjbPJjJ+F
n5OOGTQZTI8BOCOSQw1chGrrh7w2TD936dqO5n1oScXb83WZgKUpW4UFrl1DEc0OcV4tQlbXgbgE
zAvBlHidvZHgAc7TPPrZ5hy0ow+5bs6FzX82TtGVXSI6yBnyT3ZolilIrXXYOIxzZZEBZM4n2e16
mq4QhkVxikz5hmj7OA1FbP8ItWQvVADwa7Pb/m157SqZddck7U8ZPEYcICPhhTPAVtX8/CRz8ZWC
oECVj1OoSIFKPRNVrKPv0EULROwRsDzRnqdvS6AMNvpKTZ0Y12xh71IvdOSNM5OxAR+W72Frimk2
RBGMSBWfBaqotCSDjGo5bcEndlMw6Sl0VxNtmpxgmNAgZeCqF+Z/2YsEL893x/vGqB7kLB+/V1aE
xz+hquIt5spZvLfSIE6PndYbNmvmNU/UcaDa+F0NdGdywRjESBqFbpnB2IjGkjZLrKm+Txb7g5fZ
+GUf1GRWx5/+yd7s0PQpfa3xe1prVxHvC8vbBwy/vosacc3eNWPh5s2pyNFu3Zb05swLWZNh69WJ
rePHHsx1AaPwMfmmCiu67KgfO/wYQXEnqMuTcU5MsdjXA6lBjVrEfYtL78GfR9/zsA+Mg9Evtbkw
ly16cxQgtW3Na479bZ7dFJuBJq6Koo6QjHosedNS8BXMaPDvFrTTGUp+Y0fwoOXj62+8ZzpMdnWq
UYU8zv8P8ux0QXH+sXlWvn1QRidRJWkUqL46vEYXKPfkb+eoZIoBZBiQKGSvE/zDBiHKntPTWnLX
JnNknnblQzjwsFpQSw4SBaOjpvzEM953h/YwvThpJUKzfnWY2+2y5goPlt6X3RYwn5FUlDnPYQ1F
uPTmLb6/68MYgmAIIGKBsDNUNxwZ4gOtBYL9O4R+XkGdWF9tsW3950aBC18dqiVMjeybFr7cJosd
XwUI7fZSeZVpdSAobPXDB+KUyhCNeaaS0P9JnXUQdNqbZp5NaZwuh9iE0hxm9FMQF8IfvoJmPn2K
DyUD7CAhbJ+ImeofGpGIY6I/T8K87ElkZ83Wl4t6GT1aH2MnbxgawG82B8Wy0R65E/IyJw9NPohP
Vy4Pa1DTY7JEhqjYKhNK2lk2hVLh9BEOFQ1j4muklJTh9wWIbv18wQq3VF2S8DQqkflwzQETLbSw
5SknxUVlAOPA690+m2/95zRieITbKHLVjLNsb6gtMG1+iBqAVrH9OCnqfheDPTQ3kygMQ6BivK5z
eK1RJkkAdOtYKDbjGCr+gnIjrfz309KdXSP+jxo99GPVjWJG//MnfWanWcpcHA73ZEZuEbLqsgy8
bENOKIJYwNC1im2vgoQv/gvU9AC+hPfJsPi3uJTJ7hqnZMdJ8a3XxSlPa1kef8muyxonRaevj6Ne
Jjsa59NKswGFl0i6ttFZmC0iBcQRLKKhL4Zqi/lhHocEStm0qLiNfrMch5kpG+aexotw7QVSEs6O
ywetH5fzFHO/r9b2VT87SIOC0lpJxvFg8ngvcLYqAMyYJ2rk1HMTdMIbr6IsNgkV6xtl8yYD7+Bi
pSgqOgZWx/MpxRQnsgbVROdkYBQTXHoVUBxFexSWwkQTGj34bUDN2A0DTlHa1Z72XqFynW5iVMVC
X4NL1yOKKaXOiiYov5S3o77leU2u1kz8CHKOZ0pWkOY0h+QeZy9RzOfIsjde3CGSwgnzb2NKkQQP
AZjF3wGUd1Fzu4EewAaEexMNBQKr/XSxK9cg59+7/mqsv7e8bgIm4l9sRpZWXU7+PQr9XLKSARVh
KFCUgiZzor7IYm26PDv5kzyi80dKjYEEaw+GxTuAmPPFs0YrRKSqBk9b7MrQ9fNMJbXNz+BQbo2X
DqluG6s4BUevvJ/xM7ufi/JSGlM9sz/YEHqtfh9fhFk9MDtLDpcOChXCMys28ge3LM9PCc5LDJ0K
JVMc/AZR2CeVtU4mz69ZuYjBiHYMTraZpsBvnI1CK9Jc9wXUbGW/pnsnk+I+57dCkEL29v47wDHj
EbLRA5TjhsH+FhTVOL6PSGhy2Gkyd0vq0z9o808i8lo6k6Y1q7OWYhHJvWZtCIFozn6/TEg1Whng
WW5RqIRUdVDiYvVfr7DTwAeicl8VU0MgQXlpQ5OUdudLnj98Ls75V+8vvc54dHj39WAHUiSbOPMH
AB2vifNt2fYnQ0a+Yh/M9hwv8Dt7VpJt2nNjlaQe6XhDGaH01Z8aUBOddCxs2wvEtsIJsQ0bFFEM
ITJjLwq5YRKcxhB/cKOrwbV9TrfuhuAv5sXpQzrk5hL4M9Eq1MxlpYkXcMl0XG3Dj15TNoEeNjFu
ejNbd++1SVuYzjUtsgWr5i8zwNzmyfsEbyifK/2U0FTKRNjpmBfah8RySsEeTF0D9rbNySO2NtNJ
SrTH25xlMq5crS/ueYsu9Eeiy0SrcQY5LAYgG5uYZUX3lqvOWHLrx1Dq5CgChpn1EouD8xxuugXY
PCXh5ER572cnuzxeysA7R1wltn2bOV1D211jrM38Ynt0iE89tiUWVIHaJ/9h0KcGTzRfm/FwKZpq
FYWpmqfA3mk4ZAS+CS4YzP//J2VYdbbW0CKJQrJsPg95eogsYAaoyY6CF3jsjygCs3JWNzKOKbQz
WVYjsH3mDHRLPecvna6aIVSe2bZHHrX1semA8sDeelBls5z9BdUGwV3C0GP+BCcXtFPICjrPMIcR
ELKd0QI9lBDtSEDbuRgjPUsbYVOOwlsZT3e+iCU0zGZ/GrUFf3rvZgcr5OOxyaFYEkrZd3OuRW1c
VShlPpldqEKe2uGDGfCo7Zb4XEnsem5SO/mKdkixraBOLhRBlmamxetJcE5DJjBnndsfrQm/Mbow
1U6rMWZQeDG5Qhj7YT5HLzo8e6csFFbNb1RXMaz+K8EQzNVayCO5euX6sUPcT06VlMWsXD3nPTJz
F+ojINEgd0tVvR1UOu/9LqTagO7eI1hW7txmFHqDG4mCOtkTWp1MheWRM/Ws3DjJUysj3k0Vroa+
l3FKsg/eMIWQa64iJcM8R946APCtkFs2at9kqRk6ip4yQs+JKp8nSGjk/DpVj5pPT8pG2Jeao6rc
zAfG0zTTjLycQmf+NGVhC7+FIxPE+2rogNJcmprt2OSOxr4I+lzy3VDNdny+9BKVDlxMsDslrIBK
WPYiiNy+Cz+QBuoCVbB4g+fWO2jkyV3QcS0M1aRhQdXGFBia3EFZdZfOok3e5WDqXgEljDNVN1sH
X3OAXub4VzRjQbCfaHZqeiixknIIKRqTImKHKn4OKjyz8VX5gtc+uRwfuP3tBjAXmkNKrSs1Tl9i
Vx6h4V971crukgptl5Xqv/XTp43LTZLJOn034OA7cV5DE41zG1nl2Go3M5zNk1goFrUL80i/P/6X
M2wZ0z3qvpT9Jx3o1PRqmjEoHKw/G6p0Kp00ow0Kmvl+8brSfNw81VhbDo/usToHbzqchPTVdb6I
FhSMFokVHidfb8iGCwLdfNjlIbyBmDpJnfpClrZdJDdcCQpG1LJ/m+4/CmOlE3uz4d8SC0nuvgK7
3gn/oL9/fnIDiPpMBfPUmeL8sEnHIgd7uss2QlMR9vJELGmHWrIH0nZFprtUqgGRWTq1tJTkGb2B
haARCiLL04nZXFbzYqhNjGvtuMIHhMY9oxe8y6ig6us1SUl1BoehxESMC6QO5BsGsVIV+rl5SJxa
uK+bb7abUOm7Rt53OAbW0dKd8ITB/y6t+Nb9EKe4RplDW71be+2jqhDZIhY2qn9dZrEp9HexvAL9
eV5j1feAumuirTbGNEhfctnle/FApa/7txx6Jic1qZHVf72/BlmB2NcHIvsIjtOt68H0iXq5TE6O
3HlZLC24Kl80U9hAX9Ba/JfaNZ9HQhIKjhom+hR4JmI/sBxNo1rePz/Zv03ckobvU+TQOXdfxTRh
VKcae+kdU7lpBn+Q9TdzHoANh06Ytgfxup3WOby6zssMZvkuxr/28yzDlRibqD+WMd+pXxw8PlWb
jz+stOiY4D5sGap7ngo4jibHb8+yYtmnQ2pcdPyPyLvk4PZRdo38gMIpCpLyRh1pyqwn81SOl1p3
XZHrj7xsVVk81e3+zQ8hyJKJgD7oAtftZvkzy62EJxcq+CoL45pAsu7G263AlqrHpZZAfeLvIZTC
i2SIYc5WE8nFf3F/8apSxx92aez/3eDPshCjoeewl3UBdgQRYQWBZOIxDZtvMc7JobDlTun7XKmJ
CqsaB9UeVQ7XYR5psZEj226tbTDqzBnZtOahjerLGfFM7Wzhx4SwDBHmMYv87DGqqj6Tj4wVJK0u
X9bvaf0BFSkIEwHZXRPlf3RWyfwo+2txkx7WZsxoDBls6M7JCpEexhZiaXc/1CsH1eHy2oXqt+R+
Vh2bWBO+W//ow9kMSDjzkg+fK5+232hoOqx9lskN9+qZ2YrNw9ZWfnkWKv3QE6qnvwVibCpMThCs
V39k+WJ10BaOOvzjbAN94VRXwOqMTgRFe0Zi1WZbm8ub2UkD7CwgbOuJQ/9zKwBKidpcOS3I8Kj8
ZaIOTmpkRpyUhzgXC/lc2e2X72SJMCCPkWHSKv55ZFXCYqjYpCguw8COPFMoxg7RbR76mqiyvEqi
pMeSjOGkWxFgVgBFwgyZezUsocO/h+Kfvg1y1LOA/nooP//m4tRsg5U037ZMtBy09t3x1yuPJ0cV
SwjgJPD/Lmlco3sP3jwfdA9X5jbU0WPJsrix8RGhLmC/u6ywIbyaKIcF925Lln8zjb1EJYu5AStn
rVq1jC9xoSZsLOKf/hY2Rh+EzfGEO8pNEf8oVA+qWex9GINWjiKPE+dY1sR3m4YXxjNHMykPorxQ
aWAoo4e5gBfp4mZhOxQJvdWIxOlVjZZTYXCjGr013TgZiaN846gCrEfTKSMOaRUzs3kJigLlFVwa
ZJe4lfOjeWcNd62/qJY+QtLLhb7D/wI+auGjb3R7hysB8PMKH8lnhesErf2X2QJqG8dogSybeAfv
RfRiUDspxmLOwA3qyBQPbrDyiFjIK6JBWLkqwAwzQLTHjFN7WNkvVp1x8tS8jM3u/WpKYMlYXqsx
mTc5EGJTTrCThPXsUKAjehD/VE8Xw6f1lT4PjszNe4cESbkNRyZ/brYYXb0TdiBLW11LTLmLoijw
xRIFA+r0Rx6FMJ/SGZ0CLUBL5uyM0UtRnXi+6z+YAEnGnpk1WE+cSGVqnILjqKZ/OJp+JzDb9FkI
hzrXlJT0LN0nYoM6I9i+54Wsg8qFpDBdVLvJ2QA/jVyXnV7wOEhsXCfq1ma/sec8MFOBJpirF9eV
Gj1XnZaTOxkRhhh45bSl4/KpRmZyw6BjgwlCt29k6SFve2YGSsQC0+gxQJiqUkrHCYMPgfXFMYF2
X/LyZ7nDHxVvvTweQwL9smqCrWDgKGnWXY6ggHUXLE4O6r8LeoLnn6JT3JgAxUXpxAVeP1/9K9ae
MQS/dLLq2mbKK0f5AhsjIZwtQcv6GxqSs2G4X42ws+CCRsD3EeRdMUaZN5pKKjxPDJNWMENvCJKt
GjC28ABZmDCEp51hy8ZdPuzRP7z2s0viRD4whtq1NsllEs1Gc40gPHg+neC8ZgOuqFe6yxdWbLyS
T27HU+uX2XO8GB0rMseG9fKHflZ8BEMyw3MOteUN9ivVc2LgIlrd68nXTUFdOfykL4VZQVlpzpCy
pm3s18VTC5P2Dfpdo18I0uk9g3PPNA8gCRtsUdNMZ9Y7R2ZM0sCco3Yedxn+gtxqbROwp0IMmWTP
sNBizz1dKHJ2+rYu8bGqk1my50qwExwIqtOH0O+LLEei1isp3iFlLulIQ7e+JmoQf14OM93R14VM
07Gk3tjOqV1WU+aEqemB3AhSOE2VNeULlNIq05BwXobG0P3wc2Ir+S/o9z8fWfE9sOIwEfVEf7cD
XFyRi5nO3y7C6eXlWJRh2vbLpjhJ0cS/odj0zydLC1NVe/svYnJaNJGmhysFYhdLG0f9lwyHthtj
N3iTStkjVcwCJn6iM+UVRGTVdSlmY9WLsJYEQ/Cawp0V1swhm0DTwr0lugi0qGzyCRrGw/h28iCg
rbgytxGpExqkBPaHCbJ0y2nGbwsy7eIJ+xNioVJHexbu6Yry0Bjh/0Abw/VaWRXSdGp9hzkvB6jk
k7keB2E6yQI3X1K4ja/bF1+NLacz4E2+NtQZ9JlqE8DXu0PGgZNUvR59a8Suyu8rtoO35UFf0RLo
ReUHGPpLVgU19DQG9mwhzLwd0AY7Tn5M9ah4tYAPKDKN5vvLGRCNsEw/pZpb1pXWNk30vZN4by0e
FGHRsuyeDnRoFhBHikIpZp0QtC5svi+Cv3+rRq/TdYTVOrtDwZF3vCOCYzKGZiqC+Id4H31mZuCT
ed2I1k5zRPcPEh6auNZpROhiB0zSy/qnBpaKomdUza4n5L+ViLKRRln7ncQN0ypCsAqFPSafddgJ
M0fAkIsyu+JrkUlGr9l8+VFwU7BYhxdWS1amnFc4XGP1y7oR3/uN6Qgx4B6TQAYkRpZPEb7TCI5J
Wp5+2FdG2rhZuz8yUwgSz9LoD0E1fHCdx7GycAk4JF33V2eGv1YfMpE/u8t6EJvTTyeteI5w9w9V
9GUx/2YZSkL316oj6itn4+ggU+wW/pX7+G4rnwWL1JmB0g+bc+b0kHfV4Mz1cJuz2hPFbJs3VbVv
helBwkLLWoWJtiK61vWrq/lgdwZVUEfEWubuWqBLHa82bJMVUldI081R8mFK3ktF93kqbI0kGpto
FDsnpOztUHLqvI5//eiKXCLXgeXGI0qErbaWFVNFHwM3cSK9U9pMoVuAnd2U+sNrjZiuN3IkOIsT
0KELKmLaJLrMtx2kawn6+kP4sAbIv+VpB1wzna1OHCcZdBMf15s2W2lnOQ8lVvLYY6z1fFG9+QT2
D6YJJ+dsf5zbIIFuK0TOghAZaoKR+bTrRjbdaYmMSCdNZuN3G+DlMfO3zz93U9AUYzkprtQVkwrT
ym22UpwAXkMoShvIqFfQ9NJ7LKAAhOJH0LyaBA8Aiz5yy3wW/RRAURmwnJSWYHUUxebe8ALqHRZM
P8On4i9a7ZoPzehvx797RBMFsxsvl1955DjW4hG2hJWN8oPocn5urXUVIL+AkM1QIW3eWE3xR9YD
+OgGOXmVmfgSw6FRpRT6sxCNnZTfvjD3Nf2cO/7V/JH+LtfAB0bGpu10VDMsTR/dnAN+uuMNcUMg
hv3A89n9EcJaEgMIZQDegr4wptiUxQkZC2bUgyFJWW6kZzqiKfVFYCN88TTxFWSG8X2P7A+7MS3q
kNKgzMWercpPkbAf1Nn+zoVDNZMXO9OTS15Wr1ew1EbhNb95lMztociQ3Zb69606yqI7SC4tQd52
ugwm479D3v17Bh3xyfkqA0a3WbMfk5wnrY4yNS5BcbWniVhgShhFbgaUg0znSocIwhfBzeSAEauX
KBCLTQN7gFzzmMcni4Ha5PzeNuyZ7NdF66P+hyVFV735PRqeRVyPlw535zCdMfBoFDrMxtPWPwH8
etRjLUCRJ19m4DcN/UtQXt8/03NTVuGObfSJ+yWwqkJDf/lj+8x5IToKSQy5q6nmbUDGXynFqJ2d
WwSg9o4weCS6I0kTSdQsmMl/YMk5K1hfSFYbiTT2zqdQeaQyae2kYYdktwltvuAK8uzi24DTaNtD
xYOvWjWFSRaghhaeCatlEnXv0dyDQ/XipIBCcCNQZ1GJzhYpOFnTxlC5QE6vYg1khkxj9aff7RLH
6OmXuoy7XjFCPWat8oJnl01wxZ67lxsXEwiMlkXy/ODYqtF7IqwL5Bhf0ygT0yjtTjFDpEisTQ1g
GorLZTL3Vpo91NF3sPHoKjIyl+0F2RAHtP9GZx1qL9CXAGoOzwcOMCqRPYr5Vqk3hycE9PWNov0A
XYFQUaCuwRuwT3yYYQsACWnKkoD9bTqUxW59G22zNFmjbA9kgx60s13x8PrbCPQEuf6mh/fHO/M+
sSpe9DTc3eflHw6KxKMMhm6058ED6v/ZsbKSgVxcELuvMSb7GX6ZjIetYXDBpwYIfeAuLPh2P+BE
14gTZ5Fcqbu2I8hGnwmN1aKTJqP6RANSkOkqPri66eFY/+8MURAJ/j+xx6HROl//5AqCvgEHv4ap
4n4PKr7Fx1w62k0wGqJ2+X3Nr53I3gEtvvhR0fXVoQN0QuJZEbkbXpiI1U8YoTotCYAxJR09mvDa
6pt9EngzHyZqPKu/QCjzf3l9QpcNI8LAD6Nptxftke/WsgNvgpphwxzOlLMqawr8QRHPJgDsmvr7
7aOd6HZJTfM/XGUY/puBjBS25HTqtgv8CNJ2RINCU7fbld3LQLdC6g5rgu3dhbUJAvEkTMBUb+W7
Ysu7Z0DcoUyHejXAZTiGQlVO2RTbiCwQrm+djh/uCdDS9RMJgnHXbvHLLb3D3HZF78jtZbXYSf6d
OKIGl2ZiGF+75qbapiyiniH5RmhPBIu1nisDJy0msoWSdnIo29893aCdSDnBYgumDz4ErNTmsk08
/EW6PqN1otTYi+gOoiE+MViVUHK+zZhDjIwWkLfGQYw9qmhmJPviNJjVz+p3vyInN2Rdfsgll7A7
mICVQwCkXgQloegrtBDTaJPqml+xqaCzXiZcK7e0R1Y6j3YaZqm3iaKyxhXleA4ljanQBld4QF5I
z9KgMAVJq+67gLqOey8IYgxvVE5S1Y3sLQfk/ldjq/0q5xfWwJi9VU3gV7hYtKsZjxrnaI+P2rux
u2mGiVcU4gu5fCwlFYlJxpUBMRdhbIn0shSU2J2IF6mH7jDcV3ASugo1G6J1rzkLGwZcL7rBsYzc
q7PUsNEgK8CL7Mv60WE0DIZkcff79ZUIbAUZJpIzcx4M/Ph+ZfrCX4xCUbJKmW7Ry9p1vjCQCqMW
7VtaJGFg/3muCgqmZtqfPzH8+jVOfqyTGPZn8eQwbM8pdJ14A2X1Qusw3aIRhItQoOZhRECufj0p
3F3FV5vhfWqx0RYpuepJ5nLSMK4lEVS6FK9C0h82n08Fan8gFvYii9C/UC8H8Xd7wSSIQXaGAAZ6
PGzxHolT8pkO0XT5EdyOLAhqyLJWOL6iDNsZaJm0x9Om6tEVLlHhEfk0B5G4IdgE7Lep5xOmCyD8
O6DETvV9NCLDy2c/7F5HsSkY+OZcn8hDpYEgK9en/J6COoDfNH/HNdIAhw7obSyxKisiozZNUpEf
i0bqQ6E/UJfx6tLVJufEkMYdHIgvKunDwnYfKgXpSA998rC05CamU0tPU5xiwCs1GtxoasdnTLy+
AhVEKP33/W7+mGUqqw2/irgxh6fG7u/DnwpBuCVhyBtqnbEr6B1KBgZFp5ew7mej5rPseLYrKpzS
O5JLjmsjdFgJgXh4kAi7l9AdNVptAb+ILvHMGPKngVNI2IhlDuIQoCdQ/Vomh6Bx95Zf73IUpRxr
lmY4RHZaELRO9wBlueqHjfrRrm970REW8baO+vDi3P4GoVyyhN8rhIUN9fbNgLxntIO+6+e9I6md
ZmMoo62uS2YVbNDJXmte5ynMcTdx7M0ozF1nYq9leHiicfylLMRaFW3z3keC/GLIAQxiMrXGoziq
+oWW05KiXXgtqWskruT4DQaBByhzpgGK5oh9A5OjV3CZAFzd91LKnc09Dk3X7SBQDsD+WbTM/ab0
JGzf7/qcnt55yl2B3HicZX7TTfOqnC+S9Had/JBysvld984eGKg9dEodPAYA58Te7IJn+pVCg5go
xwJj9XX9P7eb5twO4PphVfZftWlx/09Gj/NnnD4Lwz2wnDuE6P+khIHOD11ATvhe6zJqQx0xtofp
CqQwnhzHTQjhtY62+fAiuofNFU1GZ4zRP9ctVrUvf141Ro93gqJTepF+z1teOx8qaGqP5e6V9z4u
MqA+DqAhK+yCVHcnf2vSDlD7WIXzLddelmGpK4dVf0ZDWlvwovu5m7PDhcAKHsPNuHHcnDYcHzin
4xpHiOTni63PusoTFcg/ZMK8mgOmVH8rdKPfaX86QWADXUq3kzg//VWioqbdyRrjym9pyKSluRjc
wkg6H9Uyqn3xI7mLHWpUYv1gcTHr01EdEmbBe7T/Msqaxuobw+lc6xP0QZi7UXC8PDsVIumPMddZ
UJh2jeO19zbIXN3KSbBp3cA3MyT9zLo/DGQ/8eXWEe8s7qNSBP9CaGxKOxAuQaXvBnHLxBWBeflO
RvoDQClMJGjnNpjL0W6A85+TRvCDdvcJW3z+cSIJ4tPsglNbUYCskfIhTvFqIeG3BdebivAc/ixN
fHvV8+I+m0/DyIDOHN9ZbFAm4dGuxA9wifz8eTQjPMOhCWUla2PuvD24DVAFalIC3dqQD16OxnnX
ADLjCd5CA/DGT3Lnxdi7X34/P5Mu84lSZkaQyjU6HIu432qXNyYdVj6X8cMU4phPhIOIO4uTtKB/
GiYUj62neAiqes9tw9r7268IRTY9iuU842xM/YQwTDnV90VvHCllk8of1MEfBvq6GCqjFtDwgMoP
AUGLAmz7m1m0crj5oRKx2m3sWAo2DrhXUTo28SJCiHIflLEqCJX2FkQPwKDMDE6KegaJqEJf4dvx
tA5djdVBovl1cP0GD/y2rWi6TeMdrQ6QEJ4h0/XCLGokFqb2fKbsDuWI/v9gVxx/V2yBQW4vFYeH
sOSwfHSyJ4gU0hWHgu/zANDeLCmC+XXAmmV9BTzDe51tSTrd0ju3t/mBD0fHSsBhN27YjpGbIICD
fQoGHoHr12MZc52sg/L3zgFuMKqrtbI8qZO0zDV2ue1b7HAx8twAx15jQ3Rxv4uk+b9YdG22FTh6
V93yBWtQ3aTQjFX5v5oNsPV+3SIk9HsvZpsv8ls4gOqD/cA3CCsAW1320NwPHjvgt5LHT9/otW83
Wm64yql6zoEAxVzvv4QBke8ND2UzBHosPKJ43wXW0RAi3jc882sbpVDRtStri4HHhhJbuaZkHtHd
4oJUeU+PUscVWw72f7TtzaBN04RwLqm3hsxkHyfd3nXrkOzPNQEV8m5YBR7VxSLGkhhSCSfDE+gA
0QNg05LDfkkVVPj30dUvANOg50agLDXsRL/kKq2ggmaxx9hVCgGUnMLenGDlX7maYH4Rw9hfjLpX
gf3sL9j7b/Oj/HZ9XLjSsoa/mtrRpLzSYOQvUMP+FI91tMv5cGce0GyJb6RgU068miyrpqiSUZuN
24abc0JMx9178APHoIAreHovc+YNWeIh2rSFiMJ/UazrOhAgFtpIpAyW6VJ9CwMWvTwzOdRGyfkI
2WUmwHhu2VY9BmvPPkMg5ZjMMIVedGXRtAQH54ZHtIGCbQIaM/KQ4X6FgFrhDnM2YPZMDQXRnAlL
tPCWBYzGciSDfYH82FyVcTI0+j1NboZv2+zYpRKJqSCbJD1x45p2jpN2pOdjK0ZNKKN3259Nzja8
D92whiZm3Wx2jFotnPZXW/jPvhSde5HQtNgRqsNe+vBzfr+mElM7vtFRiDDjcIvUdYca1W6IkvPL
VdjUN3tSPuR0T+MMg4aloVAWdJMBcoAWlOZmAtQqIMsYv/SIdFx0Mg8FEEzu1sjvIyH6T1J58LZb
XcqZncdFVRDq7ULm5pJNyfoCmxntcmRVkvi8LIuu4W9dEH6kALkJJk5S+GcRrXIp03gFQUSEOIAm
5g6GHF2VKY/v6Hkefq8YOmrcoANrZv9j9HQHy8/1GgIZMJBKKcrod9g7EfGG5vpR6ibKpoN20JeH
bwsQe/Srzxjk7h1xIGuKJSIvX8/CJdkFzUp+2/a7dDpAIEJ3wKOePLcedtln80P9zPlFxZDeUDK1
HFSlyAD5F/+VaKXF/WVpYw3pmxHod632RRocAvBoLaSulRrba34WLkx5tMXW5Nny9CHI7uCD6u4F
QkWBuw05cgP054VTO54084Nb02iBoOmrtbWy2VgDb4Gs49TTVOftI2M46ptfZGQNafd8nGYdzhTq
A0pJNnuMjm2++IHtx0s4HWf4MJYtyFvXP/ah2oAGNOWX2Ka4dTuAHu7jyrPiZzv2be0uFYvLsKNs
/suZq95o7qYDxNF/WOhkn20dh7B6o6h3hFS+qmGkNxetT22m130YRhTf8VJblhv04pmNcSRly5Gd
dp+YCANIP8/AthT4Mo8JNYv2DEkvIDNpJgVhxnCEDF96gvi+BisPwNbf1g972+3Df1kTVTjOGsdS
ZPRMhDFtJWpXqQNCMWXgRNvYCrpxHKtYezytFxBKOFiGONeJw1yk6kps7w4DHClW6W6MgnfXiMA2
s5vPMHhBX+Q6tEy7TdkMARfUeEcmyIqTa/o868iq173QkvJb+uix3bLIXHeoeGReEoJTRzxXTAjb
gL5fbCLXRze7QNSWU+ICFj90GcFc8UpRpaEmGJl+wgwITOznLdNaYMdlh+8n0tkRVPTBODj+zD7G
0xQhoJqLfNJBpJw7YiOOMZj85OzBuspIUt/LbzSTew/f098g+wmeHOc1AwI1O91X5EDn4eYWDd3n
sUqS7ZsCUk+yK/J6rlhARAs+8L1Ey4/hHh979ICSeJLbF8wOnV+4lafLJBNaYNkw65h8MOHdvCei
N1Tu+IrzuTwXRqiB3IhXBdA6/IfL66szItZfA7f/fSEs4kbzptDZ9jgthr7Jt0rY5bFyRPrlCY9b
3A2p+e2UWqNC1OI6kEVVqZQgJTGOdttNW7ZUaQNu9R3twM2CmaGD51zyhxkAIJpUfE7AG6b0mGqd
NUzXb91VVfwEHT/KrjXOJlY4Dhgye8z1KnVzAUpWBhTcjT59P6cYcQRhPgbi4kjb3CaWWSH5eLR0
r7/9ekRwoqcDVU9znNHbQKe7A+vkCrApbIXU2c83umf1W4Gdd3d3gdjAhmsmQcB5TXLE6iSWR75S
8sip7g5s5gsTrgNaabgAbHam9yKwON5ShyK5L/1wrCY7gJ382//x63cPlaoIdUFKNTzeFEz6dQ1b
QokWZsQv2W2Woppi3Oec0meOmw4L/wdeDvvRmwJvIRbt+KAro6qSfOk5hk8qZ23AKBs5trSsWjSX
Z/Ygyq1DAM5pAB+9KHm7NG1Fls7R6CNXKypg7bC1gNRA5zFMm1mTXKOOCygPRNh35vVKqcVeV6DD
At8tTef9sygSPtB7f55Q2nzQXVu7/hc0EeyYbvMCp1IxJ2htPL4by6gv3KBiuZS3ahG1xTU1pSel
/KXxJGJjFIqDjU9+XZwrqSFzoFP7lh/xT+9xFdKG+fQA2RNdOe3Eo+rGtWdvDerWTzppJ6vF0FKZ
ZyEZ0sVETwd9+pCebaK2ShBMhXTm8rWzHYNFStypfvB51nZfB1fNc/1iOxrJ//CHdgZIgQnwGOc+
062fmbXYtplxfb8gGaT4a85ygvE8ahs/zikwDyhg6rODzH25D4gk46BDLavQ5yWnOMmGO6kBRWnc
accYzjET9O5boY9gDmodFkKibXVOlsefBzn4YC8H9Ho0juNscdW4Fq0HYVG33mxNbTKr4nqVH+gB
yh6KZAF4xRpBklp+LrE2Wy85X4sWoJ04xQqIspZRqUB8kE2fIsMKVEYsUjkY4NOxLqbWOkKYFJD7
OtbYx083/GRl1gsBbLuKpauUBw/sTGdDhaifo4a+SdBcdgjpGcDfGcoeqVJoEPQG3LHhM6SNuApY
QKfuigm7RvuR3QJXm3frC7xfVziO6dC5th4v3MKLp4cmNjfWh0sr6fWD2wcO988/XiI9HPhltFF9
7EBMoQ9JLmbP6SbgiqhaBfVAe1g0LJItwlpJ9SDCzGjBC1so5HUdMSsv9MAI/xvNgqfo0kQkxD2Y
YtGUAjgLA6nMJMlEHJs39eqnM2Y1pqZLFvoFMfvQBt9f2xuU4VF/frr67r0sadSJ9At7U2BkcLdf
2ReszZQ/Puwm+EMT9ucpk/L1+DbJ86hrYe4GHlkIbSf2crwan7HV9z1suv3C+6ioLDac8wEEV+VJ
Phtq0Yq7r0/UiqDo7gk12EvE8aSLuTrap/dB+vEDzipsUhRfVCs3VONiN76N14+1fF2iXF+MP676
sp+SXWLU+GdN8N6pQ/A0bti1CjiURbXiC4xoLWvme1OfWR7T3vF9V6tTmDpc2MuZnrmrMWecNEf/
eJzbUT5Wf0V216rjyZDLhCDAS8P16/bExUAU3QLliWzHJn/cvsqSq9yZmFrznI2nu2FuILTxOmhn
GCYLnWwxBdoWdTQA5WlyZWnP1rAneZ5ADip78khhRm954UVV891wXKvKNVwawBAIw5YzMPptvfmh
zI+H9xt8JexDW6baVemKJw89XEfNNq6hC5MXrScUIEmKW/laRM71zDTCWHP7I+GfQm0LP2Sqps44
EhuXqncWITDTjcRutjYXkkqIDsUlYUPpwZ6N+k7H6EsfQrpsyc9e7IeQ87coIFwSd8Pmhd8cEytK
IZ3CzhyLjND2ddvm3JE2Bf+bimRx0orTbEcAuZMyxQP1i83Uz9hCp2lxbk/cz/sh5m6CyCbjqw09
EZ920Q/0GxRhC1P0pqJeBeag8wFvoD21qxMGU4RI4nyZTDu6jsVzxZ2pkSqViP4wsJgX3dHLk0Um
szdC8yQPuLhEQbdWimvGxLd6ZYtnFno2wynhEjL2to3E6rxw4aGf/u6Wq/DcbvbPQINyJGZFzuV4
INqpmyIg1VEY4GbpM2pkx8+axTEu51YLflmUub/DpSYl3EdJ9RTYYPAWVQ/obxb2cCTHVcpRArh9
R8phiDTwhdYh4sWhH+/vpqb6FkxZFe2iRFqRMgB9AF4ZQENaLgULJxBqjF7aQvN8QZh4SFawq0BJ
VE27ibexuZ4+EnZ25Zk7fKuDe6xQQJsN8jerDRPzMSATJRs4d86ozLPkPXJDr839axeJ/7CMXzMF
kT/6yqgtp6F9znanBp41eduqwQEBtzj+e32wDjbe8uVpPPxZaJdTdS+r8we6G74VwI2rO0u29XVL
O0vq7LQQsqjp69+JkA6cfTr+i4hAJ+BRja4m4XE83Nmcx53gG+WDQcqhnNlhWvxVOk5v8fcYWtcE
secR+do++0201nLgAZQdBphLe6DkB02wAlFSo8qRdmJWQ1+FhBHDYaSZ0NeefE8ItO4iAj+cuqMV
PEItve0DchhS5heMiUOPuxohUf/8n6C/gZm7hvl9p07FNhKphZN4b5VToZduflK6N4iJFH4GxwZO
cr9CSyh3RIR1r51u2ESBRshs2aXHTbykBqcuOpaPCD3K/J+lVHad7NbeWvy20UQ2sghbctoalSM7
rlXyMEd0RfJzz77Pl18WLG2DV/PznrNsuu7IkyGXICDOTWAutFq4WCzbqCuWmWi3I6pmy7/tT/W8
aVhUGjj/fbsRifVeBwHf8lK/lcqw1ts8WwQI4M058TuCJ8Kkx98MoNUAn0gKp65ZPDvhYG4gz+nD
7zNzPqOcIqxUaKZjg+F7KF07ese119tkpcDmC0oK6i64oM4CZrJHVMzs3ySmdSkbWRqSILW3co9Z
4KWFpDz2W52r4j9zhkqbQ3gtjLToYWErsOei5Y1r5SxTIRSskvWgFWSSd0Gi1wpMPjp0F0tZBOZO
T/DkPSNyuesENDizriirZi9mlOYGcCML4Awy9tvC4WQYRF773+tPYbki9c2J6/oCER0d1dinun48
sI8Kkd1GitjYnp3OlOd3SLmLUqDPw1K5S2obb9w9TxsnnIrZXy8L36kc7cSy2SmGmZJfF3KBmrri
yUB+DbOMJrguSMgKkpnWN2u5QH2wpw2BqgdE1oIIk2LljcnpRUrmeossfaV0E3awWGe2SkyzVfiH
cuIbzHS6TNAmQzxU+Op7H+i1qAmB6hhiOo4A7WokSBeNZcgaR8Kn36QZhSvZhMXVQkIfD3o2LvGt
y9GeT3Ga8rdm0yXoJUzw9blQL1r2cgKPQu3An08O5FYCA8WAXg6pJwlX088cP7fVYRmymXNNNdB9
v9lyOX9PUX4UiH1LEas1Ip8ElMwzhhDRR07lPNtfJdB5bvpQwkMJP0+aOV2FI7wPhPTNe7uRBp7F
jQtmDXULjSU31hKQpsEwhoz17+eSyzKgTUQml1/3ljFs5E8SCQ38hq8CwM0b8F0Uuru4IUA/7ARM
uWI5+DS/Y1YfxcCKCJUTUqrz6eZC8NzEGyR11wtV5G7kbe6YfHWGYtCr0UjI/QZkv/S3llZekug6
qlCQ9br256xUyEWaN2TpHa+4Vk7L+owb1W7/DMsrpCOWNGiYRvQH0CjVIriLg9KIvkcyxxFcQzF/
eKfwo2pSIXXa6Vs9sPmYog77uJjbqWDzlaDoO+nT7Ehr07WXHJDoyLezm2hWflRecvQrBS7PmC2l
bgKZmX/3vzCOJND+7mPk1WunHfECdap+6TUiHUh+qQ3DTGE2ydiD75fJ/sdyFt86ok7Ha11QLPTb
5zkogepGTx3TlkBZog42qMuhmfIKgXwtnxhkTbbj7JS1RrcshbSSmiHXdAXSPAWhdVV6QUUBTEtM
z+PJ+PKFBkC3sPf44lVoaaM44LEgwAbJ/XZVoqY12AF5ke+6pSRiM82H25SJK6p8CvG0GdON1N2C
QdXWy0YmcnV1WUMgZn92DEEnXXdCDSOTpLV+yC5YAdevMhWZ+00t5wlBzEffB5J1VKwmIVX6rfsI
AsF/x9vzzYr7PXiU5RjGr0fLUk/zR3LJaaqeyrQPPeRfzWYCsTudT9Lw3tFe+Xs0EkqwXtz8KL8v
rdOJs+jK9oUTr1VpmR1m+SfT5O8nmjPjVOfRlCZ9nUkLP8yYbuejRdBWAwM0FBnqXxMRjVcUjzuo
S56Rvfo2XTKVhCJozO0zCHtNwFeTGLb1SaIEOyXRbJFSQRnrg70/IFrutTLNML9oZbXBbyWviCnu
/DLDjY1AOYXuhLT/uNR6MsDtOxfo5OjC09jORXjQKfILZwPGSvBEifaslhukydTq6fQBa0mi1KZk
O7sq7puWEpQluwENlccZMg49OxvETnerHG6TEWHdjwgt6lVb9VQ4Xp46GVhZHDRrd3K6P0omRe6x
YGK+PkmFjxYbsVZzYU0NtHRVAaKuQMnGOx9FgNxdNHH9rpW1BKNy/1o1ct1QhvC4zFDOfgSje3JW
9Jc0qIVfthkwirVtRm5KK9Bh/JcHkZyhRD2HCOrgyFlfhXBIpdZawEvTry4kvxy14IccrB8/QexR
knyOPDfPVb8kW9GxJ7r1KRBqznt1z0WElW7tTOTzEUh/CZeO1o7Mmti6kF8xKjQYxpt/3k/a0YBy
P/ixplPlL+86D0hpRhayXjrylAjxQ+ikJKdw9eQzEqRPLdw5C1XWQePP0FsXuzyxMdMRxfUgBOq/
GHaELCdwHHpPo1UAJcOi3Y3UJuLe/9D7h6d1vZOngNew98kVNNBvieptgK9yqAFkb/iGQCH8Vam4
J0N1W7f+HER7opzWuzzWWBRC61pyD1Nprg04Kp838pMY3AlAsN8ksn1pcBqMZVWyQpyougIh1ZN1
3Fz1qLaj66OLG0PSTjPtTIRmH8eeXDP4ZRLiAqCFV2y7tTwp3MvAsf4IloOkKbpdHl5lGsaeWyA7
5ij9sijddkTJhx7LGx/EQezjRbEcvqizDjJhXifCMNaqo7AQLDD6exbPhzVt5aWGS618eIsOzSoF
eegDPLPM0yUlTyTUKeYKwTPN23bRPtrVMWzJYL4C01F+pVepVDDsAdGk1fhlMHkSn4jQ/hmFu0u/
/QUxpjFrKQOsWUHNxMuFgv9dVAtUPTLSX6NZDf3CGoJZs2DkojUEr4iNJfgMuDT7vAFnL8wE7F9j
a22p3c3oZ8u8Z7imMhKTqSIPiMHgdeMxwqaoZTiTEHlTb9w5AM+oRkXaK1q8iUZWEGdqTAG6Tqki
s8cd4sSq6LJoZmPdEqWxuojl60yu/eqrRCAt7io6GJGCeS63AwibHP+fu9hYfp4FgKv7OvVf3azK
BxOEFId5Ei0bdFAqcl73749+6N8nIbir4XtjjCTWnC73UKo3dHbS2WFDSukkRssAfOl0Pi1Omgqe
ausQs2DGpWJGj+iUU4alGO17SZot5Py4Ct4/3MLvAHyQTKPfu6YKZCDntbJFJ/6wSl3gbkJGV/6/
CTtqQxEPjLQXLUSv07ic9RcEUl6idTxDGNRUBV9W8fKbkQrVMbk8Un3t01R4pw7NTl2NtdIf+aSs
qmDoJg4hbfoZgBzgxuAcjpslG2JWUgbrvYEcxwnxdEI4wF8R+ShBpIa3ZGAoG0lIZYSSDeTfb5ZV
qwGPu6FO7InPaffciWvNAcR46i/db0tl4kEs1qgVx+3o/17DFF2vKV/UM4Tm1/kSv2CPkTC8m5kY
Lrf7+BDvDGXWN1fZUOvJPUHMidci7RhEcIv0lO3uR/Ar6fw7vlARa6XVs0j5uMPTWMaDdmCExVJY
VJO+9IkxlG1yB/gcroFeH6uYzWVat8SQXcKIcHDWTkURl8wyU5TnZ8KVeCmKcjslSatNawqZPmkR
qcxlsxfjEuWg58UTI/S7BDf1/jpP/SfKzFkP78gVEgJxnEbhbVJbxNBDcUbMjfVDPax9HEMgjrDg
bDYBMt8qoqoEBgkNi/ORxxlS79001hRuOjFbnZ+C6pY4YrYWhrBL/McI6L1wM/Zo6uyyLY27FsoH
2Klc9Pg5zr9EshvDV0pdwkg8YKxrVCiPrJ0fVN9hrGk0F0RsxSFm2mt6KsCKxEktgwmeObeEzvw5
p9hzhZs9P1KpHWR7u9X09cRuIl9CcnmZ8s1U0oQ9AoIy004xGfg4UqS3lcbTCKAFH/IX3QpE7xU5
5xkbXy0B50V1XuBW+hYjOxIzO5oUTPgkBhqmmYr6sbLlUQSVEe9Zw0KIKYoE76kliI9m1nR8rNbX
3s0whaOln8jTE85jaFkJPW96VFvrs1eYDNi6sKUSszgn7r/LoBYNJ6/PPCcF7iE4neYunm4y8ix1
qd/0if48PMhuu7yvsoMrUgNJZ0+MiDpb89aPp9m9aeHxkLvf6XmU6thgTzRlKiaQQTnULl1CLidy
FWsIOC8IN0DXBJyzDId6Wi841z2iJPfDvi4uhOluFlLOARGcDrCiPrfJQzxpKrBFc40UnuunE4f4
fvlqr4ozzGQG7tH8faB+11Qa+iRR1vydpDPWs6g5w1Av6mJfh9KXvlNuibltpTH4xvz3BcIiqVL2
DAd0tcI23tocj61a1tEgfVPsaHWsbAKBoGVA6UAhN3lzjSjSZdfdNnsm7t4epptVpDz0cuWydK9E
r/5ymkQQVNOETWpLThzyF7HfstyEowVkmC4cCFxpH4p1zOC9vcMpC8aqEzRLZuLlxZaormuVXgtP
gBjkJuYzQOytbaL4miSWhi3C21Itu5Cpc5qTYH1NWuDfpZ3aIa/S/mGoIyPlsmihHsU7qc+wH5vR
X9BPDa9mseTyXPv68ao0V5LN3s4VGZW1TU94DtHvVdbu7RAAKzxHCD4/qtQaQeYh4bXhPcahgbIC
ZeV/82+k7JHHlSdIt5CSoW2uSpyrSk9nscFNFRepWqcZiwXaUto21YYspkjhFPeSuIh1hLo7FJ0j
lilaKy2ZFfleE06z1T0Ta6VnFz2GXFHQTRoI6W2Rfd/8LKA9KgKvs75yribJSBaOio6saHSgUxpz
MAxq7Q15gW9LZLM5J2PdTnGpdzLj7Yof4NsGv6VDnWf6v2w317EhecbvAIDG+Bkczzqa/wFOkKBr
rA8xS03c0OBZbdQdZ7ObM62btZRYrz4dwz8b3L4Kp5Gz6VKXEdkKOsglpX01m+o82fx/opFfCveA
TVJl1JqIt9Zc2jVBDjbVjrHuyITAAzwMRXo9Q5XpMPEqnJ+5jnorLXraZAnafHRHvCvx9bmnG7v3
cHeFbzOj2n0CDCbACX9GpZgQKpt492tKB8UV8+BMxWr/Kl132B5nzr9dHpptlqIrJXe884cJgv1A
pd/zrSIb+/0XpDwfavGXB6EfUJBzw+Yy4s0ii2INjv1sClbLqGEexg0APfyzFmT+rS3GbAXgLyfz
rJwRdWSohLdNVt80eI6vsjlSUZWsi7NIpUb+tHEHiZAOJnZtv1cWvglNL+SLAtLeu5n8qVTZiwIL
Gz2J3AiApyHpiwR5VBaIw2uZ6uK2qqi/F83tsKmHsyKneIqeIV+yH0PCsdru5QB0Sgn+5oVEDMLI
JFNCAcodVQQAPgoKoCbTBSekARF4oUcsQH90TSJIeW5yprBvbpLwRuIsvBc7E4HssOcPACCniDOF
MkQwGTTnUhPSp3Wu5lL8wRhGMdT5RzzYhEqjyXPPT51e79fs7s926g8SgsGQx2lfMIdvB+DZWE+7
NJWTpfCv1S+Jo/Hs9/zOY6+9rEMU1fFVV3YM3YJbREHY51oJ0BubDMiwzfJBgS0iV/QzIg2bASb/
eqD1t5K5o+0kJZurS7Es4k3IkIRfksIMxYs1Y6xbcoAO3zow6F0pLkfCDU86NJbXXZIbYA9JhyF+
yPmYH5anBRLOzfLVyXBCtIQbSwhAoN1Y00q+hcpS+IaA5wTU5sU96emZ/54ML7vqSVEvVosjqNB4
BTVbbVGiXkoWBgscw29bPlmHRfctljDve7vXlsfXN4pmGGH/FxLBkQO9D3THRVeDzInxqvzmme98
uV1v5TyWcch363R57sU+Vd132k/UZ6xCTwh4NNgdwrt7F8BwrAglWcqP15aBXmygmzOpRzkxjJlu
cHuY7XSFvRuo30DLCLJtMHVkGNVfzwQYsYonAcPoWzCB2NHFejmnxMbtH/33q00hIA6EYDtmO+U/
jCkUSH0zlM3IwZKVt1Hn8rnJMl2Qx5kt1UijAjnxwAbm1wZk9MEnams4/VXivuMDFAxoLuM9iesp
LGlUCG9z0urXbQ0w6QRbfsIdE4dVZdG+Y8EZME7QyHV4VsTkY1t/jc1hWdY3E6UV1lOcRJrK/nf2
L9ax/Pax3xgpYymxF8Bsw080Nm96qnzbq9TfiC0bGQ39oR4c1E3pJ884xE1c9yoCNKarhHRkAC6a
F3n7bv5Un40bDPxsn/9W+P7EIfJEYk5Hjnt2cqVWR2BRsFWjhKRczm5w5IeXrKZ0S48JhrF5a2A3
NwXMDKDz281K9P3fvzjHl/eA5Twtb6swCIeyNoN4tSwiq6wCliGxIWizMd4ROY/7b+bcdhdLpF/7
dFGV7TA7QTZNMI7XzjgzslwqJ+kqJlzHlarddK5Q6/1JhP4vcwdsja9+lKvMoqjVZOWQnrDcu5SA
O1XUDEt5qrhbwgscnBZ9AEUY+vzxy5sDpY7LD/+xI4W7oaJU944pyqgner++brDAO6M+lmLmEYBR
lS8lm4neaiRGdEhJ0hRobJj3wgDBivqOs5qljmLlBsU7iksELm5k8+aPATRU4euKKzwnMVdYGVKd
BHKdtFOJBCAl6BgD+iLgi4UR7TNi5nBKRTPCc2zDYrUrgsDzbLpJquJRDsxD/iujOOQt+bxbrIDT
7/ruxf3LXp+OxBZkWnYhQJ0wvKUUJGnGA6dxnN5+UeRzadHdxvfvDKIVyZ8QG5+YRgHM/hsQJa6O
dVbr1+oEdPy+kB6OItEzBfOZGLU/XihUcQcXBMBUUrFzLgwcS9WSOsKDVmYTW3OM4eTqqFje4/bq
HARAdXQ9adLFFKsaRsFKsChutIjAmDVRaheCMyGqyGmCPlPJx8yxeozWx8qdxtqqtcpXFuVymw9L
rMhrr5wiHy33QAuddwZAka9FOgj+0lCCcziafNf0Hc3P5yxm8Ly9hoYXQ96jECNtocvh9+SCfGz9
W4nCGXYIolror18eq1hHRqUBlpLNIeaCXUheGpnWJD/FhQDxS9O3UKmGiyDOJFg4BcnOJ8/qX/GP
f9TA/sSHz3nMw5ND3qgKj+FaEmmp8kWawHJL8dMxg1k+0sYDeQSF+ZDkXRTtgKEOcz5LlvWxOloQ
rxqP72q0VV39xmyYbyLuZjFuqYoyKfuEREZ76oQL+8N88aGReDE3rh/Yafg9OE9a7XB9x+eaZJ4F
P6/SMwYIXF5693bDmEnjlwogEOVbV5xHjt89UOCsAOr+cMo34Hzdqub2+Ka6bIaBv7WFT6pRelkS
nZTZC62EB6o1uiBoW19SVef0zIBJZa8GSjUG4meIttQm2Pu5TyOpETMkCFf0VIFI8vCvVNfU/VYb
akfHi/Z5avSQOdL+O0zPPEU+y32hAfC0nGmfSzQucEe5EjA4jWwlIGROda5x4Ts0e1t+m4tdXllj
Tj8dhKvlo6iV8Sp/kRLoQGgcaeZaeqAtLSAMDHvvxd+lAxaQzwoPUER9MwRUlB4dhWkwb+UU++l4
WSb5QXKtckZdXcp9HIE9KKfJfwnw+9DbB7t3yhcgR7BO2X41cmVN92yAH9ndLx9ZmulCBVg8lctO
kBfR8ff5XBBjuVy66p7avvDCQKYQVVClNUv0LwjNrHphdnPi2NCYWTCVD8ob3uaiY9VsPdrMvuEg
Q751PVLON29FYgO7elJW9PfL9UCvQy1MLye+C7b77nDil+VPAWXdaJVUyONlD9Zytsrp9T9qzK7K
FWwqvCK+UKLM9vF1XgFBSIFsuJKpUE0HOohfRkycZ3isGfs6nakYud/M8J+KUvLOjuD76GJVgRii
5o1fGfV/L4Ouhz0U9PCse5SQw0p3ef2GoENEDhu4Ggjbxh68gfqmd3SIuLXp0FCryH1ceqgs5aUJ
/nN4kh3yGwvWs76Hkiky6AtC3NVaAHZ2eEqA9BSKmEyMgCnqmDcILFrK0hM1aS7J1HV8cjLP65MJ
TsoBSNm/zVMQcGkt7ZCETSre1rzoh263ufWEc2LFAm0stJPFZxzDwqr/qahMcABpiXypFDbAO7aO
hAT4U5Hf3G0HT29PjcP63RcYZsgwI+DgtHPUbDWlyJnVCM0VzdZbJ1ylDv+Ln3Tp6pazKkPMe31s
lnA4xjkFi1MfSl56wteK75tTSHPLGJRBPyR7m1bhchznrAKoPqGZBBpnKAbeGzhNd896JuaE7J+b
iahFAiiPfQ4qbMOBRgib1yCk/uw/Kut74NGabhNGLVBQsMJktD1Vo0UcVSJnEadBoQ3hztjSzgdL
qGi24aGZx8e4+dbb9mqbYjJckZpjA7BiqhReuE2Bx/RBoWDSI7IIIkOgxuqVUfEfAVQlZ+WMpacy
WkSN4Qtc0e92+UbTmT+4ayL0CEGhkVBaWbNW/r/8bxZCLxjk/2hF9Qg3Rk3YJKoMFWZOg4XFtN7j
EEtakI9Bq4of5LGKnQr16NMOglYKVasWltHQY+dLfZfM15x+xLdNCW4COg54XTWichn4o4cC6SA8
CEXlBy5ojRLVOCHcnZz0py2/IbEZ0XRpKJqofiYWYRLt5tVqg6uPVCwp4sWu51y3fggBJHW93+2g
NWJVxyxhhbOxUYf+C0m+DYaSzmE1FU6QVRDmEoCJtwk1J0n7XG1KGHV3mRwF8pY6x5uSoNpjSykG
s84jp9zjP5lHPcL1INok56ilyzcBqBdasfT5nbXqlwssdcndc469WA715CqN98ccophz+u0Mkt+z
/mrrOK9t1DZiPepVOPGUkgiuxDyC7/aJ87VaEZRlLOmL3AuXeSQaqwy72kcD58Gj83KS91Em9ipd
Z8qY/AklA2oBEA2EEP1ltjNLlGxdAF4N97HeJ/mHSOehQirTr0Jw3hqr30ZtH1W7pXv1pZ6rcqrF
mKJuA16dZFdRz8BvgWom/I/XNGpT2AmC/VE4jOF35UYpQ3fa06zcDCCnGroMR082041g6fzq1PlH
0lfVg1M7gW4zgHXCL8SbnPUxUba+wGtPk2Ub7tgaqsh6K7z2Z6oXnXbWT64+Oq0GCUctPu7yU8nf
ozQXIE7YsF1GFbgpiPeEx8Z2pP2t4SJfqKVG7xvm60D/WodCzCA6eiMqS6NMfR7CrV5NY1ocJ7nz
6WOHaKOBSMzDFq+TBK7IB2KEtEolG51NEyAvC+4HuYFb/Avxxok6UKjuUF3xmRXUs7ZMjkHHXMFT
4DGE+zwOPnJ91UixmioaHZ3ho8pFBtAzAdyUgVYTcaxxdZeYfOIwyB0X5LHNGuqG1gXJKFemf3w3
wfSaFEvjlH6MH4UxvWjapYTa1FQ3h5yLkpb/mqt/ru/SDY+s9QrDKtG9HFjX0ahz8ZTA6+bH4b03
n/3Nv0Fo2ghJgC4Cr8UpZ07rpMy2of2WotO4CSGwHqNv2fmW4J7+DSIPOahDZgKbfeDfHdQgkuG8
fWFCF3hj0mSlJJ9q5k3yXLd5XPbxS7ukhDtQ2hnCfPFnXunTx1Mqxh8o375GImu5H6BItjmuOQb8
6DKhRWJmZnZ+EnfQN5uYo/WjtrUnMj13a2SpKmUlJhWozrHu3d7MKu0SthWZnSkPO9wZFoY+QgED
kUX4fk9KNDn0BCE7l7jjp/oA2SpniuRPikRji/04KyPqdezlFRDuW2JYnEuZT36X7wuwUsNdYvEf
P29KRdrbDTCUb7zbHUF6Z5vFqCsc/2w5l7gFkd4oS/D1HaJtovZCB/uRagJ9An/89Z9GLc2tiJOP
ckZcouL+KgsgxgDkE54bxGzH+9SYEXrkSZuDNPe/PwqRpnhslMHHzHGuocJdPy4ih7FJio7g9Yo7
cCyyTJhEeHg0UleyPNXPFHhenzWVtp4U9GXvgkpgP+SDZDd8ZNEMVHkwyluvT2gpRyXMDY1s3ayE
YQ3JX7DQlbE0/j/KZZYdMv/y791awKUy1F3rzhTeMbjA4KcWal4q/9d/W6ANZ2yG3GczROL84qQL
rQPu10TCCsvXjiwNk0NtbFtHfp7+b5fKuvUNM27GMf/+AjRKL8XNJpIbiw1XBGrmkC03zxwQ2K2S
uRxL5ofBwgQz+MknIbbsADmsNriNb/rLK24ckzsJMZAnI3Xpo2bRRH4xIe8sRsXiBn9iwpPK8wuj
BoEYOQjV8RlPxQMrA6ZUcqJT4T5cjXlkS1u6uQhxKlVqRPktgEyVQUDdzHeQbemEyVBhdD/aAZ2Q
4GBAPpZXA9+VfSeGJw0IJiI8V2JNjJcG9bR9JIzU3IMQxfe+UZrMZw5s4xlWJrcA+81POhQNjqNA
Qd/Td7q0FEN77Do/VGv0bYmqYWDDNKuQPRl3psbqJw8YG8OlRAb/b/7TLZuuuVCpJX7kDDAb9IhW
EhhbtPT7bezQP+6gcxE7WXuPZYn2J25IM2Yy9iUFVt6eNqSuitZwq06bj5WkNnp1pAf+7n+WDzTy
EZBJYOJNOgyRwjl4D35Ih5nabMgbipNQ6QUzWKgcda/VAID6Zi5X+0o8VulCYNOc+wFcjRIavtOo
bhTJRV80MK0qqvG7auj2jNRzRvdQ5Qpkh8AlLpNz8rMWTghQ/eFuQszNU7MSlVBQ4oaiF30shIpA
s23M6y5pK2dZqKTrhgH60exbNFNowjme6I49zn3GRdMG2xxrdgJSJ2mdGTzo83tzZsMK1Il8KPsf
Myd8ZxTtbE1RKqTLspRh2IcFWp0Vcd+2dyDopSarIpBzLdXYkNOZhV2zgZ3FfhwWkTK1ozebk8h8
Ax8DWDW74zSY4JZ86TK1D86+c6L9bWauARjPZZ6Ui4bMremW5q9CNP/kS0qFyyKWHRIGIdiOXIMw
z3sctQOA9z9W3N32g+P1KBhHUpw2xEfPl045s0KgjuR8PfZIGNBut4WmOT0tX0BlI+bhLN8LsleL
BqImV+cV8Cw2Dm0S6N3mB1YEDhAFrjsd0ng1DAx8IKzleBQS9uFstsIxctIIr6JkGaWgpWaQo7qn
hwdLgELoeXLa3XsTb40m3EWmnu+6YQO1QdY8NIY/EdevzQ4HuTl3XR4Ns2ksX3XI3RFT0oSopfWL
dYOCGt2HA6sxonwn2RtPY81jwaqgfpFZ1zD8VEq+eyBcN6wOKDhbo+6F58InDKNKPc3S0vQdUvAg
GQC0HJptrSzhsofofFCa7UU949Q7VwKcwtaErSkeuSd+MNMdlWDiGydLm9e7m9Z5lig9171FiZty
InWOQRDiHs6LkrPd5PaHMm4cFyXXt6SaMMYSK4khkBTGaEL+lukwMUuAyp+00gBIaVZXyVA9pdgr
gWSRFo7o0i37RIVS0zqezhQINnq15Nn6XtNU92FGLigVGkErvZom7M4pif4drf+efLKp0q6AYVDz
nFnAMH7qMnoXz37kUMGG3YnnA/Nqg+Bui9QBrNDg6oJ/NDFWWBQBRo6hpQz/0UX5lUK8838UvIla
5lOZpd74KOw8FnCe0zaXpuBJDZvin8JDo3GCjUiZVWDcJrL424sVBTyTGAcgB4dgvKMPnxxN8UsG
E6iW7NPTZRHGFfqzWpAspnkLvFI3uyEWeQ9iA5vn7v+7b3TEEk9nDmEA+7kO6CrOK2WeZM8wx+42
Ip0QFiCCumbKPMdHg3Y/47eBYrbciuzMzzCKlxi7Sz1WkizHXPnDv5iZ9fnVeAtvT8sfd0/OUHXX
Pz/JqkHtr4YA7BDWeNsuW7ufObtcynmFuH6vR3Zp8yaJRMEDik64pLQx5EUEDw2jLttIM2R3o9Ts
26r1bLy8QBQaqT9q0S9CO9YO5HaFW3x/zazx9qNuJdi6ol0LGjZ4nJC2gcHXBlatBmS/SQih6a2d
yLeRmYYmDV3D0B8oy4o7SZcuDhnq9AMdsWFst8HDfp/Qz1ref9klhns/G+I0aQONrFIMjFv/7yxs
oo2/sXaizmtyFUVr7qRYpprqpyd98GY6QwbhNUjMbyMvDPnek6gMpM8RFZB0px5Qmv4h8TJcAfwU
zTPSZyFQhrCPi38/Pf2zDMrduy46Gw3ktNvk0AbKfQgnxZiuKOyuLar3SsS+KU3WfXceVRx05uAL
/yFbuyg7YKxIri2LJ3E+E53mfpE+NDaLLkH1lKtRzsI3zeaigv6haRyaqpRG+Ai/LA3YZgnwefpD
jo9miRC3vimFp/tlYLhHEfSWIBj2YvNuGbLN5enkVnDmElBo2vPE3QeX5Dw/R4/Ms/40kjc/cVFN
/jIaPV4L0KtZFnzpt5gUWVh5rnNjFrz/0MrEWWW7KiPLutYaNCs9p/n33wsrhqdUPo3pADwB78Q+
ennk4VZHsfwAfemBEBQwDwN01oE2lAZaUsuQTMRzeeZ6zxruJIOnVbH65X+3QOTyMaS1RFHl/bxC
dOwiOM2vyImhY75RN02AV9y/AQSRoEC4ZY76FGx3eOxo72rLoqtCtRui2B1bNrbzC1uV/65asZJL
nJBo9GL0m2R6qnA05PF2kE2wYNqmo+ZUQNKrH3g/BVhU7eQsZiKqRLQysNK4LG0g/NLRlLXG2LID
Qu3TDSDH+KJN+j1hPbe6DDRfYHZDY7I5zXTa7cMQeshb+1PTMzjwINcccKx8l0cfI/3kVVWs+VcQ
QcaXppJrdNrS8JaHXChrhB0J1gf8Dn0xGW/S5evVOZ3Grwlj+BzQtutsmvOOUrRowBX5VgnIR1oV
Gm4UsBlawwEBXIAG/ajmHd5fMtn4k4TE1uS4uGilI3lUZKR+cCAfx/zehorJaaRE5M9ZxEhw43G9
fyzYeI0DVVFptyd5xNxGoEWSAzjmpUlJAEr8tXyldE6BNGWHNCVOBRwTMRM+CNIJe54LlCP7hqAc
SIP+o9m6ylpUZQ7yy8m67oOyfQIX7WJx2HTiDXbzI6j82D2O9eaeuuWiP8R6i0U/TOP4dYRLT3Zg
Z3FIL9vr8i2tqZlXjoeM47q8O9BCvDuWb/7j+xQRwnQASY0f3/j4Ku668cFEGcijmQzpjrxa8DJt
F8DjpYdfbN6dcpi2BJdWLCRbGnjvQAuTvw6KEtPyb1v8iM3MQ7MIVG3j6ZYK8qJgv1y4yPyJCKLy
Kde2/psRfZIqSdY0mcPazJZP/IKw4byNPfOG6I62eX9tplsteOKMgiaTj/eVIlcOtJ8IJz/Y0U2C
c4+JxHsjY14nfNZX6cUPbltcpEGWb7D+2tA6jLfr1Y0jxNedgjl50vmZ/dwBYMpzbvmPGfIrnb7a
R2LJKekoI1fQmDZ8uO7GbHGPM5/ToGhj6RnLz2KYAajvh1WAm8F+AVsMdEcdXtZ9MC3KSI7e+Kx7
qTS4k1L3AO9vGmZKw25yb2nzly4UqiVjY2Lg8yehH/Udigal5RML/mTZEFfR6gwrckMj4XFfMw1d
34XjV28i6XQZvi5GJRtaSkcUwQDGNy5jALNcD1u+Yq8xYeCrcj04KYcckjSEVqJsQsCTCU91fe5i
fart3yu5batA3t7bgbBfQsHb0lMkw29jArnli+lCO+Q/W7byhuo8vY+Zhr7BZ8hHX3u1etXN8Tas
/pS1/HZxkkj//TwfJJmDEONBVdfTIQkR+YPmb4W5eahbi2ThkdWk6lxYrggq5Jn68ipM24BiXOal
Xf21hIuncqLGixTu8wpvfEh82QbhaHbtzxjTsFtU69WJx4sgP30ZzRYhaKqd6zzhqQSfYdBevwwg
hNfmAq/THl2vy3hHsZSm9VEd2QTCytwcu9Z0iZu5tK9bcTRzxWZ8emi1/0U5fx+xGbkLG/v6ECOL
OWUxHypWw0sSFAKD3xZ0jnI7LKbvgyfQQMe9SRRUQpLOch2AXI/KMXMqSAS0sXHQuAhvE7qa+d9p
p08CufryMVXU+qCiQ0YRdsQ8XJzoKuIAya5fjUFPSzdlwNH7cTQRGLPMcBB2guyPHvhHjobaoIDW
XGr+B2ciQyLEY//AYuW7lUs6BLJKrdMEN6gKN5m5+mTEEZ0DdN8PokidFWUjaM8VGZY/rJrPpR43
rd25QDdc9IEYAfRIJH8oMBxh2uLsSSHqof0xjZuKGHvaHy9efksBi7vCUbfVS36r38BhsPK5xNEn
RFnKCj5jOSIfA1ubD0SnC8ZQrkoJOVBQT+GOq109qS1p7duxqC+B45vUkP8TBfpSwL977aRZI0c1
mjI23pmyPaMz9VvWsV2VXA1ueiYtlvKe00uFGFzQUQ35ZelehSchtBs+YTowCuFwaPd/S9S/epXl
Ep/Z7D4pqSEa8Gr0QTKKeSzNWUYMBaOHByZ+QC/ZaBKML5lSzWW47ROs+896NaDO3kyzkBWaDxYZ
P/SlmXlrGHaSii8Yan94eDFXaCbkz74DGJqgRnewJPEgdB1fDcwOqD69w5hZL9mQO/3W4DCrFMYM
2Qp2VU+rUCmjsejlzdnxMbWn18J3Ey5trPXPPSf4IIzh1JntG7TkI+1F1NprPLlnwa5xzDiAWssB
eAwR4eHU0R2sbd+bGod4OyXkjmLKa3cFATDuTz6Iev+9XxnP63UgqYRf5js1MCjmVQYyFk6wPUFI
9xiCOLTJgIZaUQ8Eza67nQCaKU7alqZfbTVfb5Y9LzgjlAvhu6skufMGDnKQTxlieBymlG+MDGcv
vW707javEYQY3F9XWnUZFgEAJEy8BT3yuRKMhWsbRMSZfFUvTYVEI9u6OUoLsWrkxUkcPpaIzof8
id7P2B7DcJ8S2NSaQ7il38WXqIfmBk7jN2/l5CQBR9RDXsnxyKUfle2+YDRaN1DgCfRpv7Ny5hou
qpLly6atdzgKZOcgAUy1RIpo8ABaQOYaLsPPDC+L3uZtfP8/l99sJi+SiADCmLWueQWqigivShkT
nl+dxqKgiMDl+K89k7SUcK6o7clpsmacVYIv/k1eFZ6l7CXymtp9ERnRukvw9WfPreiCMWhhOcNa
54dlYFW/dV7pDrTl1yVXdJln3U1vYf86yZxJbQsqdEVL5weWfY5QT5hYZwZWZf0b/2cZxXkrUBWi
9F3YmHtiQgYb2yFpDaNtrufwPyoix21kCjrfuIUQTAKvw8IZArSp3OiGGIWbow2LRX66PQ83u69v
eERNu4uVYXcjMpSiL4GJz73UO73QQD2f43df6m/ZmD6eDZ+JTbgfx0xSQ5jIXpyhIdYs3kRLiKT0
L9MNxAoY74S5f6cb1TsdwwmYjH61jn1ys5eSG0Nr/RyKkYtkl69s4aEOIA6s2mdKAhUDlw28JALk
bJ148d0gR1YEsvBUQC3S19MVyrBRFEL5kMlzdLu00/RcEyTNlNFQorBus2pDpAizgoR5njNaHPRE
ybtc/uaQ52ctuhv8nNkhRy1SFLkWlD3Z6YoP+qOSsNJNH6YqToVw+zcBgUWWmiUWJgSY8YUQT/Nb
0PKDok6cCAJToeAPD44vearfFTVjanNG5asqKmqZO29RmsH+bt5556c9gkPbleMhIbbhlOwAnZK+
Nop2CZgWWAEWMu7JB/zLuXLXiR3B2CvUrePq3YR7MWXJySPxuheqpeG8sTT/kuUMUr3r2sLxqogX
7AROqGkvdhLMQ3uMmOdERQkESkGVosb5sVtrcmG2siBzAJlcAVOlWtWeCbz7UbwWaZDlYRE1vs0H
vbmznHzQchMzFbYlvw+AbW6kEp9T43/SD/woovj1ZP4a7y9MD/f302WKWa1MuMVkPSmDO+m7bDM5
Mnt/LaoWkIR3Z1qviTFe3Wdq+YSnwo/KWl23WdRMKoM664d+6BqWcn625BHYD80OxMFKqpFSkcBK
Jj7+43jaLbRlcuRxZXxCQ0HIkTrMpza4YaAf+IzgjRJaZA5qdQKiiAQ5HniAK9+mXr/CYYymBaKN
X3dpcI6qKdgJEk1VTjyhaB8p98Wu0ZamtCJ43xMzR5ng4P07X6PadqSkNA6eCnqV5NwQ8LDArdSq
0W2IKw2dyuk/x1RsTWpSbVkduR2iIAx5sksnI+2AF1J8D2sdMWr5TEi5EKqIsQFoAKrz88o0k+JH
EhzGDxdPsGu3w4tYQZJ8DYR2f8W5eUF/8serf2d2cGnQ2Rsd6GzniPjKnVKEHlzU2/hp8nNCye8o
GLV+QVMiJMtrhdde3nzulTakHq9ySFlbvUzUkZ6i4DM+Ov9Jd2r0iYJ8ZpmzSOU9i4SAHCzOGLiy
jn/To6X4zD8MftlmiJk4dREnB4CPDgwivXhHSKrbu4Xq7H5v6XpFowMFC5N5BVKdpKBfIf16AtA6
bEMTSlEMuMPw9RNY8z+pkDbpTewIE+I+QgpprRTqjpKafHrhmMVGTzdljK2fsxo/1uZrVHSYwtVu
/S4BByGR5ZTO39ExfN2zEz2as89S0MEFOJoCp28gOMRA24UGG4qxLwbmxLWjVEueoQ2IXaPSZmjz
e7DNy5Vf+iZI0B6DdYTN7blYs/Q6nbfabNtJJQG3umbh8Cr+iz48LYA0qCf9TPid/cjK+nUlyzj2
YmYf+pBr81RB4IimAVR7L8+013tFzP3w2+LIATI/3UYTtTZ3B4qCRFri/dK2Bn0SvC1chnfAYKJO
x8dlR80RH0FsIxYVnSVh95+PxxbZe5k7A6pmNX7ivL0e1yjdqZUs8awnCjha505ikDcll2IC01kc
6/52jzPsT7nmLKU9niuvSCiGCUyI8bCZOsf0cygbsKH49JLi3XYZlQFXallAaWrAWnIOypqiyECX
iHkkVLabnwYtpGFSA6fz20Kswh/avPjFHh6Aw/BEhPYXP4ezybCDjykCtceY+kcJecghTgtZ31Am
jfuY5Ur60h8M+f1b9nm18gHO8J4SqbSrUD+I3g4Joh7/SDB84RQ7IewlzrSGfj8U6HAQTW3HbZWO
dJpYUEpdhUt0e/cATTrRd0lBSOfVrkd4b6sHEmAfm45T93X/ov8G5DzOhd5UXkMigBY7zPYzL6t8
fwrcGlNX4e81fC9wJGTkSOTtHoXdlqIVu2CzHz5u6CXBIWinhjMqvI3dL8JnkCFaCv99Foa7m7uQ
94AWMqujkX2U4qBOWlB1eTf/DvP4YqPWJk7tKgzNhzJzKiqvIAGDeBVEW6545KLgXGANzDIKMYQn
WO5OMgUZaMOyNN8jvxceldUF6/ShVZ9nnI4L4WNDwZRhoudBN8olMigvNgpk5Voq/iVBhBztl1EN
sX9Zqx5a/fNaAUDMiTWHU0nyWBqGUuK/G5aLRFXZNiss7XHErfz30WAXaIu++9+8TngJUGBV7HZB
AYDHwiPkgBslgglU0apsagQNXdf84s8v3JUBawWdeO5K5F1+aWFPyr+GwlEKdI10X4r27rIKeUsx
8Fkkq3IomNAwsoW2FdCcPLsq6v53NuAzP2ZUFgzGcet/rVbLR6CepHP6YUK6EotkRXLPkVfXZC4p
6Db1CP72CtvttaA0IXeoxnnMniKRvFi9KQ0BXlVOQ7FVtOgTy0bQup/U2Gz3rC6VUF65RGXO8T1N
eiZIHStRCRNJ3abKFyn9ITJH5uLVKdDxMT/l0alP6+0A5Hq0ZZsXT/NaRIjzY0Pwiaw8MEmmuKUu
jUeWwyYomV9eUn8yNaIpTo8DV5Xk2FQwxYDsnJxT3/9GjXEgcLjgnbOl80myxiDTBhf7wLeDW4XT
36arWVyn0o8latUuDZSnK0l2SOZ5EquVnuQaOpA0LbwxDR40zvpBuXADTB7BCaN8KDwY57w7m9E6
mWYiCKJ8NVkWVbgjQ57YNd3wLK9EAdwumNfoJ4LNnwc5IOJB8XQoFVwV1MV2uYFRYSwt/yqhYXVV
rplugY6Xa+ubXVyfcqPjKuDFVxJ0VANJosZX8BJ99ax+Q7NY/OskOpamjtvySSuntgO++om3m8U1
fS2yWjgbNSkkJj40K8jrwo2hn0nGDC9f3k93vw8ArrnmXgd1tcoQcB81pFvs3NVuXVacSMQLjfEl
/lfl3bbsuzpHkfhLUK2T34aj2P7joojPl8vcd04kyaERAVqDm2CTM9QT8/nW5JSNmOITiuS45gT3
8qPJKS74HZXW4hamnPUDe7bzdptJMC5KydKMisPREmxMUNswQB93FqCi0cmhOp+/nkVrpk9CEKZd
TF43avkRTfczuaYGeIXT7XsqrL4zRFYrPwM1G1JUhRvEoVoGqpWZ+V+/X8kJkPaVUdep2TRlsm9r
7ACvL2S/JDSDQa06Bbwh1aqRHgVsV4bsxBoktKiDDebwx9zyH9IXS/NxtbOmyj+6o26juIjW0f6P
oLFIP8E6140iFbDTBxUgANK8P887aB41mhxcf0hVrC3b+WpgajaBlvtp7hdNB2MZz2SdGJKiio7n
QHd4lS8ab3BZg7VYKGTW/1tx4znCt2/ldjuEhPB2devj0JULrVwnYOUMwCcmD8z5tMSizKZ+YDI1
LVy2MMxhWxoGvfQphGaL7UMxS2O5Gm9kcsxEkLLi8mSJT+P3RxYRqjbNW+z3nPS9fqReOICL3v3L
oRWvKnsjHJRG8oAfWfvTVF0sCGZAV1zfwHwJzJogiVKPx0r17bLG7t8xn7vjuL+li+b1kY2NTBZj
Uu8TxlYDf4EHlOskjvyV/WkF63iMQn8g9nIzFckVrRpfCdWyWrX9KF+6B0ogGLkT1GzNttghkKje
wkXiw3RSqIdigo6cFh1emUlbNFJ5zL0e5vR1FsM0Z6HmWmNMZiiLgduzH6ToYbXo/r/vFML7ZFvj
6L+D62ESb2bvlmdFEDwfgGpvDABJMoEMVY/tI/JHe2QcPoaAkmfjgea4VnQLJUiBxm09TcxCdPcZ
a5CXS/OwrE9jNmrRt5gycwx8mFqFf4PBf+GyzpLPNqLjf/mZ+WEtiBHq6FQCutk4zQdYsza5ASTS
Li3EBPjOsIMZI/9Ods8tfGvpE4vtk/JW5bZKc2Xx62MFXe8JUGwax16KqSE6BzTSbRY1j0NrS4QQ
EAlrbJ0VcS9UQhvLy4AyBP9twdfNNvIMMAwqKixaT5ht75cRkpe4icaVClIA/Ai3YRBPz3dAMdGP
G8RgnaoaQkiOghuppv4lT0E9GHXlN24r4Rnunvr/pokkoTYnsIVhKJaThoc/GpnhbDihHDT/noPs
T7WgkoHToxVW1cfR8+AywI5/ftCEBlxDMBbtZt7tzZTQ0OT5jUMHEhlHM+7WRIxmY9PpJJQuemu5
pv5+YBEnpcPIXQz7VpGHGhhPOOxs1VRkYNGjLeiYw1fTV1wkZaBjX5hkmR8be4sYVbVnZcFt0++p
6wwGiwBxGxyxbWTFqU6aM2FSwnf5fCP76qBDWm95m3dmvknbex/fkC0CNzThVpQ51kYhX63bPwHj
mLj/dcRFcNwCO1VN62GtRT7ZtZoz8X1r/ecNZ6zn8IT+GzwBZsg80MBN65nYbv4+i4bsDxrPXI6I
cdH8bfka/UpBnkmIfQ9npBb2NC67jcXE6Cu5+BF5CMR8JSQy6rd6upeQ4ea51Ai0/hecJIwbjb43
b2jkrl7flMDbf0hhjvyZdcLeWAVskjVDDjpf/dDnwfE0u6/KnG4uawi3jesnIU/kFZ8U4kzufTTZ
LIfwwwS8himKY7zFr13cAlB29/zLXZ8y+F+SS/CXQeu4uUjV4lzPIQ/4UZXRbIUxbV3TNAYZdc1v
KSMWjKeLHGyLsFrERWgNotWwXkw9Cu0uh3Rpkx7Y75cUogufxtCE058nqHQyWfdwgmBXZhAIE6mC
zB6/GChWRphcs//6e2CUPxiPG2KREyk6joFOqKNBTg8GqQ+6isvVuLCfurycS0QPCdRkUqYA74y8
0sHob5QuV0PojwOZbvkAsMbJdZIHU4Un54KYlpD8Te77qvnqBZ1spNnDfEgHks5xWO3A9+6qu3yz
5AbkAAShq43ZR2XRQCKF2+F41Dl4JkhhjG9ox5/4uI5uTN62DEV1D6FXQp5Z/x+cVxZXJZkq58yj
wMEvhTYveaMoUyFy0VyJTKhKTBfadR9noUx9CeQBb/fWSsBGmpZhsCH2tBnGBEB42jRX/DBDadgX
Bo+uOdR4hIqZhx9F3T7eHlTcpZaQ+nYW4P26voXEdGXjcasuiN//u88/kZ17chE8H9b/p74bDzUN
Yz4d0Gli3WREDfEYEIkNu6yQlvuA9SLahUuI652g8uAksLYNolgtql5K8l04oXon4fXvpLIqrFkp
bI4/VAl+cMtWbzc8BBEfQRAR0pxFQj/ukCb4Ud4uVLtG0e+W+1fsejpPmU6jYr3jrmuhIIPcH4E8
C8n3mAcDs8ZX3Gq0sVfk7wIlmjgZoOFfeD4qAk483VbG/XnflkdyYAFkWCSf4CTdtpPYVf+IgdYc
XSvRXaLLutyX3W/5dNnuWvq8U2dXK6nrF9YX91IdV9ictxx/RFXTlHyutACFUCF9oHzEU7VjYUtG
KPo1xDm1yHVqYdREP5ih0Oc60pYMpqAS5VSeUf2LCWgvi/t1PlvXQZw/kxFz3ggyK0jhyCGvwrxi
RXBz8xsAy76RPqvJT4x67bBHdugPPewBKUTBEkIrQdYECe9EsbP4zQbZIDD6viyEH/f9dL6h3FvI
K5RnTjVBAzf93y+bnY/UksWSc15ZS/EMVoqfjYPlSRNJleozLQMbQwImBvi+AjZCAweHDeXSQZZJ
ZHV23m7iJnk6B4PwtFOMEKU+1SINY+t76s6YzHElWGJuQghN70x5cLikzMIh+VO2AeD2id6kxhfe
4JELQZsxuqFJRs1HLb8YgTfWwNMWp7V52/F0SO/ZCnLEZvtqnNLRdgKMpmi1ilXL3pjMwkZ1IKRP
d97beg21PlQ7TrYqz3zMcSVbim4hB2plws834FtG0Li5aqIFMn2BPV4tK7uiOoO3btgb63MIlf6h
VFnGwWYtXK95i0cFWsuTscS4U90bntY2I6evR0OP13xWN+kKXXfejflTQDr6Dwd/QmsBa0e/6AaS
irqMOnsNTAt4OjzuQj9kNyGB3udX8IXI84eHmWozLqF1AFzzGhjKG9T14ESZoq6hv9dUXDz+mWzp
JtX/qb8JJnO7tp+iHSME+75/gjJOidqqjC/iXdPX0ykgRRSUp0xTs5IwYfiSJTQyg0gv9jZgaQtj
jTfIHiWUESBIR+F4PvefyGeXH4PvmVFhOseRd15Ad2faSxltyNrTb8iIqEDG8ZBHzy1SqVkIBnI6
D2LmStWbEXoXfR3Oy0hoEidC5k9xzDiJRkT8Qf+JDVNNfkmSXVgg3ityYvR49W9xfFnr3zX7MPe8
IgyrHfJ/nn4N6BpYNsjop9d6oJSVxQZjoNq3BMnruT5I9JeW+PI6EavaeeKRnGDHnIR2RVajvDP5
M84rbSWydzTvIzXCufaSG5K0ptqhugGhsII11H5Lufh+aK2jbPtfYgaR0ZCh3OpZ4kMx39yQQv7s
C5opW4ZC6g8yBn4XL1vdfZtGpnr5QsDgLaxdMUldSAksZa3ozCuVTiRk+Lo628bj8TrkEPpiMtM0
s30GNtMY0g6sL+ZfrOQiOkmXNKxbJVodXRPSuv0qnLExWwA5rAo9NYeLgz1OIdzOLY96WD2H0OnW
m/Zirzg2BT7kLvTyRit6lLdXoDRa/CJk74BZSPXg5j6IZYn95SxKZjlA9ll+QBKAREmwcZl5Rz4o
Fk19gqU8ob4AeTCsKENr0fCBK2I7Qv/gAPuQoNEi8laVZkI+EsFhYiytAm+3VYw7pw9ZVqZ+gIOW
F7+bwqswm0rnwq5BRpKTVMCKprnwxM671u3wOEL9EQ+i/NU8Vke1m8HeIPzYLzgXMCjaGOt2ZwZK
DK65yHYOZRUb1jQ+TWtyJgr2IEQE75mjPeE7jlXUwBNWfzcrJQruk8rlyQ4hZzCQ4p4tWysKf27q
wAJ3ej8ecTj61EpaHX6BJUzYYI1LWeNcN0u136SbBzQcf05lBY7SPVe8NNq998h15P3PT04nb+Au
jh5wx/qZ8aWkJ+Gmae00ukvgmzLpho4H69t6/9NTTCjZv4cNHpTYz3YKb6i/RkaT1QQsVz0XDbb4
q/mY8DjksXwEEi9nsAVLoGxnqj7r13oPWWFqenROnDT1mxKDf32ltIWDsuxoBHtwDNwsoqu3t7p8
Ov7vGTavD62lADaWIRLaNQb0lNWfJyJC+XPfoBsJTqA+8VsDod6T0MBadAwxaxX782QmMhN2IQ8x
Vnh50l2IiDv+OSDFP59ETlZkG7hQ11gSO60hgZTxzM9gqbXVAgd3awMSgI4ZhpF2NIocSBvtbF91
x8TAiy0AWsnqbSomWzgvUFhI3dEKBhOL5S9pV5XTOeL5JC6pUpOWtRByWHZX/YabGQ9HQ7ONuYOM
FvXbO/2wpwmBZwsvcIuYnl2mNX/pf5YHdYQDDl9L98aw0gZki+F9AbGggT27gh3B6mWQ7HjGhNXp
J4jE0JhhoQ6TXR172X7ZB4Bei3DHIYluI9fSj12ZuYZX3jCUdc3N6kSqHrLJzRegDDR9jbTTt81O
atUZ5AzwvyFwYwd+MN3+il5pgp0ldfMGD7ER1j7JdIw8UDrR6IIs6lls+RULUg9vI9KO/bSoQc6R
VLbY+PEj4V6n4JD+MObIYCENx8A+3XHwGmN9T5yM0MMcbDrLBhrD5d5IUyYXhZDWF5vOEgAtw5h2
5qjjzjAM8mXwuREohR3yPgeQOOayAjYX/0k/t99F7H+G0RT07qBEJ6m86e+g+xT9bpHP0ED5SrUu
+FDpSucPPCnlyBzqKFTBYzvvMSBzFpDCfI4LQUpBiTIvSalWdVi5XqeapvIdomZPMKJZZbquNqba
4IyZCGIJxrHN6C/dUWkvSTj6iX2dOQvk6CmenWIxXXT/vUYwtZ5omtKo5B6/szkFdZSWbl3xYY8p
Rf+O16UmFYnOcPpbPMTG7UXk5SN3HImDiR1JIhZYsPc43giSqA8p8dqjWhfb2122sy++NIjuRblf
s8hdB6oOz8+zgV0lcBsfKBcsPONrZ+qbMQA3oM25AN0jDxMd+Uq/g3qcSmIz/OhRbwNCWFmxuEJA
YnG6J0dtKLRv4pA6ECUknnAjZ/OP8Ck+9g/g0Q2yEUXZq8bDfZOe+39XuMJZ2SMsb4ylkebAQHho
aqMuwnQXN0FB0WWwUkVBuPH9WoBdBhM82aPqNPP/1mKRO28OW6bRIDy+9ho54z7xAlRHfFkSZSVV
XB4AfMpPUPKCs7D/rBBRHZz5ocFAH4oqk16Qurf+zQjhmn+hswvwyb0hiU8gDiXCc75NLtImjbaM
fepwsPlRAvU95kYZYKTOoom4raeK5skG+oaRGv+A/w2EAnisptskCJSgJjD8GY510mPpvYg+BQJl
ucfJmowIEEZC5vEJyGmHIOS0RKUC1P4UcNCvaQ6/AsClM0S9yGG8VE+rYTYCWCIz7eDlE3YHOYRJ
XZA9rFHI6GYGjZ3c+D5svGJFyErOJ/v2/wwcdAefIDMJnmJw+bUwkOY+3yznlv0x5esQPwgzfCOh
rQks8XgccT9bgPGPhoh/NBsGEF5hQFxO4YSU2KKvsTDrrHsTyIfZHAU/3DStQu8lm3r+qUqRvkqY
zpSWxCbYy8vYbCWoIZkUIa8X9h6rUw8qldkaWTAnN47n6webxNUuq8YoMyLMD1g5hDV4WQfr0Um4
97teCksiztTrpSPy9tzuDu8u+Qv/NZQFcp2GrMTq0EFSNaiQ4Fc+SrPwtVKxiyQkZ38rtzzfVfmW
1qhPLfDS0GeeOxC9dfvY0dGxliC3XyiTdWdLW/FJWC2dRbpIFEYASnv5O9Vrks3I6xl29tVT+g9C
59dmbPds6j1IQuoxImvsbmepGKhwunnWFw3CnbH3vYLmQSYCAdEv5tM+Bi1AviZuOEZjmMoRvSBu
DFoUhHpssWA7gZFGkRxwivR7t+p77YmtJ9X6xXsLjUjQmkgOiNuw0WtTQC0OX1og+0LKJDanbHOa
0SR2fvaA6Y2DJc9ukaBEjyoP9tbrHfYAskvUnAAmLHwMGl7eSDKzno2JzE1asMzSzb73EI3p6nwK
iMiENdCqx2uIB34WgetQAPuphXHKNBDh2QmUPoFfhwKDxwGzmxY6CLGKlMJXYht9Jpsvf7YiEm2e
n400+KFL7nRVVR8NDwfgRMAjxibC+aMMs2uOnjVNdY3e9AECJBF0tIuLWaWfTkoXv076BveFZHq8
irHTynHe/NDMhznMeD3rtWR+MMSKws0KemwLt4+sNk/dUAclTNxRCL01Hzxt9hhIO4IaXVwc12fa
4Wn0J1yl6iBWCRUUFtd05teVouQixgnnU//QYtNlAkAVigU+pW89My/OHtxff8R7vML8UlsErv7z
l28zdzqie9Qy4B0S/jKtSfOV7Bnse2XIRt3qvFKh+6XGh898dyeHB48q3jC0jbGqzI0pTl/YHBnO
HNR57IGqc9/8OzaqNzd/Mx/FCPTATbtOi0/bpkODZuaR49FY+QtpTrFDQTP16aNy7JtozPjFV/lG
G+iOdAJQ1L+oRqU2uaYy1RizAZILMmuUT6QuVHHQMkgxHSjeQyxIeQeFnc6wIKGRaGNXAo4NF7kY
M1Qs+na2hYTgbVatOsMFtMzkIHIu2BfvZuDSkHZBIuOvDPBy6d0XFYFiLVcBzqNjfOm3daRLT+1p
YGesRLj62vwa4bE+Xa2ui31vVJZVPuZd46ab2/MlnPAaiNFNP7oyweiJYLv/YRwHohShYg1pLlBb
ZydXyya6e97GxCiT3j6f2bTLHZqomWBjwAjuUXVCx4/YFY7ns4+VSfuC6F9VEJSaTbcTfeeAzNlX
AMu7NTZBv9dsZ4umJx7xh3aKj0PjGV4yu+SEpCG5xSYgNmJHLL/kWPtKDaUizM3/N/uBEtJHRcum
H2LoDax8a/OatTMYm8XVLsHPEiorDCLW2x3/CmFjH1xrVlWqef4d3crWUSOFwTVzHqwItJiOxMF0
sYDA1wJ1Y2ENDRgmVSvwqvVHoR4A+rrBKrQxjV9FmTpXN60g0KTWxx9q3eldq2MxbAZAGmwEz/ww
8+1AhI9OUSMayc4L/SmhSSaiebIOEN/5zjs2Wr0wBAdWacN1pHB9I6F7ydu68sdaTdYw649I4+VK
3VRY05HYSHd1qlYp4nRNzNKGNqw3omfCMdqaqV76UHKdjCR7/AQUY9m/N99qJtBCrVPHdWmh9s2D
5goO6UprdQvOIQXoJiSnS9JfMXoYzDzpOjl2hnBJmsq+u+vXqXjTP+iAy4IZjjq/sYYK5zRvNutg
UUZT0/1j6yAE3CAfBrxadIizFQV4iLDw5OJK3D4I2+OATbE6z7acLeBieLt7tmx8cgmygzhszQU/
V/pEVLADlqO/eI/yjNUvGNITttHB7Gn1JQaz9+iUMUM1a69jvV/seyK0+IXr/xAgllSg/5CxpzZQ
S0CW9i1itLG+NG47d0sZzC7GRzhoCj6BGn3lK/5bVC9Ad+57Pcriwg6oxPLAgmZEiKgk11hA1OAo
Iec9InSjCuYDiswZO37bYqd7fMAVFtdSBZtzLri4DoyBbt6i8B6C77MCbXMadQM2I900gBhJXmCB
XVy4hWY8Ct6zCJRO0sTCz3HLnUhtAmR6VVRxX1jheiNfLDdw72XWnKALp/d5KPEn4tnkropC2PEa
FJZ9McxQR5GHI/ozI94jQ2AqUa0Xmw20tJPC8WB5lhoLdOVgfmc+FjZakpLE+l3Wey4e9yLjpPmy
uLa8wxPDlfoseJ81qGT7hSkTrnUJSqOOtVT4pIvV701M1ZNUumDI9pfOL4Usu26L2EifWA2KPj2d
FnEeorSY4pZusumQ6qni5lCn8WEh+OC9nSvR310Dd95eMXc500Jv63SSYmOf4mV9BQj1y+jyVRem
jxmF78GmXpNogzBkWTAmzjoRJGbh+yXyvcVV7AQmvg8q+M4qrbioth7jvd+w1lWNsj159HQG5kxY
jArPo8E35AcFiz4dZIFCWOrf0+J10aacSlFmT+uU6/jeTi8q9SevSRHDmh/7YRWwb5pF5PjnAYfm
9Pa68eoxklPaoS7A7Haf56B8Np2/usFldjWLkLDoStXT1y/bjQvAXOq8xfv7gfxLz0zpNLjQJNkl
5jJO2Hr6geCkgqcFXleI2NWXg+4snw7xiT4b1+hUxB5I8dbA9+fugtBKvHWBckyEw0dznnUwByOR
RqBG05g1wfh4cfI2Q1oIu+5vlWXUEDf/30U1/IHrh5+/6xK6ZJNP4/hF1oGCdFHzl8DNF5RDos+7
lNq7vI+W/ziAALrl0IgTphZMRuE6XWlYOKZ9S0Ee/tpry6gQ/Dmr/aMkap6ktfmOHBZA3Xitht+a
KFztOM8dEdtXjSAA6hwz54FFYD5aw5wOqX5ZFwGFjt5IB67dkhwMe4lii6DP+9sAwbhdOA3v4sAH
VbDQHjFZr0XN8U4lhHwYP3618jjk8x07dEhJ1/VpjLxOKHaiMdVK2pOnU/19mGRJ1pLUDfYaaIPY
pnrA0GZ0+rv2V8aZ6fTgdtVx6TnHr8Bro97u/X3LRfSUCoicG4FQ1Lby8AqqP5Iyy465lbqZTo2t
/4otL5s42ASHEUUR1CqsVrQZi3uY8CzHQMMzsCWpWef6rGcgV9dxYpzsktSPS12+Rr8uC+eUBTft
aZgRkF3FdJEuA/5jYFqHehGpO+6OJkZuKAy9apSSlgWgkFj2pYw5kvrhQjfrDxfQ+aM4VtTaJNeO
Unbqxrm7lFaH0fyZNHOwl6PYvx4wgRfXxFlPWG7u7/KeFV3/W08MqnfHRMtW5hkm2I9FqAysExJB
Vlzbn4akJNg/9WWIFSkZWR/3uPvgYLr25LL4HBcCWCyUjdrM784Dkrvz38nhDTSP50bmdVHCjr2T
2t6XSqR8S7xea3VbEZav74yFX3UJBanmUDyJw3HAqWqbfx8M+i3HfN3ll5tsuOgrIIzfx0WF8/MZ
WerPDY1tgdeepaIeAYr9Vup8xA4db5+AoKKEOOmWM3KL8HvDEmuKim+1D2wL1qkyTEa6iBhf39IA
ReF8+/WihDK5g8SUwcXDLYokwImpV2+yIuLZ+LQv8RHiR3JURS2UQfLzYLNxs4nAALssxczZCwdO
iT0OLtBq/YsLggDGw1EsL45MBYC3MM+v1kJ8+JitAPuYjnBb6ZKafW/HEoZOJqL5fE2FNeUL7Upz
UM4hpvPUcA/xl+eUVj7p1cdDSUoiWAnVBYfPDsbUZVIGhje0WhLKPSjJTWNKJUmPJxHgqffiJ6S3
CGDcmjUsnV9tTWRcWChTNI7TxXX0NafkQln4nXjxNwwDrXNDo0L95mC3FxJWyxjC4gLR6WxBvGWo
oNbRuYCYpA0ZHK+ByXzhjUKnsjmVbeYaRxo4xaTHaPXEaer/kx02rdSKujvrvkQpeHQTRAyOLYXq
0unaVXw5Fnza6vgoGEaxQeaG5Sst1vrQ3U3TSXV+h5ARnUi7GSYsGwp2W7c+AlPDxp30hwcxsoM2
ovWvN8eh2BmHiy2Fqz8u0Iw6joSQHNTqJCEnhbKw9eeoVuF7qrk2Bp6hqAHHvXwLg02Khn3oXLoq
Lwf6ODG1f08FGrO1tPbyX843y63bJGVJ3wsinX50Tu3anO3EH2DoN3ZO7HQ1q8iVQhW3XDdPWY71
fuUzv2J4Ct96J1/y6xHwoz0KY5LriXNKA3lbg51yxU9SX0TjrSfnCBuQF7Jpg5r3pDpUj7Ko+3NW
2Xw+v/Be/5kcze4R6DvarmU3TbS7y2xhSc2k4gOMsk38QqdMVs9o6cFHf+6iuAdnHP0LNyv1qesw
BIkTHDxeTL96b8Y9Nn37dAjwvgxGxS8s0DN/PZuwXJOSxmJ78B5sYSmuNtY+sNMZ5Z3/lsLvr23l
na+bO+SebHcF4Yuj5Zt37VKBqOpsg0fn86An88J41x0n+jhfBEwKckgIofj3BehjP67+t5RVOs2m
ZU6dTmUcnzkZT/wCuJWnyDrwWk/CX6ZoK4mn7E2dzRYqfeP0Ry9T3XhLJv5hzuuxgl7IgJtglvYb
MttoTUNUhRXxxjDYgVn3u9cC/Chuzmhrcy0nmLtoHu6p+cO6MwCOrkbmw0DTRNMC8MARQzcqKyRZ
z2K3zYcbEXEdjTANSlPOOissX6HTf585uAF8K4ARLYxm0dgk96pmbfObkP+AEMSGA4/gUYladWrk
XqGOHhf/xg/tnXemvRKI/LqrOaBDd6ezsKzidn0U5yarv3UhR67aH5cZ/quneQ7yCGJKEyVp84+/
XWN1q99Yxz+/wKnoP1JiGwmxrkomhA1GrHbfPYdX0w9o6KU2p9zW376+mmaOpUAsDxKlpt4FXkQk
lVLtkQXMDkKARWw0EfIkwUURXDIVV644+ltGudRk2VK4U0LoG23JLdR+5W+SynHJRjrQQHkrBBKJ
sjQx0y4RHzldDBPvtXoW7VvJeVDlO59rumyTfcP2DMED6nTBrppc698BxSUr6qQnrp5Ie2aMw1Y8
nHeEXgGJElMIVbKZVjrxu2c6O0ngT5aBw06/ZhU4piEqkr0DGcsF12sjdHIUjysXAqZ4Q+UG40yF
u5v2sV1aYxR2Zao8C/dCJ2mSXhjrIOCK6AI60nmIpyQCaB2gxQb/LFTJg5XyqJkSuv04CLl8uyXs
1JC7Sfc9GOFB6eih61gi/Vgt1sSEvmtFvIiQnNrCyIgHSBGEX80sD8HWGu7w0QOnva0rtGciqaeO
Owe7nBpzaEY7E0lzAwU03vnN910XQYrCXcNUjBNc622J0lm1s60swFAGbFbJIf6nw1Ca7X9nzSTs
SpVN5Zf5sLQkjJucBSlvSV85gEqOdCNGDx53M0Y53nygkWubwIUPhAXmWTauFKihFzjyvx3QWnUx
v+jKtPFJ0/Hh8WEljG6W7wSg/+M1re5CgvLxgcf94o9wO5vdMN3quJQpG9KSEDhZt0GmwJ4HJ8Jt
xNLiIZxUXYAFkvPOFj0ET2Q3URM57q7P60uzHc+W6+ghtylCGjWxnjQMGFWsbH+IB1mIlkWOG6pk
kXyk9ElUriNEACm7A4kY0utkQIxS0NuT7UOJwu0lHwdV5bO2Jz2mDZXxdL0BiR13TB3KYH774MfC
cVgy4x2Gpm0AW56KqvNgYi68sFhUgndHr77/Ut3gEtQO3wOCG/vMLA5TAtRUy3fRJ8L9zAZoWvst
BUDWC0CmhO1+ai0MchRxIz42NQY62Y427P6THN23lJYiN+YORBC3ruOrEhLgcEXN5wkWGoen33ip
Ku+GHd5ARu6hr+pJgEBj5G1hmnFX4yOu16YF97m7PDhCI+F5b5d5UlKJEfiNDTSE8hlcO85WLay/
ro4oFWOMmddtt6KPyyTwQFGVNYuN+Pyupg/MNLnDTRYp4Li8KrnZBoOL3GPk37GgmR3ujv4RV1q+
YoBTyWag4PVh4M5kNZGMlGX9yx5eWvBzJ9mWbWg5udHnU/8OF4DUfoN6MlXJIt44uNStKzE67/CX
Nhxr4DKqpxb08c01nMMLMpzR5jxwB4LgXoQ1/eElRp4UuqkSGtOSM52Jp7w/NgrRdfQD9wK6R41K
guvLGZOWVNdbWLLgrdzQoZQKDBtpEj+j/TPLfWABv+DZHZK/cUPlRN/aTdeWIrZmXv4EdacIIqkc
p/U30DgU9E09Y01c/bFVqWv3S3vY52/MwNp+fhnUHvcRrapbMIJDgzvciz7OSTG/qtNsj7yBMC2F
qd5bFU161RytLwtQ4YkoFsgs6N66UDNnUVE1dF1hwAlRpN9DPs/YgBEtzCz8u6PAiGlmI4k+aAU2
uLK7L6O7qG3vlgisi8rgfAx8Rdx3eJiDvH5LLL9mHs+RuQkpW64iXB4FEnlvN64CDC/MTXnLuNoA
BdFKLPF5d/Ri4LEGLG2ce7L1bGvL3ZnBiFjTzf1x+JUNqcOSt1/uEvSOQ7IxIr3fj3K+pGpQMNUG
KTeFMFI04vVLlpVYHG2ZpDsXa3+HR2uzzkyf++ORbDus//pJo10aP7BWyrLW/MLfUPRZ/AruOh5K
tyj90gTxjT2X0Zo4MGzM4vcWJ1jcKG9o5b/AI5ehvPBd7pZve3wYl09MLkJyl5kiZ8umBzYgakyi
IXKAgJIQXRY4pE25NOBPXIzQxMshoEcKmBzvOigNKrfduMuzUzvkVAr/m18MUVb1IXVULJBOj5OI
M0pCkQWXyg4CUD4Zfkb/YQKEomVSMIcgn3wZk4A+QHSf6XOTJ7KK9ktBhfbMzB0pNSzzxBobuY/n
yFRRWZBohLRVT5KpPAuIPOEcUFNp3npkPoPK+Hu77szIXiPPGfZumQqk0iPk/eU5r9IiTXAGWbk8
Hpk6xCuz5MI86Uq/GouecxWvP6mgmmUkCd8FM2fW+QgPp/I5ZVYPW/Vt1/hWMeyH34HdAfGAS8rr
ET+Ea0rzhMZqzCtP74nCi8KemmVA1xRaKm7m3Jc1h3a+ZBePtmvfIurglWnt46CXqqfLZHXMWLcN
AxCrBUealH4o+9Vf6gbZy66fSDkw943LZCOWZByM2wheDx/dkN74JFI6qqA0+xShPJPh5Oi6nKKJ
XoP7yg2CCRNMh2joyRiblqwxvWxiHzp6Hin63q0qtDH8QIwpDBB1+LmZsQ53uywyaiBkqormOwi/
Qw52T+yGTyqtHaziszYMahCy6UkBGY6Dg1b9IdRc0Jf8kfKqKtmUepOMAZsVtoS3t+klV9ajwFpW
4sWks9IL9lPSoUegyJvv/eykVrIRITdh4ECxUBPoa5aiobuaSzsl1nwjnQsZpQ6cuOfepx2HSiFC
ISvS9omjKWZ06yWhpJnWhmyTlIfp7kP2S21hxlZXbrbLKhkVib6Fof3PoQ0UuNzNkVIUi/BhuLGc
YxiWP07eCpReRmS1SZ6LhkJfgR/5KCCnQuovu5NMroBOZ65BsJE0Xtka6/F3uL0cR6BUP6/VodDW
+Mn+iaUsUrBcVUDv1ZFo66+/4DL643KAym1k9f01UeMuFIJIxnn4iAd9Kyp8bMiGr36YS4/zho5j
6Wbuj+Pt9zDGPhKy4M30r5iq4MZ8FcQkZbiC+bhsMDmHaNKZCNc6nk7EOh/SKWeyZrwa0PLgiObH
Qop9RnIR/n4D5dyb0MhrByiHx4T6NPCmYGNzy0QeA305zoWnJRUZ50tJobdcAI3V4gXWri1ZGBt6
43z+MjTrp2TNcTAbIWibIkDKzVr7QCe8x/tPN8njHmzaNTeh/tMO5xEneu5cFFfhFbMpiOjB2ROb
Bao2/i2kqYhCuCekn0eT08oVtiVUAPLzyODdUKiMOW62dCUu5H8FMOnNTwPKrGf+84ffJ2dWVLvE
QIEaHIyv3873w4mK2j3OA3WG8FyxYe//FdOrS3FRsrG1JNKxxSsyBImMsu+y9+enmpVMN7LejdId
slxUpxYp+/anMpPATlEIws10Zc2vkt6q7Kvy+XtsMitCd6lxqaznwYmZjfRXsKs29oEysbsdm6TT
Yc47UvpfCXMAqDrmWdhKCay/QNh+JnZ3tdASjBGXUiY8OZK5L9ZT0OkglOXxr0Fy9U3lLx6GuJAA
1HMSpWRB6KV2F6ri91bTigdAg6ihZMrVV47OXRnyYsej0KgcGZ/+gFZXKKcFNZ2xF81hRG7rRdX4
09D2UaZa9pg1EB4e0CA1Sz9knXc75/H+QsrJt4as6AFh3rFJyeHN81Y4vZyg7cgpbzkiOIMK50rC
+EfYtiQz8qwNbp1EC1gTe8pdCQ6XMVrmAfS8sLbcAEdKL57r+asWQ62Uj+SaQnDHhZgRypTpEruv
q+ll68+oF7KIz81XwQY5X34cgD4jk/UVEDZumA/aX1ahQFHJUnYu5ChnhDQ03WkrEAA2Lwvl0H+o
SqujxvHRtIcR2GDe45hoX+1K4MaaWjyz6YoC3kdidW2oXPZw0oGHj1KeMuNttBwhwqY9qrsR6Lov
o37roIdshA6OMSLwiBDkSm0BGeo2blvbX8kA2lTOgwPswpw5WGKIL1MKvxQcNuE7p3YwqQKmbhFu
kKndWi5bhVstr2lX10eyZgEhmeGl8qIBIyuDrKW0bUqMy4sUb99JZ4/8iTOrGvYLntP8kVTA3vwp
n/4CGPXskhLdrpaEhaHeTd5XEexHzKnyQ5szBKys/9Oz3htIlD69yNpM5CXK2UMJaYCbIN/nPHhC
6OdbGH2cjCTQhuhfKNEgElDYlDAc8I7AtgrtibZHBmJNVbVjmep/llGReclsYomjp6zM/nlWlUa/
Mfne4af0qI8RfptQAN5j4duPo5laEZbJw9ZpcqlEtq4URefTEKlLj0PKj1YL8Rpixmt5LJMpxxBg
epFCdWXHk7pBTJMfzS4BeKgvw8YsWLDMhw8a+1ECBOQPUX+mHA9s0GrG0B0+kaOqPbB9A18jWj2F
kyUPO+vERsQGpOPrPSV65NXCTUR3Mt9/2f5+bC7Q4ekB1G57P2vknNn4XG/tuVO2eIzTFk0Y5XL7
kvqslvsfbzT3G7yquo3HonYVDJnewJ8A2NFBIe/xePK/XlZDNG2feGmYs81BMQg4B3NlQGKBQZ9v
aOiYCFnCd26fjh1ZkrPR1904/lZH11C9ychHt4M+bF5SgPffs1PM2DjJd8jmTjalLsAB5INVWjZM
+5SXHaklYaUROfMDXAF1YawbyFi38BCredCSUsUbzrmVXEB/z3BcVbwtOnXQGMGkfIYTE9NTVt22
GtbOD0QwDVRZwPqmucv+7KTrhBIDYdplDjXdV796gUNWYQU5JAeddvL8PSO8quk3k+SfqN3V0Gxl
Gp9Yx44flU2JB3df8zUZ+2qTjobI7Zq7K+lgfSmX7sinacro91GJk/NKkciz8cbV4n0ps7aT5FXh
8Vjbg5mOR/voE61GWJ0Z83wgyB9cfw7xDymLYUsQg+bwLuVAAOYAKiQsKwrtc2urwjqd/htjVp1y
rw/LSuFySj7YHcZsMnV1m86NIO68npWv7rV60/vwngr2gP6raBiExIakcPYTNp/k0gIcCMT5NcKE
+tpPQ/bxHyVoXfedifETe1pAieVGITmH3//nGDAdulu6JwOg3JzHe+nxtWsQJJtV/jeeeQVHx4kZ
MP3q9IlpQIXCvR7bWO0vQQ0SVvxEnC9/U4ztNekT8td2x9EPw+bqPhGqpFB8OoTRIQJ8FxZsZxSd
L/lt2FGWDDqe8mZwX6SF+FvUDW+pGP4f+H8EQOhfgy9O39XdySlUKXzP9FylxepZRgdWT24neq1j
jc/t6ZnVhqUrJXZzPM5XeBgNpU0z+syk4zg+pj9EseFYECcrms+7Y3nO4xlmnk+XA3xlc53JITXd
JHh5h8HRh6k4kVKGpG69rFlzgVNqKXSYEXhXgoeHwGF28C4VtGQimVXeLz4N1uchnCHwct78KuER
rBUxCilGZF0NcjFWujqVrqcsEyGtShT7gSLS2JsB9TKMhQRebkBbkABBf8FPluM76zo8BaeH+4Qq
cpzMRlK74TJpvRLkUs/DGHuWKlZ7dby1NU0uJXv/YKxJUkFXj68/IHBbyZZZUJl1MwxN2Lb3aLSA
ZGXmRx0+7sJF2LKVwwGTwLFMI78NfgyYc9mVeUa25chLkwL9lmnArITrF/ofwnS9rh0T+CiFgyE+
XNbHf/WoNB17l+OE66wm3lNSogPvN7P3aTNmqKJqDdMWenoZhdV/vlyCax1OXxuU8sf28hEXt7Zj
JI401p3ouP/g5XG0WLvXW4x2CwQcpzhssrEskRmpi0P5J23ntz9HUZWFQVkUJMRnxTUIretYbSTN
dAi6KqoLDPDmcMmGmyZzf3C37qzG91EBpyzwJGLMvMaNG3WndktK/b+u5I1SOqeuxEu4UY6bMI4l
aZL0n3+SCmaZVpNIvjoKJQnpWvlkcz80RrsFM2UwyIbQn8jsibxV7EB2l8sqhL1ZVYXfGU4K5wyu
ECKDFmAfQmH03crXK0yB17mSBQVoDVdVPj7QgQavX1Vx0G29TiuM/w3sUypEgbrOi16lRzjKL0yO
v8BXEc/OoredWWPo0EfAFgl2b2qLmFQ8pwbFoStJa7/oZTy6fiwzS5xr5LUOeesP6Ulmx/UEBegv
7G9jbyNZc5Q+klHyIj/lrK8z8BkNRL0HFZXDr3Rh4GnU00CutDw3P5yJCA+xfXvLIRcSnFiUsJlW
6Q5Y+bit9grj0g5pDpU/iKq4jwG+ah+A33xIQ/uruZfm6bZZeKICzqKhxkr1Z3J/1dQGE5q2QKYo
fcwB+TsU3rRhLy2D0SZQvqYT9crWe5jYWRizJbtKk1r6QRXwe+ZE/4D5ppB0VO/Twt1tYJkos98H
Gk1Pvy9fgyyZsqyn6BhY6zIBDRZJcU+oBP0rjlggXXYkz63zSQiiuVkoH7UxAn72ftmBMmNcBIAD
N2wU816ARkZRBFzmHVWfsbePFnPrxwuLRyYjdJ9G8+Gwka/R1wtIVh58RbkHVYDtoxOYJDK/uU8Z
9xxKFq6v072hykuNqB2pM1ZPXOJdbVntMSH0SKDGIvoharf63qz6S5u++dWkqhU0m5eyre7QrErQ
sfZiQfaCklEHfLPesn6U3W3yjzpD2MkFTTl2jYpo9Ek/2X74Q7hf36hJfM4LYBJmZ7y9MZlU9Rdh
+Xh3whruSjB3lPMqeOOIVpuIZBmeBk5a7i8wcB5RjafZMUoyXlZ7B0wM/l9y+hhGFWGFio4GVIYq
NpZDbirmJcf90Ce1oonZVFqu3rA5mpPwF/KU0aQyhu3vZldDi8FMACheRKIX/ObMSsnfVf/W85EJ
OFzTa93eezEdmvIbBPGS5sjZrx01Q7EdedbY+aMZklMRWqeTI1rVOtMsydg/i03TNA0f2oeECh3X
S8jLI8F7tCpY+YB08aqIa+jWhFp1cYwQqBRdbals15yRHC6ozEog8xT1AXFHUyFN/cHVoIz5Axd2
pxW8T+bsVmn2SQmv3TX9ed0dUgYYk03B3vKsp+9Z9rPIM0ahy+7L+a7mV/vpNueitu7vzcA9tqVP
EBhDRQA18loSNFLVFGnxLgz0zeXTHTed8Shm5rESLyfzOw99PqYKiA4szaPuUztYc3z0Q89T5A5n
30hGQBlnpMPwEunygVBrAVVoGfsXwdBwUSB3W58lOuc5OV8DPl4Irup8QotcK992IUbSKyuC+NL0
/vX+PD+V0NNwx+YmsbRTzvkUm6lZBqKWQg31zPJB5EdsdVpqPBCv5Xd+dqmKTvfTRjNPLhP2TQzj
Yh1rKBrXXCiJ+AWXybVgrV2UEZq1BT+4BLK8fPyHT10JC0cIkw+o6sDPF2oN/bfujx8mGy5U4Jkm
JwtNsPnsNFhpLbIgt1E+1zZdgsTFt/xUXPJXgrr0GegxfFxxYb62F4HoUHElJZYRi+76q/fxF7Rh
1EZoTa/a1A2QKTQvzFKjsJgw0DIM0Pq9VU5DHuNlRDm78chH6dkfzuYkADmS5Bfe0WfTEGEBD59X
uJg1XO3HQbv6IiIReaGnVC4rPSFrFZ5sWSZhxEzeu2/4poMHa+eXONmkG3bj/y57Ng5XUrnqv6fa
PjOvBOuhWE52RsFJ6XdKeIYBcw4slDoentwk66ATI71+AmHrE8sJGfjUs20PMgxjlDmJEnLdgVpC
LfKOY0wc1HkpEmnxzNSLU5i+u2w2VBBfKYUud8s+QjUYP/BHSlrmizR49chwWNr4hrKLOKHKQB1j
Kol0Am/lnvCbPV7uwH2WURguiFCeAAy+GAR/1eoNPAgq5Gzcyi5BqqFRSMcWQfyZKaVXbOzwlgFs
TWoV2GCu+cnDgmeCLqY0zY+mKncWmSFYuhYflloBRmsJ5V6x2eHwBeBbiJ1EinbyIa6HCr2KBWo9
PSYMgKmoKrAIr6Sn0XI2M5VwVf6g/g+nJy6qMIsh2aLEE6bZkCLJtuXdUSAfWNgLuX+Nfzhbv4l2
PE98A+rg4LUvqWDqofjX0EOFTFTTwGBV1v1dDWOswqEzefjWYQT+tQLJZvTu4FE2+HMgXxuh2qJd
1ZaQu4oVj68TiKJC248YuI2NtjkuxBC0D2IEltLTcDYepsbDhEVsBAV35YwOC8r10gB5INtyXLcB
/MrKeDU+TAztyp8IS8JJVXCFpJf49SkgzKhXaJz0Dlumm8JAPrQkJkyJpvtIjSPsR5R/ouan+i2N
i9eeFv774QqjXV5UUmCph+iM8uH7C9v7SwpKddZjq8l7OvSOX2GqxQID4mtBaq+z+KIySRyDzrBf
7FAL1LPVwybGv0fbJ4GE5VkrNRQtj+7s9UzXuwTEuUyzvosxpH2ow2TuvS4qWe7Q3UjP8MpHLqK4
XxEK2RS/U2trJiWTRnyvG3mE+k+nXCk4n5/hogwZy7jqBJq/28xFhyBa8T9cJ2ujgD3hBO/aPdwO
jiDiAXzbh6hyVuC+5r1YO0+XR7MsjXbsXgrTDE69ErN4Iw4fxcFAUeoTXB/7EsW2ydH8Gu4VFvxM
zLg48f5CJo/rxKvvD4bXf8JRJYw5pVENvQz+28yQjiZqB1IPkTMHfwlymj0663q2i41RK+MC8ilq
A5Xj9UFI/16vPFFjaj3ma0Wkgpg2xBhM7hgIl/jiRa/l7JFIofiwxWHLzne5DaQAG/jb8pPMUVFK
cK797NmxwMr2ViHNCSKHnAMmfp0eaNclLHa7I4Htg22SnRhSkgkncS5TxJX8z7WoHTvhfRlnMF12
xqzwqdCsVloi+t4UWlTXTbm5ZzxWMOQmlvqL5kLZjofrQ+pNvJVC3qo/CwFy8m2oOsw52jRMWqye
gtmrnv6shBJF6iy8n8a9rQQNUw3Sxc/AcpJ8HpVywKJew7mp1pC8HTMAGBJKffFp2UF0Pk6Jfnn0
QD9wPJjVH+rRGU11dmWgp8E7++kBFP4pvq48e+yuWacHzhCaUELPsh/k7/3MVQ7CzVJfkV1Cttyp
NgvNIkRs72cxHosS+F0pgLE2UP6OKnAcWl3ISdd2C72xkkJQL6rzmqAFRN7Vqj05jBfhGkmAxNlD
s3EW+DV9IWwuujF0AomYwJk9cerVhNJ12um4i6z7z+0MDg3JXjYjgwxbMV7UorG4MZLv4VLm5NxD
uFmlt4Xl/NFS6fYlViu9EPIXxfm3ZthDzPOSVVwzQckOgXZSFvjVvmQGA9s4GLnpwSpSf1ffNpgd
XdU08gDa5i0T4zdHPM1buzsXQq+SsBYbHSa1FkW3xJp8wmgR9WtV7RsHBEf4o414KHmRRQQHEFm1
EX37+geAUzFbwmmJMEGyDX9dgd/FUAx2Urar0SoZg/BOEZ+4NoEA8J2DPtL24LPFaJoU24mhPCvQ
CPLxHf5SyBvl1CQmSGNYqSTLffjQ7rWnp0XqJLGXyhNTKSGFMsu8IC2rNSJShOow6wSWbd/A2D0X
gVYWeaXkIBuj48uBS+JnoXv+JIdSRRx7URFzZhsYrRZaLOjZeQiRiKzZYqHh3Wb7u1Ws75NRUaK3
ioX5KWUv9oQQ5B0r+U/AKQItB8LnBMzUNgPOS+VnoVSligoM6p5vJ6vdwnMP+DSZRlnb0oi2KNRQ
vbBiLNck7VymyXOG7IdgcFx5cLtPSDk86i8B364mTA+LRVKdU5NfulWCdtQqynK5OCwTW1JchDMl
qKVEKvi4Xgqq7igiLR2jpRjeRowRWDg8ccHlJBuOGavdO7REXI53YQys5Zw+YVQa2QrdqX1xffe+
92aqNLTBQUiWTlzDzwUsA7yNrNzDEe6Py0A0yGi0y24XSg7K35LSiJfEL6ddC5w5csdJ/MFoFr8y
SvS5W1EoeYsk9+xx7NfVqxQKl2ZSVRD8M67oWq6tvhamXHndwKaGeCI4I8VnEYf+Lw8fAr4ninI1
lxxHmDcrLks7WkcSG6zMfSJhJR3ShrIIszxuDu0nfkbgcVCAa5BBvSzWjMeFmAKjrKHliOmj7QYr
sTuD8vi87WfSJHIlZz6IT6oYmhn4bC5vzGIb2Bs5xZAPHF4+Bb5ajXB/X2lpz2IlKljmLsARdLtu
PDqr6yNOFVIVOeuGjH8NdUsmW00u4tier1DpwyhMzxaCqkbBOkBrIu5Y7bi+aDSzWWUdMH22plRb
NUfYlUc6Bmf4cjMJpfAOUH4wQXpNOcKY7wPc9HyPLLyhhi3+DedzKYaf35VbcLOd2rYHDwAmY5Zm
l9mQ0vhmxOGVWaYmxzjJEf0C4EyeFYN3/LKfM6q/qNRSkhqUcdj98+nQg/EfT9kjESJWpPhgZZq2
961oJDV6MxrFGZ+cTdqugc0VQ7l8FNZdqah9fjOW+CbppQzJNjoM/10nXXPHC7Og71nizOaYfk4n
05KzbQoxTavorRdznQtq4pqLGLOKktkkojyq8NYTCIx8c8eMYcvSpW2Jx5caVDAP1x/fzDEZEhxR
PIR/78xnIyECeD7m1pMXueazHmguR1FVN1E1v8SOaAgo6Kytm+Aby6x1Os6nCbaUgAMkAHwC0u6X
ULMkS4NBcwH1bqTjmeLfhqKHbsnEN4lErDlpu+nNA6N8mKj45SQwtOpu4xqOsRq54pQyjHJLLR7D
NZrI0YCOX2kbbYn6SD81hzVs8ZOhhxCF09NVfnbeglcTqq2Miosuyfn5VFMN0BUjxokF0x262Xo2
x0MEM1bcH3o3oKZ/MSeD4n1sKbOLjezwtUXQ5NT4+UAuLHN8cFOtEnx/wGJb2vlBjZj2fd9ozQyk
TRPwWot8GmsH7gOm99Olb5LasuECNqcmbIaPpt7KmBO5ISu0/LS43CXDl/JskKf3eyVZ9pX4YrFU
PChY+kIoQQpRMTtRKCM0aoAyTJioeK2XDg2oRoKlpLxpuQKNO1MVON9L9OlQc3EUg4HzVIL1o6CU
6CLdrP8BP5I1DpIDGO61r4nuep9Ic8nGISdPdVT1mwW4IF27AQVbSZB2FMxNGgW31DZHgnfz2W4+
fW1EjgI/Aj3hSElZYZOHMXy1g2niTG7+het4nzuZE9bK2ZN5ziCrICIipVeHvegtTW0hOqZoblgL
uysGNAbu8iKBQzZCJGVZUyTRGlTBrCcBvN3pS1M9PgbduXeiyx5LWLW53c2GVuKVzzJz3hRRlFrv
xKhTJmspZ10PYrnuwijU2IUhO2iaO0kawFjHHhVvlWJBesITaLRKiaq6Np6IIq+kcoaxtTnM/8/t
FAPsi/dFcpbEnlEUSUukMZcF3hVuWd4A/wF2obYz9aJEhP+bIDdEQi2GbSTvfXJ6po54Cp9Br/y9
JvWsvebzU4mE1FYyyOQi4vJ3CZjRLEqVTS7sDQZOje6Ice5yyzm3kCu+5+8Nz2GuVDuDP+LBJcW7
kwP/aT8bfVfgc/VqhPjQye/pQ80c9TpsfEwon2QVRGpWYC32tImrhlf8zQDLxc2O8bEzVp6i9D3F
rpDxJNnrEckQkh1Nt8DLNfonrhBydAPlwIPPK5dedHdqLTxjcJI3A4vtBBn9sDySRJ+nlXji2kk7
inl7KsZiEkU4tGIuzMiHMY9O7h8MUcZa4QRRN2EJFDafoVX0u/DDCnZp7KuMlJurE4VEnD5Z2eSy
EAvVvPJCaspSF8/+GUQbPVeB/5TasP9kbdIaHOlgP8CqGlu2qrskLlqotfTl3YxWVhrsJpB+QWx/
m6TkE2XPsRXsvZasLLU3fpUUd4r8p2Drs3F3b8sqO5OTMoVLDuwMuNa8lcSzLSGj+9zuQnguSSF9
Epfkr5384bfYULgr2EwWeBcSMHR1mB1noBphDKqyFyOwXwc9hzxig1N+BjICnsuM559TzvF0B1c1
MBPrq0+jGQqX0022AmYiBB+FfUgOGZ7Pq9y3xivXKZZD93/lTPmbqLPvW5nO2vGnJB/5nzbVvMES
Fw2KcCI3bHwng3GcsCKtNdnSJ04UDXPnNUyT/pmfHi/zwoGX/maZJQQ4E1E8oP2ef1AkB0IMhSte
6LnFb53CzaOvRRf2QephuIX2c0XejEopWDqCDOT48q8a4qJAsXq9AV37MUS8NOEgDSCwVR0sv0oa
pp030tOmxlnltnaizNyMbFHU8XizeQKbWMy1hBlU9Vbsam/k9ZtbwEh15Q+i5mPuT0XQNcSvj6Ah
yvQDXUWQGEV+42J4gFulh7lH5oZn69Lyj2lt2y2ho41b1ZUBkxanGyRHxLAxyKACfYt19i4XMt1o
jXNmU2KcBck+34cVtm2iPmkU/gclkUA4fh7hupDhVV4mWepbD+noR500EkKYXZFjkXyxx2ZOmNde
Fq9Mcgqf+cf5jcB1KztKpJX4zZC560FhoP7aRMK4S9dycRsR742KN75DuKoNAG6zzAl+X/L79vrk
bqUm2BmGQXIa5xf3i7sgNN1hWDKu44BWR7FcFYC9p5190s4RF4w5ftnae0ZJyKTZLieykAjN+jSN
WGeupHjuNs+41w/NrNC+aq3kMR2/e79Qlk5Jiw3JZgwUNyDoqJXlx18KidyhKx6AfzmCV59Agab7
v5gsi66VG2e56pi6WfsbjxSr9TP6SVGga3CWwt5c2ax3Y/dLVTkQ0/tcCidjDaBxhy9VLAYjIYt9
FHUyzxX7qW52n63+98j8EON+I7Ji0oprkQFiigt13OxPRU7glD1AJpvo1Il9bEBOHVYGyTNgt/1G
xb+l9Why6UuRlyLsI1jccMWMNLXfsZULK++s77la/TEmfbl52w/MAHvCKnblXwcOr6SxL/3bH/3E
h6JZHo2PrpXu3bS59G/DFxeN3mInd0Uj98UB8Q+S/oPOFi1CMJ7qIp3Ngo+TBIvXk0uWClh56tra
L4kxhrWhfGmd2gj7Q1+poQ7gh5PfDkHi+26I3N9qmoGuJjOHvFMjtdT3mUsbpvPB3YuqrxC5wEN6
DlL+jTevTNy1SLwE8eA6YulNbniizhf64Spyc75SSL7HoDf0bndybfaYqP4yFf2aNrmfI7NDa4T5
ezgdaImrbU95GXOSsupy+vsXj30TulrmI49l9VnKlRoE8I1dGQzzbbdDolTiBipeD4er7aBFRdig
kPHWIQOerShtNl2ChUGV0iQ7RVTRIUngqC2vOLsVOfMNU99eW62ZdX/JleFlC+xStOV3Cfx3Aq7v
VqUMwyf1wuQ+lP72tWukgNZhQhvZyE1mOe8K9QiHzbqrqL9kSz19JU3vsF3Flfpw8ZoUf13EITN2
ifjlivxxcR5E6MG+Hu4DNRzRGE4tf4kFrg5UkRbcFHdDDlsfrm5GtIahG41F7MVtCcsYxeHlCLZi
Aw7iOGAhjNxarnLlvJpLHyzVBne7ppRQkw9/KMpBkAubFFm0w4AEYolthL+zIlUqJlgZs2M1U8mM
XUWBL4NnCmZUBOzwngb+uRMHykU1BrkvFT5g8kA6JWKFJ06je2t6gZk11nX3cOJg0qKMQ54dxgoc
6onGUY68i9LVGjPBjLHFwSWQ4i8ZBp+TMGuqSp3anprAXBIF9icAaKZ+MmrSJ3jZwW76aTkVyYdI
2eiszj5SkfHQUfWfauXbs95iMzat8ClIchgbhl4IPhjE0rgPKz/BVvcwuIoBvOMKKgst+NTKzyla
SmEmUY3G/483NbSOW4PUtvPTTj20GlWD7Rij0wC4CEiaEBYcjVYj7EuoczRngQXEDR3hKh+65G76
g/GxffUVG29mKd0trl3XhR4W7+G+ybaYC5VI3jjNygVHgUIxnI3gy0Xa9HHMdTK/Wjq2d3aSwoQB
YkNJ0LPTCgu29WHJSMcpLvzdgaF8nPJ/FP2X+4eOsa92E+Pthkkwx7TKDfFzMMzYXvAUdK29R6mR
vL+mQZrxA1xLp8Th1mq/A+v8EFMlbb64+Hm8/YS2bwYwWj7RfGQ6+pudX00zpGt9CiGVug4uYomv
DMqJ/IFQCccEWLd8QQ94zfHSp5SLUA+audpVfUr+61nlxhfGQinqCBAmG7Oi0T3VfP1ge01wKVHk
9bwAQ5HlBM/QcOpDW6KL89oTb/i5XE9nXXNlc7Yxuxq3ZCcvfQMzyyX56oyXHMwjyS7E7Wclx4Wo
/jGe3whW2DPaxbfLT2aKAD8GZ7BGht2a0TeQgdj672zggHHJQcUcsBuuCbN70T6AfZijoBBNt3FT
4v6be5B9yJW90a4qfeud5D2ANR0ytwhqlH4ESshaZWNeaKvlAcBfpicbsj7P3REqL0ZU8kl8Ef1R
fn+jYhOXz/AkpgkD0cV8ixZOwDJ5UFW590FmuXZqofhyw7iciW2+jKNBjCXOlUJgU3/JQxHWQ8nl
DL9o8GbplRVsxGV3nJ+wCnUXGpenn6tiCtkwdFv48H9SUFoEEWiaw0zhfwsUZYZZBCBiqSFerKm2
wmLe4YJo/U3QxjQRbrJXwPhw16CJBnAoBtJ2ZFa0MK3MxhvMPq6Wdl9qOuEH4fqrcnv+T5RG6kgp
MMNGDIagtHm+nxi6glV3ciO4vXg+GJMirk8VkMuv78+wyDRumpDoM0nj0+DhqQpWTo+mQ4z1iGnT
CLsUo02NkON/KNeVumQSCDGAURQTM8RMwsrfCXQCcBOU81LvsQdQL4+G/bvAdR3LyKJb5b/KYyQ6
GZfchGEJgoP91yhHlDTSAZW301vWd5FypKbQmg02osekqdF/rska5hnzW1zt/xnFJKyNVLlEqgDu
phphKGoXu7UJ/QwH1ChBC6wA4Y3LIZdGA6FDWEhUjMxwmPrlOpDj5cK8lRKR4AxmKVX1UD/zAvh1
lAXz4v4nONnC6rGMC0BRApMNQ/12KW0ZZWQLvHv1HhoM+lvIF4/pmVn9abWk+MUS3El1pKw4FlD0
hqzCionwTfh2UdPftTW2kKV5EIAsLONRyzxmgZBfU8vy4Lu0OktazNhmrZr8VHcXZMWn9xQKLyeA
8plXPJFg1qzzm9Ey2osNTwA1leUfrVLw+aD9L/LB4y/5Jt+c44ibRFRxAu2Kyy9R1VG945cvUuUI
u5n9nVObiPKhhbE0w060a6Axr61MvK3ih8ICtTuDwEL1h54WGByQg4fmiIJC6tK0EgSqKDGcjemK
KmQ8YgkQ5q5qPpd4QdsA2xyr+Zqpj8zsco1jY/rcDENNa2CSj+LHVAjUXmLYnoMeUb3xqR4hSlVO
0y3ElDPwT55lwsJKIo56AlNHAp0Y7Nb/KBrF8XzhmKfQ6sGH8vE0ruW4/FGs4gYCl2Dvt9iQoaHl
SLx1C5W83onXYr9TtUFobJJele6ARZjFn0Cqv7Wa5TtzNYm2IGXwI+WK6HStBimg3fa8hbQXKCf0
qJEWbcjwkWjId1vVMssqbma15Y8pGIbH9kMtx55yXFCD3JPK0jwNuPCCio3qvP1J4BmwJov4jfHb
cnPk8K+qM8zNgr3JX0Wwc3YtmXcfxCy78uT4qKti+g7QNDHPkDixZFtkZQR6dy2nZMM8xgtYpgwd
Ld0mdL39NKXSJhXyPNNL5gRr3iqOmWlhB3m/Uha4oqmxTlbxJ0VjtoXJWlXSwk4+Mt8ovXeSZpF2
Egdu/GkbWVhdcB3FRCdL/7xeI6JrTphFfFu3OQAlRRvLhS88aYYKf2f+X5KdSsFrmd63vtkZUXec
EeyFfIOwmBVnTcdDIpXv9wIMcFtmUNwvMpiKkmqqzI/7uogFrT1Mlz0L31xptwoqpA6KdqmTQAXy
FxL+Q74CTDqn3QyoM5cVi0LObmKsQA5J42Gz9USvw7lkO7Dhdh9i3Vz7EzQoRDGwf8gr7895z88Y
MpmOS9TS45+uqiS4yWxT2yFwsB21HWVri2MKeiKSDNgJqd1kPRGpI/s7gol+8EHWvT9ptVfMvBpe
ELEWtyR1E1oRLETX0CYm1LzJIT0sbRLE8MQ+hxAR0NtQ2hC50+iH6XqGx9NwBFCQtMPVZ6lOlhTw
E+AlRI+zGGA9yp+wWBtxiiv9XiZlOtDGn375PnLLQo5R8fFj+pnMd+4t97b/GQbqmhRvcft7T/r/
eClSgHzu1uiCCXgTLj7a7lSVG0FQgzIdW0E+ed5VC2GwePCOLjxu/tpqaAxdE+cELzXqaWg36Z61
S/hIv04gwZoJBLuhRWhI/Bv5aJZD1U+SGNqaEtDDT/Qo1+0SDaT6EUrK9067vw0016dBrsb1TClp
bEBNftGxKXGKpero/tfWtdKlSpS3KUyNuqjP/iJCs3rbDvNJh3M9V7gLGmAGoxi9ya0a9E/+sqfd
DhcyPDZAuny1Q29MXoHlcEQSEu9Ou1prYGlaqyCraZ/0cLpyB9S5uroyItlkmHfR85UXvbGw9MdC
pWuLTbgdEydMVrhe1QoDyQBW1fJ5901tUuqiiPMI5L8AYkYGpGJESq7FdvVeEY/7dxUio+jT7ruI
cD+pxnP2v4q/wWoH2uDt5YKb5ctX9X8qTJ6WYzccUt0yq7GBrIMdNN9Eh50MEGwFZg6xHIOu89kc
naQ8LpdIavGesO2knDtXxHvaF6FMWGvwy3pvPcc05lNiEW7xQGHcyl+2pUj/QiYa02jQS1xVBj9F
X9Q4/3xzeZ6XMKxs3GWUp40jn0576Kq8j0/qTobZO+wBnAO2vv+b3c+JdqzhtZ5cXYiOgBfKr+wP
AlESD+HRE+MTHhoPaR9knf9o/3b72hFO42F7t1fn1jh4uH5x+205C6Q5cfRFpZOCS6vrgjBPzgMr
PGzHX+1y60i6r9lAZqycXwi2Gdg3rTbTIcF7/p252vpDc+4VHt6JMjkv9UbAavFYRI7sn93z3FHS
4MCxx2Wc643zbVvS12oL9MYP/fg37Hl7AiICj68HPSNQD4YFP9u8D7em2+Tt3XiKBfbnpYcR73h8
OI6zQlMtbaJsc03MBrEaeYqDdRwaoJizXWaC/DFWw3fTD7EquYF5ReCxJ5QnGeWWbYFCL7mmnKt/
7RNN+sIplXEQaad7GlkwcPjU+8p7UWnmkgFYOmQ6nKWgBWCNtdQtYvUl6flVeV2mUG1H0YMggcX8
ExS6SwsQGIuhGo4LcFp7esASaSy/2UP95BCka62kZRm0dWAtn7NPwR8APKQUQkzuffelA/DAKkBJ
L0qG6NNGW8oRN+96EjO6raCrOKjgGR2BIsa6kLNd+cHP8PDdNiVJ3wT63rNvnRI0udNiOl0jY3nn
WoMV5QF6YRROYFUNSik/eH8QP96YUcKAy5DRWx5bsb8l+cxqg9iclog9msUJljoG+IoB/bgipMgo
U0phcLPsldMdzD99hVhexjM87uSeWtUJIEnATYhgh9PTl/etmsh013vrLHxR6qZELRlPy70pNp0B
xaqyW6decB0HZas4fh+Jht/Jp5q3zoJqIQmwbS84fRa0s9AgT4VOx+wnZbXdpZc2maUSnTaohZ9O
HYxvEN2Jl7A2pZ74wSZJN0reqwCWUuFl3HXscqmWQDMVOhO6SG1hgkqlOojLgSBEg7d+3ZOwisL/
6Is2YQUhjFtr9C/KtvIRYK0b1HTvrta20WmS7kIHPne71jrULgyerx885gjvLylftIcJrUSarimq
1gjw2rvXszMYPAbk3BgExC0KEdjX3JnbO4ZYeLvk2QfnDTzjojBnC+op9X0tqS7M0iyGP3kPYRPS
g0aacd6iRzXcLeADDcxBrCNZCSI6vtyhfkArr+qoHgSZ9GalIC2AMEGd8Yy+MFyfo31XG9klbfvk
SyFSF+solkWevQWAP3TqpVl8kq7MLxhyXaJIluaOZyj6yrnUpwzTUODIRSjbhUMdLXan7YtaBqFK
WBJ1FfCn2bDDS8692VxrdAURW87R5re1Fgb3/N+m4iB9bBawhJwjRic+yFWz7szUjLF5F6JbCAYA
j4yclMj2nRVhZ9A966wn9Bf/gSWRq5Sh8fl/mkAm+nLZfH6n96OL5Q7VNx4pgSEDosBJ+Nqmsvj+
zIfyj2/1nmEIPG5f4YfaCM0sNBaVP6uLDLGPPPCx4amqYXx0bIU/7QnGMrr0WZEi5tDJbRddmrUU
1lS2FjVoCFjlAgiVnc5eDIJkfluGirWqbgoCy/RjgH3WdGD+cUElyEd3CKLmg5otmgdj7lgbkThD
erHWJb+6Ukqclor0J2euEl+9TNZR0PLwHRHkLiQqfsx0YfTdUjtjV2rTZWdVldb0Sj1MeAWP/DXS
XHBZ4jOEBSl+O92d8Kz/lVENrPDTCNK/5aAG4WSK4JwrUTv2qHvQVcSLe+Yg9ovUXU6PPRBkLsxi
PyN1XmzKUTF5PHae4L8cZD6NBGzNqXUqJ8TuEup64a9x86XA8W3UorCk+lrOeWGTH9ax2nFs/ynq
r8XSz5xQEnlz6IbJ/rreSV9E7on7ZyTVWV3qCs1gVzOImP8Mx1+yEOyMnZ/2MJuOgoiHw6TQWoUd
SIF+A6VcwX3GMlJPaD1MfdAkQX+rlDM7P4aksMDFfUVV2/RNRoh6O76cQhpXdLMO03YifdcIa8bL
r02P9Lred/OJlADBqMT9EHIxFpQc8+xtDSkwfp1AbR+x5hwx9iBlg06JEUUqa8pu7+QFQm2NfyOU
3uHULHAe0+FDGe0HpmoY5GV5I/NDgyCH526wDwg+ADy5YTG+orxQ5/ObbB5TSye58J9l1bwV/BNb
rgtu8Nkxt9TtsyE5llANAfB3z1zCrxb8nx/C7CWMJHTHIuDStN5htmmiB43kOC8a51/vDRvggUAt
CYD2KFdP0zuxJZh4fHXEOMihvYQGhDSvqep8GQoq+hAkm9qTXcdMIO2O2qIuDLuzYVduOw30Domb
Ojuasjqu+GyaE5M/lJWG3PSwdPxSdeRaEqRCFu/6xp3PXvn/eM3qxNeSTjfsZW7bLooET7201gyG
aregXBaGb40WCPZWEb1zhQECveWcYYs4Y6q44rhPbqttKiLleoKhvzp82f5PvFwn9fbCZnwhlPzl
TDPSl7mGJUqfaQd+gH2aYxy7/KWEmWpOuPhpgi3Jo9dEHx4ASlFNVcSI9kfH8hf38SjoynSxvLBm
muWkraQGaFqmhwsFr6+Pw3Gd75dM3/qYg8lXvAsG5B3RPisLWpuKW7/rY1ANOJD6EZSh8DbsDsb9
ZqiBr7X3RAGubvKxD94mz3Bp9OjhY302uNpVveKicLdmFaOL0fL1lp5AO6erwbvklGNEQZSwWJ2j
THeMVACgOt7RJSBTfHUgd23Gh16Qm0Vgz4KtoOkSAgE8NASXsH/r7D5BJ5jIlRslhvLu7VLMgynZ
mVlWMk9wtcUNTE1XmidepdY0HJZ3DOppBcDC9jgUrAhxk/7QdR3nFQz9tYbaUihnC3BCvrA3DyRd
TvmwhezZlr1NTN/uWnhHb9ztvuSTVtdM3T1hiehNHGJ933W/b43BgI9B6LOEFVhCaVcmSfnHIxiR
4LDAl6s4m0F+6g+Q5B1qT3gFjSSdzW8hOnmteUJTm1MQ1Bd2zgQw2PKEuZ5e8MFaJEaiPlSI0yDy
uonzVwnbr7H456cWyACksAh0YQYLo10v2Y6Sr2UbVNMXYC++IPJhHsI6XVoj9W85TqfpXtTvHTcT
7b9c9VxiC1w0ZVaRKxhpqFWLDFmtRtpGhekuLjdY2t4cd+pOBaApe6m/QLvJY6zn1GuCYnd4HbRK
hFPjTGTPngUtFTvHUkZSHcTGzses7lnwSatie0ppkL8GV3IHMoniSmfH88NpzqzcAuGOG91ATwYC
H0psryqGs4jToZd7/MpnU8bk+qPsDFGqipAOBj3QX6SUUd2HO35ZJYm4SqnsvqmFmMRvjaYisiSA
gFv6kJT+M/4WQy05iPAt3D4DCXn5DJzgXg2JuHNMxOofhtOniqdgQCudEp38PazEkM5AzMNQ7/xV
ER9M5PaA1Ixhx5oznd8ZDRT/YWyqyXJN2uBt8rAraULDXQQlVh7kdSIaH10fNyLMrbljmZddF3uH
ahDb2wbeQ/B1C+PvW7ZUFXVcWRYimToIWIWH6lmfkwsYwKKAnOVTI0+L/8+5jXDfKttx+cCxoVE9
BkuzNlbvXkbfP0nqsfPA3Phgr2BVwjxvUNPB1JdjDhg9fnKkAibO20X1HY0cMdQ+6Yu2joVo/wBk
beysT8GWfpKth3wlkK1hI0J77KgrrW12oTspQuKn8Rs4GpzF84SjMfOPKnGC5fchty+MXrZVe7ul
O3L4+TfBotjw+uBfYwZ1Gzr3RsjLeFjVxyP+y2v4luuVcvl5Ctb2WB+YUZx+D+qYifGrw1UHIdxS
nHPdtYN3EOHgTMVmmtQk58B058lyFEMe1rJXqFCtKYdw+aB4Q90LO+bSc/+AacJcCLB8e3yLbUmT
8AhWHU42EYMSPlLaEzmJPjdlLzw1o1frBR3LGj3qK1aGR8O9Q6NJaag90Gep+aQz7IePcECAOWu9
kv5ddIspt3c0+fqTw3orfVtdCl5zmBuTHq9F0NMwNJhI6YDTQAhZCyguX82ECgojuPMw72CYfHBe
7ksg2ehD9PD8HPqyO8ZRTeX/rIi2Ralgy+AATTfZI7XiStTJd61v3p9GE7d2HG7M02us1ahU2647
1mi9Cfr9FsZ3yk91RfphFMlWsPUWOoSnhroK09xSjkmeZ5PG8Y/P1oa0bHVl2f+XyFPSM90El9Sb
sXORIrdR019iANrtGP5NyC/pJ18oWrjw8Y82p0NiELjBM0WhUOovhaNeMj4sP/ineoKFx35eJtjG
HZM8OU6eMr7MgtyH7nUQDy/19rdFuDCN4Pfot3GTTmw2SbE1F7c5FQBhWRspxqi8lP8PgI67p3UJ
WGD4dizq85NsuBf2AfW0SzNBIC+MUghi3UpW0maEtK3wOty3gk7LOdY870VZ6thdot9ApohYQ2nT
tRKSoDh7TY6wixbftYaYzWeGPXOHGK9RxO3D/zoZwz4W91wnUg1Bw7S9L2Lp2iPT+yjrgUxJXjTZ
4lTwTEmpj4GGlOp+MZUfIakfEM+dgGwBNN/GJpk63xbHHxp1AIjKSg1Ch5wgLhkFv01Chr/IZO9Q
sAHn9pV/ngNgiFQW/IwfBYLReX/tnIBjsatBR/ztPDVnzHWmz9rTkoM/AG06b6jre5LPqdyWvpAF
2fg9NRoHifm6v/BgjpS7xHY/uOXMpFrXREmpGDy7ZiOcjmFqFqMAOSup+PH6myMem2/jC7fjqZfl
xCfYQbU6xrMnKY2V5+XkYeNjCk4wT+puCHW2Qjmux8JqTlXoQUlyHhyF1AN3zb2j6chrxoLozpl+
Ou3fM4hzZdAs2kYPxX9c+yGz77iTDypm2ndcnc2VJAyF984Dq7XY1AfzFU0vRha4ue4PhaAGQ1mi
7FoVkkqWn6fJO39aofbLVpCnHIXDudcmcRCAtENy0fJA7cD4EZ8Sj9t4CKv2Vcl6Dnomo4MNgIQV
SjdBhuZ7OKc09B9bhfROShlXesQ5RJOqD5woDunXf9MUYYfYRKAjgnSXcRikqKj3oKdfC6IsCzhe
JbAhLfMov71pLHFfm9TKZP4ISPoGSU3DWbOMKY33Uydedsp8LbI+DIDeYBKyCelIBMEn/d7iTd5d
pr0v19To16njSTDPI7K3ijdFOEJIxkIJLPkxtzDW5QvWgiBPQqyj+7VyxfRvCnSpPyEfp33dhuIl
IdJu+jeauGMHrW7ngfdPAsRpG1HDTlqdpjGJCLw38Yk/ovD+OHvZV8g9IR06Voj3KEvY8VfcQwv7
jjfvtWQ/m3Cg5yL3/o2mwTmnjwEfsh8VtsRrSL0na/85agIBzJYNCcxQ1OO3uxEvzhJvAeKq6Qbf
4OP4ee/dEmM4ERbTFpQb9P+55RbcqSOIGkVA80cuvjwJodAbdxOlr/Dt0L7ZOVq8+bUVdcEE+f3U
u6m4wkzM0o2efXNI9vLVzPCuyis5P3xZjHTYz+5gZ5Wg8FIwiho6oTEu4EQ52HbqJYX1AxK8N+ep
lvTI2OCScUwcGpuCCPk8BJqAaUWB5jP1Hy9V7cdnHvSW0f9yADS2soCPKCo+2xI4TYWMmLMwsc12
lkXT24xkW7j01/I+HHQ3gjh7eGb8qPSenL9UHTK1++BbstXLoiHv5Q3x88BbSbqLite55eDGNU/+
Ph8PDC2gFhKTanmdOdYQ/2n+AwAdk21fnLkYMK1K3NeiUX0CyuNVjM/nRx6Sf1ALKuAlCEWxb89u
8U6Hxh6cQbRdPTnFLPnHUUjEjb1TZI2uG/YfsJfXsf3Tc5/rBllY4YDmvNel4AhBbj72AJoUaRhT
5Q+HzviYY1cvtHPbWJ2rKEXQST6UiZZiFItVAf8RUJDvBgu4jLwKJny4pCE3Aq81Pc1Ue/ADMS1w
OJF4lfk8qng1Jo3X1y17NaOBNbx7PlZr8Zixnxa3BZq+xgYPEP0Ncn1sboy895PBb0ISrlv06Da8
HHGsckibMe2s8f5hwOtKsRLnFPUvA19viQwBa8n5J/g9kf4zt39boayuENoqS3qxpkWWk1lrWJDf
fer/UI8auXp3VDSCJjRv4VmDd0HVTb90RI0MAjgGd23Zb3d758DIVUQfvCNdAlaD7GYJwU2gDOhc
K5y3R9RfMX50vdDZF/LeDzqFbUNGdDsnu2AlIsq17tdB+Q5fsov8e5sSmpo71v2jyIFgbRQIUCqB
D2JSboSuscKjfFXOGjS+q11i24des0KYf9F2ucrPnEwfZ2NHnQ5k7+3gffMVvLww9yut+LVsPhoU
uphDeT/RgAVisRiCbWluHfaADILVYqo+ipJ0wxRpP0tPfO8HbdtSPVCnz4fDQDgVsV/z2ok32ujc
jv8GKM4um2OOB3H5X1UPARIPxoulMsUVSx0YiEANdoEU0INUSJZ3P5JNnE+svKZRKzmubfFusu8P
l9NsWC4oNXoB9YixKVLyENOFTBbEkmGZeYZ1xSIR1kLfSrA9UBh0CywT2VtX7SVmER712iq7nvUj
kCf1eP4KbE4uz0IAbA2Ze3LsZb36aLpX1ZYmRQkUH889fXU8JmAPtKAt67p8S6BSyufQ0DrJh3bp
ZdXI/6LCoWFgItOv6FL7q7xcfem74A4GSaUHmJXHOwHbBoN5N0mtf4NaVvkSgZAM6JnqymhVfnVD
j+jJCSsAJzqUF7tTXt2geZD5EAp7MI2rjsrF5oeK921InCvrw+vY5jEoxSBgszo2MVeO7XwbDXRX
CHvfM9YLdFT/dQqyx9chjIsR8s5EYW1cG5lFmloo298hbG3JLp5/tBFpTJLO58sDkzeynBWL72K+
2lV6pWTFy4SFEVGtPT29uLGGw+VM+YKxZ8oe6RW+DUcc3OAdUaVJxV1br6SyKQh0soR0Xe2oiNJo
vYhYM+uboFSVQCQwjog704hugPjnSyYQ4+7MONvTD8U17W1DVX/MJyMoaP38G4wy4EjYRRnt4acR
vcol7IJ3HEHSG4FIdkXsbliObjQkq/WlCXGvyGXib+0VSIrVvfea3QLIHW9fhCJkUb8oMVv7GrCg
hIkUdWINnjXryiBSAlFWvIYobpEDKvNv/SISWNAUzJB5/CZB3MoDNmcTzVo4l6H4OfGU4f4sBiPC
vOWkBJAnKJNlaARt65duO6nP7nvD2XwEIoydVjwC3l2qt/QdtGYP7F4mUDbT+t7mIho7sE3DHNki
4a5+2EvYh3qZgKGXBHBWhD3fPuppjmLDRfNUlVGYp5oGQ1h7Ek3T6xY4WCDJu3mKXUAGBgtUtV+P
yIggnnVOkpgr2D9zJEO0byO7ayyDBxUSTgMkNAb/79LEuJkVWeUBsFBzHcTzSqnTvgecj2xcm5zN
OnT4gfax4z7sZAcmh8ZRilbBYxujK8rDaF+3UUcbjv5ynpSoufeTzsL+89crMkoLmjTrkPPetb1i
5JGdjKXywz24hSJk5QCOMW41J47HFHP3W2q7CG4lM5XHya+uWRQRPztB7+n4FbKatlRqq9hK3btP
sr6Up12SX0+8uysJoqSF0xHtnqZphU9Hsdg4AHhP4p6Aa2c4TyDIR3oe8f1GNMhtGz9VeosoG9v5
GLqG5lSJNIoVdN0SJ4ezOPuiFn6AWgTeL9cZqGDsgI1/wSXTWFoKCroL0bjIKz9zSF50yYq4wKhP
4qhzElQrtaldxRenS6OW1Fsi45hdcffMq6JhmUMWGUw11rybL3rLEs04EdejlQtemv1thK3Ilaqa
8JGZc0ED+7Dt9pEYmPg8AaN0zHDlMtrEKhI0AgkICxd0u5k4QQd331QF5eX5ox9hOR2PFAX7DBMT
/ro3XRinQxuMOoZo8NybHaIFlP1Z1HW7oZzNTtVgbjh3g4jJOO3OuFk61KJsHJ0NIJVPvoNeNAbj
NCSyfZHuVO+I/pcdpbtBe1r0c3HFwkRQjLdX4cUl4Wxd9CokJwslWTsgHFaYA2gbWFtf+LnJE5nq
ZT0JPlrqlfYhrxZUhfA8M5/kJ01K4ff5xlWkAFNJAdIniYLoXgCqSJFxEfsY+LRyP/AIMLdXybNz
XPkbuzPiv4cuQZ3YUWrSNyT50ZpvDqG0xOSXJu6JdAXuueizrShccKhcPyOG4nMptn9XSoJtKP8p
SiBSTMZ821cKT//2zuL++nkYaHuJ7WmvGtUr7jBn0mHee0F4kbQGw4CxwAWsO/1yA+89h/QH/ECX
zYF3zJCIY7I/sYY9tYWzpa2Lxt4+YYiMf8swnHeTbyYdLjJyFfxpCWCReFbH35WanMKMmcKFgV5y
FxvvvrucWSHmTUW2Z7fB9HWiCCG3tjRv2JVmtgg9I3gqFFOtWxo3XRL1vDvW7YN2NC5OrV8IJu3d
1mCZ+dB4JpX0vOgE6XiAMMUIbOvGjr8FzvpYm0ghUetAD7aUPAPeEUvZTdKTzc77DnXam9gcSKMQ
Yu/FNSo7SRcHWY0ykeENoy15r7B8Aq33+3BAm1VK6gClbaD2qai1o4XlHYgWOnOBkI7yR/YUHwye
02xX3iCh8xv92GTtBRSyMRSdYUmANnFvaQrWbHUEHtcAe8Z+PILj6e5L6dAVvrq5nT7Gm9q1i48X
U/g+diJyDZcFEYE0N1Yjc4G2NHHKn6gIkbtrlRgufrgO6cuB1KMKHa4yGH6lb9UzDDPlU6w5Me2m
zCELqXdq8HDQ01d9Ua6qusSRR7KenuWWuyf9DGJD/T26g27Gi1j0MItq+luEVMuBHcWRko/pY8vI
YQUXOzzgwRmvz2qQg7hGXBYuKb+EDdu/pZ/THSNfHQgNvb69vf+Zo9Li49Ib3FtM+yISCMJQ/1RD
/LVZc1pqY8wHk+5ysk6pmJDJkZLnqJR3sONNtfwykn72BCOmHH0s3UTLF9eSJqQ4y6L3Z9LVB3OB
xyFTVKruzMnuyBlLsx9iCb7+Y0a8YOCpDkO9kYBXS4LSjX8xPBvQjez6r4n+k6zdHnQpVeGKXkPU
E8nR4PI4xyaPHEN32iRwHYYDYLDinIuVnUDCkQomVeYBaqMQoh2dskP1Rc81GOk3PWC/T9gtF6hX
OZSMVC/KmSBUoiIyv50bD9sX/fLWCfdJ+n8qtpZYnZJp/KrJRRtSTomFmV4skO5mZJaHRMVCl9t5
Ku6p654ViE5dpMTSYAVD+STLpPGZ85BNeF1RFfKM88fmit1+N/8E5O8eMgJvhE1AlVVlXn/FMo8h
EXjMJdYYbWtcau7s/NtrOX5ToIhmrZyppFnRbfU0bKgSP5yGnasSgXtwfVfOZckg0zCQlqp0ah0y
mAAvpcj4/BYeR9nLejKGr+gvOGDN+UmwtNmQNgXhrsqM1EH+bqhe4lmedMu67zJ44yERX+r6RaEF
piRQMYNL9jXG3WPFXouQy33tVPWYAUg74HC8i7YOuuj9RXuZAXm/maYM72+Sf9C1/DifE6O0SvQ7
X2C1LQ0GB/sBLY9uysgDLsfR6X2YoOq9W0IaETjYJxETF9zyUQaX5Hbhc3x4nUeqmwj47r5nGNKv
Oa3WPSXAwhIIJvIuXaR3BFdImIb8xwRXNG4yX8JFaoTKjB0brf6M9BxRnYAbwNpZh+pAks3LN6q5
L23ZmfAl9kUwZwdY9wBUIYVWaJ/6nzr+qlhCtMn23KVuvPy4/+1PeiulRsz2ZWrDn0/FHgoNnLmQ
ju41Y+bkz/LVdnLnCr0gKX63FNdOKdqXk3k7S4M6E6ZvoZ+1zV/Vyho0aSpQZvpGIIiD8OeQW6tM
IFDzWhYbAq0SrTwiqlww1iXW5sTj7rRDbGtydGAXZCviH3KxHiwxMbd/gH6d8/cGVRlI8h6rur+a
Xw39jAMMgPf7YaNnTR7IKBJ/tYntrfVYU2zYgDNizy3vza+UnjSSaYrjyyznQO4avZ/7vr9dCKa/
hpv6gbq6gnbJgswLGSIz1fKfepE4qM3r7U1Z1Td73EePescchxC8RzYIqCBxhG+KMJ+yucv5ZSMb
QceSZbA3XB+YVALjM7PrCWnFUCIhc2wvHRnUKYOK7zE/oBe+WVNa6BG1x6VpYKtZWduM8vikjdL1
3yB7x7TxxIjokqeKq35bTCvgV82RqKLp3uhBkRRQFDf087gxseYZVio0Y/qWzo3zJ3rNEfZ0Be7m
/yPTYUXfq6nA0mIZoYnSwlPIVE0aVvOBsH5N1Y0PgZqLRJL0dqS+gGc9x6ivlHO3EMfwnJlIHNqR
o9PHlZTuNuzfrRtuWSvGtxtbNapxnXeyl4+gU0ZEuiBC85jAh0C0j7iKPU3vYHsRUpwrS6u8uWfy
R14TagFbN1pf8wSdHvlUZ1dkIOnfQvP0jRggQXBXeGWektLRpG3vYRE4hbpDYLd8esl1jy+n7xW3
/SpfcpSOHtLG+ltIXkJjrV7oMlx9uxJRsZzf/uupsTLE3UdXingFLVawT2bXtVTZUix17MZQu+xV
/tSDRfgqc9I4Z+IVqVUrfuRcw5v2vLYyTvtMJSptbvt6Wu6ufaCMb43dTCcBFhpNkDuVZocqwzI6
z68eyiSBXb3FlOIh5fKgm+FsddtU7OJUnNoEBpSXAmF/27gh4fXTow4S0HLk3uUg6N4ltQ4WKbbT
Q4S9LLQ6oHRE9uHvBEsd4fXOy3NC+Ey/6OoeAM9aTT++12E/Xmk14TQ6PdQbgixh+uFuTml0ydcq
hBCet7MmrLn5KM/zlQEvsF0lZ0ocInrnLZkGCquijvzIarh7z7HeSDhqhiLNP9CbgmvC3aaHbMcI
GkAyMoyCrGbTiEtfeguNxEbfoa3qPIsJH6bHMgYVKE43nRkIo6ex9Lufz0FqG0uO567muh2ZN/cF
xpnvgZxPzprHSHtSz1QX9IQBUYkBHPAMPWaUqDMXP4TGqgoTyn3XJ2557VGMtzyvWrxWihS1v5XV
PCG+OSkOl5xF9ev1Z2kpslRYopjFkkKk8uVc126ra4hJwTERBwgi0hMN059gFjfvObGuMt/XYef+
uAim7igWyLF2c9mqPlRYuWXvwOmnNwdwRPGHA8biZKrPyf233/lnLAaS8Muy/awIT44d5PwvJDRY
qxTmrzg0uj2LFjDUnN7AdXzaT9eJJYaNQt9PPPl3Xb9sMA2+RrKe55OggUZnZQV2atp6Y8nyYXsX
HGaorN6iuwQpxAR5xykB+2w0/pjfQlcM7dgeHj2zOrw/aQQp/8B1RqztTw3M9A7mPYhNXoI2oIvh
Da8fmG0hvo9XL0yrHnZ71SlyEmHIJRgHi2AaNO1rrS1YbuJESRUnopl5AvSXs90SyCOLGEtxUilc
UiC+w8Uo8Ktm4oqZXVtPz1HXm1BwZWpYeK53MZKmQjga/TW5/q/e5POF5BIK/rZ2Ao5tCER7nght
ZJiTt4z668pX1CXR3dLdTIk9NsVX/Lk9ur01N2OBKH7pmpvlD+JC68BPcJCAxz8EC7tL8tfvDl5P
mpposr7tla3nT1A8wWllri/sCRqN+UCCXD10Fb7KoQ/q/x9rGyMTbzYCapegOFyEmvrbIyQgqqmV
cJihgZxzrRKyv3EU4JC6JLD+N9p09RDYqtSo8P0gYUX0Y3KIcoiTKG5AYBRvb4o+8Za+SNhnKrOl
i3zx1AUrPf54vVH1TjZ4rYM8DXFS9JGZFQk8NrevrjC8C4GQo76bNy5y1ijeBa9BchjQERdU75yX
b5My2r8GqH3rx5bST/zm2gnjhCurdvEjoOjVslDaQe+mF58ubI5Bm6w6RiJx4UNoL/XrfTkn9fN2
BEEtm/O32S/SYKrslaEQeegyNam7ua97MKpOoyEpdmk8zYhmDgv4108gES2aHQvXUEOVzE21eMgt
+B42b3laf6bc358NQ7kwM13TWM7pPgGskDanV7vk58UEMEKrbyK3PNorN5BjTYWpqHGGzRczdDQG
90Xwo/zbZgdFytH+5flZ4aLCPouWPKFiB9n7KmfNA3UUchMN67JsQVAZ5sIUv+PZqCe4zTTBtygl
fV3A7w73OSgEG83ui2qCAxb+uBtj8f11lHJD+9gKT8bLHa/vHZO17Ke4Th6Lr/08RnpJHKLrL9Q2
nXr2YeJmV/bcv34PCQALcBodioVYPO0f2ZyC2eEegT7YdS6fA2NAkcMGQPB57vtjN9bVqW8NXeyL
YtEZyPNBXF39NV1ggZLvZITXON6yAIcjugtJXQHaJGtmju+mdkCnkV56Oler1ek9T+ROt5EskaOX
LtIWwSSnaugwxUdZN3XD5EdcImm1uEs+lyf1es6p2dhStvpbmvO1XaoB/w4nWW24zjR3vE0btnrH
LlljYizZGyYyOXy/ia2WZM0wT/NYv+yoUWpz6l6IJjJJvyEUBsQNFIO5ujcHiYGoqcAbt8uocIKc
DyE8O5acOp8M2CRh9R7ZXBEWWLhBIazM8nNrEtyyD5pWhwks5WT4gmDVeAUZCOP9g669xvQekXTi
wy4MdN9c90BVsQvQrDmBBjc4BON3cB/0vtvshxNVUENEktSq7rxOE5VHtI9jMMqn5TVXW38os3Bc
yKKDp6Fy0mkchRZfMSANbOQGpGaul02+J/d0hGM21Vqqgbcn1iTbnwx58HjG4kahbli+y4tIPRBT
ZxEwVVsxUwAuxi6L26pc+rrR2e2oPRmEnMC2KTHBitGrA4D3ww9LlTbABimi1biQ+XEJj17I1bjC
6abHV/cR9yUCfl+8zseRgjffkDwewwNrOClr2BetxQLF798YGE35sktzE4is8HZuK4kBDJQMix7V
PHrzfmhS+QsP8ps7uNagmh1/uZ6nUTWvqJA4kqCsWXCbKh2SlnAKfcyBLAEjp5qyCgNhgtwUho8J
R3xrkX9ehxPl1No/1MX0HV6v6nW+9244PSmJGZ6/aUEJ30X4BRVuIxRSuZgtl+BgN1Ykp3/cKUYE
dVYOhKIXlxpvTtKVpvXKQ4IkjE/xrn4k4udoSkg9ecdZbuXRO7PtM7PXD+1KBUigbSXrsDqEL9fb
ESfvrhDzaHoNPWbogUn+9yY0gWV6jnUMGuokw06vNxbKt5PXFJ72EpYXCVnEgtAHLK3cgRURAHt1
0zduJ6D3Bcv0OY/7aaSXYBgOT2hpGFY0+kkO/Q/UwZbaXdx+pmGC1xIx1eNFE4VVFMg4/wqvQv2a
yiJU80DZPVTNHtC5euM7Et57nksLX7jSgioezr1Im/p70IBeStnGzQkcL17RTi+aWNdaUXtJpXK7
33lEKGn3fBynERa/jpzQAAYP08lOzhU1w9z1ZgrALBl3k8QQZB3p2u0+hmTuW2FJu35p4r8KycQR
mvzt99f/hpMHEHSC3xdx5dLG9mw15+vKYIatfsTcNQ6bAlphNyzxyC009VinibbbJR6lI37y1uL9
NFmsXpfsZ5msZ1Ba5F/nRr12Q+07mHvmcfV91Ee8BTLvLZg4TTbDbDenQGGSBi0CJK9G7Zr39owf
J9NpNQiOIQVo4Bdaoc6gqOrLtumWIAWCADHV7jdbPy2qzvVwVp5rx+w8yjYOMlkRQCp68GtyzpR1
L5IQuF3/jiRAs0j41Oxb4OlXeu/dQkCjdwqXH1Te63XmzlCDKHPW3r5aLJSFSc46BYLQj+440zmz
hrrZHcEi8rAcCeBFr1crWizZ1aNImoaDEaAYZ3WB7Oh8El2YHAmsJAUmhDhp9cPV3NbCh6sDUiWZ
l+PeSW05wMw2WPoMYhMTfOv4a3bAjb4hxdA2TUTwyzF/AeeW43FL7BokiaZUpQYrWK71oTZAhdOd
yDxPw1ypNlTp9EM1FFeVvqKPnUV7pzcEW0ZmT0sLBK4YFm6on4M/ArYNQcXrfmg8oYZAAYa7ejxC
BWngI+Hs9RBmwp2gSajhmYUUTEPdyvZg9vKYa2kzNbxGj1zcegK7BUi4EcIXXSamEg09dZPNkPBN
L3pdsdMPfKjYpo5jU3JndjKii8Nf3KudH/A8amc1ZyS8i6080an2TrqYaXEvWRV+XAborn84+8Iu
1+lFBDR644kwDqDnMlJT5rfgQxwY8nRiOAoIxZoLIKWMU1rki9l6e4iK+uidvdEdP+J0Iq0yov//
TSMwmKHJ/XJKiTZ7mJcQvMbrpuyEKzxQTgvAkI6jvhwmlHvPVnyRqHl7Ehc5zz50t7C0QLx/7Lhz
RCtB5X5dE3Nj+O/Yo+PzO6UV+TFcI2uB42kDV9TaHtJLvX9SMHAktuf4BvdREddkPXCrRJ/CVE1y
peUcwdI0z1/6oxpzhs/Q/OWxcgDChdAEV3DMPBb11F9bbm3GhSj+VDiemClWrz47NQmIRaPEUAKy
4MUQ3cwcsPLI+lrhZn9LeZHxmIX23a2luMFXUQqfihC2ANkK9+LXbZ7nTK1AFemsE8rsMsoJLSJw
Dv2BvzWzIdkBithyvzKjbz/QIuVxJI8humh0692M6yzfhLYMbD5uHkQvzFMsAOpeBs2NP9JRdvdz
3b9hAdlkfMbL6FzRb4UqiDajQTYec4OeqdZTLg9ydt1VpJxaDgEPYzMtz33weSAtRXfaIFGdu0yu
DtjKz0rPBfnX6WSbzaMCkrn5NkUhs2JLibOFR9SXHUaC4mCyiE2akU/l90YHu5kGKzMzqNhk9U+w
FJJU8if79gVrUhBmQAbV44ZZVpEBIyC02hW8i0T4Pb5nWcyzZVw8asTchPISMYCpujErzaRNCLE7
IiNUMW6OrSwDENvQrV7sZvNcW+C/RlDiy5MPnsKEbxrr78bexZFRGaEbQBpJKT2kcvah8FLszk1s
bq9OFeaXI/P1VGMXBYr4U2Bf11rzFvXT8OWYh4xr2nyHXaDf6XaOzKGF3w9ZrT3cv6dLVwl7hrj/
YrdXTXJj/Lbz8Lm2XJ9xmiVHkCd9OftsUMLSNLMzO2jENXlypQvUQrZqYGTR2wTl/Cbs+RpJeDL7
GzS3tViDR7XkUqQM6YRoDM9tlEWlVkHYTsTvCoeZROQVvaZ5VKekxHjr7UIy+6Ap8Qsq02nMVcRS
ySMtlmSx6GAJ2uT09neEBWkC28DWLngcJ4VeTEe9nCuot4/cKksYWsIuOeAvOXiNvZsD+D0mxg3w
XEI6ffXydSv2hdrLotghKG2nOza/CBH8E32M53+oyVkq+uLybQ9bSWpju+35QBmHGYmEoNeEJAei
gDXCVU2ojHmIC0mfm9TxzT0Ljzpb9Y62Ttd+JNfEnWFkk2NMIHl81WLNg1Zyz456z5NLp1QUKTNw
Yn2X2IZ9W8zFCxNeFseYl6k0GuUSle0WLN1Hmdl9M44VrccxEw7+kb4IJs5N0erjT53aWqDheOSX
/GOVQalU/2J4sGrq8G3oKH1rMf+5v/Qk1yVSkhlvzYE2VUpCHcDPufIJvTm0d1ewkgj1jajB0NMV
AFVWItbFiClRXNO/ozZnsuVWy1gSCI6FbRoDX4BIfRkyl41d0maHPOs8eMCcu76iLslh6LSfuYg9
rJmGvjbxDzfYh8uxNhHcGgQgdQPn5tvyCQOgPj4zMKtd6WlPM9SZps0z4I6USt0x9j0FiydnhPxh
CnxAwBmmFGOY4sLb+7lmZ+aUOrjanrkD/p1hyWvX2P0XIyco7RZZLJpNzjdJuihKsWC12eb3faJT
UF7b3mwxuFqIfGwTVxP0nfDgQAEHzg901ScCJWztJ+mdUaEeF7KTLCDpTTfgw0hOvyQGAgNM1pUa
u0geZRy7Oh5gCwxHDWef9zUOMAHVNXvDJm+alsW3I3YfcviyUlHkG6jFIpvGO/XF633iLCxfYn19
W++YaJtby+KeYvHZ2jl19b+SAwlhoE7a4opXfJ847w5TH7A2m5ejcPrqGjuuZe7XOFLHYI2KzITS
3JhdKDsMhaEoxXL4fOs81nQ60EzmbdtW8COmrTYWTuhO2+7vu5LetEExKAi2bM2YFp34aPCRCcvb
JeQc79zR7yMugv0VDmo3+u21S9wfiA6UT6qfXuXctYYagloK8amg8P/QQ5xYz7XNewbsjpW9e7N4
1/ICEug4r+HsqM+aYHakycZsqpAIcSjGYTOfdIwgT4RFmnA/PLN7vyitcOO1HCZf1A9dHvw/sdmv
tJpM7/ytv/QvriqiglJqmg10TZhRa0NfZeaCt88ZShBv2bJbwV1lnruka81ExYMpXbrrGDm9cwBp
nznf5O6idn12fN94TrmxTrnfusly1qfbXyVX3q+hEQFvYt267oV2EJ029E8Va2rLEuLbrtWEjY6V
kBAaSIZc7wbsF/8SE3V8pLFOc0BvVSTW5okPH/JxYrrljgkKOKe8TDmzmB6jUWzibECkTrjaT5Sq
lAGGMGAkAtfgx8DPlfX9mcNR82NmFCX/rFKswecDoze70TEtoMYUp0+jTNxdPlOCgQ05XtUpQicl
j3JnSyTZK0J+zTCLZzb+VHb7cNbrV3Yrx2FtZYQOp2kdA+6ILZ619UcUDhZcRgSpEWRPFgvcYgmF
UI6N+Ez/Qy15/E7meG3me4WWDh9v+Z4WfdHzvGHvOh9V30HrWdhSNW2ovloy2Dy7Uc7/xtfM+eKM
lVK9u2ffPsY1FLB185U5XiwdZoBdnQTnc28sCCfWe+fBavSGimgDSluCkU/CUpT8cIHj9I42n3SU
LQxUPwU0nfqv3riIuT2nDYGiCP8JlhMBXSY/vReV5SUTPtyMp7C+ikzGxlgWkCMtUjhwCLa1Kyit
v1oXcf6SfW2EBG4Q8cDUmdbQ4gCQIGm/9Zi48d/ZdCiCPMQriPBFUvu1nShHpoG+EmtMjZ9ntGew
r32NH6OkhzknQbhTQbQm52bDPkf/scS75dELdGrEltGJ3CDCU8KJA8FwVAQh3yej7hBM2rQMoa07
YHfragjIsRGpYVqySk6zDJX3xe/BwYv2wYxmXoMnf4pkrdPZSgC+Paa5eHihbB/ne9irQOls+oHh
HjoBy7YEgcYestLOn7Wl1/Gm32ISdlh7hg3RapK+5M+wPf2cCvoUNvvBZXMBJCrs5Cv+mvLrPRUn
44LN0nxyLSZWfvzSCeQ4HNAP4kAXLY6o6RT7uniYdGdHP6l1xHpYfAERHC2Pfc6CSjHaMwMF7l5j
5jV/CyFDbQ58NlnC8iAxhKzxODt9JjpB3qHi8L8ES3bQWjFItOHhcPkvfjvKrVw7woBtG0CKTtUC
qKNGq9DBa+YZE9iEqPUM/WyDqGHvqnFJW83JFWTrcyF8513pdHciqS1kCmJd1yypqF6dWyMabxwx
L1Qxh/hqOr2/2wi9tJ2bzKYD9R4QXB5DBB/t2+dMxTXRgSiRLHn+R/D5WyS2vWX8UUmatfOau7T3
oMi2+oDyKQWzXvt8pVnffUPWiut+4Ts9t7ttvVVnpCGcvoi0a9OYQPeCeP6nUZxxr++w++YuulnP
BJkdC/od5Znyy3HnHShWGOKmA8vQB6VCd/Ie6z8mN+NU38e2Iv+bjwFkWpZreLHr+Omip88hZCqk
5MQBimdp5PXvoHXvnLxczJPd00oBGojADcxaVf4aw50SdsXVrbxbU3l/0WQRM5FLYUZiy7OnB+Sx
b50Lc5P5mf+v31t9xybtlm3QOz+Qr0+EcCQT6hgVW6y8Wov5LZbJBAIu8e7HW2rdjYwizI4cdMdb
uM0BZ6eNV9wWTb5w8ErI9/FwtEA6SdjF4avITEBAsJTGuod6NNAEUuYozRvWHPsJ3UFtFi4+vvBE
rXryb/phEAx6wnYLM7ge4hRjywjBaFBmMGUTe6cRFfvQmXLpxAmWgPDSgIh/7fvEoYoUeDdsDcJj
ESnAcw3J/J4bNwx5kwUby8Bgr7YlkC1GieVhckhUvTKxJ3FWv+6bOJtYATfhuz8veFHw6ybGRn/o
LE83WwffN8vyIBM05uVnR9JOqnmdZsI/4rorYAOQTxQpiwW5e476tQanVvN5RaoFWh2WOuRHmBNY
Qh5KCmTx5980LIqI8ZmsQDEAbKlYlfgToMoTeWbK/aJsCYwA5UEfyyoMI9bDejNW/4RWNc/szBBP
j5TQUz3p4X1QwGSEAk8K1xBvV8EBEr50n6UBtS7JTGnddTHZKKeSsN1HY+2YDkZZbMVatN7AqUYI
H7tnvuUiZjSTsEoMhcsQNyLMOt/KNypXXXA3srxYX9VI0ESRPG1ByuuYRdeTWOywkIRIJB/tafxR
LoNnq/dhnmBw9LF6H5+lq3OaH/VaF/t/9cW2f3TjLPfqKWrDGPgjm67NA4Cv4+5+K4IEuwUoPpJ4
rlsJ6ft860oOC47E4Y5KN6B8sPCKqFxYwmt7w6Xa8y/0yvjOGEQFj0FtEwYsH43z1834b++U/rCL
JBKETnRZOegg0laB7Pg0UoQVZGkZ6UACFBQrucWZ2p8L5rZ57KQMvvVk7JfzPcZAid336L5OfdaO
b86r3sGXjIkCuZ8sRYB3zRN2PTFXO2ZqQ2MrWr5qeLqcGP2t63vPHW3267gZpQ+2ugu+u8284+/c
qcDL95zbZsm7MgcZ6MYHD0cXsvzjoH1pNZ77HF1lcITZQefmeaWkQ7cA0THl6t2sDGoB0ExLw4ut
3vmqNtswfZxTqAxGe0b5OoQMHjwIFqGFVuivDWLWPnxU/uI8s6p1tsCnont9esUpoy1UtvTir/Rz
GdDR9F2ssKhoDsxpoJ9OgSSFZBHFLeFfETbDg8Zf8EWggk9RaR1blFcH8Vs9qcTpggBBGiMlB3ZR
fgxLcYI2v6T+cdsuYJ8TtfmGZvWGs/a/V0rACrNxTvDlS+4LbbHez7b3mkhvq4sC69SxQZugCulC
SWyJlF7QWxeRf9qTpalfxn52dqswT/6OZRUkFatekpAzvuTBaUCbM+zAhOYlJUX9nBzjP6kWelp0
WrK0EVZR+mMmuyzjDm8uNaGVAL15f/eIPC9bDZvE9kBxFztPQx5iAxfwwJLWGg28+S5i/zziyj52
fDkUGxZIP2oPqHV3toQXoLsAxRLktpG/yClhZFpHGMgm8a62JV8qOau2bas4gGk/gyx3vLIK9fBE
pVqAz537MzLSY4J0ixpPGGhb4nnjUYszppoBdKVyrvJMrYEmOaqZvQck04A6zLXSec+pYP/40DlM
Kz32KYbqnwhOT5+/r6m0HUpkXBpcHMpR6vhf6KUlMU321oKWR0A7DZe6kLnGp8U5icUv9u8iSP/J
a8hcrtINf7D4LZnRzbXK4XpytxvUUkrbtkSGS9aFoXCzGn2HUxlHiynCpcP9MSldjEmrz70pig1L
q7nApJtLbUJ3pZqv+7T/Cw/1E/StgQ4N6ysSSSJoC9/CoIbJbnUwr30GObT6t5yCGgPL9+bgh9vK
z4EyWSRbT+8nK1L7Yi7aCaHz5uUa27HUhEpfA5gubq7uEAC0JoxnNG9PDdmZzUYkW+gJo8VhK3KD
lDLlXovtjrPodwBFQKpUqsaSDsMmNymihKbRf0ElqcGr5ITzMq+VpMHa5ucIGL27VNdPGdfcHbzC
XqxZnyKaufS66Bchc/mxn2nP67j/mJDIHTv1Kn6LW5dHTjASYGR8X+z2Tc1fD1JOD5Veec0NnKJI
C4TzWUbh+ho4r146ZUXXigvB6rRzAxNS4Pe4E/mYTI0n3YT/nqfRwUXWofGFwpnY2J7Z9KJPo0qa
14tWdO77ggSw8ujYazRjEA/wWRYvhxCnP3v8uTojuXNE6eOM6dSHOP4r9rAvaEsjvj7slpV9OEvD
MnSdnkxLxMvUKEAHAwAvMKlnrC7Idg+mbfmSNlXE5E87zGzpJkQIOzq1Op8LZbpk+BiT8W7m7RIG
x3Pgf35MhL6NBfC4Avjyaq9zvgf/x0I8sqY+LHzckGTXgqFIe1/SY202ycqE6BzV2Qi85WEhup2C
K3nl9XBqbXYm3S1rWTxFC2CklsL4LimzMTlv1cURqUQ5GH6xVLKVeajGqOV6N9FW1XhLzUI+/IcV
ShgDr0fR5UvFhZsYFJKDghF0DQPu0t/9oHzDbLuxTdLQUFajztTH/c4dxj9oWo4Dmt8qt2S9ZxUX
hm55FKHyyCj8rXH3mrDlljfquf+V8zYEAf8TGQAAKOUfYHNgiY6PCQzkVj+Zml5k0RlRhfXChDPL
lJ6CBPD6X0+dHxxk8V8fHo5lU2c121xiJuON6kfdqAvGTLIAQbecNoeNFi750+Y60n19oXrbBZ/3
S6/kZTkOiSQunbNV88QOcexehpBsHI1etcS4Qq4EZ5mkeKr8aWZ1mMAsBc+AiyjAN6LrA3L3eSMi
daks/XnarUerfrfIFmkvIZVKKJJo6uiuuKWh8Vi6Mz4yyEEaqpiJgGw0Nc5lkMyr7B18viOigRkc
P6xN9SRpQbnFk+SbNJfCPLYs2CwCw+eXg6Ff8ITxdvDNowx1wf1jZYkrX7QiU+OwCk7YuXUHejj2
mxSgxuDW+iUvYSR8lNhUU7D1lc6f7umBIgfjo3tphMqsCuSkptoUcISCzyOdOCG6x2BntrhFVDmp
oSElslNo2N4gvXPXgo2p9YPIRv5v02pfSsPJVVU7+DK9yEXNdYVhFPhhps3gfl4PXwPMYlFASBan
mpYjh5e4t8gR2IKNJw5XJvA+lQ4imhok6vlJobTNrh3Cc1kXYjfv2pZyflX3NPE1pkhCbUNZmGV7
9kCHd5Sm3VWFXksZFJTfAZ3cuJLnW6g5Ffb5n5AkQVd8d3kKq/t4Rri8OH0txxbcMcMNUu86kKK8
sY8UFBflcbbyKJmxxGVHjEOaYFQLRFafz6Cy1nB1uS/XhEYc2xtWVVvkcqpPPfzYWQOqr3c5Yb8S
/o2Mf5heVslroHUUELlhVVKK2gT52qx5Qdrg/j8deXaIu2QRd2JN4oYigYietelSANUBIVQ8diDW
T2tUI2CfM5uZvtLDnxBJsaO3kTsfGTYz2LyI7juurBpkbBmjZ5hFFz/2O9hINTJi3AYN+K6XQciX
K67pR3laV2gFYPB6icp07q1mX4Roz7mti6cNxdi82HLvdqSUWPbzCrbIBNDD7DIL8hYwRi3jXRTM
GPiY/fCCQ5RhoelmyLP4ZVxvv2kijWYI4UdF51Ss1//pzIigJCszJY3/i2385Q769y7AShgnCAbn
x6ju3ZN6PwsiBkkFtHqCrPMf/Ts5oaYEMm8i+ciIKBkQ6jEfSs5QpsaUevoxG6uhNqmZXV44whSJ
YeJSQGFmzo/+ScFB6fTyrDFHg2qf3QemMlY3JuymLNzBA6SIhMn2V+DNg2NmJVeK7GzXq4odum/u
IHzCyXDntc40ejfB0ndJ/qt8YgCX56VPCTIiZqkryMLBCQzdE+KhU0jr390AqAThjbR4VTqIb6UF
8nsnl0md+TS+T8GTGW7ztegibRDztwHB3yUxvcC+jayhqTp7cImqhjgivxfL/rrzrjn2OD0feE0o
T2rT6h9cbIOXCIExqaKNE+bQXgROHT23I2/HuZ0W72emUZgjrvNv6vEV8N0Wln9bD4grvE1k1bbC
tUnJMTkT7kcpcDX0UntaFHfC5b6m695PGmiQLcAR6JXO8jNS2Woa6dF/o5mNlECXd/3XXnB0SlnN
Y4KryKdIBCNHVVpTAoWMKb7t7sLL0KYnrsDUct+dWgTjfDGfNv6gvdJpkKoRSk6seywt68FWz6RN
Ro6dWqeNO22Ch/8hW2T3aEvn66twtODrx3wymtNRXI74BPLtWeHvAmvoRYivckvXl6xtwGycCdQj
wznLxL0xNrEZkhQb0ByyxdEe6d0+zqeVw2FmyftpvviM75+W/5vLADsQs7Tcrf783p6aOFuo4O++
/F/hMGZWw8TsgnvYt2ECWxW3lqlJdHNlvmCoJLkOVNTtv/coWITV0xnWCn6YbvuOCsaEbQfSNTIu
QnKlXWz+LhUvm9eMfVDNGmtLRkFLs5NeyqmsH+1snpXJqRunJ2+XY7mEPvyRvNku1JGv+ZHeDpVJ
RhiywagCtA/JqB26W+A/WL3yJTB58rYvhnFPNm5D9naQM49OO8At+XfvQdKafNAVbsrLqATXgXFp
b4s3lM3YFGEuKATzZvzbTkJQgKt0n8miDReIus4mRYNI0vcQQLIY5cIWCkT+YuJq3MWqOHs4ZyKg
VwYcfXiMGLui9A1wIb43p/hPlDtYB8a950YBvvOCimDbLfXLWhXaIeVZMQMRcXzxfmkbhMwWTSf1
X1J2idjfHoCatfP02GjT5Rl2mLyCjTvNDvJey7cLpTZpWJNaH0EK8Zuqi85CpEW9oIWf4msfOpMa
w5yKkp80pvfNSrAsvWMRkmuqRuIA84Zdaaui5OTKjDG4ZmfdOL3zql0QtJHmJekjy578ee2iGQwT
42MV7Zl0xF0RQ7ZjAUs/W8efl8pGDENRfpa4oWpjGvhvOAfuIbdzhsIDTSGy6DDHANmTM9opBINH
49Y0SebRLKofN3ZVEEcWvPYucTdTAV+5Y2vM4oj6IkYUI6pRcraMeNFOMQ9H/X0fcmxTgz2ZcVDH
hrRP2bGeoHm1ZykKQV2g/1XzDI49ZlxrVlloZZFz5AoIaExKUcFgLTWvSzme0LUBnwq1gYYANpa6
HcJmHzxpfkV+I8ZT4lYnkmd917gYjjHjaSMqocXdXhLuHKWap5gfzMhYHCp+JCesOUms4t3XS6FG
LKF00PrAlTScAKWphxPLyo1GkMjIwD0iPWNxri5oC06kZnyvWoPpsqG1WaCTjCVqRfw6IawYo9un
WJNpTuS78Ovq05f1Vqy9YTEhZpAURTSqCC89QouT1h+5XbfYYH70qsS9ha6/lat1CS3hKAzdGB2Y
nVNCMH4Da0Bq6QNOsUQdhx1+BySPC8dHS1fSBo71AmTHAK3Gaa3KvVfNTpgBFgr7zQnEeV0ftC+b
MHKu6tWFJdGi7MhDw0+Vovb6PJqetW0+u+G0T/CuH8gLBk5wdXgItQ25W0/ilFfl8zxOLTaIWPfT
h50C4637NaXzeJvVCw3K6WUOSa6YwdSqoqIY+/le1l3wPPOR/mfk4dcp4VcYv3pM+vMKlITDNhj6
UbSDXbrp2Ma9i4QIUDqIsd9G+zfdz/GWli3rasGJnrLcB7TNxphLyVePpHtBiEXHcqw9r0+7jVMT
Bicz5MPPtVz83yRAIE4u9wfDXI3KMlrcPCwzRxOj2albfFvCHHboWFP3lv0qHA0xIim8mJn634iY
nwrScek5Qm+yOc7a/4TOqT/+ERntWc1XQgUkEshPtTBCwJEw7b5l5tMhZ9Xg+fkEPv4iMPRYkRyM
0+ZPevGNqThHXzmIy7kHNUwSM+lFP4muaC0gaTAscK2ZypG3QN1/DPMAFwPmShZZvk/BtJl9VqTV
AgIIHjMRD3HciZADSpowmhZyhYf1zIDRoN7qgTPOnBUcMiB0M1pd43Bp0bSPFCSCxefhrXtvWgZu
JbS8KsQYrRtoJKIiDceLd7rTG+a81shFSifm2QkdYm8XBeLBKzUvHhpcl8WLZ2oaSEIfHooFqanc
waktjcIUAuwcnN/T+PiRwIgA3l1fxKXvZ4XN6fblV3kDqmYYSfioQPR84X4iihaU6HKec4lU+D3F
TVsBCzQ540IoHoHnnxnn/lXdOlAbXBPXTtNVKEsV34NaXa/bgrbwsw4olBGXdDd4zeikkukEegaJ
GxPm7CTgQSSfZITFs4LktaLOdPRE2kplQHod/Z/kBAP1thm+DpRXhcRPWYo5sdeWpw/Ufdunboyj
YnMIpTYovQtlBrmFxor5MdnNf4ernZbloRps4WdnAVzUNbnXm0dIuL8uTWMD3CJv7+eJZfG7mEc8
5HCnoheNOzRf3+hbmKVYSEbzNMCAJ+1yP6UBZX8uDjEna6UApVxd98J/HERCZqGdSXAV/M7LNc1a
IW4Nh2pqirGCReznZcDvmVv9jS8FCvUg51j865dcZTyqHV46tRFPm3cv0Y5QURY9yORgLUMbNunf
ikAyKy2FaDGxbwQDBrXY4TTOUVysYwh81Fz1K+U0HhA7/dQhKyRWFYIVKBJnGFvM/w2bLgWykUXL
2DNCnPNLbjY4rmN5+Imeql7samr4iJUxT3u5EQ4szIfqvcxT4jWWT2st7vEQdQzZK3a2HJWWtNhv
9cOfgI2busZjjzz5TQ6ZPE0Hx5ea/lcrhT85SV+Z7a6S8R51D8VNd3OmVMM8+7SjYfRBJhO6QE+d
Oo9CzU/pAbInFiIHeBJKK4h6urLs2bYUynDq8IVcGfe5a1WAbHo59jaBSuYG3CQfzyF0qPxprQf0
yFDucez8SIHR+ka+FDAp2bXzq8FV8ZPX50ZIQ6A42g+6ybhFDNsokPjMAVrndkr8GNYRBZ5rxJSj
QuJy/NebusroL0y/5RWBeJllx2FiN+N5xlxvQltikXdk1ttpUP6KG8CzK8x/sSmpPVEBKaMAwwd+
M8w0yMo5VuqzrKgphcYtPw+Ax43160rcSphEHMHmr7eDPdCf5w7dmiRZVxbe7WeuFhFOs7ncy/na
4KkQZdGvuqUnUciTm3jiJIBZhL9XtnupNWsKyUgfuWvIcn3S8+HWUDxaeagmOYKXV5CLeCCi1ct/
pIA7Ys7KkRtlJSDqv1f50gLp2VN2iwETxcnmoXhYJeZnFL+3vj24NVwZq85rQcgUyzNT2zQN1OYB
k1D9aOGLVYq/cuf4H96RBktH1wVhqoOJvkNfEwqrsN6CdGoBowMvKElzqBoHFxizKWhW5wZQvnK2
RqLDhZoeiWhxHDRw7CTjwoR/PQ/Gi+EQV+bmIC4SBWWPM44XZy6kf3byBXeDdTu/mIL4E1IOGhcU
WXZjNKsQ15eYxXbdvfNfCYyAi3CwYth3EslDKld2dygsBwUhIdiebS89XLh41nNKluF+tPWS4xqz
ksstwnZk8WzBvyESqGCt1Sx8DByCGEvzDC5C0kRg2riY8nMIM8+WkUptD6yJ09F/R8ZXdYinic2K
FqSRbXO6ZSaihF/Wizfm6CySB4X/Jl+XfgDk7NZ8WTr8kG/74m5PLXTmSl/pPWREFR5dnidyNTFc
A5NXE6KEAQFSEcTbWYoqH0/VyhbL+ciKNSKHl17A7GiJdECvu8XktuN0PJuX2LMCPyciiZxQUDVJ
zB/RQxvMFPjrzUq1/Ni9keHp36Th9U6v07f2LKEG2IJi/Po6mbRM98i/pJWJvNkpQ4uysUyxq4sY
MeAXlGt6DDzMPGD8jYckxIp8qTvRnWUPH6uwk0tu2ZczrdHpnPhYojxIrytDg6JkVeU9bYTZXUEj
JhJyO0cWqnTHTPHX/SrPNNDlq3889MjgGNiyz+PvUjXcjUe8XIZWeWSOLb8diHoLhpCRZGGeIY7L
j3hE4Tzd5j/U7OIrmLOgBbEHPUa9iK0O396nfkI+IYraZ1dMIYKYawLwIGk66vCUdkDuceP25gK6
Fc1kicqy5DIyCQDcH3eEiz0nh4WnXqLt668qfeXOFGOlgqX//n1C2pq7quOTBsJyWAHuHJTXlHm7
JGUZxQ/CU9OiLSlf2s0jG9ShSj3WVn//TRPq1BgwiNdLjn6Zzbnf50sHTt7+NwXZqEfqdjEFItgF
YoEHJdieitiL+AJPX0ESRz5qSFdEfJbXVGNPkA/E8g8hmTJlRBVI7Ya3N+aWS+k/8TB/FAXPcz9D
5qbvOXUPLABp8c9R5TdNY7dHCfYAk7+DDqvMQ7d4QvsNNxxff0grpun4fmh00Nju97AdsZo5vVkh
j4EzWZpJXeqCr6hwbHF7LqcVcQGGVOhe275n13//UlpZSkAHNM3W22tHxT2/55aoHolWNbVP6SUH
uE8SzSgBIryUv5oYwY/7FyhmOeEK5D/8rT1h5WsOtg8E2wtZOz6DqhHd6gljGf7qg8A/gxo2PQaB
Lc7/13POk+79BfDCw/D8HJfhTxToRLrGQ/K4i69ehbT9JrQVD3mhYTulnHJfbas9ot5h6rmxCrGM
7J0TgKM1iuENgfvpiG20hyQNdpd7NJY6zXTATaBpEh//c5HBwQNsnLqmh8XRO3xGODP9e9hsaw6n
5Nan9E+J2OgS20X6Iq62TCB8MusWqbk3fWvgCqfAxkdNYt4+sk19NHSMJoJ0t2FALYfZKdvjBk/d
SKZSg85owDlQ9O2QbnmO8HUUeFXu8FfjjmlbsUclWSQYYYZmHGwTzTF/ducO8PPyb5DDuSW1ooK2
cuSvIy5j+0nk26zwdURTbY8+2rZY4pJBsHaQSKX/6aMB07pUX66XfEkd3MRmsLjhXvcTCzmVEXt5
3r3lzUXtU70+/eywenH/rn1Ij3ktbZrstQ/eMRs7QzytTUAbml+54UrlEbTizIBnceOhPy7qN7T5
hHOjy+zSGp/lLcUOpEX0c+bQ+R2spqfnwWbjdbr5WtOIYImoztVGMxhUSPQDFtNfEvNLb09tBnPX
ut20RLE6LmeWMfHRk0yYHvBY4wg4MxxOOAELQDXxJKoBovnXfYR/Czav2LYYiofXSjd742aLxHiI
XZgNHaJF8qBSLKZd7xSXWLE64QTlVI45HDXtyCUGJCsfLKvIqonSDFEgIMd09KwlGAcoDsXsBhGa
VnmBZjzt4Y4LcIIZhAeMmBxTMmXsIhxaYTY98JYajp+8OZ/CrONLR/e91hj0xWrJJTjXs6ENtt88
oIPR0PrqWGsXNONfyWWfxQmEYvcc/+IGm+421DYLGu1YUXK4Kmi+dIuGfFBhzkXA2wv2PC0TG1F3
4Lm/r+1viCHnsRBOkvMT4Egrh/zlF/2dj3YUpPIm84bjma2EOMsZ1Psv8itgii0jO5mUrvZ7+CxF
CnU7rMWHFvUFCDgYhboEA1ilOqgiHv+vtCPnr5a44jTe3nVTjbvCpAWpRYp0+yjtqSKJHMVAiFn4
Kb6E0BgSNox3wQbwhjrWY/AMW4ByEZ5+dbDcc7TVoLliFk1snZpn7fRLmH+ExMgO4XzpO/HmSE2n
uXgj8sXUUAuwumtW5gPQPreMmOn864AYGP33wfArcv6CgVmTp40K++UWoJvVcSycqCW3pKf/UcLI
J5+owhNOdsoY67cbjGrucHZxcyu8Lo1RYk+ALx6XzXOgWU7alju841gqM9OV8u0wCtHKdKXMjdMT
8dqy4yksJK4BUvQSPtomWJ9ymmTp1NqnWQ/L67OxvXMUTED4PFAdi18SRxUlu3dpUem4M0RXsflc
F+I7ahQ2uawHx0aCCnmzsr2AgcRwvKq7CelLjQ1VmdXpbN5hqFFY/F1VuC2F+Ue7yhIw0NAPFuFB
2XTh86mdZO36eZWiGWIp99PuhWzW5IaIGk2gWnuj8Es8LvucWp7QttBn3dyYcQqHWztchXSi3X5J
HwVI/oXkLOv4+OFC2D5BJ25e3drwNNuCZkd5zBiZEA1N1aWVWwQ7/z9/JcuSOqOggUe1m5D9zusI
3ztz4UMOAZ2FFy7FPempNxn3pEI2Pjz4sxYjiDXijXCf7VjabLSUWFIcjF5epROthit56I3WqLgW
h+yBfcVnXykaJtmG+Xplu+Ql2jjHY69YqVfwgypoEOpTWXKuM4VyADJHLHn43MSAX6PHQ/x0XGUf
tZzqhFm+A1k2BSQsCPrKCuL4xfAvOXDACtcXlBghln9Y3zcmp1U5OHvFVaFpqVa36CZD93/fuZJq
NeF2d5zYH3uNLoP3RRdamIDxpoxUSqrpkvBf3ddn+oUqXwOPzch9OuJ8s9gvao1v5CDH+2YMA504
PIkuX9atqVAkiUCgH8w9jGjFrVEkG2uU4YNsNis/dLwQlTD2H/Rrj+P1RHe0pkZAZuoqjbR1NwpL
8+T+XsjC5Nb/8Trr/tvyPvILKvqEyhx5Ts8j64wtbuF3B1xk3/YERxSjR/j3i1pp/uRrCDbrpd9M
eidH9DUUdK6DCAbPb1WLuBYcMxBBLJhNJO/CuIqaGWD+WGUOdu9URJnpJd8RrSiE17QbcH+pOKxQ
l2mIQUZ58xtDTqofDYMNcBQqAnqbst5AQvoSgG/9S6TOQQTB3JrnlRR66EOtw/HkRV54t5PGghor
xYNeEuTaP87Jek8RJHDFmqQFU8zp3VA/vjfhJ21GkrAGNDXQsQ40+a0MG6GU6ANmIhgJTA6GY5sc
eDSwC+PtsEmCMKEha96+o1Au1tFhxGoUuQ4hEWAHrKq1rmp6Eo/yd3h02qTsd1O0KaAvWnZEpvaL
Nx4L/V5eLPdzBKq/rrFQlYlvgcIEntKA+K81/Bid9u95GFpCq4lgq1Ux4d9MjPdaBUj6yBwSPLaf
QJFPGTwz5OqBa6NJVS1GxE3DVTkUjM39rk6rhn7FDuHFJLDnJfVt17Ugqc9jsVOgi86W4oyhkRGp
DFk+K8iKQZ9qs31ljpVwyFolfWf3L1qduljBHV4l5o6CsBh7ZjjitILRosw4yiszG1NerR1oqlW1
G9aUfxRzBhL5u6j4gF8gCNrZVrXlGPX6PeVny7yddtHj6czIsUONyaVShN7vQbhm9CHl+85v5rzU
H39cPUD1p4HPF1YIyfszVPwRP242vTfm+tR8L2MZ0J51YVhjbzZHnJMSwhCxnKXKyOa+oIJxl10Y
z1z7XqWmik8DBk5LPgd1FwGkEIbsJBUryeM7n5aKjXTSFzJ4P1tkMnCD5+EmhMxrEb8D8fDvp2dE
jM4XVWP/7M8X6Ids7toFz9tilm7JLkagaEuWPxeaYTyEpupg0HAZRZoMhN4r6+4BcNnhQKF69Cy1
Lv0jdmH6ZVEaEQIXhOwrr9AA2R7GyLC5HEZgWw531zMpCjBK1Lo03ZoCSGva+TQU1qgPW3ShW2a1
peAMQXG0Yy984QM+ap4YybwSqsUs7nWgxxLcGDtNxRWHE9+Uo4iHlaMwt7Af2xBTuxiGGDd5hFd8
8jPBrz/K1oEC8Mx8/Lv0qMb6Gju2LOAD7iunPHrVjIr1bW+hkP4roGJbDghRimrK6jx7j7xipHCy
C/9lQ8veN7CzQvZQQysxOO1INHx5AE4nsv29zhD5L3TpAzdLnbjdmZbSXtzCnWuJxHZQzktEV9gK
ARRTV73gOVu3m1/9iCt55nZPWOwleSy4fkIeA/HJPFgfQAG2PREjYN9PjDPNUOf9uEej4vWxyjQZ
DJjtL3KqsJNpJuMi49Y/Xe/Ul4J+zIen+/k/5ezg0QmEuyWZ74k0yaQTaAmoPPYnWdBLIfh+8Yd6
lndKIvOW825ZRFhWMugHiGGyXS34XJnCkocLYTqqRVCDGlu2zplR0NEyZZ20LDYLjOfzmxKDIz8H
+bWl2LBfzSh3AwhcSpm1i6bb98BSR5U4dW8AqPucGN8S80TD0v2wIWlwJOji1AMcVFIykV9vbngf
YiTg+Ypf0AJrZ6NACaV2nEdbuESj9DLs6N3uOxbI7FePN/zkhJYGEHUEFzFsa4k8Zk7eFwuMrLEW
HMkF+ljvUqH83IYG962VmAUmj+k3HjxqUanEHurU37ZsAJeJ60X0vbHKHBGnyUDyiSeEjyZT8Z4g
HORKeRrjB2+mQcpD1qHi2O5s4D2xyzy/zO1yYfjJtj5Qty4ZfzoU2flZa7xF/kpcKNy+MIlXph7v
rUu9TlRpEkC9kxCWI5BkOSmNTmshEh2oy53GESYAQUpTnVVUV6kW2YS1ZnSrs/XO91Q4vNmRCY05
Te+bSuaUkNpV+APsWi01vnTTdbMARB6E12JDcbFsOcfNvqctD58GR6eWFdbYznkgviynSH+TrBXJ
Ll4VA/9aRx/ostxGNWmXtISvmmbvaQ/ck2Q0qI2bDM/XygbZ3QiUH9lTM3QVB+drgTt/XkaloZTd
nEbkJzNaCUX42EqqH281Aq4go2As52TTxAyQS3GStUCDAuiCwCxqK1UYsVrK5j5g09+w1+bdOVxi
n0EYX1NHkNVbf4cSwwGHMxBTooNi6BQvYdAPnaZhpJtCJTKruA5eGxIF06Yt6mmSqtHmKauuxHOv
6ZTccMQLOQET+7YKlAiMZR3R1gCSJXOv+vNK6cSeeKvLixW+AT/zpTwX8Xo4kPzucJcgTBZ5ff4U
/ECVtXnUtNccGqoiVwdzqop8PqHR47Rf1e1L9VTmOpbuC7ua9CK0MGPrqdWicgvcVcpOxgWPowoZ
FjWZsz64hqJVqjftUWjGrretBu+Ckc4NfngnpZzScJfc5c0qu+cJjlynLBnEVIv0MtCfLnZ4mFSv
3MPvJG8DRq203UY/c/038ChH/UhyyPGx5xToJKiYyWPH3p4RD04/n8LFopYxQITIH1fdWwBY8zur
xt3LQcZ748fppnzjHqJsQHNjKZArxfv3BqjhTlKFN1YwKoHSKgw3TyW1qmSWypq5rHNd2btJU9S7
ks0AL28e02noz9QzgNrE+zdtIJmiEQrTuy3RJVAl0++XJpDJYatbFdpCk8lQmuA3M3+x0imJIUNb
h4WsMTXk54OZ/0lSEFOGYLb5FJabk4PQMUAQPtF3jcGsYiydijUW+m/MOZ2jQedD/7SYR29oJmq7
AlDnOpk39FtczhjO1K10iBh8KvTHSY8XIAoy5B7AKv2KEvnRlzCA6db7YaoLDiRUzSBQhcys3yxp
daMnSJ7UBmwLJdoXFj4pRtSn3tMu0biHrzvYl5VKWeFsLwgrl0Tv2YgTv5Z62npoZYMfHgwKILt2
rIbc3aZkWvTTPKVS1+ThvnSn1hiNS1NVlgDF1ucayr4sb7+LnauZQxxiSZ0094Xlws6EgHOfD/u0
qvfxARBjgt3cQZjS2JRtwTtlpK2bj6T4IYHLLO16nNVLFquz5YSGftJpAKHu8EFJIL/EHPJKqAWw
5E9CZ+mL5xWJp9k5Is29iAyxpeST2nulJDo615pq4SWGW5+dU3ZqdJ8CrElM637zFtdgkTPH7Lwm
IpON+iWLN/qF6G8JgLrKd/hhqqhu5bMDiBi9sJtZvipR9LaREhlm17kq3xkX7v2KnbJjLdFVE+LU
n06JL1wADB4Aq/gNJQmNACpFVOGb75t4kwi43V7evCrvn9bqoH8GIQX3gpRw84qiwT2KigVl4v0P
IrZNof6wjzaIkd2nj1z7rhpxOraYxE/kQasWXw8GteCF/sIKvuhEO56c0iJ/WvMiUCL4fBboNhhK
BvKkHTIzgXQhghuGd5tUBnFaBE9Jor8AkDq0mZkxOWWQYNcuF2Z+uK2G5kr5PPcd5JVStiPFtNVR
sURm/JLzT8F+BIyO3cMLqN0dHood8Y2YSg5MAslAxEBylOj5aw2DPeRMI8+w6DBs8FRfqa9PUlsb
AJY0CkjDEKpr//5+Ak1olkdiZ/VHwztwYF3SWV6FCjHWDnrJh+kXW6LNOzWdJDPme5BRjtqUq7tt
bBpG0d4UoqFDHt32lqyeCgx+EAwyNV/kXFIuUovUU/IDxUIz8wA4FMQLIM7HErZMw0+Dt6x5Mjas
5NozR7DWVTUPHIFpYZeTY52p2Vp8IQKniFz351cK75Rqk4DzE4T/lgNErWb/oaZQrQF0Xmlv+1Ri
UNhJ6JWCV0eEVWumTI8GWLd0YDAbg03CwNPDQObAgG6eQajR+V/cl28ZHvlTJTXttsCklTNHjzWn
SrmAxIgpO07RFP0mM7txeyFC7ypqV9F2Pwvi916ivvM6K0rWElIFaaedAHYW6xwlpue8RHwIXAMc
pjEIevPInu9zZUwn1oKxkhiauv7rwAnNC4yakGeELDAeELNXAWUPO6IkzXuE/pCePXCQDK5H4UY3
g7dMg5blv7+Ii0369W0LqQ1O11bxaCs/xAzq0qeN5S+SR2KhsfkHl5DynGPNkOiDzlD5DTyibddP
ASUga628AW/fo5Cw8H7RG9diNKC7jIw9/DqlMX5Ic5Efv+xziccGU8o8tYBz7Y1iPcK4p0Pe+qzR
rUZuHPZi+YcoVwGG7mpENhyLJykwE8OYfFNQv9DbXQONxa3dzk9WsziFVB5Hda7zxpVGLTiS7UeN
LG8uqOVY5iXUoNlfA51z4s+dpIEwh1wwo5Q+Bih5K24xRvKOvHyf2F7PdDIEsyW+sx2c88XFwJMr
RFNPdaCSVUrQX4EWwOG0Om9HWGpt6eEMIXDZWuD6srgSnVkUC7cgNTedu04fDWVOkWJiOzFBMCmG
KSKCz1XQd3qmYdiUgBAtpkYdNmG1Gc9tpIAlhKokTrhdsqvWutEJ6cTnUbw8S0WDOVV2sJ+hRxqu
2mqscnCK8dbcaFyn3Mn0XsWlEVbZtv6126t+hrKVkQwD1Sd0SvX6Y4rPD2IWDp7zbnIXw6CmXzCi
RV2j1jJQR1rpaskydyU9VaLDXOe79K55WtpFo49KHvK5+LU+pMDhWQsu5ZkrxrqarlM3xRcM7sDf
HfmVFupmW+t49eXf+xPlz2pAnQXzt4cAo/iws/gldFSIHIF4KlWWkrWECiiU3zE10PbbMHRyzQYS
pIZPpwNeUfN8AxsT2E4DJBzVzukgywo1gUlztbWvquvk1wXI2tkrxubPMO/SovXtMhdm3OecQgXp
iANsOxt+FJoKBo78kdd/HWd8mHx1YyDeIr3xan5tZtMd6pTTAMaatl14sOn/esPwzz6Pd54p0K5G
L7YSJF+94CiAFnQFWEbZJzPqnVr/B0L6JnL4Mlgp/tp9Bxyce4gbDiC8WS8526kcuWwAtGQHGdRF
BdDedhdiUNbxXKvzLEp7KI7K8QPNoMsbuq+aGX8zGCLTgBhFY2iLT51wSz93gjQfXRPlwPt7nl9W
wCAW0xOn64TGk6RG2Xi5mx6Oi/AdJCIDrArNipiTq8tTKfRg9gF/M7u+vVLFX6ancHYUx90LEYwO
XLi9nor6oiFMAtvvqOfnpsbMG/+Al6k0547qNWlahvrrH2Lb5itmbc9tGq0kH7FqC4C4aCY+SC2i
QW5Gj1Axh+vB6SdDWkBKz0ool7JjsO901uHx9CqWwnWRqNAsaAC1oMtdk38NtYEPC5U9a7qvd92V
ptwyjXXh63l23857UTnQ+4Jj8p/DGG1eO1wr/Vf4L7htI19jiqft2trK/Q6FDLaa+lGjGMvC5/eH
aQuTcbjDMHSBzbzHruZr3bgYXVKD5F+1sTn0P4JF7dhy1/RePx7x51gENY+lVv2YzJ3d9KVwIhFF
Y1yO6aVJV77YxHVDAiCOHi0Y8L2s5VXXIolU6zGY0qMdIZ1gBW8ix8gzF2KBKloW/o0kFOBwKFGC
9a7EHC3KEpvpFKoT7hZYp3FVQSKjrsheL6H0JMluy7k6dFPkELs+qMFkWjvWZGobADdfgmu9HEbQ
hV/amfghGa7fHY0yYgTNycji2SCZgSsl6991aK+iT5U7Lvnzx98E6Ya8wfuwI7gluWUErICaXjZ/
KXHH+Ikt6PRpuRoST0Elx23UnCuWBqARQevK51Os4nRoyV1mjGl0qxqDnHyRWCCrhBNjPEaSgrsp
hZ9dqepRV771OAQdkd3qViNxpPMxfC5mD3rREUsmYFQ9YbW7QBfga9lyCnESKnxiC6vRWdGcW3I2
7SX7z/hEtUPhe/LC30asW3yp/KsVrEKPc+CeNezDrSYU7d3R60178rZ3qt69Fm4I+I0r0Ud30H97
L6b/RmyLFdJGGxa3VNLoNgoyztXLo41pGJGeWyFINWLNhG0FMI7eUhLhwj3nWY9IZUkxSliHGKUc
GJNqNQAgX5fLYBw6OQtmlwnLxD6KExsrGUv2DLfFv/SLSqXWI5HFIEN0CTYVH60swDXw0PGVmitc
4dFymddXbIKgIc2wAZFsszAhXkTrPi8FcOFUM3tRNerfOxfzedNjM6ThxgFRFpea9ZEKX5vCkquu
jN2SXx1fsei7zlpsIoThOz56u6Kx+xFLcvUoeQIjFL5C4FrqlPx8GIxmpqiaJoY7aRvJl8Xhgb8p
FRcE3fKYwooHYskHLX4QkWz5k5U/93AdKPDTh+jmbTe6MRmdMRPN7YKsPkNX/xo6HUoNm7IG1Yg6
+uz/71mXD1micuhhF09Y7RYMjssyiLOJ34CXf0pWKGelA3ePRp1IdqBMxPesuLM0wMjkGNVgOL84
793UXUOze2n9wDpuqJfBFlOFK8AZstx+yhgXdEYxfMs5E/Acitx0f3fe2Fshqxx9PTmfbhhLSYaF
6wwhspIQ5L4AcCXPfNgAn2gGD5ki01/lXjjUAyMFDbOctDnTrKd2hrTYBp+q9aiAe5TvVAvhZt4Y
+bNxAcf7jH4BWRZPlzUB+R2T0+C4rzF+XCKN5TJsRcW/edoRMiaT0l7IiCGj3BrUrSG+3iRRGkIG
6FtvXsoT+SSc16kjNoOG6mrriObbSoTPsG52FoNN8nj+V01f/E8wIb/Ps0va2VWPshzK79DhzE2T
mXMHfSfH+hLLc9QNbVh6e21xoH/t5esidbmVfcHJBq9bVXbWVe5IJK0zMnFNO7ugQxVLObI13NMF
VFZrjSNSAHv31JZwMOMCi0CxjppM2vLKGfxSk+qs/NmIhNpyOaGEJTmcysQ+uBXXwgLz1tPzuWF1
BpTheB75B0aktojJmlgurxxu+rN00p+9UtDnu5B7hURd5efW5gc9fLfKcndBybOZZcBnEbSiPWIV
ZsbbDNU635KL0RCYahNqJrL2lRc4zDm4JTuBqRlsyqMZNC18ooKTz6ku+rlxJ+M0aHnmlqtTYjZ+
wTe/ch5ghKegGI5yCZm5jOOewLV/uJ7z+s/jK0+Rj+I3yCCiBtyEYPTEllDbyd3NmUOQbikuuHAy
thApOuCLO7f99q5Pbs7BwhU5y1k0LxXSimhoGtgneSst4JTpNo6iBOOkPEVfEKgvPz87ZzGUybSU
+PvoGkp6msQDNsOYvngJzPaafOR3JVfKTsuQTg9TGrnvnJnuzAD3th3UUWTHfktzlnfzR8FonUbI
XVWq2cXlApvcHfNkykuzuMSZti+0AUOoCxJ+v3yY1Z5M2fa2DTWnDuSAhb7iBfGGAudbGkZBXt0T
sWxPpsL4Zpdpxw/z3KC4OIxDtGemOPcpRcP+0Hf4Xpm3bxdOlkv96eWgX3yTs1mNafMOMmRDz9QU
/Ku0Tn3LzEYY8of7Ht0YOG9UznM0Xqf3zBTNehfwSh6tjv7wuoVemPFG9uFRDa/K3aOEgbWp5Fo/
n6P8Cr0i4UgPLfLD7BjKosmvZGIyGV1192NKnfWNlLvY3PLQMzVG3+8JLGkxZMFBlg/nCwSW8INF
/t+ubuu1YaSrDhh5Jq9RDIzdVRV8go/jQtEc0b1HU9WLZmmRvOXasM1jDL/VW/7vqs49jCjkda5C
Ur9+YTYjuYm8qBI46BUWVv7Lxn1dQ3VJ4vVRIBS+B98iQDtEkAfx7kc74rjxPFsmAfXooRoNdlEd
UaRWCAhngSO6QcEBxXS+YrtVepWgI9BGIMEc9A7BTHYITzjmZj3tlAX4fnnyDakYgzV2mJepgZSF
fiKih9UG9k8PJqiXHs0LRCBmCliuarMH4YXpBoPlEdg/2sfFikQqD0xTVGkj4UWclKkI07d3oC+t
cw4j5U6eSkyNmKXXx0EnsUk0hfWl1p0gbtqw3w45tRN7YT+ztG2EvuSjZAZDmB9i6avvlYVeb6Y2
bV4N0IUj2lD/9fVRCQ/E+Ci+/ApNZVN9KIAOjshKxdV4vmSGsdLv+1YdaiTD55bsQ5smwiP1Jbej
BTTS0+2UM3n2V8uJgNCnd7tmqPxotvHVryHNCP0npTGSbWeV+Z/NPjzHaQrCSzYwfSngFW7b+Axe
7VA9YbocMkGS/IVqORN4/k+tplDhdhtbAK2vj8F1E9vlVUlvdGkjjea0g7SKX+zNXGBXL8b3ZLvu
nMXxGQizEzSFY7MlBqrFA32xlYr4a7BJCjmz/HNhqyRC4G+sGUgLANiAhb8VTtecmfszOqUVMj9T
wzxh7imnMEmHdzYaX2CVRo9RjTxTPYx20Ng21XRNWMR2vgx/1VHPcgRGk3qeIzngnIhR4Gi2/haA
wBwVfsjE2pRuyLuVmKCwxH/+FfyAG0uGPqZhBKdite5Eg6lvxOcEF4QUOA7z6AMShD35zzo7V1q/
nVZ33c9ibMvLDKblAePSRdkvyMX1pNjMUx479nT9nE6vPm8jXF/Ze5o+zQ7z8f+AlezYOduUhwKE
2lPajbUyI41fImiG4VufMh5uKfR2XgMXZVdHXwCKFHA2fpMl4mBqpD7mvF4YQAqjMKnzy/ujbcj1
DB36TVyFKLXATb7ML+uxTHAtFnTzf9/BQa+BzbWcN4vJcZqDiBEMu8pzziXtdvqYUmiPS8T/wq/i
Brh+AOQsmAfXdJWc0gn2JxMmwi/ohZ1/w7ElCbdBWCFNZ2OELSm+61PULo/HkDYjMARPyzDjP7Qh
lvp4jZIzK02KKDQ8gbfdbQ9suUCzPKaZn7A/h++epGYvtZFIBX1uRNWj4QU33Iz4UprQVV7I71uj
tH+P83+DJliSxLUrMvQS/TRtZPXVcxZHXEPE0HYTzH0B5eVHhjN/WKTWuatWOgSTtVIvKOuMhDwS
pfrQ5D5np7CzWeeKRFRoWyoZ0nBVXglH9bFWUGS/bx14/53znVxIw7zCMZOjDt2VLRImPH3Z7DGl
VYnD1yiZs8K/hEjz+0DAsnCLcZVAFtMLM2zhco6ojivkOMjsEegIP+hsnLZL0KoDfIy2P1lp/SSF
rhMe1HY19XibARHsauhVKZ+nSb+Wa1HPcYyWFFWdCCtAxZH9V+E6poTZZ6w19onmlRuGGzlOstk8
+S4JvgrzzNn9OA0lRQ9w3BzV/W5EC7xam94TzmIuK0+rJjcxYFU4QZ8ujwxk8O/Bzd9xbAj7fP4R
FUN9MU1cSS4CNgZjz7ijv8CWoPWsMAyJKfxZnKIwCSl04d8oC8cFuJWy0E1kwm6tFZEH6SZHV6HV
Isj/f57+J3p6jhKYf6c7GSmF6D5hl3XFzA293tW/3ztWjq+/k0qjsqWud1hd2Ec6u+080Kf916H4
ff5qX++NDNSQQRrtkcGfKVgb+ZnNhAuuzzhngwtj6evj4uk464g/lkwS24FOyih9v9JwLUCUr550
a05Q+1WH8mQ/0ksK0n2Wkl/9lHYdU4+ysYVp4J3XeRHKFtaBd1SX3xUiuq+ffvUXOEqVYnDIChCu
gQBm6GIPXlEnMDlWngUlqNU2wwLgAJU90h/tCgPNEMoTV8u2wcM7NCXILhmsv1iSyU2222LMo9tO
m9iEFraXJ4TUK8mbcpctrMU96jy9NNn2/j3pxb7L1Kik3ub1/IkeP2OkjTCr0JqvfwYl784oKXPs
4DenyBn09eQJhMz2U1akpR3pwU7c+vzwWljvwMV5WpLC/aYDVvgb57w7JaJMqYBRlzSLxNjwkhhs
G065hnvucmtjydhqjgqHMnC5QrTmTqYnx7wkRK1OK9hN67FHw3MPeRMuxcUbuhJBmN+aHnIlArCD
/LsuRd0vQYA1YjuLqL+oSR/TIuYFw2St7GBROW1nSdgCZXam7lU3ZTyeo18oNMWbgwni7BGSKsm2
2NjZbtsUWGRhFJ0fHK6/TS5Q3k5eotG0X5P0lDcxkIM4WoOXkQmwChxmJe1CQP+MmNEMEIfY7PVe
f6/TEzWplOTaamwG7AVWlKwb08IiJ9JTCzePcBEH7kUGFWpzSb82r/1M8E9UXgG/1BKQfcoSC394
msLg5zWon7D7n1hpWWzcj751WH8HQV9rCG6aEOwETCDqXB5q3ztteiLX1uxGivPzMpem5qBfJ0T3
Ccw+jxXiks8pexBu4AujzHZsF/ohxU5QhXSfM3UaAiEDtZqB06B82/HVxKc1qhUDl5MvlEPkhVPw
b0XBTSEu8W+ReNePgUTcbdk+JAhKD9Fg9XoqmUXu/mjm+39SZUw9gmglOXL13/ndGYR7REgkfe+2
XU0nH8D8h47pa72fa28+LG8UIC/gnqpu+YTu9oJajhLFkMkG861hgz+j6yCmepbNEVAIuRvP47Vy
5hkDhluetLOjDtGljfNdX5/4GOszF4rAZMXz2cpA8asBv/qYEUAirLnmtiq4gsq1Skk6jpZK5mAt
9q+z1CpNr7BH0CEjFFIbC8h//e3ez7s86CyS3USHUa8aKx+HhKwXBBoIE3SoN9E0U1zE9hQ7GFyH
7OQ/uqCfgIpD+fc8BPSr1GpXHx/pmmhwF+DPh9JMqmyy9R8F722zkw8dxeC/ixR/ViYKIPRjkDOL
vqXO234ybvOI6u5OHObrKbZabNlESgf5KEq6B1XiDkRHcZKk0066SQPIzYFhF6miKFo2vF9eDpLS
C0yy4QOsEoI7/ThIUQ2Fx8ysnWsuqIyS9uisEv05gvWaxMiiQLpbmfB+6XzHdDO89Z2HGs1ui5qq
3+FkZ72rhxz9MSD6QiVH9ugp6T4KsyZ43xRxUPy2KaioPVWv9MLZqCCWpaUauNumBXHpWzH7SDVZ
7p0CV3ZAPS11KeYdimNPeazhidWLksSazLC2zV6Ige8O+EXNTVvuroyPMd0jnLcFSFMD8OOw3kWh
IN9W/f9VzzUugSKLZUoo+bi7Y+5QaBje6gT1fmCFy+s7GK8b1w+155Hvq4QSf0xfcuMwckX3Lqp4
MBGBothz4/vR5ba0Sn8Hd+krNCC6SoFMOuTqh/yvAGRQC6r1IiVe/wB3m4IvY57Y68YEmzBi305y
w8k43qsiaHH7huFumaSMpkgvnRK3M5m8E0mYY5JWMvzkx1XvkD7hY04a90EzYRntQpEpsq+HC5Am
Wsoopq46yltkEsAxI+zoSs0wCPVVGSn8v7n0ySmSYa6uJPzSfvOH3xkBx07/1OEMSW3k3/llY++6
Qpt8pA1b+v8wn396e07eiZFKis82eAK0++o9C5bIiQ+FOl/7M/pOgBSQq5P1xu6snX/bxgUsS3yd
e/QATGFJCMBfvmtaMp9WgFARWFvF7y14zXJqMn8KVqbS4iYR/wrzTOaJCfe9/1Q5LCZfYn/p5CKe
g3iJH/cISvAvwbXTgco3ikr1y55+oUOXhuMo7UqyVjO8wjEDFruVb++mwPW4etoCITy97/wf6Idk
RRVru0cwogbwTBIHHXkjdPUHRG9aTDrFLyPLNVbG/oz6KzNtvyd4dt0I/d5iAqtmIrdAh48Fo5ho
HlYFUOGzgj4w1mA2Af1DYTXJk/qbNjzqoCltCjq6tN9BhCa+tA7IO0LBAzb2YOC5Op8JhC79uL1t
kjshcdcNjxcBtP5+Dc24pNkh/fnVvzRVoZX6KPLXF2IeVUUW/aM4KcYrPz92japhbkmwiKhbUnHJ
VebaFUh3fBGLSAd0MMQP7nTyaCFWXp3CgbTGsit81OuEGtxhWG7ybRukPqTXx152kT96qIIQk70q
PkowUCxY1J5vxA/RMC0CLtiMOKeQtDKYDMRqqFQCSlVx5I92yE18Q1Sgqk+j1mSrd/X/XmnGcajR
9Pmhws4aGy60fOGgM+KJyBn/YATvNqXRELrtl2Zg+aEQyq8uAcplQIQa13qFiwEF8NyljIBLmlKV
jq3Gli5YpKk6hVnjxXUIEKg43751fhn9Wl0yLGxDh44JM9SiWKR6rBX0e6/fZx80si4/gy03ZEaM
6GLH1s9qpMl54OVzKbnY1LyGRFb/by8ZQTly8vKhQOoomcC38gKkF6G/OZNa88DDCYloFkan7/0j
7swIAv0akaA8NTAKBjJ550BaheUhm9J5uvfC7//N4P58iF1R0r+UZHDttPj8tttK0HbM9QaLYlO0
GkwdizFhwmbI/bc9tuZxvWqwFDZGJ2bY+c0PIpwn2/FUl4XqvJk/XVDgzYGVKZ4B6I7D1q1fhByH
SD9xdBVVerrAN9Ww5Xy0xMpHFbSR6wSsB1nVbcSI4zKZVt7xBD0WJ4l/HolfZg7Wi19qNskyhYo5
clWm9MjVf6OYpV4Sm9Yie5uUkqN1m+gFKsxSJZDxPvYISQcpEkl0JD4UtPSDHVBReTb1y6vCqZhG
xMMEqnzTfzy5Qq9ZeFvMTd5AyrGBalh+E30+6IYBE0kWx7JWSae2CqvNjym88I85p6QDRCE6I/jr
WsE0Edh4/qUTWksPPbt5NCxccqswcv1DlEUAROzf8ZutyGtExPR49JhOH2KSRzd9z8chCCKPfERg
7RAkJ8IoKbA9qqOHtUFw/F5LD2lq3I0yVlfJCPO2orp5oYVVjh8LDz64BAYZhj8PdG+v1Ok4FgD9
bNG6TsagG3W/qPTOPtanZYR5d9paRhdrFRHVbTjVvp4fqt5b5dI8XmWPoEVtyer6KzmUKDTUwYP8
TQK1vP6IdpCuHxLcRyi3jIcAuU5TasrD+LhXb8+sqO76Mk+wFXQSIo21Lwj19loAA0hNrhvKqgWw
8qJRG6MCASSZ2TSkLYkhosOgui9MKHICHQJhrbj/AcfHFEf5BJlF46Z1wWuMZ+IHjTmNNjCOMM4D
o7DMCP3r06EUqgDzbl2CjPRhC1eAymK7Giu0ZLzXCEsSEA+hGGqdvZrKfN0FeC0JxFz0A6zF5etc
YSAkAj7GbwIWoGXNdgTBoYCc38QczOoQ0alaGduhtGHA4hL5+0uEp7GCXb2Byv38+A2+3IHG+pqY
g3RE6cGuKDA69xfVSbqXUDR33uOkuXBTJ/nCFjudCqD6v7OdY/MKLcKUaxWYV8KPLjuyemTOeAG2
FY3U3OdVpb5qny/dyzOWn4LRYxJdltLjT4RQmKMg4SidhV2Od5AtXdWaJwzhtLGATqRX+yALWIiu
RHAikV2tf8VO0seFJkJ3XrzX6bK/u1zFuUeyBa2VaYPSkQLLjoHXsH5wq5z+rZDpxsq0dTwTVokh
EeH9dGm9S7c5XuQ0FKxQsrRLqdTAYfrbsr7CZxkg/ItCIpl+0yYx4peLG1ctcu9zvI+L30O5+eKB
8cWcT548VEqFYUfsAC/XYEvBH0sPL51a6USHotbzIVsTmiEFfOpCGbaaHzemnqsQzXCph+t7G78Z
Q8VvnxsTDm8bMmUINA/abHnbb3cDDO0A01duDz2lyfL0PjDLP7tDcwwHOJYo9NusiV8QD1quW28k
pnwxPHz2E2rrk6BN5/Tl8m5hU2rRyXCmJI2r172o9kcDznRmVMiVPpow/rndqYEIHRgFEen2biGA
VYqLcrzmUvYPy5BDsXWpH5RNdGWsJXJlrJR2KTUwekXAK7Ft4nXNrN554uBe441tVs77TAcpWf/3
KF+nEvhlZq+eOjBvYGdV0IsdOX0iRRtcTlhf86MDrOHSQIsO8bFq4JShdyOngx6VZLOxhz/SaAkH
R6916G0FocO97HqHhTR75p+utvLjQ3ZTZUhEkbjc9dx/CAfCLbdfhb7fUMoCYuJ0tNysDWYxgfwR
ZK6whLMCACdGtOsT8mVO14VAUaxjM7KFjwK6N8QiAC2E8d1KJlOnocfkY7/aCUtHIGblVFWt7vGW
SPKXOal/ZJSKgfXG1LhlbshvJ9aReUn4rIRq5dXT6ImF1kCyv2iiAfbkYS/McQGd1ceomoSsrLQy
DQ53lC1+qbzpXQLJhclMRHt5o0vqamugmEOsp8Z4w40oR4gVViT7SqY39ZB+O/a+t4k39AkccDkY
yvGj3SGbk1AdTobN1gZY2K5aUnjF80YBbEllwbg22UIKU3XaBSlTLkHhtzpq9tXaTB79GkpyQ4b6
JdPIcZgOUP5QsJY236sS/klXZO0iA9K9xEHnE/IJmafNR9f+0s04stNnMYySxlmFjzgSSWhuQS+T
mMFTdkle6J5lZvFwqmcMvKnw7cSGk83OFlp8N2ceOWGbQESpgk4UGsmrX7sbJ/wdktWaqDRehnZA
WZdl+616QJkhoJfb7ZLJbcmWnCmR96NdhuR3xgQxQyQrSw6TucPS2i/Pi4wVraodXircm+xW0pVh
fvGe1WVrrtYNL9Poaa9C2oR6W+sNIXnwBdu19XVm3a7jaybR+azlv+juqLqoqK2W5uZXBWu8ch+o
aQf6Il26Gh248X2rEn/YJ3/55V9+SNCLaLuST5RkxFZNebRvGZ5qYcCbyUvPzP9BxC+aVH7GqZ+2
Hc+AB2tH9gju6uGnItGONx5osSSeQ31mwA+jGW7NqsLhBWvA/4GluhvqLxkklhS35pgkKgGeN3gm
GN/4QWBGY4Q4lEyf0qxHqoqjrAt5FN1mHMfDmvSe5zXELvpCKFtngVHX5DYXb0ePtGD2rur/HkdX
NneOexYiTjKTjz2tSlFyS22gO/yrjCUj3rVwfbn/ZBYkTnlUVZcAPGz3KoOSLTEraa7wPXfvR0fJ
mPIoMHXYa5h1YINgyTwNquA5C9JrYPmOzRGRXqgjtOkFxbghenDysIwLr8dzkrEfO3U0YU6Q6d5K
G1mP7S33PzTXOx21QgbAhTZcgRAWBuqyUbQKrtHk/HeqGmDA0XSA/M8M05x9eev7vLwnw+hTJgHT
6wGcHAaS0vnf3UmLfG9f3S1IvZX0BjC6z/lO1Tboxn6lSIuQYvY2cmy1xNFBiv4r0D/wyccvi7qx
31Y8Hjr5RzGG+5FlCl+vXRQfcvM7gcvwv7Dq9gjz1NpxNxNAua6Ns+VAInCEIVsK1lNN11v0JzB1
HiaTY9bfu85CNlM5jByiv2SC1yOUFIbbCIAV2Hzl/16tald72/WhtwY9yTpoeaNhefF7lP7jCV5s
zdH/oH4YcO0A7GznvxQdxkie3sw6Kg9k6v6yZKprHycPcCWKwRxrqoPo9QaYe7PDzu89sitjIt1s
ZKZ56sKNYizmDhrbknmEoOn8y75UIFnQz91dnUTuQCVcXElip2ISk9GjTPCAakba9Korr978Tj2m
wD0VE5yYJRhpDvg4PG1hcHqyljO0ktLdzW7Ptv9mbpbf5OkKjp5CIkUXkYLipmo1zjVJlh00i8Rj
Bz8a095MfdRmfzw2BEfXO+5Mm1VXoyObETCGV+ylOWyA/Jpq/RntjaxWJXEUoMCKb1cHywTFnjY9
yCgTY41J+Aol/Q1KGVEOwaHQRs34NfXRYUsFxv25HJuo4Om4AxCNWuKuKDa+FUYUDkQKsoCqEnOQ
JMOIV/8NN/d31iL4+A4ZUapfcCVpzcKLBca47toMD9k7ctNSaZvYOShE9f61WX8aAvYlqoKMXmIZ
pbnHVttL3QciIIvIobHxkpxtNaWV97bjJy81xTt2mLi7+LbSRl/H1MC1CeXxPqQSXMcVQx9Rp7XH
MaVBwbnLFtvUkgssIjwnixfM0vZOaJdmS9/nQMZ7D/0EW/QWaG7+7qtFRdQiFRSnt9dK4cPXEiff
rYwNygVhrR3yJVU4W67HW/E5UXzn+0iKz1pFuhaNSDrcRT5CbGrVgd238en8WAxLr/3nrIwR8pnX
rQxBgG3NbyHKfzYErpiWpbOtYPDQAd3OH9Pp/A1IHj2AsAkQBmCCfdAU4xlvNRFASpXMF+xBmCTe
dY0QRkyCOXIoYPwp9AZmmVYV5svOhCQyG9bI9YVAYf/fXznz0noa+Q4e53pajVWpHxkhCz3Y0i6G
B36DU0ggm5VcvSAY/uECV3EsY6NT4o/a0Cl0zajB+tKDxkoVQhf6CHBK6SgRDk9V1rJ0Yokd3U0V
hH+Itaa+aD1xQcOD9g3RG42LGabeYw51RQ/22ShqTCVWrRdOrjo/IMyW8fX1IgPsK4PFNGev4NeW
0y/lTD0uxjhTWlT6jKq94+zdJ4K9MeXTyFi4tu51Q6rmrgitgVF4qQe7QQFie3rkMRWgRqZJNjog
XadYARTNUGgTNRRwB0OWmwmpbhC0Klrf+BjkNDCTYrke5XIwgY73rjXnDBIGNnS3OhS14vLDiqc5
NMJURiu3kmESppcfYouMXczr+lrXcImBJp/0pCLilYcAj2KGJ+swT0w9uGXweM2BS+XlWGkBgFWP
eTYp9eaB6bTOxxOiKq18XwDs4mmcTBUJQnFKCmsrtm8KOP3VoXVqPBPALMRzwJEaNiKNW8l3w22L
ipSEHgJlDxjXMxOfgCViubIPpBJgRMBB0DFnpuGSprZjCEQJANYu3zmJm0UVXYWfPCy7OC5U/d9j
tDoNYX3fS0R0XsZZEVl11W0GbmDQ2mF9NzvAJYQXsYW0sDbAdKpmKIvkrxG+M3vJCuVCtyZbt56s
2YIDmFS2NiAHW6IWxjoEpKrHsls0lMtKSzKsi4GqOQfSGg0AHZ5oJqrFXYgwDZ6v4J4KTHF0tgo2
IsxVAta6TH9SgNceUpjL1CAMC87sS/gec4Cf6sdW00zMoLky4ENP16a0ZuEuVg8ecE/sFmqOBTl2
WLec2+UidG+Qz6JRzf0kFAOb8gbeDowQG7I42g1KU9qIUFqeXoPpJclqmE88RK1WDPSqG+dzkbAC
ZnptTU/zGRgP02kgM+wfaKhTuTEMFBLacEidsNXHPmtV3F0u3A9llt32mvjXdU2J3gI1qCNoHQMm
KQMbzvYGNL3a8c8xnKl1QGdeUI/UY3RTh1lOmNUZGFSENphMA8RGcGLY39qN3YTc4ycrs1kfRzRh
qTDrKhZl7m1Mk3qxC84Q1pELF9Ht5Jv+jr9iBjU8/YwB4ETB787wWqmoblX6Pk6nRqFja7jsH1T9
nFiW7H39V4vXYx4SZmFm+ipSfFUEg/ZOQArtoOKIDOpzXCcw8Oj7MBq4WGqFvOLvuyxDL01BP+9s
IzogJAxpGx84p5IHXUlemoh5erRZDFQ/t3SlanE07aCYHqk5S++bJMiEY2cm/YLjhaRjDWT6ebim
2TcgWQ2jpIPM80NHQOfMXm+7Xq8FfvfJ8l1dlLNlea7GCkuS8GDRSsGGgSRj9afkCq8i7U/glT5o
ndiKfknj82COvf9mUNdpIQ4OY5r9b+wZR7H3ZtDPmk+WNmTcFLRDntLPygMSu4s9u65wSdW57Ctp
SIqie6J/LWis8jVxrM5Z1WJWU7ZJ19ICh+8f2gJbFRQyl0jcDvZEwjLnRBlXuHC+AM2P2NLi6mW/
/F7euY44Y0kf+mfEQ9jkZflkLk3wsVKhYwju7xYT2sK8CQXKXVDKMWkXHS/s1cmohdW/xjC5g5kd
/lRSfxAIsP1rvqxBGhTRcw2CL2Baa+wrf3AigjjDaeZGwDzEjY2/6h5JHvxpfkVqmeLhy9rs7t1f
drmr+m8g7NFzlb4fVn/nrgMljBEWbZrBohZhJV+Y7zbK0CZjrzMOLJWkNnvSNhAGFWerI/BUujaf
ZCkyXAK27p6tbklALQr1hQHrT5PoCzArzTiuFkCCOuTiBQ4Yi/B/N/ztQTwnqW85xv2mkn3kIuo/
8Oo3Y3EOOa0zdmpv27aCwryq0IiNBF5Nue/EfpXB4hJgeEmw7xQ3aVJmgc7N4hUWUQ0bRVjeOTsb
ytItmuBKsAvx361ZbDjBp1wvzVWKw4k+HIKBcGzcVsqhekn9RdGni/qznk4c8NuUqvi1bl2ANKG4
R9yLiMYZP+e8LTcvuX2UU0hWwUp7kZg2+If4CFX5UzFshHcMEdT/F+rTjWt/S85+/K8Ip2Vrs/Uy
dTR5rmBuq8/n9FlWrbv+z1VUG4PT6OgBXCzR+abXljjkfg327Q/v6nA/A0EQLaj/YGAyHPoxp0aY
K+p7B81hL56h4n3IzriKSfNIHkf5yPsODc3r19FqlsUXMmo9i8yu2xX7hUuiSZh8VBuBjdMF/Sbz
nnP9L6h4H99oIwxorZt8LPmJECn1S4sEQgznTx0zyn3WDlpggzlaLsU0NKzG+Geyd90LHM0YtVJj
QJCEaTCOAwCEb63iuPfCkIORT2ipDMr5qT18Tlc5E4s9OL4ZNF1AHpan9w2Uczef5qw3wOMVit7z
OiFlO6886NNV8sJzRrBULLajzYSEs4HwkB3aP71TH0IQvTvviZEo/HdZ4XNxwvpLK+D/qmT7BERL
uUocGpefmOKMs4a7yHSmMZP9ycEZOpemNr1slip602VNqtD/pUrfBUHCEwc73HgQ+v+8Zm2w29pC
wG5aDPvWIvag7n8cLc/spLUgdpY2UkmZIuQHyxjE+MmwA3Q7qUmoe/ogoDDsPzXwMvTHBB/qwOft
ulySAeNjM3DWf6fJ+wPD2NO2X6PG7eM4wyuoB5p6o65tCf6/itBOTjaahrqs3oAgicfXZWHbhiaT
M0gG0fAz51kGIi4VIqGnn3RJRXp7P0VzpR10YBqDlppX336M0G9ZywBnJavc+0+Ne3sPFhwMomOG
vkE9vdJyifVdyoaPjtpKqLNvY7Y+3mnNyFj7VuX22GA5DUxvdks2uAzNNfUQxB4KLi45zAsaKnme
GmsYEPFqSFCfTeHvejpyGiqPzFoie2gFqADnv5IVBOJqeNsh0Xmt0osKIKEAJ+WXpLuSdg+JxB9c
pTP0pzQfCM64vIY/5hXFtT1FBtbP/Azht36hvZVi+KvmDz6Gn6wq9DkqTqSooS4fkVaIDTurDKOO
5leHRwGdgghFK1dzYHNWDvnZlYyUNEYExve/bF5sUAhYLwhksNJnPiMpEnQSow1/lJ9Uz6UviKdO
chLOyuMkoY5kxCHGrOUIJS882kse25t6Dp1IMj7G35ZSCooVxpFS5tWMcd6VoHBy4ziKX9Jd8bBX
Iak7o7NMJrA4Q5ZOMb9HmFHabZWFP3XgwaU+B4YMLP7H5mfHRBQF+VOpuYBAZ6++z3cc5ZOke8Yg
4imLg6qDwmGuBmeOEMHPzxE75W5VUUe624a7GvE7O7F6gP0IRk1O+OW/Opmc8r9qzivuJrexiMQP
qaGgfxukDmFJw2Alxzuu9K7mqu+LEUEpKJmNwOdL9IwUdj1SbnrK34xdIhznd85bPrenLQWbEwDG
zbLVIJN3EI3n0oZFx5gvaarHQmCGe24Uavqvf5/Z7iPNUeyfajT+9k9ucfXJ02v/j6/q2U1ZNyDk
GiDlCMMVktlKIdHC3/P9b9J5ya364ZS2hLfUJ8eucye4HQ/1+opNG1dq4wY8KDfM4BWcnRXqF3wX
TmSr/XGwH7UX3X+tcdz5YfNZHk1j3/QeGmT90hiKw9oGmRNhW9/OiE0H9vRQxhgeib1YN/BrSv1M
vlvGt8MtfujMIecCZoTs3ezHAcGb8ZpUyXjy8u4tkpJRllQsTuICJOCab7DAdudIN+rK00Cc0Lbz
rfTu7qy/fhfC11lZ0ObT0TN1T/A87PKoknExujbzdXStbuXRyuR6lNrvmrm2e6fBCunSYJewqX51
4DdimIj2IGxXXHNsPtOPzesmKO/zBpTzh+4ppcQMI6FLJxFd8RMVIaS4IuyFHhQkmdqCuqQlld2I
DnN7FdHnX638e7fKd+2hb5kvcKDk0zt3FZ1QO2rKE6eZjVb7Kurb5MP4Kb9f4Fiz/YzCJggyLyl7
2fQgZUVt9sjRThbA3oN6iVY/hSd+aNkTpYvVNLFGF3LsEwMrlPY2TIW5MGDO/xikm1/hASHI7WsP
r/2EHC9yOwCKhWjHxsKhDwTrTgXS5i53jyftrWQlMiAme+Ar8z7HsnXg2XH2/458ePGJSpa4S5yL
UPlhQptcNSLGE4iQwERt8+yeUvP1K/nRlQ0i4v0s+aCSeYRDUmPnd4HYuaHikZtevlMt4PnBDSZm
ZruGhTmfcJsV/N2iGRKIMKjwzcUAdyx+Y5rzxWYJfLPAGkqooPAQOyZaFotw1LBazzrJPB4Nc3Gl
+U/N3Ao3mpqMH2sJDVS9Daw5Y/AExTqSHRPHtB5/21q9ZHJH1/62pG4q8f9OXOurcQ03ZgmdGIX4
VRznrM20dZgjs36pVY0CaBQzT9XUOUyTVHg6dCJgPdiRK+gXVsO/Az8T7vWSKCEUOPqSpQcLqnmg
oYEkxyHK6zn/vo88Sdy0pCiqkowNSrlgg8GQQcvkGS4G5wmw/rl8r8sNyydgCfADVtbBPtgrfh7F
ZN7ohpRuZBuBz/660eaA4tMEJinpBz4etPEtdWcRub1I3RAm3Bl+VI7eObNteb8kuhM3KNLD/rsP
+SuA1VD72NqqydpVsIFh7cP3jkz+Eu0GoyyQhZtSQiFW5eAnYl+iKiM6/DrXa5yV1wlN5wKZDkDA
aYZ666LEU6KZNMS2s8XI/kHLSYi9gJvuw4vIJcnJ9SzRwSPKwG5uSnGEah0gc0Rrb7XnsQBUJUj9
HL4ttpCLOga8ghwHrogiCP0D8PRtoHwkBuC+ntEpUkku00o7c2NwlGV636KdUPSwan9yIaZblVp6
U5aIMncFtp5eZQ/TY/1Dk6FDsnMgc2iuT8bfBKZengNxeigvFvglDgKC6s2Lf2/Q4uqho/nDJQBu
Ar+/MurP9dfm4w3DI++qQ/WqNZOc6KIQnVdCBySFzjvuXDiiFvOWlXJnE4wJHPFY/ZLVtAmFzuFV
iqH8JUuLBCTArWn4IF/6Gu00H+iBFTyVqDpalMv3AldTBSDbWWa+O37rp+p2qUlBZosYN04FE/Qj
Dbezx5HHNIdU5wcTQCfMf4r3NDXRq3RIUJd9aJOqaRAQnYN3PjAiiM9dbVu8H0yOM8FIZXaUXeYg
UaaHPzAX5A9B0KB6BaPLfbxtIiMiTfRrrivYpIYyTwpPnC8J7O3YcXXGi5QFrYBkfW59+SwL/10M
OhHz0ZG312b/uQq9pC/lTnMz4hwWjgJxwM8gXlQv9+6gXapNaOuchpZhtMyHsecxm73UkGJlrVFk
2YXZE39YvvNPclDomohcvnglT+AvB41KSAn9Z4BK0xibcHbg2sfE94Xlvw+pNnyUsMGLXxWK204Z
L4616JagsQWRTyN8ChuVslqmHf8HQhudZSt9BTz6hvimJ+41W0QCb78QMF3pBlzhkQwZvk/GH6iq
hz4y7GBl8cYvOg9iX2wi0n1vRGAGNX9N2+iM6LMf+UDKz+T6ATBIH8pgTHi3ce3jEKhWlt0sI3xK
35FV+cj63budm1QEjxC2BSUHEMBUcdkLPX2x+52l2GdQKaCBRkK/ym+t4mL4SGwxcm6dDl65i6EB
MI1eHgBBPDdqUYLW/u7KrRcsqncxcp3vWnYFx9lLF3eKbxchQeHc2+ETt7sQ6j7jGjt0G0t65DHT
IiOYUb4+84ltQR5rVyCbT7Q5vwRPrBwe6ZocWfSLrVaQxtMazm3qMmoIHG64op+0QGJ7r3pk1v3v
ej2qHJfkdh5pmDObglhiEfGX3o4rV1NF7IQfcPiWDuIkHIF/TpFCil8Bry8bxiPrQKQ+lQjYi+ZT
0sjsxnlpfRYQjRmhpLm11up5sjlC0Sj4Z8eKQQ2W3J90ISWsr+L6qmVh5IVONs9TR7Te2leZTnCx
m8ix2rQDtci0lpTbGiTPfMKBTQChxq8m5fETXzKbSfmZW91SERheMgYZi+y2eag3z5o4D9yHizpP
BDMQv7vmpFrgUSHKM0M0jz0flgMiAVLB10K+s4WkfjQKBOeWdDmEKL1+2bm1NK9H8KXj9MyLPRs1
EOVIEEeWqagXeDadLYJN5ykaDy571h/hmG5N6NmdugJN9RsGBaJZU31xa5Aa6q6znDFpfcSHo+1u
b3ZIbJCmUAqMnAH3yxs+x53wp9qOSE//JR7Vc4j2YYscEiM1FEHwszqjR3MpphNd3KxYInNEso9y
eyGVM6+i4VeITsxJjD/pBApAWHxsMV8hrd2OYk6IW1Vv8F6aegHuHTpCWimYHivMcRudEg27/Kcw
m7SRaYSMBZsZhCHgMAjd0kQ9r5VgV20Xq+YWhehQxFzsriwvLkj+Jzup+cNcosCWApp+aqSIzzrv
YcWawCfXn/dRBk98Uz9RWmzGs0UWjhomQadfhcdK8oQcj81F28AUAQ6TcXaamkXoM6GGcZOJPhGL
mukU14iw3vRSHhZPnZDp7f1o0r6fQJV3d1vbhdftdqr0KtngunTIHhN/DGU1c5hVQ7UjTXQw8hTD
v7zZsX0i2K1RGwCSWqh3Zr28T6hb8+ud6gx4VbN0UEm4S1ML4fW3dpgEpwqS8pfmuTzN2lJD0SIo
NcvOMg8An1c9FmWG5HWhDYEtgdHdDJaaKUiO2z53HpeON/xsiNCpE2QPTgdpDTXeVi+PGKjAnwUO
jGWV2Hxpc+m2UqaK490uw1KGEgav69kngqYAos5K8pZgKZULKiOdQhWPuv6GA9g4lLnC3P0ggD33
eGG+IDD+iEw+kts8kjHvopsBqrk6ialtDMkYG58uoDDQ5u7zJ5CRHTyMBQC8nQyTBh7gz+DhYbUd
jkHVyrmvqjpwWc3VrqOdK5S4JeZwf7HH/5WCIc62wwoKt1POTTYyxYVYkkwPqd3ypGixeUaCehf2
wTm/S0eBXytdaZqChgfxeVmLe4dNU5OUgxfdRTO2TzcEmgF5hyZa2TOrw4SK+LLnXudBfSnBr3yr
0tS26Lp1PULLYCWJbAUG7agTJtHIORNXJ6GQPrE94QSdNcrjcU1REz9v2u3bnZgiXQOZTR7cu3BP
qaGS5KmexO2Adst8WPeFlCMryshHULvp0gWAUkm/qiJuTH7Ci2mKVjmyBpXp0QdCS71gAHxJYlnj
/FMzS0LfpM4FpeKka16EP7yC5qy3O9CSRXv4/xUfh+ZkpxQseXcpCVT4N6bg5pOcwcZWnSuqHOoO
K7ySlWvCOe1Y2e6iUliTTLdsXr7dQfpWYtTnan+hBo6DoF0qmHSklTZc6s+/SaeCBE1qekfco5ff
UHGUvL1gsRw+u29v7xvZUb3sJ/Qdti1isHJik91XZsEsLKcXZU3ML6jUH6/+1nIKxs9m7iRs2+7w
O/LS7E3jHymHAyjAVdQXvQddE8+zeo4LSUFh16m41UEoMOBUA0cwS92wz54N6YSh5mPozEZZYE54
WS1x84xOXK23RCLTUB/2qdCumXWQsHpRf4ysYaNAehufDpiXzdufdNfzMXlNIDq3gYfKpjehO2l2
TqLaonOpgPGuI6sJLfvG7msFeHaUAolzqoo3cYJSGduFOb1LP5A2ExYqk941i5+cZXBxSS8bigrs
2DTm3WsNKrt3Qvps1XyalrXAbeIu2x/EJEUR89cWIRG4nQQbnxwZJFVZR4SwKoeVDZ6FRXcgrK16
OQ0uyaMyn/xtbfzu0ITdI8ahbkCySX1culnaIrBs5kZ/FJLqTZUNapDRSsZLFQSoQlcqfGJniIdS
8aj9BxH16W+plaaaE6Oj7EnS/UrVBuaPUhxGdNMad9WZvEAETlpcJQC+/Uw0LEB9tw+dgzbZMRva
aadocbFKKcQYgzQ4l6F/M+o+d6wBM09sPY47WiAtS7dD4/UU3wI9DMV//29+5tjCMkc7G/tG7wMj
1YX5KhJ8JSeWArYxNgIN/hcIA8hJa0N3nKkpgL7kd2akIUUKMD1Pe4ly96NsKGIGALIXFD3snFpc
hQJ9EDFrtT0Mu8YXRGB7em5R/u5FXq7SqKak3T6wJ5NLOSGSVQgwnC7PNJCCYo1yf36hwzpMZEwX
FyJQQ6vP5DoWeec8GdYKrAO3p8xU4BKGVhKEYjV/9slmZ0BD6wQ6/mq27mXa3Zvlj+azzLQal9Hf
mTd+hD5YQCsPPxjk6fWoJ9gT7Vb4u6wEBFkZ1FmSx7XNBvX/iIOaT0pqv/14RjS/ANep6HLn9l+M
yYZGng7NAVyNgW45VaHpQRJGGrr2Ix4+9IjDkCRH4YXuas+Hhuzi47n++QMZOAu/x1m8fcnGHl0h
zMeG0qqZHs42s/pnDWhHHWz1mH4+xU6GAK21AXzRb86DakBm00iUboHZ1kEB4ZxkHz1Kf8B6rc7p
NcSNklkMrW/DAtToHc501zlYYFs/rDCS1BGX5fcMhroBysrLPEyfZemwb6cOGeA5Ch6tgMFzicd2
7XHD84EA+HJZ3OIPI/fGDBwzh/iDiL47P7WoCJq0nJgGOMfj3ylsPQqy8RITspF8wEecp8SajY+C
9vUtVJNrwNhXJ21W2Mnjm+Oy0Dw2upvBVwMKHLdtVHzlZbq2TIe0z2QNZNU1os0hM64u5tFrZpDJ
h2URTX/IuUGBrx5AY03fkArCb/e52UfFlcUmHsQURcv9j7XqVR089qB6xZyIU9e6oJQexwi9PKLW
qf7rZfFwCaLp2Ym8RxVfqWu2fA6aYG1vYM75N+JjJCPWYmLkNF6UgcfA5fgZxNht210k6vjhep6r
UqDl4KIiqhFm23odk+TkqtFwFWKTWHqCk6hGns+e0NetFv+8xum+uRxDsHbQe6oe6xTWuyiUgceH
vu3UltEzQm/nnOuTbJfmaugb/d4Bt6f8H/eJy2GcV5kvPHNo/HjEJ2KxfG08GnL6T/hm1ponTmwG
lPvmUFU5QAB9NwP4uUECd1YuxCsIwEq6lCqPGHI9ldJ1ahyeJlVM4QR1XqAy83EVe57x6j7oLKJg
PMqqozCqYoAfLwfpZ8OYgJXtysampsVLzQPdx1Oq8+aqxQvyBtH1j8S1UJV69JzH+7rB9OLpm/Tl
e3hmix9TtteGrU8/VEcrqlB8H4nH83xjzvHA8njTEMMZvBYJuNwWQ/fK5TZCgh4KcbJG4trtQDtL
B+yUCTsLFrCdIVX6tGKM77O7+h/aoAw9d19MUDBE26EevSi2D/8rwYOBI0Yvaw8+QThKywrtxmtb
LBhi0TbqTid7DM0q1yBeSPTwTZgYBVC+r0sKOqDB/7REoBbmHy6GZ3SYPLS/lW4IxZ1HOldWfHz5
s1A7DWiuWONuM0e9zjxHRvQs4GvKaYbZ/YllvT5WwiXSJsXS+NXb5LAQjcaMm0bLevKoEs4qwZ4S
lFgzxMm1nYP0+5AwcsW6d/U8LANDOPXF/wqZJAKI2D++Bi62SqCW9ayawmXeKcUbJgJSc6lkvpcs
lKsZn+2Y5yQSnI/9Mz/B1m50Ykca6jUIa3FNuU4AEuqC8jpIOxbvRbHst7mLCzWQ920bBvIvPg3+
Rz0Bl2rhIddmDNomlNwxJAO3VedlkAavyS0+D2JGoAskIQo15qxwsJEuFEL6UchuR+jzumbq1Ynq
DL3h797Mjc35WuN4nPo4RuFChZKV6t7vP2cKh+B/FujikXJent1tiGIQLp5Ka0faEZYnV6QAqPVj
nZdApaknS2sHXlwtq0xpfFNbQwocTxUg00rFPQJB5EdN4dUPtz806pkhwggnkRp6zgwgqqp/apAj
Un+/dsSy+gUKtVgSfeszKluCWZrI2XomQstoLj+npYyVqv6sXBoQAYgAIAA9+3490MAfqDEixVEK
pjGS2H/5nmxJH82DgaC9vT8JPS5idUwv/cVbjc5oQida32MhvcJ0lNk2DuBizgkJ/rRFKropeX/i
GhUMZDP/TPw9med7KrHfLEtX9G+hem4s4EiLKN8TzVLGvdZoWUWKJs/rC778amxqvhtUqwQxye57
05WuvpPr7iWWfTD8vSRAmmSLPk54szEW7WmQaXRFolXVZVr59b9MYKFAglNIHzVBfCg19hjq8wsf
/BkpDH4EBn9mVJxd0qibn9ha/5lKXPoU3EgCdLPCP1nPnv0tbYPLv181nMFZDvG9mFdudMD3Y+tA
dkNeLxkI0PHXxmufmzNwJf8DypusDWYnJtSSzPejwOcxx43oPSuJoN+ReL+aS9R2/C6PAEb2oWRF
M9d78ZihDLWBHI4y2NlmsROlSNHpzCt+le41u/bjcL+2IQWARs1g9K5IB5TvDt0JpxbNILnV+gMn
dHnxj8LVktMr4GYfISF6AzD3DsMcQWL6V4MqXfHWKpLPlCVREamEy9eJVBgBghxrsAZkWQmjMDZF
in1F/fnSm70Pesw2DicHiK4+DFbcAIvtJBh5aGuoQtyi5eQEEgCqCsciG6C1riOjFUCRcN8Nh0cc
bRAOoNVZ4bPlPNZDGVu0b4lvG5TIePYaUb6MTzsis1UpRT7xGoMxdyKptU6ig3yi4/zqPcmToocb
hfgCXEsuXG/XCkK6juilnhVlb3KUs4MwRutLxTVqljpgUOdIKwv3EtxVXQA2v2b05tD3RzS9SMKb
4LrUiAZQhig09k1pCGqwwCPcKL4wSFUsfUkeVEPeMwk4kzmp8MveZxApUQkx2SmX+gkNEt32kSVH
qNuTipUy1gO69x5Q6DCT4i3lSH8aCfxTv0fJfdtnW7nhM+OApgDX+SiuOxWcMvHF6f2pp8U6GUOd
405fgi7yU3pvnU/qQZG3C6oRIMP71DIPBCGgVgMT1F+NU7T8+egy9MZgkeYr+PcmCaJU6FNYoCvk
pGWz0cCTXg8HIYj0SZjQijjfCbv1tq4naAnEspf1Dnh2Nk8lCCmTNTetQWwFtkI23d9TcpskYs5a
is7Prx6ftOF3glAfMgxt0g1/BRUNCZFCJuGdyaaAwNBpgTVwdN1AiQQHYbQu0UVqFi8NrYk97jh7
Ph3aaxsEzwH2XBAHyvYpPgxxtEf6D7id0oWmkvlHKxDtMmfOMXeGhxB3NVvjJlRH8VMSvYCd4VS8
7z+WMJE/WDkHYsx/Y7n9t0dM259+4tU2UecyRvZI1xE55F85RO7s5Wqbi4rVqqwIJtbsTW+GKtJL
G1XfZekPXyQp/FrFtfy0jQ+gcnL960Jbnylwh4h6Kn/Qvyi1/jx/cbi5r/RM8kxuNu6i7FR567ap
GYgKAiVYcpGnu3L3U8Nv0XhMJzdczKOFYqzF0Wyn+9ElvopgZsLHjiSV+PBvYSrgW8SV9MHISMzE
mF6JlsgnXeNCB0ZUYqBjtmjbOSblR5GHokwkDp5IDhZ6VcSFS7naVKjxNcEcB/a9AXsthkLKsVgL
sfracj8u2yqOG9n/QaAuBZd/lTzB5C3KP2hUaqrmafj2/DhcwLeXkjzz2CtJ/DdwkKBKrWCkWzFX
l5KL47UZqoG9hWrbgDoWT/Mr5HeclXHV1yBXHW7Cc2T5ihiPlcJ5BnPcXKkA7QB+soPSgRJGAMQZ
BeoId6UOE8qUT+EO1EiMSTiBeADS54SmEMqIvFeSwcff91KaVRp8vRxZPPjix8xZ8wqxZnhFuPzL
+NtjRf4wnMuYPxLrbybYpr37+vrtYlHyYEla/fRVqcqQjuNDDl/BRp2NZTkZN1XSyx1HrNALUx3l
arv13gIe1ga63QpBMcqrqeH8BpdBko6+97G/EPyKBFQVxXSev1zYZFApvijzkieWeQ3ZimD02O+Z
GhIw2vQdJ4hrLpvvvRW0DXcqUT1Uxi7r0EFEPnKZfmQVX69m6+c0XyOimkq2R9tyBY9OR0qyAk6n
twIkJLyxmowYU/QClEGbNq0RqmFBLSW+QrnN0O22lzYmd7A9FEpkp2k1WTXeRjoG8M9GYGB1SBZ3
VC2QLPxKq6uursG5hX7mqMuabm9x1V2Zs3yjtkYmAq/JPw7QxehcUyZM3FXG//q8fEzVcfw9g1i7
QuFXqatt6G6F4VCVpstbJLshT2U20lUwH7KlLYol6d2yn0zofYPrgHsHLnqMJaSwdmemgsOfJSTz
0HUIinOcpW4eeWywhbhRZdy0kua9b7m9T/5Z3IhodAlty5gsHCtXnU+dVRoAo4qSkI2rkELj96cR
S6NQteU03XcY0FxDamjN6EaNf/einGNJYSHbngiLaHlvweKCMEfUiCHiJEc5EUQKCH5ms/WMm9UF
nuo0xQPM7eDwybC9KH0EmK75VnazEYq0vuj+H6fvqdJMbknvGyurQKgi5IDEnGDu5HLh+RmGAkCX
ACf9lurgROTte6/oND3fIuUe4AND7VDji3EPW4llkpV6p/OlIfJ7h7oHk+vnp8svSN2eteQ6y7fI
JHs3G7qSuRaadtYfqORjo4k5m4CLxw4X+YQkW4sOEXI92/6Pn+okAii/K/XUwESm0Mzm9ahaBESN
mIOz588ozOwqYiiVgfHXIoWbqWgLSfoPsua4mxCPlV3QR+U7SBo3W15QvcM1MLB8rOJD1OtTC0sC
ltJ1UC8HM8HLIVbXn2f9JMLfdKenA9dYc4HCw64TGTG8HTF4F9IPiFTHw4MAJjZTXrQrCbe1uikL
xj1XlRtrc8CnpMslE3t2GJxlVKKm7l43GqUXVU23slO0zRSynix/U74Udep2tNeBsuwLwpgfgHOl
EiUCeFcqULWaicwvT1GTOuag+SseuBi0AJbOm+Qzxfxf1qkRje/hpWH2oxFqFIPf9nWOt4WNS8uK
pknu5knpAKY3/kkmOtQvGR0dnLvrC8qpqSYzk77bZuk3rWSt4EBYTyvqt3BoiSiTzGU5XI8B9v2A
kXmEpIbkUAPLS0xf/mjimTShB9yvbtkffKmec/BjDS5j0Cz7JpYfLlcyZPadBS3c2xGa4gkaYhS4
3xidl3q3wHzpjmaPRI0FqkNmvVLMzucx5lZv49g7odW9gZvjvv1zW9T3ck2zvAsLrTcDzLzmSLJs
8jlGtpeWxzvio9jA3VFpO5KVoa6Zy5DBugvhJ8boVBCQceVGmo/nWPoRL/ZSbDiCyyqJ/t7/0EtG
Tkq2tJGPfovg2Z7hGWCMO/tCcibZJIddDbizo+7SbTsxQ1antqpXio1Z7iXrQ0cynJeszKuSMt4p
sUTZ6u5+NYHOYno0QJU3R7tWCcm9PMUqifeHQT2BLjSfBIyHAl/nyPscDIvDSeMD1Q4dgxgWHj2z
qKjQ3bb/CdkcyvbnnAloCU7bfLAiv64+TkXfennGT8WFkLbPsWB25pMVRQ4SibprXR4YsSwTKuUu
lzAcUOqPCD3QxKB9uOVBBVxdjaY5iGfWgLHgoJKriHikcUIyhisGgByh1I1dw1SfTAtxVd6MRtEh
OqfKtOCoSKZj9LGr1wj6m5NfJJnFlarekA8pBBQmNAP17zPeq9hOkL928WIiJpGxRRoRp8ZYwd98
3NPJW7Use1A6alUN75Wm+dYP3o2wF6qlayKDjqYS69US+5jHs92uly+QaJT2An2y55RCSlvtUFol
dFSIHvMXTMiN8atOVrlbGT8/RaQHwELPNa21tseoAI27sEZMHqzbvqYgACF4nOo8UxhoGg3zRtwD
SBw3odUfLcjSNFa8O4Q/zaybl1WQXeLhFXJ7N2oOHLQ1Tnid3o26lLU4upbx5MUKdcs+FuOvK2/y
P2bexx9dqQJdXyhPThRLI7kMfucboyqS/rct0xOLxWmXeZGfgz6+dR7sdvjXLARtKrNeO7CFwEG4
GWg1VjGR+oeZBCBYQ/Zu36oqUQsvcIZZJFrm8vvkSCZchIcYdspeDIxoY4OTUd+dpF6mrdTyJKzy
pX/EELYlOPrjsL1SsP5tDRhuJMZzzgW15aIxfy8p/LmI7drme58hJDdarr+Y/uGjXVX2HWRih/sG
Fut1zO6WsxIJlSw2Pc9v4TXy66U1M69lu/mNeD23/RrXNTjNlI7kDYwvTKX2lxBiTm89uzeToQeH
AfoF742hCUfcUFgzpuw2dsohnEYBMojN5bw8aH6yRNN5sMvBTXRMte2OefLI6R6sbOoc9IlJem8+
xapYU44FUPtyINL6lMGkrv3r8vS2Nh2+PKIiHZlsSUdLHmTD3NRtKDaGoL50IIZns8HvmaV8gaZi
U/o/xg0sLi/fr5BISffkGoESGK8KXPtSRgRg/z8jfOrrwG6NbUaPxpsJfq8O64YVVvcBU1A9bVZX
8xOrwoxai3ecQZH5sbQwc3MG2dYV0MpEHMjKn556vioaYQhEVxyMlmpJz8j5u/jdU7gEFIGoYYNI
Ig1VPrV0lN+3ri3R/jJ217yAuNyHn3OUcpPxVmbQ+RpmzwZ3M3KE7qoihIvzpJuNCYTcvH5Qftgh
LBGERUBMfHTZBs2vIXmYXG1//qDt39yq/hVe0UbEf9/qsLjLTm8clieo/CPHaPKR7n6JiSUZ+QGJ
fJkOh7A9GbfovjgS6RsXDcizWCSbv7iX296QI8aU7N2gUj8ithNHZQsmNwtiERMyyDPDqTg5L4Rx
dNAhY4bP5LbnCjh9wKvrF34++2HNW4ZiTIkhMR6316yARNdjHMoF7h0waWABOBxefmtGuH11h2Yb
eL8R0jxb4nlHRhE1H+st8hClnfvaa1xfKV5Th5+qCt768If1qzCZozTxyKuLOL132pci4xpJOKT8
MCQTsIHlh1Yx/aBfXc8CuwwkYp6DnbwJcxR8547cYGLMJ8UD6tAEhMZ5LGVP6lCRvc2BIdEpoEe7
fG2z8p4tQEymcLB0ig5+RarL7LyF4Uh6GN+nVDIGFrT0vrSfBio2612Lmxpa/ePnkoqQPzSlI5Pn
CtYX7K9LkAWS9iUngjDb/YMlJjZ1bIGw6zX4Df8fUjgNec9ySLnMJ2uYqwEBjWoFDz0NV59UEoSy
9u8S9AuT+z2WAKgy5twF6McWiQtgwRiXte60HIQH2VGVGZwvCYKVlW+g6DBZceCNDUX7DpvhuaXj
i3N/kOojXIaMqA32cJXfbIzxiRX47JhnMm3yOEZvrZ3ddhkwaWwqOZJz4g+Q3eQONnFwwiZi+RG1
zty7HB9MSDzVvbTlwCEq+lL+AClDyO63r5eTjT1sTaVLMzCFjflOa9XuB1vlQ1m5tGAg7cczj5BU
8hK2cZE59fN9gIzKxR+3ImhQd/Sx4q55nDXTw4DKjNP5TVJ/aS10xbyqyxVm8A8bq3LSZ82sNK6b
vbZuWlozGVw3cZj5pWqMjmmhzhcp6jcSWYpVvkdNa7owUGHcsx2adr1micXLT6bwEgnFOVthNUYP
h47oWAKyT3sb5ifjAEOcmmXN/NqOwN/FPHVArtNY7jwBzM1Uf6vD6rw9V/0Bfv4EIQTXliUxn+Ar
OAO+oawMFShoX005fYQ+hzHEZ2FlXFi7OC7L/dz1vEErAK4rH1vpEsUKalF06psl6Bbq4Y4kTYAx
+P+ni7KizxDHf3qS9LdspjZmI1qHseG0fJiOu09pdrgc+NDFDApCLFtEmEuWRVY9AaWqDC8CETUH
mq+yPLLWm21RuKqfI8Xy1yotLp87g0QSaTP8Q/pEixscNRxcUcDN5fkmphBmLG5qQE2Ej4LH4iMC
ZN16Oj42QvHHpXqxq7Z4rEWmYEq8yyzA5h/BneHyTntgBBT2hBYyT0sSUtz2KLjxfeBT1NfAalBH
/40yd+XXzdGh6C/R0lONYPb27DoUi/Ao7SILJOiXejjiAwwCAb+ZryYHP37/gIZtRFDWrgfGfSZ+
BjRKMluxl9NlqmQIIv6BmtrPLTOP8IuPD+D6yNypxG4qV25jl8v8f5Sl+/U2TnGfcXKJvVGomijJ
Y5/0zjlhIE4Fz0Uxs5cP8ecgkdbakUpdKBnjlI8KdB4W/1EAaalEFpzjaWwRVrbZDNqX0VD0I5xK
nwpWxiAbEdgO6BygoS888X1cJ7FEtAEKzxrPmNTbC0ZKfRIbVPi0IOyyDfPc5y32h2MVl/yU8RIK
AFeTTFag5uDY9OPyXwNL3ZiEmpCkJruDiOMq3y/+wdYVpvraKB42xGQgtfPHF77X80xpfTPl3ai6
KPQZRDSiPCDOB/CWTUlLWjNnUB3gJg4iAHFI5ObkDdE4q9MTJFdnfrym0ElibUbGkzHSSQiefwmT
1Yt2HY+ZDN1q0uWVJv2voA9QtTRJSUDHetJVH6MMFoR2teKyBc6tEQPphHTKgnig40kryMewCMyi
GtDU+7b6VO3vaY8voGPjMMiZFv9GPS0HWoJMUHujrE1v6MuybePpcyRY9etHkM2hNpwhMCNQUDet
mD74ODEk7YjvQ7hWIN3PNtuOoViWx0zeh77bwscgXWObg8h8F/yVhdEhiGvP5Qz7HNc3gpskmD+i
2XiDndCkpLkljiHK2RpqcMotSmeyHgsJD3sKZL0GpTjSKRTNhVQWjP2msro/umtMexNgf+6jL1H4
hkWdcBv0rTAnTLOU9Hq8FVzjmoW1yvXSIUsIXR/9hljkZdDJuS0T3iDNSrfMCjeciuoCesg123ae
t2AgIL4+nXS3RCCPhg379zNozPVS3KkRwwRZttTmiV/XH1nrwcbEUkdGKA5oE9kDU9d6JlAPjsFn
Zjb3aZTWGzdeMiiqkriIrNpkDRzBgJD48Q+P7RpCvui2xNXWHMYBXVIrTUZwHhlA/4kG/K60BJzr
nxLmhCMSWGj4DhJ/+cmYgmpFGHst43ZMFLFREAzRLVmWmKWmVjU9V96/KOBCEP6yok+kOoZqyEHl
rWBWWEKTcvchLBann5QQ5/eIx7C1xKhcsL0pKe4OsXeACXXujTjEJKFPT5tPWxCcgv6G2sfOXnMP
+3RLxxZKSeN9fSpkCPd+p8F+Z7hnLSdMH2oz1c56rkQVn8sL0rvbT4/GLwXcpYxsYESnDQdg01gv
gWZVcW2skZY5BSjjrcyw/Su+tOBlA1/N3D3xqFzjlRIq/N32L7233UwA5RjAAHfz3D1MJ6VwSdsH
iUyRgU5LKaw6FIZpjLVKeiROq2iAKEMRrqNMg0a4BnC/VrPCItt/IC5BQ7xfKtOH9YEK9vPagPyy
oPoNgP3GodSS7zARjTI4+QZrn+6C6HVYZ0wXaZ98TIbCVGpeLdvVVRFhGlUNvc8j0dZe0I3arEuv
qAsK0PW5W9i5t8CZ8tjlIeV1zkHAlMp1yGAxXKpXxt6+qEHX7Sf4+oYpsdkMjiMkc0XKXxy9xs2F
w739JAbsVWbQUnGzsf60vVwiQTsvtP3BsV5Y6gBQ7zv6is0a4hRJateoX7yXekQuFy1bKZIcHKc5
TNRB03LoXtNAvWrV3HP2J5f3Qb02ajF1BJ5rrhqBPU07FmofHlGUgyHFPoNNacWX5T85GOZIPYU3
xPQ57gWJKGuhkwYl0ExVTdDoefkcB8Xpv23R6uihLhd1VQfQRh4kxEJ8DQ3EdPShliFKws3uPYzj
Zt6pzo48EXdNHZSRvCPXo7/rbwaFLjbrNckS9hGFdgYRBk5znhNQISCKjZ010pwEQ4jPAwuX4qFl
JemugzloRbbSHxkP3JPQlIwLAspFjtLOdwle4cMQlztWXM0fDX7sc5Q5DFyDtZYTdMTw19CH5rQO
RcrJmH6hTLjHs6j3a+KDz0qvm3dP3ApTW9RU/TYt970W+ri6ebJhuhvTKDBq54G2QcR6LQBUdmyE
J8udqs9ps8S5CnR1JQhmBpEbAofVsX+9BRb5iSQbpwNAmCAZAounnBqMtRmXGioll2qIOXrDyict
9a6Eh/zfZ78BdDEj0zdfCuuPYhI26+TC3Hmxv/e4nY+oQo/gsNbIkZNK6cOcURKh5px3NOLhzNuy
Xh9T013k4V1AvLCWDqoEhraMPh8RnICBWH7s/jgVwIcgYlA3K6uwxXFwiN1N6gipCqhng4mCNOWg
FIRwX0Z4xBFvr4MF4+yJ0gJmRpv+A42RyT53X6r77gCVkQY2DJUXW6OEIB/56/1rxGmKOlVgJ+WH
FtvKP9WuxtBbdGLezjTOoog3tSfp2bYPLTYBM+FbyFCWMi7o4hCs2mSs5rU+mV5mx4EEt1HRt3KR
ynW6FsaFdpruJ8Cccs/KVRkiMkrwr9o5gNF4utWC3Dlj+ZVi4nG6ulz1z1C/dw87Ql1GBoxt0Woa
tktbiIlJEUXjKqMlmv9SmY+qZajvClXvSLhwLORQVcmkwQglyrGxZHVJGWtQbEYyuXVpUq/Xl5uV
7//g2vRszuCYidqRUTQeEirKqrTyYEcsuBFCo5gYNbDCsNnR6nLP0pLwjZj5zMGUmfJNY3wfy+pu
PHT3s8wmcoiun3XHw1D0zFGvdXpqjpPhbJQP5xEBk2WhHFjNQ/wxRirfXFBbpyRfDDhBzlZ5rdq/
IGN90QwsGcoQft0A3GMuxn9mrd4KR6LjfHuoMdtwsgHzeiQusXmowluXuqseEPFNWJaOPkJekskS
gXlMDY/omByp1TA65K99x7YrQ/xWxqndYP5OAX/TdJ05dj/ktbCHIZ6nEt2QhfoutSg6pWIRpPdR
QPdgT6WNZCIPJXvJXrVWi913KXNOPnm7tAom7H7KnOE49rISqYs4KynaKAjpcNUGhhYtzur3CbQc
s1zqfF7SLP0xLZtcZeDx5XQbeC0oCs4QFEB3UW+fRTkfgWRy3FpDMNApuG1km/0M0grJUDYezjor
Wx3pLQsLkK7lVgHs7XnutGRB4vGo1SxXqPLUVOBs5HWbbiexTG8caStgi10R4Ywp6uq7IS+QR872
IINl7o8PLv0LNmGIU2ysZrste32woJR+GaUlBXbcvpK520o46D35ZRBiYeMx6EttS6iljLy39GqP
POazCzmeG3LaNg3xOla9eFwlzvMncxIFnAhkGZ7IWsxD0LqudhJn9CUXcfdzYYqzvKigQIiyRe+z
t+2SZMoL8TK06V+stZkK83z2sCpBREFGKEaYFnEDF2Mj01N/UMAT66sDbBioEEcmqF5CgyrMaoju
cnkOaTb8IkfeO19zltPoeo3I9IvAbJiTXGYY4vgVVM4O+KKOLgTlBVn9WT3o7rX2rOrmQLnhOA/b
ByLo2iTfyTQpUbkMl7nj85PHL1XnLoFNRZJu+NZE56mXVH1Qu+OWEDd/uCevKPcjWx6sykWMY87g
iPvv33I01JMGBLH2SW1sZTCAIVC12e3Jwcts50rDaBQzGd/tkZVs4pJtNyCh7xWN0tVfQzWM4gEh
J2JVMSsLmNSK/kI1SuPVRHzn0Mm7nAmdklU+qT6GEj5ok64xczsBue7PxFdpmHcUMRAOTjLDebRy
ulpDkfEWF+F/Dq2OQxIV67RAzfUFr0QKg2kLcwof0Y+BMINdl5pLj0SceRdx1qdafN+uRbL5gb3P
txLxV1Tkwv9OV6CuY/GglcCK4HWdKEgfSeVR0HzMaZDftqBFqGZweJmgJJwDGLR76Zcw9y7vPjeH
4T/Lo64HsUJYnryfIN5sUYjxzGNowSGCzlhiIGWZeKi7+c6sbVdDWu6vozmKoW/TMMmw98Zy3MVx
8592EuaL5nKIYxsSBgpxcF+mQ2Of3DONeJP5OcIrPritEYz3gfPovlrp+VHrEDo13ZHtvNrqYHLt
Aks7KD7a5TarzMPQ7P5W+W8WpL13xbdhbNLzpJSap7JE6QiW2xVB6gp8Q+VoE2VerZNZq6Z7RNj1
joXtw7fQNcbaBCuNG+sqb52H3kEOZqjelGIgVxszh5A3lRXKxjMDiZhngfRyAFLlX11yazkLQ6wB
xPEDAnLc7w6gi+ANzH3Wy8fvs2rjNUaw2/t8DWURMlkMrh96tPpYZsB2G4P/FEP0T8iIPzo90A1V
nvy4/QJnrspWaxjPqei7fVgS9f4PlxqoZQOkLLS3s/jiwYMmApVoys50qdTO4Mgwtc1FhEkDsP0l
lmMya4BxfTYGVNe1FadZhSfbjiYFD3zZX94fH985EaJE2g2EjsNKFmnRLiQMAQSsMEfsdQycQaJB
+zhKjhCJMBPVJUW8LHLCPBLdrzcA1ZMml8R9q3MK+N/+3hrrxlmCNMv/38f5fCxinaGH6/EM2D20
slcS/u1JRXncBrRUg0LBCdmRzmawMiqVMu/Y9w1UUg1NJcNYzhwPLsX7hQ/CevsNT31N0MTLwlJp
9lqL9XprsCHB7i/SsNd3yDHHPuhNkKyi7/7V7Zi9puW6rKu/sv7Tsc4N0sNmnYyiH9Cggbv4m8YP
IIXTfXalyobwuKALWZD3jIH3n5g38300GQlCC68PESq7CJ8Om0nqwY5vNKWRgk5LKdbzgq6or8Fp
yJ7WrCsesOGkhow6nU/C44FsPpPvS0DX5OuEgGJGcB56r/Ot2rHjTOQGLpB9mE1yJMUN6qh67Viv
pm+pRXtG6TWHoZFagD6PuqWq7G54RNRdgbxZ3DrRsLkTCk1WPg2v5FGidERG/focXEfihQCjMSaU
vhk/yo8i5nw0mslpKFXbcf+Ft5Mwbgfm48AMpzhGC3hNwDCrZeQvqc6HCscXLj09WjTK0x0PY5Zo
1SNts9htIy4X1U40ODb4ZjmHB7uQQmrWAljGJVfcmsTOTQvt6xjL8Pk8OQZ4GygN2Gwnl2NYZ9zw
awrZsV1SHGMX9hbz6QXEErQ/Y/sUHQe/ispKcmhQpmcneD+t2sXqRosruHPoUVaDlKOthV7z2QTX
Jz+zCXeeb2MqXxcrYay6NfL+IbQzRrj/60jcuADiG/2k1euqRjLgGgpRj055Qrf4mpIc0ANma0YY
LkA6Q8NP6GZEv29Siam/ps70gMp41a/pN0NkxkwFSAe11QnibsDaqC9ZTo1N5gGL/OhVvfmMMUet
xr23LWoBO7GbwTUn4YyMVEht+BF6iHDiXbsL2AMOLeoaOPBacWUVx1LU0cjiKVPBGuyvO+UZVCQc
MKZIfwiBPwLGGPzwRmS3NOHQ4FVP4g6IfTD+Vp+AMxB9Zxt4/2nX2RL/yVEKh+bbpvuIYH+prCjT
P7mO7Pkdw6kWM2etkGndq5lXr8aCeZECnxd8yAhcWgksTgbkm1YT3yvfOpxKlVPhqPO6DWc6lq3f
EtUqKvVp/mRxr2t53qe3DfC9K5chfWwqbeWxKfOry4VerYExNyFHWhKGa41/DT165vN5GUwNlzSo
HwuunhXGjhpaAMAiNY/iWyomiIcStvHy80HJwlhQeAA7NjaSiSLC1QcJzj/QBxFQTdEepBNr9k+R
oILrsbhh51cz3SaBakLPtYaUW1KoFyWmHd+SbQFrsQkfi4QmjmeJM510Wk9RdDKb9omgyRQ48mJp
nQ9i1qEz0D1iVOvomFy/sGn/E+0M2XMYpLPLb0YUTGipYiOa33oAa1gT9vmv8YdIGUfR9jjr78t0
Bom1VuQY7hcNuuUqQs/1RqNgyUsHGSi6SWdUdpjQ4tPt48u551GmAPDDzmqOqZ+R60/URelQbWoT
I/h5g0OF+2Yft7o03mrLYqNPCplWgu7uGFOOr/A2L/hDm1I7XS+GBzdt9u4AGVKXaNY/8NHLP77X
o3Y2SZu89QClsBu06riO1optq0T7HENmQtJtt9kaKGJIxeO7w49tH1e+eVWJfBgUX0irMQdt48C+
gwE7GRd1QVBMQEo/hiLVrofMGrGdsq86KRguUN5aBq36xROCOlka1Zpm6A2lEUSYJCb5rJMySjzO
ERBd5WaHuUUjn8PgVaxkN70OJbUGwuJp19Q+S0OrdH2g24eC7cmZ0a+BweZiJ1GHZX18Z3/+3NR0
2ZvDJELb8E9lvDRI3K14cNVQp/OR5pC85VcWpcwU6Ys8bbmnjltGLGoJpcVYQ56gNvOkfNKY2MxM
bW7KdDMMep2YuCx+r+mrmAENRp+It1L0hV039I6DAMeLzF2XcrC60RihggPBc5xWsVkzoXosUS6l
s99eeT59gb9CatwK8S2MFqhMSDPQ7E+pBo9YzH0nlRCll+GCsg+HOUYDUaOQgDMLwesRKSWtYOWw
C61JBuzftOvuz8VVKP5vRMDjpOfJV8FO4vj6PGzog/RcSWuueKhrzacKX86H5qdHQL6GGnlLC1mk
tWJi5OJtKMZKnNDHg1Zh6QNukGv8SUISqIPwtj2gR3xalX1Fkt99N0JUf16ugvfRI0jbY1Jl+6IA
l/Ue7YJEBHBkOHy19voW9kgsPAJeUU3JB8Sl6esaJ1ylsdfDUYcNUf8L6EJH0R6iHDLvBhokgSrB
P3qoiRxVdvajTv5fIRrmairjzxVYystyEtU5MeG9VEnSojVqAlqokNwitkrQzhHsrk++WYN4diwr
Go5xALhDt7wRRwmsldqRZwBFH+9vmMyyF8tXUTgSI6AW3gT33T582Zqk1dwCtq4QjP0HY2FQtshK
T/xG/8pDIuzxgm1ZvDdxVK4HcU3fphZiakNMznicZIw9z2eA+mEEIVy4gJ83SFkWUk0UmShAZdGF
X+rikRh42g2NyxifuhC1K5Re+bRWLT1wsqut6FOQ0WwV0KrC/wbw4BY7f7Ada3VUNfZ50fmfoCoC
U0pCMtxXmcMFzC7yhlW3LDgmCwKM7CZg0GO5J2A2YIkpxo8aiVjSqh6+nVJ7lNZsIznZz2qEHdui
0yA3jqsoCPrTBdWSkAcJPaZnD2XAmEaERahRM/cVAxkaa4m7CKSZuJG0bq0lrEWe9U1fxSPgCx3z
Q4oqicuxXhELtm+CwQGwVDz2hpe++0jKMmIGYb1JnuqMxdkaYlLiR4os5C3yxSZzuV41UjsU79J9
7g2YJ0+EUBbHG9hbhOINKpFOPvWvOjgJfVktqpIbcQ2peznquzgGagJy7F1Q0q3NGs9LZqvJxDH/
1HmU6CVnN0X+uGmof5AfHU5j39xTyEbFdsC9IfttdZ0P1GiwQbHjNv/aso6NftDAGAqpwjl2x1RM
/YAfzy4CsQcfUuAPxHb6emecHNOfOwYZyPXCMrjkKJWdtEG4qJCvmwI1E8gzbn6dh21FyWHf9spS
pfEfHENEoBZCr5Yziy2trxYItOTt8Lndga5XquShDhTc3feStNzDVV/bvLgua8x/A0n7NUB3o4fQ
6Dk1msSQuzwIHstcTeaLurR9j8kiQkBRWEbBVFPI20lcjt7d3u4QirXQIGOZll/6azqbdOQVl7fC
tOCpBEofjepJRCyb0Iqizb1ePVJYPK0oa5tGDMNN7UKq1J1jscJAwp/4tPh4hR7B0Af2goG49VPN
uzQjexSR1EMuHZ8MrtdzzoYgjeuFTBLa3gIZ9B1fInX8jxHn3UwzLo9iSyWwbVpbrpLUGHDix84y
Bq4/K5MlSlTM9k5rEijhl/3MP+gUB9XhQf7P1KbYR7sjF5VJrUAeYEebZh11CxDzeZwa5i33NTcd
I3NsqLERCBTLNWsifFIHOWkI7y0wUxoPXbaUW/rpRLU099l7WpGODdEWQdKZQ7gRc0yIC6nPGquM
u67caoXtnkOPufJpBzSEbwiGRfzgPq8cHs5qWvpquFvwKAcyPIL0fYLFyazzeq4+8JjxtYdjQhnt
siaIQmcWUrQ+LYEWcck8yK33vIkm2WcBm7atrN9pRZRDSiYWtGCj8PrcZAIiLAb1VXFoDyUdf+Un
T8jVYQGXq/G2V6D5ZmiikyCnxm/TjGitoYuI43QaDtmtgMBMoeemAFGDTdehYFFGvUsqbYiZ0Sxn
U23rufsoBDS2K2srI8AERv+7wrodN4YZci96WWuZwTDUk5VxTYRz5V1hyQmjnWu/DtSVSWholWHW
77p9DelmtF7LwwNoayPHmJzb0qjJ1uPeAnKIwRSy721bLcbLaTUaq6UaNhQWBhGock/ONFofAXZa
lYSIeZfzSsVG0WczIf8wVIO+RYM7MYiAUb+lhiMtdeKLfdtLr8PwV27BTALnue4EMPb6JLxfKiNm
TcOw+93Qse+oIHBkc+km/QpKQ/K6kd72Y8SdxfEU6l1gFxFtyD2QR0qeMu2Sr3gXcV3DA7wXPrp9
+hvn9hw3CAJ8EsQy2zgGb6FAvAJ4vekBHX569p0ObaWUBHy0D4pyRFJ8+H6718d8sV1N1VHJuWB5
iXJcIBz+geyYk7/O5Gtl6Nr08Qba8r0ciX3gMU+FSYhqmfvan22OHQDD2K3TMSvBu0wwDRC8QiV7
1YLJuBJgcZ1yVflTTGJSbNMSxZjZnruAgUWmj/TgK/UlMrmkdXlQZcPPSB3iXr7HNoLor3kzllKv
UCTuOIpoTgj4psNLLb35JKyEGOfHAaGNzvVVDM8N995FbjhXJAa4exxFHFVl/nzfMhaMT/cT4UAA
XITg29YZ69HTTyudq/cx4RhYINGFNAlfjV7mOY7wZ8W78yNFn7abdaQ+CFKtSod81R587oInohE+
pFBsUsLw+AcFF3EncgKHXqwenYQw9/DKr76Wmo73c9d7uWdjJ6LygtxuwaEcMpPxnwNqxGXhiYYN
YrHcEnrc7ZAXPsGPvAVin5jA/PeftmYLr7sS8hwKMY+Xksw4ggHDRZk2wu2z1m09FA2PFbkwZZDG
0x2kTTbxwIGaoBuGr/n7NAunifOaWUKlIdJrLbNxVbyZuLHdkIqAHWFPXYrzrwWC7Jpc3c0sbPAS
IU3hpIoqLp9QJRYJmKe1sLJj7gFaPBss6hSQeZLzHw1Ogz2ON/mmlg8wEH7EzPFg197bRwm7xgqD
idh6bCFIxuKavvVs+LVd6h3Q4KSpWgFwKJ5+3E9o2OVolL+qUUx7xWuoc2s2LK6Rr4sXxazmTy53
9qi6oiWwVcICLr7UKMGkYqbCoOPyYxcpigo5YQWUu6nsAOML8Ghe58u38Bjgn/wx62lJNzLZfmrI
JUReilZJAzKaOktTwE8p4IZ9u3k/bB2xaDa2184sEHjTJZbOMgizGUae63Ingt9wsZfwri+xyPLv
u5vWPOpCUN9V4u+1WrdcZIBa8BnMamRSp7jk4hpqz7HcQ/y1NJXOY8gduSWidTntMS71aqUWDR8G
nUVgHIM95vifQOm+CdPWBkcScUYizOtxr1yabj7XtFxXnNiHEMx2iFyRqZRT8dvpHbbscVblZ4KW
2kT6XH3j7RVrdBrfg40MyPn/tEYJCndoZeOsF4nEIZgQmCosRZMTqwMlRiK4kU0pkVcyY4QUd0mW
pWWKbe8rTwmWWBHUReuM/03KdWi+lccl/nIGK56qPNrJl0Kr/np6Hp03bVCIjxhc28MSUnvCqf+/
en5Ff6hqT0PaXj81pu9/lPdJLn0VDl97QkPrsbB7iOsZ73/60aNJUHk14+dfjxgvZ9ZdHCmeFIPp
tnLcNet6aT5gUxXy5vDFfFZUeSq6ZbD3pL9r9Kv4xNP9DZeNfCtTmTdXzvZZYke0Mvk6LkFBy/zj
HFwXyFZH68Hn9Ih8uIgxQMDRkXFKoxoCJioeUV0oNxdd2IpOa+yRnF04KNPSTpxydT7QoFfvnNGp
bXquJaDDKy0MY1OMw4Ew2GZ0hw8qmZwI3HzuJgQ0VsU+uKVUgseAbpMb8rff1dOzv4gDlB4yaThj
bOOAp78h2T8EiPE58mmZcwgB7afvAixZ2DHTu4A8IZw6w2nlY+FbAsIqbciMk3AmC52CXuSWTd8C
lC7gEoDHCpraFxRcLoqavk2d6DeM3BAGMb2AcFOzZ3gYha4x31Gvw699e9g5xDzYDCBkQPnpmZgI
gmDGrwt9lVbgYcEWyTnvaBI6eKMRyMIESf+2Jo1A/4nGdPbbRyH9ATKH1tTofxPg/ygEF/uiXqqB
aTQMvVNzD9QJFh/GEVmJ0+Y6lfoJPxqLK/qPduq+YmMPSvOOlyY48mmTIJpyuYysUmvy9nX7kih2
ZK9U0wfJSnm0XDKRIe9tttz9vYun0SOrDQo3ae3FEtd9UrzSt2tiDk1u7Y3tQqtSGiZGrYYqA1F/
yrQUGaIKo1ey4eJYGQkrHkAN6Bsaqq8mKT3t0R64KIv3gDNxXpggVJMuQfcp3sGzFajI9lhvzzh9
YsB9cYoswC41JC+aATl8ZJtY7gaKzy6oQaZHcZOLXJNPibkZ7MdyAW6/2ry1MZ1BGG7b2Fs9WTve
c6b1WsSn5n6tZT92S1ecZCU5EDDIHXLS+c4e9WPr+xjELorQ9Oy6nXrMYV0tDCvHCVKVWUBdu6vc
yRdVFL98OAiaGtluF8Wk9eAbESZb5hbY0MH2NRhPRzIILWgzH8PRjdyGZsdgHJto04OoUjLzAJvi
O3dWRWdkzTBG9GCTy2YP8QsvNt1HhUTdRyJ1I2CygmB19WCkDR7mCAn16Kx9P3xaMl/yUaTzpvAk
dp/B539kS4AT8AGzOPtW4+qrTfhAoVHM1fJkMBEltDQhjaFhvLsCpGVPttQkMsTS1nYnXi/pdlDM
Gq0yRtmQYFi+KA5ZqAYSm97ecNaRsvoTzihe7/5zsRny4jgZNezvW/iAYVliDtIEedwZ0pj1CmzL
iVgG6Xh46JiqLXpFN1y50R2PT/eUVHg52VEaSKar+RtSJXTU13lq8NO4e+Ai8i/9a+Pyh63oZEHS
EgiS37MYt66pTPRymcDsgEMPEHRLBnsFmkuVjwfnOhcufD2LDmFZ91Rbqt0UvCvnEIPVEzAWCqyi
SonxFrNaBLyLIQKkoptfpJosrkl4i9C+qRXKbF8rTc6Iaj34SEV2Vc/F+7DAtBkwaORk8Vsrpuul
4JdkiIkmE9FM+7Kh+POPR525sTqPu+rQ4B44WXcbIPOX6YCvX3HNlw2OtRpTUcJeYJnPQyv5Y7Ua
loBc57Yx9VjBjCMrmt87qShHZPFPNWwqIf1noZz/abu0fAY8s0Xkv7lSkhTikYwYgNTOks2RXOgG
znHXz91fDCQXmw1An1G1lCRSUpAb8bu2MjM+B0zt541dUzqfS/dExzdcMt1SQBFd3D8/OFoCoI/j
edLB6LGxxq7dNjSk1SGUI4SVoGfofP9++ps+/FEgDEupjcNGLxAE/BMeg58Prq+X+//zEANhPfIn
M1HMlObqPvl363Xg55r8UWNWWBm8YSxVZagXg0/RG/LlYU4+G7OFqybIRxli8nAvDyBu8mVf0ROB
cRNSlPZiLuTXjxPgmOXI/I5gzIYPE03kQ+nBQYq7+zMVB0FPm80V+iW2DF+1cUb4LgG3VkJxOcnm
BE4jn/81mOgL1iXshZrgZIJkgKpuJNaVKxSI64ysRPhCoH6Kd+8G3aXSEZdYfPKXwabgQYmoJCUJ
gkJsXiXRlHKQxjFmzqP1WYfUTViGLNlzMWX8W7IOHq1KwJsTm7vctUqiN9kTv/hlGpQYL45bHefm
Ua7cz6z7LD1tpx+YqGSv7qaqQxUwgEenyzC3l/tJ5O5wuDoFw+humuXkVPxveDMuhR2gyy92FPXO
MdiYMXJiRddh5j2RJm/W4C+RygRPmwa6+kE25xFKU9Y4ORoaaEmum7+IQEACwzP9D1RxzpfGrDR/
dVp4kha5QpbdM8vDoNRES20RXJofEr6qi5710Ev5uDwT3Rtt5laz53E7wW4IlN2nD/PLxWmn98pF
u7DRlANCB2xkWM03X08MnQuicvdS+uKcz+Ur0mCmMijLjW8z4cSEG8by5IPYakMv3q2b6/oUKzkd
guQ+s9ynOuWpYiNy+DH09yYWYT+NKKi3oADISwj0vt0+A3oI8hcmYTB12FEHc7PJkmTOzQ2YONRX
IgTlThlY+JLDEAztZyCr/d91HXK0y3FvjMX8XoUsYI0TiLeDN+9VDvF5tXml3oiR8RBQPp+bbehK
ksJ4mg9yL0VQc0FyeKIz0aZXquZQkz0jDON34TAdC67xu/1JFP2IpFIsswVaOQ3KSZMHW6UJthVc
YXjXJ8H9mG7aB0QDa/yGW+yQ28w3mNBBxUCzO5u1wcypXPi0yduvxmBmGMTKLqUQL9Rg9/7EHnCM
g07UTcibRLdUmnK+yi8mV1KOSoE6B7ry+mbGkhQVb7qVjx2AyOQ1qJcmJCnX/MdWOAeJ7zb+Q/cM
bQsP363mapmL27oNoFptgf5DTJvQGWqq7hpF6yL6opiDr0Wn+RGwg2zeReSIJyHVskfnJi/HisS/
wKnxVPKPuqeH7HU9/mmI6kOF8bMWJLWhh2TbFdOL29hUoqk7vHHPlePqF+Uajcudb/C9BAEqbzfF
XZfHOr8y7YKVj91Zz4aE2FGR+4g7FJ8V8Ixi6Z9dzKZQnOmbaS+g5SZ+l+g3QhkOPGZ5rRJKq5fM
hQWBWSDLQFZskDZuj2V7oiYd+EX8KkH1KVLbDLftj64fkx2Z+QELME7IDUean+NPu4FgDUbj5sPx
ReI6pnTi3X8vzTp+w7s2H5Xh3rDgRTglQ1mHZw8rSKc5HyggiAP00xBGMj9muf31GEFsj1qtipVM
dxD1P+RnL4o3h7pVym2UupByOWSPF8W0MolZEw26G843pMoeyl8aVNkeKvdmAssMw8NuEJ1yY1pH
XLoaO51xg9axtNyJEtPAxL5crl40ZXiezMGyfJfJseauqIDUeBKYMUAX5bF+Jalq/CCdgNVa4ogm
pGrV8n+QBPIWyWAAABOSLZ0eRZnaz3Fbtovo3VxNSKacB8H137tiu6UZWDPcArRPJ90071o6vvEu
D9cw/+ky4Ks2uh9TBXHOiIvu9cjYhHV9VYCOeeQ2Nae8KjdVNijQyTRq74ho4wodNrR14LMjr++D
aLMTwy2/I7r/iJUvlDwAtWG9ymoZuXBpULFzLzbIcs4H2iUZq5ydLRgeBm5iV3Al3WajYbJJi2rC
crPj/V7h9lIbVWoSEbKBg7PRbM2Ny9xwC/3an2EEkmFfxeHLZJFJkpWs3vACYFq+lCpMuRbSC60K
JLCjr2x9YyNP6Vw3L6kCZimKjifi43sKp5xvRVAuTKQ80i79qGU/oXSeU1LPF8IVMqrV/JeIDqMY
7Cp/jjnZv7cco5i1+AzbS/JrN9s453QJwS6dD6l2KWQfpxVRXrT8AtGENPgvd267pK/4nwJyYRnd
dMVATYmVP6Toje4ib9d7rqitS5vm6M3yay4c19rSXKDhSyMXPGMHn4xsJCtShQiCzIX6//3dyQ8C
57QF49F6KDlDzWesi/ZBeJzi3UOhkIazwyx1FosBOohQ/8WVxzsPNa01Qb6eqUP8qdPCBtiqKvPW
SfWSw9fKhOKlmagPp5SS7YAmpQj2NmQfSo4Zv8/7nCKuskhynBN2CfP18auJq/JwCiccyc0qsRNl
EAqObjvPt7mK7cPdD0HZcy94DKkHCpS7U1r/hdaWp46TbMoR+f6XLPPAAaDvacnJ6Sp4DZ+nu7RJ
HnlKZI/z5SFQPEaTV5wKM2gPvSVs82ljHHQr1p+pCoNgfdCR9prW2NMUbnI8tFbr2krPpvBZpIAN
Ijww2kKIancFroKie0ddlxZORhS3dDm2ppy0BNl3h1G8uhq3lIJr84vKhaM2IGw81phfSgh7Fbh8
a4RRvZWeEWyhoz86hx3iFx6U81Ot7Y/TshryfB6g0wVLW6tBBmyv/FlfPHSQYFF42gxCo6MiYbt5
MCTm/3pV21Lis0oCu1Vm7Qb4q7M0w8+uuqS930FR+uzLxbMMJAQPfIVxFW2u8kl1DzKwumMST+63
ku/zD6KoxvBNq5sxpJnuiMZkYl4V7GMRVEccKGqjkZpnwlxul7tESoRbRf0L+mPGuB/URK92rQRr
WNEScRc2N6DoJqQtLqIbcREGKr3wGBPW1tvvdtqU+BYC+CQ4WiHY4WdBLwWEIb0Odrz1x4yhBa/U
EXP9Icot5Yxbon4KZ/c6Y/QRgp9s+8zvhBfoj3BfJmfveR/UzxNm8ineW4BnF+rXYp5tGiDp/cqX
qVhmSq/N8BrMJxTeUC0Ru7u0dE5uKqe6T60XVK/iNmqktPVkYTJH7wdLL8FYOX9b8Cfh+J1NrCuX
8f008np2IHEVfksrOuwc5HiIaUgwSJbk847b/F1sVuX00KRVqk5t9/Mz3fPySOsjhOrdH2DMQ9Kb
WSB58HR7G1JO0dK3zIT26g2gxoXHWcV6iUVwm8GSiEQECOKu7TjxHqqFRaqJtpMCGORI5Kq1l+OL
NuPIT9cqbLsOxzc+nAjYgXLdGwae+YFXi/+VAwrCdfKayFhMWE1mpe0GL1hVo2b8EIzNUdX3flP2
v0LCPZS8YTnunMR555EjGrSi/D5Ek0BvhIZzkajtxbUj6Vp89rRHiu4pHT0qwXPh3ZR7D0+hMkmn
7R79gdNVqW4ziDm6LRAy1F+urwVGefgXIti41s9QQMbNtirYKC5tSwv5Rah4016A3Sdigw0boN2i
SAHwDCWQo4RG9LWV4Qtwj7VYHQXMoSjnnavfD19LQa/yPsSqU7pl6KBXO73i6wtNOsd9qT6awwK+
3rgQtON93VTIFgJP4rwaF1muhnfjYIKyyQKK+eoqG2wRdeLOxrvR9oWjtROtGAikfunb7iWy6P9f
d0F2C9Z8coQlJL6lNZXWHLSINQofWnVL20siCGV+ID6KZZz5jEp5IHrg6LhQmqeCaYmWDmDayNeu
NqbGDRPBciSMhLhO96RWnO0PHcLRihZ/Aq33iMK13KFlriF4n/qjAOy6D12IaXlSMjzYzDBLFk++
GifhblkMNfcaublBNDJWvFjk/XWh184bGaK1j0nahvNL9z9Gc6mXlxW3jQppFX8fRcBNLBoXl006
OmV/W/LCJHll82/K77ZMXAQZ+xDBUNcI6jZB+16u8wLiI7cDFbXkTTqujmInZk1Qq6hbMM0qUJrv
CKqIIHiHJaH1G8XJMLJMpGuAu+soJi11uFokDyFNjIVH6BnSo5pgDzgnywsGWxjR+1iyoUrGNw9+
cXkkLTL0rxpTRhPzBcQO0iAyiNi/Hlymuk8DA3AZTZnGcBQys0sCBfDpcsh83+QpXWzxq20W4ZVB
Cv0UzuYirM4dI+8kkSFTKQaM+ED72xvbSXLEAJtnx62Q4FNh253Sj74PZoOHjc4nQNOnYEYlXp72
2I1E3FadxWsVlEx6Nz6QhqrLmzAPR+gZUUTbEPFqdG0XnTyM7c9sKnsgc294OEDpdLRRH+dLHh/h
jCzvilPpr40ZR24EgSCRDKHhjBPZLrXHGr70FiHfu+4nu1fU+1ADYqkbu+GY36Fvi0V8C1SPNAQE
X4DYIoDKoS6cCu3uIU1IdSIR5FSrpxQ8kDvlv5K12IHlXTTUjuaJr5ryHtjnfMPbnOfn0Kcp4ERO
5uDumeAurROrqbmRHiwK+//RS3iyD5UXs/6jkXaFVHuH6JxglxBvT6YscB8+qxoFTPmvjwTxPuzE
Lyy2lZrJImF8uptljOO2UA7kr3xkaotoCjPExKhYcCKqa6HRAdhQyoyvM4QbgdwOJ4T1F6NxJrO5
Ufd61MjtPrWGXk9RAOZPeqLL0BmXhw50f4QYr982kQWxDMxXDxlEbgNGWU4tTU2EVDuH/uaLm9aM
WFTaKF976ab1TYp6li3h2jh/eAT4qiRKG82deHLijBa0f/1KVKRfZ+GsXUcMmlNycZPgafhMQH40
xp/dsC1Iv0LiQ7MAMU2fiMJl+euhgrG+ECLh4Ak/meZZmhnhfA3/W75XSP/DkYQ+9UWny/3jNgr3
Di7vDSyWBw70uNeqUTKLdgqJYfoTMEYxp5pF64GCjNiP13GvfrrsPEWia+B2PGb08BAyDUiSvUgb
RlQHtz9ZZCpkSsjLVRKyM5jxBEfm6IP7rFZ7MD0pXSVWl3klILb4cKoVkfjGXT1CklG74XuJ9EwB
SM2oM5RrB0D3T3P+Q6w87UtDhX/WxHnDgcJhqzlhsCLP8VYCY4jtm42sgSpq3CGS4/eycVt+w46s
eY8C+2WBL0CgzugnoplVnnSCG1Nh7SRyiqlPxOuPjVMduL0MD0klGmozyA7dAFKnxAmIn+miNtSa
/0ZdfqQllUQs1brRCphRPuWj5rwRWPH7zF6/TQp9Z/8J5cbk7uR9M2VTY4lGQ0wGPAjaQpOcc6XT
ciD+nU9YfQvTgi4j3gDGwuamFW61ZDD27BPn6S/xFMsVmdJkpj613jiTdE040FkJotlfeHx5N0JC
oBE3vPSXOrihfxNYdOhLOysK9fByNjY5i15PUTQPjUipezEZFF+whN+TpFAvGHsqh2XBPpg5yItp
CpoHrv9Vqx86EbX7ttV2KCOw22vxW/OFBfA2624yBQqDfsp4ggzAkD/L0S3YdIyLjDfCtsB3bOhT
ztJMsDJ2xisDHdQ8nCOlV3nrnndwj37HOatLaHnoMK5GEQcwD9TIo80iIrrNN88A5gnA+1xTZZfQ
inyxrzRPaCCpjQfXiRP0UJLEkHcq7cBFGnuWx/oG8blnCvUiDjuVq91uc0ujcvIkWNFT5CNTaWih
jQaE22eOlJyHvyAlan1NWVqyfWtmSeYOWadI5AkrSgnSAewax1iMKodRYuKm97MC0UiMQhGDi2Oj
PyGOdvr0/0I5J9iTEUYdOa99TGEKaxhw33ztbOQfCGE/ocwTJh/lNvVCTyjE33PS5EhgibKsgG0n
CGFVaa2yuVU46WAp30pW+ABCm5aoyBWfag0/GjpEKz6ZNvdeJpQ3WTS7ut8k+1FU1w3pgr1M2/E+
v26OxMzYcnZVY2p24sZPQsSfKZyK64MUQKQB4TJ81B8C3MgfEEMbZR3HFYYfS+3WGxFL/clCTXbm
dlZCYOxAm2HQb0TYQStv6iC9CSr8kDQxJChLS/OGBG6rURcvi1NIUlgeyP1HnrDb874qmbhRo1PY
YoFFO26+kI/ZBs4AidY2Ylhq+YAKYW4v8Y8lIJhOrla2iX6Jgq65KUmxC8lKEACn53gy5n8F2rxT
aCBhc/Ne2NVBeKB864EM3pyYdNtcVsTnZMEspGjhw0yTipLNOfx30gNrx4M3tLX0J8Bkx2/2bxQ7
fmOkMNxmdEwzauWAkOh0As2lwm1kXFwKE8ztrg9xPAODM+5C2bu1+1/uJxLBxy036L+b+VaQOYCj
Nmu0O9h7oHBpeGx3BsI9c3vYFy+qPJ5tEYXosG8pjcxsTdQPJZjtWxSp4YNfQ+hN2tH6iMdw9zfS
YPRn1BXKe3eEmq4T0HNQGqHZ6MwgxFOc0UBjpq8TOB85ygpidjn0FaPABGZ9eUmbFGvsFgMrhEte
X0EgCVexT6kJNLvSZRGPIdweknQXoEm/SN6WSBTFlz0uNzoBj5HSuCtXnKi+oMjv5drQte2krLdT
QWS1vsLDVtWrHAp0+lhfwTz7NuVe3+mt85uKlzbgemBXx+59ifFItRMvSenUgjF5P+ENSCQXv7iq
Ws8RbtW3vJuusRBg0oE9ZDy2MiBIXyJ5THh//wlDXvdXyo2gpRTenFUHcN1mR3qyJ8Qa9k1ZoUy1
0dfp0DK8f0DFib598c/dCjm+P7DdjLDBzWAUSaBO/m1PeXIWluxW0+XqktDgBVCN2eHxcRYf6o7s
uXtBYz4QLrH2HxfCjCXttaHGPbyT9YrdW87+cIpeSwziwnqFusSP+rCht5/QbSNZ/7YTTrx+KfDk
5/QwqDaD/h+S+PNTQcbxjI9kdVPd7wQafEdHK0ATdrWhAMIriAAZIIa7ouTEV/uMxXG6UITgDS+q
yB4Rg2Y1ZUxeVmxg0I8yopFSkEBP2zRBKVuhQQ1o+woCb4J7SPcEEaQKGhxoV+pmPy3i/Jp7QNqM
licl+7XvkfENLeIru+Epu6gAR7hud7aRKYa0/wrjZAYAlunVtk0kcD2y9eyu2UmWYwfBHaN5WpNX
4Xhu+aT4i/2VWWxnHPSSyxCaCIeu0LiSLunzzDMQmumJ88kWZWBdyWXGrzNNYHDGBJrmaC2JwhMM
tjKwiMNZoKDlBTjwWk488Dk4KA+gq1MwWiaAtSNu5mq897RyS0gF3o17LEu6q91ALcjPI5+kIJPs
5AKA86t+LiHo/NZPm5rdgx93Uu9ZSlPPsFH2P15CrKAXiVy/1kO+L565EUTAtwhwHA7w8TV4gzet
rcabveS2ZOF8w95hOHppVNcYpXYSkpMRklKqRhFdqDBcyAC23x316o1XCTZ+Q5VxYzUyf2IF7Boe
iYu30emmBPGtvPLV3Sj585USTVq82OjmkF8iC1AvlX6ZJRylK4cjTTFejZ5/BvkpYX2T9+53meQ7
Gi640A5dC6G0r6c3wZcu3HO1yRmTdcZlsN26+aYDVKh9ekd75HnuPj141ryiVniP5pdttJQuOWBW
cxpAL0/097pOFI/uySlMbNGKujbhIFx7W0CvKLg7Af2GYrLmz5RUrAzOQ2va5oON+9weTzaYmjN6
f+MfgQHkjHXZeBs9/n72o0HVENMeBnu+dmOS1hu3AbqzHVGRHLFvUSasIM/FX4WAr5SFrvUiR7u+
ZBBxSNSHPF4Z4uycnGBHEzjoAqdCiZwD9jNIfHZRP1gv6vJIL7woyDOMs/jMcsZtuf1Fsc0JcA/3
iFcfeNYR2Sm/8yHZ0BJ1VIsVR2rxANSJdpKJKet/09NoidpJ74a7CJFnNh34lz+QIEj92wbFOzjf
puGJZzKZrQZipWMBNw+GF01vbvj0fGVx03QWiypqv/5UzN47JW02iln8UhrOeUlh26zOpV5OZzXe
64rwNcTbhibZB6+kIClADNnLYX7Wcwk/8vXxWeMrGzw1mtEoq1u/UimXvF9zTx56nJVJtzCNsNOS
t5NJTFilLjFWulNAJuUoPEMnjBY2icOm7XIWn5waWIVjOYkml+FnEOdb+u5UsCiEj8nEgP5xqYka
pzkM9GuUYJSj6WWlujYKxGMBNHairgWAf3dZXXr5sbUScVXQ+0hEdSQYRIqPRb1D0r//7DqeI636
wQ9aKDOy0FTWDfxr/GjZkvI9yNl/ryhIBMDh8YbXWnLhZQPXbCOpoX+QtGgBKI2NXGn38L64F4g2
rfQc/ybtfEvD3vsDCsYYVgwP74xIKEVPNg5iQ5w5cWTt3T4db1joujHsFU1P8uUetb0lXHC7VC2Y
upv1l3EuyB942bvMrlmeNjQsZSVKTq4LngdvtvOI8ZIMEFIHZ+w5erVCzg609F+FljpiWYpc181K
gwopGC7/IIoi5lG+6y99qKrDYkmqvTP9vWu6ED+DmxGkYvbS+2RWsctvEMCAOAYBaOzYMlnUBRHJ
IL7oydAkiq2rdDhkBZ9OrxhgXUMh/jI1A+FOB1KQjlC1rU6MMp65vDkfaq+rmVd7VeGWt7sp9dvz
Z6m7NoDdgWD4ZlOFFD4qaMKcmrkCSrXnVrquY4cMkdGM0BaxMJ9viKdzU9Wxpz3CpbvV1JtUTjgM
kpYTjo+IJ/f1C/lIeBnZWzb/gfZe04kM3kifT06l5tWZqyy2zz9tZ792hPLpdELamVqSc0kgxqso
TBRmOi1zcQ9txhqkd5RdNKoSnC4Ads4tMQaPdfEOuhl7QWGWIpwxmCj7mP8DYt7rjUUjbuYCHZYB
6Ajymx84JUFdB9V5bFoUy2yyPHAXgEsJ2MfXv0JcrosjAzBmKKjA1f2iPelgNgRLwKB0KMvp3LBp
MRPTCPX9hQN6LvkmmSDpzhOqnGO8/5dH7UpGtlp8tROUtVhMfHr6JJq9+xa0Xbr2l7x96MgGwzGE
wlXRvEnWT9U9O9qYf05qfMC8ofJTFxKPKsosmYFQL3jMUAMC594kn9qo0pn4HxcNZMM1aL28kpR1
ztUYQ6zxX7QdplK9wGjpnwlncpICOdutI6mt/lMHZW+qbhztOSDyu9f9DZIDPkr/mhIxbVxv3/MZ
HVovgFiCDBmIeI/wqJyV0RFlxeAXYcYASUWXYRzYtYBqb8YqCEKDEaPkimow+u1+yeOuMzzDLg3A
iW3AyXvGySanPtJ/cP3bHQKzq4z34bBfloNYAP/Di70oaOYvWcNJ9hxMR9t35yStaM0QVPgfF1G2
ql96ULjnhAT5eWFRjXeb8UHAljqyUZX1hVisa7hZIxsLlj2i687XG8KIQ5M7SP5lw4i8HmfECsQK
1cScOjj7aPMf4FJPSx7hQpkShlpQ43zLkdV2cec+f9PuuDnJuyGZrzQY33RdONDoMLSl5/AxA9jX
QI1hQVqf4HhcvPkgwAT++hrXFy/o2tjW/bc5AkpGrUPWWTc1aqK5/+rD6nLsjWh3sBw3SQVhy710
sDs2eOKZfgKNFAS6xMjOisde2jU/fGXSxRDWsxRmB6jIxQSkwfD8RtSyMWW/fCY3DD1A3MVFcXRu
E6baJYFY4V1DGDe92did9xhdv5Mt11axjWyAg3Vwkm1LTvWiQ81YrKUbzwILImYuXIIZLRru+Bzx
PpPQwwwCiskXQTuZaKMkXI3GqQNftItXmCIMaE7hHVPPB31CPUYWWkZ6YAEMQv9wmVXbsGTrOu/q
giEiNlm02Ny2Jdz2kWoBQ5XbMExNlsbVh93e+HalPhnsT+PR83QD6y8n/hwOpmf9zBmNVXjKSM9u
gDu4oBoN4LgamDGyG4Pe282eqoE3anpkaTBLevvrjm9oxqfcx27Uw5teFhri09b20HJrptIHybAZ
/mXSJHXAnuL5buvwcmwZDqLFHCEFyzq+e/92N+Ix+KkwA4mg6TFZH4g3AdCxxYLuIo88MIRTDkPr
OYa/k9EokJ0FVPNWSJGfVbeqGhgTg+yiENrppwr3O9EQvNa4hImfKFn0lKTePDKoL65rxjcriVOQ
xSMsQfaQflUwAkRnOqHMxMkccQXpsku7KM08/jDZ6cz74Na7f0n9xTmx+doHHHa2DFHJ3xIJwQAM
pVQ7hMnOs2C0MGZGW7zsWp0hCxbRG2AkdTg6i0ml6U3qPNkdpTYQMNPhJrMvhnH3n50GkrS2jtFF
07VBrKvgonGaDsLYmZ40dUCe6OusR4LVjqIRBGi9EGZiGBR+COl4PuXcGrTbfjHkiigc8kQ01+B+
B72eVGrIbGCFD/JiCB8IX1TEg1W6ZVcQLFpjiUihg8cBkCY+MJ38zovE39o59fgZWCpyd5d++wTl
I/e4KpY1GAUmVR9KwV6ElRQJtSd3Um083V/JBVmwQ8KJJpV6sMykkm5zT4z0wf+EhgD1A3diQS1D
day8Mvkegcv6LGrB4xRtupaPECeHSV8uLJGy86t9z3CWX1z9wmEWCAM6bAk98rQh0a5yViqtlJRv
xHhT04SjZx7LW4Q4szeVPm/Ft265LQTf/2H+tBT240lrryhP6NJYDJj8xJ1ykZscWzGg6fgOvCXZ
QFovj68USbuVelqte+j/njTZtzjj6IIu8ns0uE5FflY4Ln2W3YLmDatL7AqpDcVr2aXBagHaMPBV
V4WLxDQU8D74YjuUF5v7hUZMaibQWx1pe6KW0O2wn9eeqaGyYSKjzQq9JwerIqfrCebOBQlkIUD9
luwXIxmoRQd4414E5itL/xqhFezwklA5CIsb5SZ1ElsWboc0u+H3nUhD72zQn3kBZGIZUZoyWFzQ
R9fhQn3IufWXOGIG3VyKbuD5IF8bGoKwLlIGBmjk8X8RKN8H+WL2QTX3vkNMKbiF5jprPzrtHcr3
Itz87B5pHGlz/G8/inNxE8XITpccIOrlpVIGxbC91ZLN0TA4seOAmGCWDfYXQeCiMmuehYwCEgSA
arzm1C+33z3Vr12glpBQ3q/bJ2f+czEyqOi3hvMGBQBZGhWhwWTG1EpEJ3zIFBpopIgzEXU+NyJ5
9tq2TLi86oesULNyvzmDxRN0iCDuHrndHt/+oh7Pt+bbLGve3NSkTAUB2jcmQYYQItUIhE21UA40
/2pF5kibONRG3KFgfix7wfAvoZ92A86wAEOy9vnke/5Q0nuV+Sdnx/2MaO7YYqoR5dF4s2mS0hDs
k3P6wCbDDqY5pZwIHZBkZqQ5p13XtF2JhtnaaZTQKamHn1Ew9aOAWO+MgBqYncInG9ahYSlonSA+
CNV9UZ4/whi2fs/oaxHXdJbGd9+hok28j7MmBPvsFa6p6zjiinSpItu0gFdQ3LoOs2Lpd5lTCNEw
OqL4iAUxl11cBwcq+iTcsKeYghaX2zZHogKb3VXs+9nQiEIjGLCIG6NVuGWVF//hSa6S8AtWX1Aj
L3z3CPKJ+CeGsvGQ1O4Rhgb70/PQuK5TuLABVndTfBwmoRaUYzDSQnBSYGSSJz9qCg9J6wVHSnXb
s6Epc9msANRsi8NijlWZXSexaPqGL8KCCGlFpMhEF2ecKAT34l8MBZTkU5CB/c+ROsJvOT7yk+ol
pGZQWAykC/Mtec5JjZC1TA9I05lYWcYluJGEKGlWxzvAtmuCTQq8cNvlgOu/0Bzlb3n7Ih4wEPRz
fVGZS7NedqagIl6wzCvSD19GVxNiXA+C+eAdbQY1Y2u2xGEY7KUKcnZsgoCZyTs5iSRCfMNzaIgw
nD28r2gj5cGfKtdLQSNc+Gls3u3Qm2RyLyWlDd+W1zLBIYRlQbzb+WI37efx7+f1WOGLabxCqheu
y/PFH55AdmWnVjWH77p9oetmXEY8TlcA4Q3ZbB0L5u9E8hxx5s/6hUbKM9NDCCBhoTJvw6Z7yXcD
TCpRU7uI0nxOS1zZGJkgY+Ufk/yv4xJqOPybvpvS2xGxnMxMqZNgWYqRn/1dnCIf5LCt+Wd3L/x1
ecW75CPEdeIIeAkaMgOzuz9h58ASmB8IhQgHDOpfU749lK18lAF6/uCQ6EZIqWpXcNaRy5ssV0Ro
iBmrWJ41NPwzIc4BBlp1dDede3dLHDGY75RqtsSDToWQq5+QqItBWbHR6ilehbKzc5W3OAxJAG94
2jXdZkI5bKrkLDtUx8lzR+X2IkQtJ08FuAVkSyHBIDsbuXwXZiAiGYyOKVxDDCmUSGGWskZd/eDu
/C8J3U+f6914qWcjQP0QQ7k/qXGPvbQxGfPGkP2w0EpuKLnC1+MEAxzDbMhnYZDS3AjgjO5z/CG8
ZkyF9PUzKlBVkiOBFN5dkaphOjt6aAgO+ku8Jwiy89gonp6RoENzt4z909lbFJb9mLBA4XpyhO6A
tV0W9hI6CnV+Zl+X1n2BOuTHH5AftRaSGnWVVYTAmay2PPyqvtzkkWtoG4Ad+JtqU3E7hEikoKJi
DjHOvuN5OUffsokxv2UXOLWxuPs0NFFmMzRm1F8+OuOizJ5x9bgK5XIIzUJ8dC0EBOR7g/SMAnQQ
lTAuG/55DLSqvG6q28gnYXZL3PLmv6xy1XnzV18MRBb4v6z+euClu9Rt3FW181IRRCOcC92aAOWB
KUwOCxef4PcEuFc5qn6PvrqseRcdAmSJJVyKj0wdnLvA9PJmpsS09Z3pgKz0mZIt/y+H1mIOZQ5D
zi5vtzgNZeuiwb4/oh6izc+GsIwEHM/BdMFP4TZlFn+52vN0nxWV0E1mh52WClyeivToKiX7GyCZ
0gkdHuz4ZJ3Ch5ahpwrDwrm7zAklc6Ii60Zwx04rbXf0iTuRLlm3aaq+PEPQ9GZ2hG7vcBz24miL
SCxTjOVXHaNPnAJx1cg6CgMzDRBTZSDyorMYvqBDowEH0ZL2hyCMOVZ23nXeBgv+X10C6BvQrGbJ
79cYTs4fsglzpJxs7IgMNOyR4VPARBne6aHcMds3SESiwktvtwxYcUcrHopT8IXjIVqkUc2QzQUD
PvPx0CrkbVX6XN6/N8rWJuKncXKxPD6H4UdOIf0zjMlVjJ203vYI0nU5Ehz6MbJsGx2ZOgyXyVMc
DN7VkfZbo7zyb3s1ZfALkU/CrCQmYxdQpbIYoVThBWk9zFKRCSU2/CCZMgfK7VQRO0E/lUfm5epL
G8crARJKDscEUDhFnStOJx4pDzjrBkjiDwvLB/Qsi+7kWYF0Hv1LrfSCp9IyKA6DE/CAC2O+ex6Q
rRXZEXkKEROJTo/f5LWP1llQ9KXd2EUJcgxGcZJ4wEEh38wopXfWLc7c7En5y4twpAcb44wEYGaN
X4VrG+wWOzJ1D5DdvbqqDSfJTQvsEixNgA73wYAzNCJtgJDbS0rINoedd843w0iJ81/QsgCw9LXP
6Hokx7n0BkVJiqU/+Bv/p/ZuNUolIHNCeCVWqisbVC9qmb9KB4zpu4bECtrwY6MAehzFSkqK2PIk
Ek+AUq8P3/UXg5C8MoWUZc+P7NFx9IhbM3to68E+BUVlB/EGT5JEubz1KPkc1m70QFC03qeNPxjk
2LwcBEgg3U0DRIPLei41XOIjWpPx3aPx/RUaRYUrmFGveGICQ47p65bNcmH04TIjAF9srKcXuXho
bSzTEViU/Pxw6vBP3kXqU2LjN2sVaHeMf3y5w11XGX6s+aL8eEf2nZpSr5lYFzPf7QPJ6kFlKYgl
88GCYzHOd25a2a2PG8CSJHvSiXQJmT9aLelCPXWdGAtD7H5f1WLXDYywT/OY2pV7axltRsuMbhj0
SlFsAGzDBIEgcCb31Ib3Pwxhl6OTe3D+aVfZnT7wkvD5W5w7yEuI9oD2eGALM4w3j8AMMQ4SvO9w
axYWxi2uko4OjzpARszhJrZexnXtwqjmJswwJKvL8e9427DgzCx0Tc8z8Q0ZQrFameczcmxobXzO
ikJQ/7YCHUEEAGu1n9PQzCTFxAuej2aoXLmOiJPGCCfSwtHe2arlXU1UdkkEfv9/9rMt3i8YMSyG
a1uwr4Vzvo92E26IsZhofqPHMN8AXBhpuhPR31V/VR6LsX37gHyEuRqfTEctSvW4RIGsc7jhHlPd
Q2c5gxoqupklfwtoSgU8vl3d00YPhWc+CCTojtxeKGT5LRmfuNSutcjfWzqUbSlzZukudpWkMzMn
Q2hVmvKsr7DKw3iHdreF6uj+jZoDKNXC+xnORvL4jGqdWHI3JeVWtLgUzSWftvajt5x6tWGWOxb3
CGEcmWk/YxDw/M6o9thyHeeEl/xldNvlM7vaKGLMgUe2Z2EFbJAHH9LNxpemXbGPIqmTZAnDohcE
HeBZRCPoqq22MAXmZqLnoceknr9idFqncd8isLRDFQ0VLE9PaaCqGtSMOOpvLH3fVyAnhAj6vDT4
87efv3ax0i/bRtQpdla2MHY7z+/B9rSE3WN3pB61QRTRKl65hNDjjhe7R0RoXha1pkbSNaD9AK3u
H64UXiss3xm9h5Nl3Rx9KzYuR3Cl7AUG/5pqRGtMxeSnXbrlllfB8s+Xf7gYunfSPD8iYhMm15+M
bwGw9P1DsDLkU8LxdQtX3wsdUT10R5F2BK+WDZOX84SWIyxcMIl731JeU6nX4CGMAkVMe3gFkmCH
l4gWGsGZnNXYCB+FfjmGBXB+lYSIhuiGPiCjQahzRsBIRSwlhVjDHYFpgtF15Gbbm4P/xBpdYuqx
ru2C2ZrPWJzFB8Kyq88mSPBlxZNEtByRgX2hs1rtnrGgZPMncRmKJwpq29wfbnDzn4LXX84w6tzy
OuAdLQnUMqqo2en0eOV+FZsEsiD7uXIBqRSdkPs43NYEQ3BRPv0Q6b950ZgK/8vaskyI+sQXVO7C
bfomf5bY4uqx3+QtnfIFs8S/BzEzjSWwxXSxe7OhgYyZDpWBiMRH8/ST23ls5neWeK1p8lXCJFwC
pChwUSs98HMPgA3oJrBviSHlV/kSr067F1pjlxuApNqQJPR/fJ2V0e00rkXUUWvU14MTwjblA91k
O/7/g3OBpedhjxYjgw8pgjzMd6VdvWOb2LT+N/sQnUA6eHusmUI37OMzLeM/KvqM25HRKpAAcxpE
BAuoHOlAon8PRVkhcFiUKjt9AcK9eEKRRL93y2FJGzFgwA3hjqPK+6SMCGOb44rKm2WaAorolMGl
r6ClfEAQ8Yhz25bEMmeUhmnfds07Ag9V2hhuuvlAC1IpjAc35Wgs0MUp9jpkP63Fnc+oBftL902D
iKlqfb+FC78QTFzPp0+ZV4UcTgqv1NmNsCGtt0ZvJbzxX8YO0TcVNXhrafazfnRzvZO/9poGMBo0
/spWzVgJP9EWC4dVusftDVjRMER8kH+SlBPS+C0SRggl1fpRTyQ4ke63n54mkZQ+LhtgAozlxXsO
ddIsTpltccUsFPGODtuYnbkMiwaiZtEvJLfUHPYHgvhr8ELRftx2zKWWlgzxHVruXsfOE6E6TuTj
lPsRPrFG2CCLCfWBNpt0+V1On/e9pODCoCBuoIOBfqBBSbYtyq43GlOelc2+qtZ1jylaoD3xhm19
mlFNcCAH/W8F8CpJePfK3jMXoiqrAY9bnCwVGdjPJoZgpSaR1djRB0r56XsVIobpQhqcuQJZmrJg
pcTv3mXUuxeYiBEXPCdkwqcVI/RIwIv8eb6VahYzr6yPYo0TyiTGVPEuTWf9MYecByRzSawT0qVw
HqcH2jqNHDCR6SS95CewCoR93BsRPnNElAu1EgPD+wV4jrSK76NLUMMixOjQ1vn6ZcgB2Lk4T085
qEF66E9zxJA9PoU/+wG92411vHKMHD57wHpL1IzDInuErL85RrHuf9oEuBRmUnum19quA3NRFWM1
E7b0d5R+vXdV8OicUPq6dbjGu9WUWGsLpWaczZkNSCSwCCL1gxI20iQVrxot+ldKtW3XDpSpWDTw
jes94ZSE0vASr4047wwjwL0KpgleET6eCs/1zuCKRaTfq+xOBBAJs6m7va1mp5A1SDEQu9d5a8id
TLz70W3FcFleEPFjRK0ocZzHV2ORXmK5MwINecD9o00NI4RG+pPIi+B+p27y2uiAUHDJbQhGNioB
JbVRBN2GAXLmVFaPVB4anLyxsQfn0BF4DL8Orm4vcKISRqE7gpc4EdKuBu+9vGsACph+AsbVISTV
X4liQdhiRHdj5ALeJnYX+uNTv4XNBfGwUMIv6Tv0GcaL1+EzX4da8NpsgztdPAc9XwSauZuhYBPJ
7vgnZVZJ3Xjh+T/y6jcvON3/GqL1JvpTqsVeZjXFBf3li+TvnU/EtQ6JNzks0uS1qT3NMaFpgzJs
2aWiqorLXqXNmA3uZe+uW3yIsEpF/3GlvJsa8SttsBLAqQYUAhu2RE1zjV9OxdXQeuG+3MwJphtC
IxkcrhHKjHFE2E38ARKDiay0vzB00DzRiNNQss5ol+08nIrTYkGkl5x1I86y9NVSPyJrc2O7bdIR
MrEreJQmu2OAXs7xcz4z5BndlIm4nXwduS9rrwNrUyJUcoK3rfSo0YvQWHadDBrO3/6t1i4xbfQq
La1chybD/BU1wyqBgyzdgrefeocfAmr9jR41GVC71uKtNaDavDohDxWPvFE2eXga9dMWL/TxJu5v
dPhe0VusKYGP0PpL+dcT2hxD5xkTlEv+3EuIYX+u53pNSDyTnQ5AQeuOUUBI+92jKM3MAOx62Jtb
FzStjjSr1yU33vLWV4vQTsg80Z2pvGfbdpnXBreA8i1dlUFgRxFO3sgtlgOFbLDMcpktNVhS3kHz
KxZdcmJSL0oxUYv5vT2S1lwF99NtG5+zlDBCM0uNVmUx/3GuILfBVPjlRAcK+PHnaJp2pDTMDyf8
GVmgieRXOVGJTTRndmwvQ7aMP3bMI+facT+VKEiWyw0Mcq/vX0GBDqlY+TLlA2MOM8hZfQUuhA5u
HCpa7IoxgM3y8da2Rqr7o81AgCNVkr7bqjlPL5AHuoNc9Fu/hf3OI9gBpfv5tbZ4y4/b7HIa3Y/V
xQhLMummKgCzFnHCCHatQkHL4pDu7qc/HDIJgY3qZ6P1Lyxh++c37qh90iI1N0TJTagRwX4YDRam
8JsCq+F/povvHJuzPcuwwDEO8gPE4bxA0i4bbuYNUzIOVmzbOKV/XvdmwsVGDNZ8CghWigDkXU3g
ct7FIgSRV+5UymmmkNM79piWIUTYd++UaO9zcT2ZBnrOvirSgNvSwxwsyYfbs4LUNAG5MhAACE8i
1DlvguK7AAZJkJmb22uh9aYbsRDWW7EkqC2IYXcBIqtFTHW6byXKW2mf8U3ymCteUipjRo0njxWe
EaTuoP+pwp0cqeI7XBAFiT/rLJK1oYpr04fDI9OxmIx80z/V3mJvIDHHM+HbtS/p8rWzxL2bnCb8
7s2UzbAOln0bYd4CbBzy26zqG+BsBigCtidf2ikyan6B3vq3fSldhb2CNn7DBCud76bhs7EnkZu/
FbO927zL2bhZZy3EAwUWFgLDnfeWGws03MFpTi6m90WSDEC1/bzrAUl4FDg/F7xTLCjOYtamjnRH
cGW50CmIK/jXHTsxFL5KTtwvT5JNDvrXW0+sDql1UeNcyHPpIc+EgCmLd0hpQ4vzYKeZtDWqM6/+
W8vj0H8oBA15eI9aTJZZEMuxko0wRpnRzCNrmMwWmTmVWD006HKmQIPUZ49gZd5jFnsCG13YIwcV
243WUw2nttoFC9dLzN1tjGm0R4A8Ifn/yzknKBK3UM8ViwkTFxkvPdmjeCwh+5UYugFgUtQUNKys
zWeeQanKXGNud9kIWWKUFMvwds8K/hVUHdVfy4wW5kNiAkqhvmkPPghdkLlU36t0PI3CisuzCUDY
f7D3oWDhcuuRmSOCIEDDt0O/hPrnI96owTNAwXUbJwf3E+dKsln9ZeaMAKJur61MvoP9SFWhbBOG
zeRV0Va4U9eR6VCAOXjDiLrHNVDD5c/nFP0uuuMEth0YSeNAddUpxFOiipoapxCGeAqLGd5bBqQ/
o+WkyJ5Qo59PiPA0xeIfGkkT0W5FXaMkjHPVZWeOU+HNwyn6djUIlFmUe/cJy2I84E85heaRGyBh
dEVdvEFufjjflRQaxrCdl/EfWL+rnpG7nUomNEx97FZm9ERcRuVqETPVWkN2EijgAUNGqtAhV+vm
UkbOa9hX6m7tG11/mYErqrrt2MzgLLU6YA58GyNg6BYxqOby4E295IHmFTybzoc0yhAOW9jJAHwb
XuNWUoyBYMDyyphoXCtkENIAdE2gHhHUe6emlka5lBsGmwCysLQOuIvEJp01T5Ory5rz3vcg/UJK
sDqQiZCTueCG/alroosQsJ6aT5kxO1//BBaG59LpZK0uBD9Rspuc0aQQkGyPT2nCAIRgt8US/UKG
myP4IShr7JCR9G+AdsGyJawcYWt+fhMHzTfKdo7+hPm51cLjvaBe2TL9ENmV9qKTWTZpeEl4lt02
1YBGhNZf6eUIibS+slpGKZoOGbuRJ93S93SB1pF5ZpM8BQyvLfZi81xyNXbLSFleAN2wGJy1xXAA
gZh8nng3vLSRETUOaAgrC3UHzZ8UY14uRbITGTdBwkatw5/1A8k1K9eKcXr1Ia7IvYhKg8KdvD8Z
YhsLPgc1PoNZT7FJ7z8TSQtphRnqHkZgwpbdzwK+cPLh+dzf/LFGhUZyhZM3JnlXfbIUpj931Dnh
FcLkH5DOhlEgxe/Z3YQVnYCtxr+GXqm6vlWjD/75mFhCJoIBSbmtx8e+0C1iB8cBOnxTsfbMm+Fw
3BvPDbONcYJYNyKjUAKLVdXEYnTPn53YqetENzrCwTjcb2DlYKjcLBv509NviRrMnXMiCG7F/aMV
J+aqMW5UqKXXUJ3b1EL6EwUMna0NxTe1RBac3vRTAK1u07MksED3oBqcOmi0NlOyvAvtsVKEoe4G
xFEj7xJ8XwyxsIaHZE9C8Z6SJb1HM4wJlg0SATsmC6HWJg1kv2J8gIF5Z0fvGPK/K/Zt2nDNztDJ
I3hymkKd0isCfngdvNmUjqhGQ1NqskMdNA2O8WnqUe0+sd43sIH3R8vZX5rcRXFXZtFYc6TVt0aA
KWzyMA3+2E9nJ3RFnZLpot62TYpzEVv1I+JuIOXx69dTalc3zRCDKx9gWQNb6MvtetllSDPDcXTG
2yKbDIdfZKEnqbtsXdl79wF6Rs83Rz2H0ItnwzqbBJAJCMs5TNS+bmQwT+oVJ8DEynWFBwMx67H9
WZMSfBDpeBl63NPvnxZ7+pfA5+YgznpQrSh+w85fdUhdUnjgUAWBrSjUA6RDpxDxEtlTf02E/EdL
P8GIxvx6ozw0ito0TXeoJsx7Og1WWCL1+ogKbdE/ZvfE+SzNMhpYWSBlQ31UZ89xVcKBEHRsSOO5
yrszABugIWluv2/mhaEBkOaTkTQiJEff81C8F9xhLgjT81oCiMEw6SAfC6ztXoVYHHfl7pgJq7Ct
g3i0ZdivghCfTIIZiu+ZB/WGxVucxTQ03sbDFKO9PaZ5SH7gBtIjFFqWQOIzgUOljFaQ4wbWQXSd
SMTQQuT9RVhskA9xURMABtRt6R5S9I3IviaJSgdDV/+z2B8d76uZVg81lWQzFl4Qw6ydZtHRti9G
aavcw59eqX1h8oPGCcmaLbMhgx06ARMUceCaZJnOVmOQQr+h9zGbQw2AdFh6MY4ih8FRgdi+Wm+G
3reRjKTVLXrZsZ1TweoIxKexZDfLYK5PmXNRWl/fjT5LVmreJECRS+4h+vlJE9xHP1F0uqtzkuCz
GeZBHU0AAXbkUZcFFcQ5i5Ml7TDLWzS2xY5EHUK+MPPK04W1YhGU1Jdx0JbHhnbrxGMbn1Ye6zFF
TE0hjjSHQb2RAhkOYyBkG00X7jFb4Ilz56Rl5FAyuXItBckf3zV51WHvFl4X4VT3N+TEEEO9gCD7
9FkuK+fl6XYwlUretuYMKJraXFldIvWN/ZELjBXqS/dzHL/+0hD+K9bUPyIzrEzpNcv5DXesZMIu
rw9fg097HJaCdPdN2y+4UzBrsNx7KYD2KZmOAHGvFXv3+xhwB0nN/zjs2sG2/wwvM53b9yEhO89I
YCpB5y5IfcNg+cW996ERw1QQIKHrR6SLTUrT1usLYs8PzRYLJ7Vwud+gwQoksNTpF4Wd08DwgnYJ
4CnaSauVEMzczV/z7bPtzCF50p2NTbNQOHVRy48m/b+4Mj75ds2rPZ224SMewEvLQNmh1+RhMa0n
Y1L0H6O2CBec4apJE7OESib9HMFsphNNRtcczbdxUHjniRTj4XuNtJcALw40+lBLlRpjq7BDf67W
yl+W7as7Rr1hc8whG+fTa/iUVL6i91hNdHzuAMY+DkhhPg0YWhgKpSWrAEBNfGT8vDK9i/G1ySxH
NGseGDM8o1Si8U/fa+Z9Up0vQKeoord+1PRCQt3moeB9rFCJIpYC1ttmnQrzYZ2sJn/iMknoRlrD
diDT199DIwSC+Fa7cx0Qh8pRQPfXbr6aQKQrTtQpEt/xa38IL/AHx2BVWTSuBjR6nFTdw+Rhsc0V
SfWvWp149CbZW+4JEfbDofildExw/ijXknhxxM9DhC0IoSlixavyGWjtKmH+jBTPcQv4FusDxKB1
cNe/sqhduWyld8lwdPUwiJ9/bapAaUmUNVQbzyulWyApo4FNhxDqyZqciw9xAWRDv04jt7NPSsha
nS47pu+5ywXnf+3VZwbXAeMONaunr/wiw1jwvr1GlJaeJKoRMGU5vDQ9x2Nbzvb0SaZc81oIVGV0
jF47oJBufGVz/M2vaw4JPVuJjOjzUvk7JWk23x3d5TaOsKAP8dRz0EwVhOm59Q6kIU63p/RW4LCF
dgq6mpXIczId8ijjWRBQZgd4AGbsYIaPNWMLovKplH/xNeMiNll6rKjJT0MisaoIq4ebDBTJEB9B
0HNtanU0vOd2v2FOaGn5TVcDqeVUT2l3mo/tUhEIuvZ9KvgtvdITS49379LS7p6J5Z3L5lpwcfhN
3uDNEYOVlA6CIfuLuZ3gnhxw24+j3yCz4wSmjiJyfhMRXGsnZn+TCxLAJkVIMIz1Ay2fAaYTSNz9
Wof/LihYUmxy7zeG56jC+iOalkuznEyF5wmFP0Dc6GbOccbqyne77EvzlfP5Wh+eVTuefsCBMaxT
m9dZBOIxgMDbJxQ/8KWvQlnA88wE3v++yAnU0CmLqqwQKZG05QYCD3OteFewI6O/A+nHcSxsHxTD
XGHX2T39A384bJQeWi52VMvLfpWpKmG9gplrmmN6f/040MuHjFOiB0ptvig71hJhY3YusXnrEaFO
rXYnilILdWuZFhkXaRkCTod3d/KE0A3Mgw3wyGK6h1lNDqiydzTz+z013wtobm6sYDzUkFFhZ489
pKse9DQouiOQ0ERn2r+ZmQOV5crffndaUFN0UUT0Ohgsm4x0tonGfBpmeRBNeJg/zZuwSRE2SggN
se6foiwvdbi4S5dlsRugWUIvA5BhUKoeGFOcti3P9S7UKnqMOLNJa4vKq7aMyxqjdgn1Hwain1IQ
gQwRxstFmfFrIPZXbASxYPA+pHOyD0mZaY5e4U2cyE3BpDFpsDhDXb9SnWl2C+n+thtSlUaX2cqZ
CI3A8EzA3YoDvj8DVBYHFnhjsfgP3QX4On9M95Tbe9bod39Wjr/Y70D5zv9a2Ln2May4xRCV9xwF
IZ++2MAFQNv5tbLOrtGaSGBa1Hp5YbIMEgdYjrdS0QEFqh3DePKSSUKYN3jXfKf4zzn3NSTmdfPb
0hjUalejRmhCg399zlAyK3jiegLMworO/2/SWaSCilS4VLHYIoMU4b9btJ3SDhNJ5dJGVvKiVw9a
D/8v6UH8EjvGsfMrjRp9V3B7g8ZY+xah2oPGCSOVqZIiykAuW90JvxI+HIUCQrY2IZzvpFCRep1D
s5AqK3VXEjaVX65apmkmSS3dtYWLvDdbMRE6fRh9CzDKuko2jRVK9WEOmcn4deuwmg2uLoXBbtGE
UJSo74yOr5KtPB7VCyFIE2m2YxZ8TyThcpiBbJPIYBPbSzTaTc5AG9xfUy2vE6t5P2T87/HqkQuS
hDiveykzBG0xNdmOeu3yAajgsMBT+HcZY67Z5SUBszBFfTu4mG/tmTF1SDs5ne7iI0C6ylxvCaV6
HFGkJFGR6lTGzMFs4QHbIzd93QFPgdPZ6OMdQBFvFWkKKSTOmCLbedlPNKskW1bAgXiyQXiDCrmc
z2owVrVPNvJamFL29extf1tsjRT9oef2pM0XAbEu/ENjlqqO/npMWBkdHVW1OeF3wX1J25bkvnSm
QjgODm7wUF7DqRTviTCJ/CVepkKZ43TeYDQs6es5dGYqRF6pAzihMcCm2FUutOcM0NP5U1shdvPl
l2t1CjEjGRVniKrMtktijcAJGOIKh4dn/n3TaWFBzmX19oMCF85bpKnXhko1CuAImsOp1MO4w1cJ
/scL1atozRAbfqS6TktbKFm387tnsgSn9YIkHpRzZgdsweZA1LTl+lRpfVYGwM79hwMh2KsxOYgd
PS7ezbwION2tOx63ykixKbfOzlNB2LPeBQEjcgl6ZdZCjTt/nq+pGj4E3UflD1Yqg1Cmx44nZIXe
5gcIxrxJtTzVdy5q1A9XKLkaolTWh/Ruld8YbjlFqjZ8ZLHtBaQmAAsfNkkubZXw9WgTlRTxusW5
QZn4/rOw2rLOSblLx205sofCqfg63wkBnDDE5Q6GejBSuiEKMF3rzk+NBL3EJ7LTrh8DLrsRyYHR
2ZnR8EBCkPFnHf2xZyNODpktY7V8FFHoQ6MW8A8WWyenlWZxJloKmLdC+O+QpHYYfScPuNf6rhV+
VQC6L3ni9X2iSDbU6xzQQ4KrKCDPYPdFeufpUMoLSyzhQxVjfRepfzcVgEqVND0M/aO71DjIDwzS
SZ8aIGGUDUA8GE/WbS24jO10aOq8ZpKTyY78n89gEeht0P2LSGQQWKWxLh0UVtBCl28Bd+H6UqpN
elEdkm2ZOZKAvrW18Q4LVMFEhZTvQ5w9YIPBjLaIhNA3ekzwNUddJBxjfiDOac5PSt0lyQd0rwlF
m+u7qgTdVNwG0Fo96i9ENgYawOp/Una1CQVmE4abg+l2PdW+CtwFKoCVrJuUG2m3HazYo48rv6EF
Sdw1p402CdIt2JfeWK5TwmOl0f5X8GxAXMy0tkqWS/tG8tf/RmHtXIqEKqcqTlVgJPfc4S80UZ7G
M+QbHxQiC7ucqrbhoa2vWs4pE/kO0x1ykdhxZmgJMZ+xsAqV/rIuQE4FSviJfm81oDbRXCig54ud
awBrxd0Z4zlPVR9qkPAx8rPIC4V8XqWKcJemt14f68eIlOhkKs4eKVeneOZEEhQXZZwOGZUliy0w
mPEMRjKaTY33/6f8SJsHd6EkVt9UGfh3avGLBLujhq4qtpdybMZ08Q3BusWLNEJKDz9rXVxsUU4B
EF2/ffc5hqiRNiSlQypnMuVeshzthgbqBdcbXje801HOHMnt2dwZEVvNsn2O2E+WZnjgRVibzSOK
dz9ffV7ePMAKRvyvYqMAwo2nw055X2i3JJgtyjxF4KOSQep+v3kLp0bnZwMscuJUc90QUoSvtYGz
yHQQTaV6OuSklH4y4L7b43dgU/qXFL4FYHMgAe9DFGrIydttzUyYAvgoQstSRuOxFwrDG2ahD4jK
t53FXJTHhqcyP4c3unINr+I4CFi3ou3asS28nA4P73TOgp79FwaFi5zkjRvksKwk7p8mdoyPI7TK
5HQub6AzAaDVjBmrQf4RSLW3TazuGIk9JN/g0pl3A6EUQj8hj9E66bMCo6uZLT2k1Rp0x4ILD3OQ
/ajYRsn70/LKrI80FPTnO/RkTQlTK/6KGU5WIL9zX98QuN+QDv22tB6jNO6oYuiFv0r1oiYKpMIw
GyiLuZwztnbPDlUuQQj6MIavPbJkSmRMns78s/4CG6FqK8ygNmx4XgOJRvS5rQPGBO6Kx0ARmYBn
omCdtLK8vQ1y23CfF4ufC6i9R37cO+K4kv4GSOscXFrmdZmojmAdTJykZswliPArYc8ugTwXbzFM
N5r6yGgNPrkHR4RPz9iM08Zq/ZY/s/e3g/0kJQz9ZiUY9lKGsCGPlG+/morBpGfzL5oAV2rW2FPp
P5sPSeofxlnUyr5ln9/+3H42sA1khk5jeNtn2xgozgcJ8PFjAGKVri+Wxe/cFxQydXNzMR/UPhQW
JgsGL8mSaFPta2A5rbBD0DEuvsffNyZSjvB2qmySagFKNcWQ38XmwY46i2bVXTCFZK9MWsI6vyu2
dkYKBkT7egcf+1uuVGlpVr4g4DKb7lpMaBuOSmqfjxIl4GEEC1Q5NjXOSBOtHVSOi6FHpldPrzpF
job3+uw3boJU65rgCTpw6HdrO2sowGEpgmlr1CDorJkT474Pp0CMT+FeCJbW1gDe1No84D9xG0MH
a9WCK01EF6YIZBHyplmq6wbuOAg4F+GDt/TPOLHPS+azR3Z2W2qEhULtbwGnAApg1XCpwd/kTeqo
o3JBvwG8pALQ7gm/D6rxG13oYJfwu2bFqfEVe/GM248NyQtul3PU2ZP8zF2P8pqp37wyohe76cMp
HMiHtmCb9g6z72bl1eBW8Z4BfbLYwi+o3f2gXkYt9m1SzZlqLP5qQne55AYKmpDv/mZ3xEHAiP1r
ZuP0pfmeQD2kbkAKZXBNOhRZsHllOIQI23BRYpi2bXuQ5YcUBpMtL+LYkkX61T6ui+Yd06vy3tue
tP3yaRCin6ErWbWUXZa7p8Zdm+Lg/yveUyzCudf2n4Ud1St+E4lIzEJiZMIhwzdgEowWfKJ0hRtZ
UdjzkzsMFhNewgbG226TtDKdimCUqfRjcLZ+sCx7k6GTECaWG5JpCrfptK6MNVkhSfIXfiBgRPbu
C1p5hRtj8CXsUA+1v6rTAU2PJ6AYeqhZkvR84x1Az5xCetxSvYlwWg1+LJ66TGlMAD7uVjx9nlFt
XdjNpL0rmN2FtCWBUDGPD6Oxgq8E+2DK4H+leI0i4Qokw6trNOGLlM/yzXkmEw40I5Uz5sWBUXd5
wK3DfGdobY2AESsNrE65HdLQuBqs6qHQP05gmdjBmRSTWxEGS0pRb/DAGTyU9sUiKOm6WgHm1P/t
Bo1xp12Xr5VrOG4a7v7RNgA3O7VxiMZ4nNLncSWTFq0cCOMpLwpxPjOmgIaEcWCGI15M9+aaTWh0
EgFdtP7iN+IjZLWpZUR7HiPN++wBF+Xx/+eRp+ndOHwsLxTEU7SFVHuT3PAuaWpzEV9YAvOhVXrL
qHSri0vCWYux3gU1vGaugRDG9j+A1Gj2S4590zK+0xYXsL8ZX/V+Gz/rhJ2gZtfxXiSP+yQgfu4m
tJdbtWe3ChmLyXMbMXPesNfq3xMOTWMbpBgk/6Q66p9hfbhtK7+p1RXurr/7/8/LJx/8FuCZKDou
GP3rIjMtYZna1zt0jON99hC7f/HmZn2V4PEIkfOfaE99QGX8qBGuZHwtNInMhHrq2seOWJB6I2sA
m+hJAdalg9GTpOaJH2nBXCe1NEthJD5RXFSAj421sY68hLB8POxhNYB2VLRCi87e5tPPxbxJo/nc
LOsqYW1FT2Yl6/yx7lQwScfzNrgjcBalcKDqpxB7I/Ll/4/hLFKlyWlmfZ2VYZILOL+o3jMWOpYY
c4GMvKv8HGY+x/ofCEKWLAKCEHo+2fw0M1W7ogqfEkp+0/ZFaA+qGq2atZ0b7PbvM5KahDkBgdgZ
LJRsHlJjiKVg7V36w4omVFlQ01soRd9ZhPnO6hQ6//+PPfdbBPfRt5lZYYDwgxuPqKCVRTlhzjwh
UPRLcl4VwABHS2iYjKJe5z93iV5e1GBx8O8w1hw+eed9yC7yg18WfU2521NLIrC2yiKTDjWANu9J
NBuIY0mRMzqkj8HMaPfE6D4rpUYqSuPhMFyHuDpjccJMWUhL3Wlq7p+lg4eA1HYe2zMgohBXj2wr
+tBdDMylNWYhC1LDaEzbgoLh+oU51mzJqbulxFb8Cee+E4brXomQqmvIQkxnlecCQThnzzJ+HtoS
Cj6LVehZ1zBNmjJ/jDikt0l7uoFTwLwpp/F8IrivReOg/Ars9jh7j8tuskFfzKAsLNtalFFjq30f
deCwpkniY9aGG0hCfIJRe84wk8TbCBEADF+VEWTV1hwso5SqVTgazzI69jWeLVAWqoWYN2qnlcEg
61H2BrLlJFRunZoQxdI0E5WGc/p0MbAq0Qhc/JQjQHVSSKLsLftcJvFuTDtAtPmrwGZYdR7oPl20
iX/aai2bpk0tO8iKnI5RgG7Ze8nfxNjvA/p+rScFjGlO4+6GV0eSk6U1gJJwMYqfo5Dfs4gbC8A/
qgIeP6sw+QM3JeDEngUJSDTDLG4vR60Av8WsbRDmt4X3WERLmvlTMaLcCTpoCrEInx8yMLpM38op
By2PY34LOT44IICSL9d+zVpeiC7nWYFOpp/tDaWQp768E2AWMcBK2gZt+6aj3GwXn6BOzehJ2Euj
L2RvYaNiAH6T5q7Y6vpXZCixC+/v8nC0KdB4lC1/SgfGBwaj8lhNoapoyqWA55mEoPbWV0JoXJ1J
1e5/8s8Dc2UoCr87vXrpm4pnLO8eQzjOabxwoLxkm1vK9TR8XNPOsbUuIuOMjSfrsYWstw93vqWU
f+RBdWHVh/Dqd8Xp8h0YGopw2s7wnWeu45DiraiZjRfrn6BN8xPWvwkrRN0sdos4BR9NqPxhDH8i
Y18ZKaXvtN3J2ernxRqgIsNT/HFV0aCuaipO7ntndKXI9M3tD9LHbm9FOFHn/4ywRwMvCGR9C9uZ
4hxnVwOYiYkMrs/lEPjlS7ahKc+11yL6gOHVrJbxvDxHwiIa6baE/Kr0MIrSVb6PI9CSpWnmslzT
daFO591TYKJkgEwqcRR5eZIzN7xfvD5KoFgvhviXIfovX4OYuC0krqcbhRU8a35HKC+5Vi/e3Uvn
7hTPxa2WWjvxlYeJQfFpmkVErhdMIGXaNaoi6VeY4N7tXz90bGubtNvoDfJx46dftfGVMlXmfa7z
aukCwrBHYIItq8FRFsPkJzi5PpHGeXRpryDjcX1bdd1xs7892erhs+uz4J0K1w8OpXdFsAKdnnNl
0YAVh5TUF/l3gyWqFfVb5eBytPn7Ttz22oNJPeOamLQK0tQ02xTAV1nXGkVykuT9YdRL57VU4bj/
IOBg09tsdf/zYzqaNxhVdcGsZUy2EDwC+9HME0H0ScSWiywnW8DfvKogCumMfassQOI2T58upqhc
JkKVR8qptGZmahvch/LGCTPNFqj/CEvfAsVZOLtMnjXIXI5wCilZLGS2cWRDhrfiS+EIQ6fLQjd+
kLAXE0gn4kUfpMPXl2hhDlIOBMq3qM69ecsepfQEuukKbofmQzQwG3lRInLbjpGNtT7k+FLaR8+l
NDFiVYxFZjsq8Ccqkl58CM80t6laBeKn5AejDwzlXB6U54BwUz1kpuoDvSkt3eJGurrOuGBeVtBe
9bgc5dnEtqGXWIC2vczcY0OT+oUh+VlJ6fG126IJ7H1wEejWLkeNvM24hw54oNm/My7SH0gRTf82
Amx4JUR8yz3p57kJ07/hTrgOyAo7rHT4tJoxZQvNIJAk32iNULLFnZb/Xd/o/5Z+r9D/bEfGRPiK
Gm/J/TKYyHIERJ9RockHLavLx01YZveqWIbTWh4kMr0fZJSmn0z+BM/D2SyYekvef+v46sBO0VgQ
MZFSsCdiNm38V3EYVpolu4UOw0156LyeDRRv2POCABvgDGR0HoIdgXhy6bsGz9ZHmxCDr/6ist9C
Ye358Uw+1Ki2Dv1HX4EHQ7MyfN03uOwuStFrVEX7iWUxgOdbBh8ZKYjeWvkQOoy52HuaT7cjMonC
voPLNO5zJkNuWynnw2DHpMi515lRS6JS9m/8RPDm7JIbT4/Ldg7D8mSTKtWkrrwaREieAvJwyt6d
f8gRURRUV10iLjQpJeVD9hB2hZ79bKOtJh488UVEdoqTzUtm9JeNtNH5wFXyp2f9iZb06I3+qssr
yJLTPbL9HjSPdVY8P/Tnxqmk4vhE4HbSn3bjjsKWIaCZJpAbJXfRWdByCTOnwNdwfeWW+6aXxe1f
4aH7dt7nUY2ZktXcvoa62FVjE8ULzQvQpqeBtgZ/6hOLqINYVAHuoDLxQ9rlbCGYHG1HoyszGfDh
OTx1yu0hKcfgd3ou5ZoPWFzsj6BXG9LdWa6r6j7Esr/zxM7jeak4ycVFaUDdyJxiw7JBqJjTcDYZ
GtCwn1DlNXFJTB9WXJCLVY0r7TVYwx9qmbEfbJZd8tHEwFx/TqjwQydfQoGbT5zkTMQ8Rjska07W
K9KqNgS+K7fta4EFVBqKshUCwNS+cvY2htl7NiiRWWz/w9dv8IkjJeGdKeJcW9McCrBTIprkNFuD
+kqecP73aUshBUoQFfgaO2fTnKqqFD45Wtwhwey9tKzfUv1leF1X3zEuiuysAESbYR2F3tWuOqmV
bLIelcy5NhKEhOwOwEnVhvJNk09mhfgPDDc0rL31+JhGHjf8H+OUDQUx49EU/0jgvzwtoff2vOOm
eEaQKWVry1mGfQ07V5jLHrQioBt7O4oEoiIOcKNSs9NyYEUJF69DgD7bnY34kPsYYsL4t6ciHFmZ
m2jp1Pu3g/p/KsOXWLbfm2DOIojN2V60v7iKzG+SrBASMTJXxLJXwrrBD9EYUN1j9xsogC5KP1LD
GD1E9dqWdtpItQm/XlXBi2xxDTHht0kbkouLiZUHpiQIW1AkjFEuJ6UBcuZDuyTjnfk2uFwZvLIc
/pWssjQAAmfp+G3sNYqd5MBDxZtXj9lOzUAlF41aEUg0Xm2AGxbE+A9uWMS6NYxtu2l1Ek2dqhXK
b+HdvqEAQfHcxLktNz+DMRBTR8QfRUHNQxc36l0qxX9uYVICmUB5J9rUVW1YnjeAgn31W8XpoHKG
cAmJVn+powbNX935VAFtDcoDIEURMAYZCdgA0nOTm0cVYn9ky1MptNzjJKOQk6YZ2oSUEEbMVhx/
4BsgXd1mGSmpUZFJLAdSKFwUMTsTzqQiI3X/TQe1RirtuETUkGOSKKg3IHXaH/Lpa1J5dTAnUGJ1
i/AHQGrCkCCutm9442wm6whFI1uTOJ7tsoSjG5550oSsNURQgsbPZw4yhH6j8QEal3MYOyk6HeHx
0poqcakHuBh8AbllKcRinh8TqlITUvrD5hSYyoZKn6ayXATkf+kdPNRqqMV2TJqotFsyteJVKq21
0SDUjGLGrix+1JuUBnJNkYwQ9ImmV117yIRL7+6+nCgj8tdNby7WUQx3vI7JJ/2TvpQqIescKUpx
PBK8f0sUgubTpQnfNbgJcMMf4NvkgjNcEq/MxZdCp96ZsOzG7WjV0tD723jKv7e5hUT1ZUvlfRGz
wyz8xvRkT5kYPn8Opn76ZT/pUsd9e70H1azYXXy6BrrCn6MCP01Vc2meqizHPq3e8TInCMu7M6dZ
ZfJ7vfbbGWeON3uoTyPSnQTN/6C+QJq+rqS4XAtQ+SSXtSBCD67u4YhQoUspug5DS1qq/0MUfyOh
BbWsCth/gcPBuVnu8KqCnHNkqx6RLKtQeEZOyVdo6xJw9DcJJQdnl13wrjn9zOlg0nxep7G9kzcb
q+YGIEvAAN8eTZJGtjQW8PJg7RVjbJSiUBdmYDZ7D3aPW+Xb5hJ9iS1qQeeWT2FXmQu5fNJiaCJz
goEgQpKIObEveeTIrAauryKxK6N2gf8mf+TzUJOdaFVgznX3EJd5JfcCoH/+cfPIYqd/Ywsa82wX
8nbm1D9zNUUqa+6qPAJMTqPGuxm62LvRLXUOL3X95K48f6J6+sYFpjLHTRwo1EMjK7DwSV/b0Pq+
P8E/knYOv5cbSiJp3u+E6VqL05NBAc1F47pl0Y13sw6Z0jvJOiWHU4V/4TISnSodEwg/yNMIVSd4
QCASVPh78MpJIMXMlQVWS5j++I3p198Eaj+qmQO5N/Co7exk6ozWNq8C7sUalqsDnTG2gxSJsffF
Jhn7LdtoKtIaD7CBKeYposNhaIcb41s0xJt5DM+b5AVCDzteA+yirycTnrtDdiyK7a1YCoHz77Un
DYhJXn9axAVUdGoGo/WBfUAVrQ+efUSlTaycjZkDVBCROWZ7FBdtDLVya3NIvt0vs9+ZPLfCr3rj
MK3oTJyaYq2C657dQpGQ2Aio6mAQeVhOBM/l69F30sqq/HZ1km7BZgtmuMYV/RNyyOf9Ggg0lpdH
ut1SkYX4zLbYKpc3Pa9NF8UwwtmNC1Bvr0MnwEtZNYuWYpUVNPTT2hSBH0p+qDa2Vs/LOomLD87D
CipzsD0ux14GKWpW1F7ID7UIZkYAaflHlj05d8XrzoCn71U/f8dieuG27MihFWpfyHW5OA77x92d
ED3OnjH/UmJOjmuoP9QqPCHN0vIfw386POwMBg99JNfhnluNwyQLuacEqx7MpmxCICZag9hcole6
eYguJRwVBxEcl96MGG0xsXN08BcsOck0hwXNnpwPJVnwTU8A/EI5KgQh97mcTIP1w6hSa32qFwUi
Cl2J9JjlmCDpbuqRHYXpBLqh+3zoy8QTjDzO+zd9fKwX3NQKejBqGK12o9o+iu+mJWMwN1q9Q8WC
LBRglpUGUxD3NYakw6sPAUbRAPS5PFVkF5axp2fJzenMnX9XapP1J5b+zXZ346Nyu22ZNjRTo9L3
Uen8hvpFNOjx9NVv9Mcj8wEUnCmysJhAhGSY618lWLb5ZBsgLuCvawRmUjXuJFOCkY3dXz4lIxo4
Hf6EAhqoidVCXXFBHp4rOxdzf8B4DMxs1w0MWLJxeV5z47xUc4KhxQqFvGKwbAggS8W6yntk9Gxh
N3Sn3gOSIEghLYePvwcaI2lbZFp240ACESAxicGJCZmlqsAQzJNKlj7jaf2RLlZDKBSuodwZKvMj
+iJRqR56b2RvmgM4eJDGAb5WE8R/CaUEOqu+ctfj067m6sz+ShZdEyY6B2A42F7A0eolaPQEevyN
EeOLb7Fh7Ii0gREdGrqJZp2tP8MxKaEr17t/G+vtB1Ayp1cqIVmtzJ/y2afntsMJSLemwfbujWzq
8HU22SHworqfvccDfHs+pLTe/f+D+MV+V2ymZ/1EENuXW67+I46g0X356ZR7CCWX0iohUVI8IZ6e
VUqoMVfgC7bwN/UOB8PlZ1DO3kRrRRWgDAmKlXfvDyTNoAbQkOnxg5zSTKYqRM0MXr65maz9jE1n
P0yqi9DAxSX3EQ+ZldTu36ERCfoaK1jcDMcbYmWmTozyV5tzuc+8mOtX/NQhj3HNiJqzdRD5y2l+
BavdoOuTYiQipXbXQ75wPJhHBaKfeXEAaFi5o142AxD4iKok+cjYB+M4J83k5CiwQ4rD7FJafufO
f8LpWGTM3f8nVt/vMcxb1X1LMJsSUE4H6JzoNKPZHCNmy6pScBZjEpSt5ejSG/SRAW8ScgCmVmdP
xaLGr6W6N+sAMBPhCdinVOCHqABzh92gS8bZyg91dH4RbmjQy6rO0ttJTShHsG4JdOq5TQ91hVDH
/u/p+66WQufD9I0a7g6LLgy1IR4LryY2kLbW3nrI+FpC8p+KT6s0HHxfdRbXiHs9ZmbeWPmOA4H5
nu722c1uG8b4bJTBwy/wiEa90EEGLGwSZRdiP5oYF1dyrS14765ktqCAktfwfMvfMzSMPZXmsZAX
DllJYf+e3Ae8ublB/j3GvbFCHC6iIs++asNhdiY7ct8CcyW0BOue8R6VP+JEmr4bqrzNOMTzxJQX
sh0RMMBJ7wQu+MlCoKI9qpd5ymzfP3fGEBiZWb5L4kPbCS1xekSNuC8lfZqf46SQgQv64pNawxHR
tEVslJhXK+sz9xgj+aOr/6sezraVL87H7sEia1GKkNN3FPNR54LsNkLAUTvjbcngjiNfHsj7CPj9
s1LLkoCjtqOB6kiAf+PmnntOPuZIoqR+Z6GRizDNvlpSIJv2VwkmfrY8um0Ihs+QOE3Y8O09Luf5
NztPkcDPSSZlWTU3A+gvqGvjPdfnlvONRXTyQQHyRa/SOou6dSsLTCA2hdHMbvGh02VnbkRqWUeJ
Vm79vHRF4IUEeS7e9ybxb+bdiwzNH9Xtjxfiw2cNlORxiD0d6hPFDlWIShFiM+ljlTeU187yAbY7
MjCEREH0x8vyeF8EETvFeX0QOCebff1JTIxBS3cvB3o5CvGIgZRCnfHsqwyQwa01wEwFwRl/QP6X
w5IVqZqNtSxkm90InArkjh7t4w5kOXzx79622RXdZKymOYFJDna7chhgVj3CvwHNQeO9laQ4rq70
vEKleWDgrAnXlH+mlHtZ8hsstbL/MzWGPFDmg734ONgzTNmglk0kBcN01SfudPcR6gGEqPYrX+CX
J5hcS2WHxtgO9JkBYsOFXUG+bvCnSfiHJRA+XC+jI0QefkeX4OXND/RTvjRsG8VXkKEZcWVZpN4V
g0PNvYlfFoOmp5bsGp78adAOGbuAP9AkvEwcOO3gkSlXcu/i2MhzexuBYQAYVVtWkbsAUQctBXLs
3Jv3/f+hxQQHEwj+oAXSRhhVSiA5mV6wlmr2KYACmb2akPkAkNtupYP8Mgb141Od9I9nd6ElxQ/5
/YuNips65KcEWz4EKt6RioQ85i0DBVlIq2VcmMStyCOuT+HISuTMNTY/TBgjuNy1ll/lDXIrI2Vy
xJbzZ/GCdMHENqJ7TH43gW7965atANdkXizv/qxO96lEHiuHQ2AYXEg5tGtoQRtNkKTqb3Rgx+0B
1jQ9IDt7W3UMvkIFWy2TJgzkTLOpRZqywf3kJMpH8EOxg9AQCARq4bP9DLBZU9Hih6Mhtz2566ss
iGnTwESZWDVrxY9CazU5hb3NK8IciGInHY3MlYJ9uceovhm/kFGyxGvB42wUO49/b/szqEzqDRAT
yGHdASiDjrDoI+3/irNUO3HvCPZU1zrlZoso5sPxqDOnNyTXE//MBuiFKg2WmDCND4y6aNTP6K5U
dho1Bb87CBReHU+30JTSRNkSyfioGmF01+Zo6U+37Yn0nYjdul2cERryKKAN6jOam/+w6C5Hh87U
5xv7iNtvNrHEtoAeL0tgcVhUIshOuyFEg4tmn36ft+RsCBKsC7fboQYbQUJEjYkV447Gz0TA+g63
XTe9ps7c+STpFGthM+7AcchqotRIoRLBQSX51pylx0MlbmP4kqaHfnRmxVLcsz8Lu8DVR17qPjDg
CDTPns8LgprnwZd5YmqjP0/dBo152s9ar5f7n5O1Uz8gw07CxukBYmMoxKuQ/D4KsLfH65c1YP57
7ObvimcvdbaUmrJqF9GUfYvNacJ6D2cFRupd2zTyxKAwlZd95EyHJuipGasDtGUm+Ye2So6J5Y1V
jmxwGRUQVnftVC4kT0PJAtucAFsHZBIJmKykHnhEhujiC1qX1oWhFrKzF7bSJNl7E7D5n7jVQ90L
sP0BvvXK5ILO+QHDIUQAA7fM7dfvu6ACq2USSymgqHxyl/n/6H6fk+5lgE2eK7GG2iExPp3Q7oer
BB5gqIiymIG4iKjj9/gZ4PcnOmmyuvYSkT8S28qRpk7xVt1aXq/cuq/bRwvUMK5a7qfmLiKaD+pg
QFN/CojGyZI3b8Sqob9ud+R+KLAqFzIHi4GNX3qOXz9/76BlWwG9UknuoJ+XQLnl2dTTIS659QHh
z8DoCbt/3n8A15wPop/+jQR27X+O3an5NhxdXXRUZae+3ttTILUjDCgbsSieRA8LAfqhd06sZS+O
VA1xhQyXiHV1/SNgARxTsAS9NpDmBHZd8RkOHisXg9+5gSTNrO4tgwK8G7yf4+tUCIOO/Q09U/mB
LYQ0fiyuhw8rGGp/1VzMfGdt1b83+tvEXKM4K3u8ZxnexUveF7dVXatP+iT9lL80XFXDkA9ublIP
C9p3YE52cS+YEAlU4BzK9fIqKE67vwDO/5wqgnx1GvLQfKFYJ+Ub35CxDiflrEm6xsMlCJzlq9nQ
4fChPW2Zx1qGdrDASOUrQpT2rWVMp9eyN03eKYw+bD4p9K6DbQkWbuTmok9Q9Qh2ia3jTxLVm4Rs
X86MDBCbTMfxZYehVoYdn64fXufpMTbEh69QUMSZb/oXoZQyS8Qpvynr+ckWkF3wtVzQ4EaDsJpa
yeSr4MHpc8tAdGDoD9+3cht/new7fNeAIB6cuAOXe8iIdTwPk7RTSaCeMQC8fmvRlKgh1siLASZO
9JgdLFpNag2MBJ5PhJaN+PIeCisHRYDHKSdZT5HV2KAUhTJwfu0l82jYjsc+fYHIsN7cg/kWp7ya
AnEhtgFw/1ZPFvXs+f0+YJ8rBBx6MFBVobdb3hOpPjsRcBxEdhboS2GuUWG8i7g9mdAC+Scgkpow
OUHUTDFMSGuIgrviFCT9xV+bVKFyk6XFwZn6dim08ayKIUY0q34j3NlRwhUN5+JCuAdiT0ValOFx
l64+g+xZvrqECtBd84Dd2RVqXQyqUdT02pDPkKiub3psUsdiSjTx3UnKt00XW3E8Xi0jLEN/y7Fn
LCtI6PocuF45lS3UNpILzVSZeRdzcMoumMo01zAJ9vkq+PtQLmwhVnG61Ac8CZoQ43cTbMQz2jpc
/n4Uu+gNUq22VfsrsW0GjdZAmGRtKdFzMNEJ7UBRRCg+RIvE09ti2Cv0Z0dBFrXgm3EPUG57q2E6
0tpT2QK0MPJ/KweaieHYYGxo+ixsiTu/PY5HytS3gqwxVb2ATPDr2N/haQ+rqRZEgOb6Ze7+tovB
bbRWUefBFu6f/MSQUGVzLX5NoQ6KREJW9jFx3x+Cm04oKzt/sW9AW1LzemSkDJW9vcIW/fxGr8Z7
UFP82B4Nnk1XmfYEd2kdM5nfuDkegxJwB4zyKdIqxZaChCpHkzCmT/siaqlAR7MYwfSTowBvD/mQ
j/92h41IPoj1HRXvkUtR9H1TCfJgkeh+YMJ2kjlFmTH2j3qml+bpZH+XxD4aA1lXQRrcxCmgruUF
tIjhfKY+usOkU9PKfsdg17bMb55OyDnxQu6xCRxs6WcHk5AozqBK2k+bLb5pzbW4UaZxva28X8vP
WZJ3FXDy6ucw9/VJQLuAThFM58z75p8Lg6GIwfpYj3J3G+TjxFHUDjf4RWJFZxXle1CahF+UCB0M
j2Lgrz65do7JykaBwRJl3XOQM0LgzNCU/N40+71YN0aYAhvcMgREBWuCJ3Y2aNNVAeYRmp5NLRzc
OeQzr+qVO/doIXFXCwJCo4bzXfDqjYyvuwm0FALB2rwcWl+TAScT3pE0jalJm9HVLTLRCjW5ook3
yIdPpjk5q7k5DK2C3lzK+pBSLWRTctGGCWPgafKiNLBEjk+x1KFHYD3IIbjzFnUztLK7jV3K70sJ
ZX4DDG2QsyDxiEe3isPJg+aXrL8lFGNaSS18Ei9G4V7ERabhdwqH1NzfWS5ldUHm1mDKN5Gesw4J
qLP9gv7YVeso15c1/6BPkWz3ZLuK+JbFBjCrak2gUgFOpdHY5qOEJg8I6CF3DzI1DxhyGlHdf336
RM9Vy0YUkg/BNnnSQ3yOtGSEQaMk6lHmxR78Nrljhq0opS9XGArFd65GI1p/oQPtgeiOm3t0mHR0
9nsCMu+RUVAHmoXt6yPBl4DwVtqDaam8ChXJXP7hVtQiwRBVsJV8Ws2Y86MmUQknPwjgZYlDImml
cQUifYpXvFGVp5RtN+hG6jBiiAcvlspGXsDNRsbSEkyhqZR0Xgf1DCGuln7aNNBmJzaibkhoV2DE
hpv1tjZCFIo9riNtrxtwq7pIJDuNv7bIAU7SBFP3MQqwI64yygvzN1Xu1inaumkrZ6hpNJE9qTE9
wTEObhzCt7US/2UTa0nCKwSxofJ96bJtB2AyVlSjrKON+H/LJAaN4SYZvFM+c9WNXChL/udAHO51
TKU3MicBwORlzRoWlnA+BljJ3zNO5QfANIlwrnmJ/gYwfSihVTyFhpoHzimGZkg7LckiJ8iaaNyP
D8eeJR5yExdAlbMwGT4rQG/wfhDF37hGOh4LVyNLDcaP6pUs3K7vo+gvdRv4uzV2Vm/yQz+mEfru
Ws9pQO7hQ3jVkyne+RRI5SN3eSWrR3Z+f4AtM4uFCrIiAgv1TwabBe3XslDUTUz2BUlpXLBw5pKU
Z14VcxcZqM2l9aA3tJig/2AzA01n8cjmTQEm2Zdqn44GBnjQl0Uf+ICHbVg6pSi87m30MKjwU9AL
BQSwcEWPtOUUYs1UxIbJDHW6GJQIhB+ERtN/fFk8IVv/CbzZoJpyogqcO9LNePWzEn8kmbep/Zlz
/KQhQyNdNrzHtnOAP7IkuKqxFvF0UbNvG4O+JEJEgl0W0IlM00shurk77wjMuxZUNkbL9et3YxTF
3WIux6KQ7Fp914GYzdvA1T2dXVR6YWaZzQVmyz9kwLhihwcXu+wuOgfm7WFebDYhQw/11CO8HG7L
x6SuCLE0yA1faoTWy8BejYp7zrPvMrfbebh3d8AAW0tuWt/GQFpdb3+Ac07Stg/mWgW/1T8uswNZ
t7HWUDI0V+fZBOYqU35r+CRxWrqZD3cQ4Dvw/0DeyI+kgn0kuiIADObmdpcA+NBqDQtRP7mUohik
adm7MaLCCyUBUuqe2U8X0x74Bi77hn4tQcuhnvWOMYdnI8f0A8JJ+a4MdxE+AIPAlCJKcY99xp/f
hdb4AjPDj386BvuL5o6pIAjTXv6g/InXk4V2LgCtk2gZyFXkoFzxumBniBSb//7fSAxaLWhk6YQG
eLuayGnoSsv/iSUv2/dqJGoUFnIyuNy+a66eMs7ccJqNRhGNZIYuMHUL9gi3tqgjWIyyw7KeX88O
G82VW0Yf/kJD4nL2qwZKbiHfoSbXbQyqta1/k09G7AhWAyR9vZKOmsqhZlZhFHC3Vddnu/0uZixl
abzk12mfUut8a59AE7jeya3YJ0XiFLRoAKUliqlIq7zfMYPn6Nh+r96YtAx45UHxpEozEzIvYDoN
47YGzuUkJegy8I7xzJTi5LIu7PQAvmVvxs/UB/fasnE6ZAZj640cDDjgJ3q7yLYxha9PpSG86kSa
Fxk1EGsnaEFnwRQxdKQdTKERCapSqy7OL7FTRHJV72vs1QbchwGReTRsSAzWNaDN35+S+Mn1pAtJ
eM1XURR1hOp4vEtq5uDsEGCdxpzr3uTFI00T/XUVj2EFuiaTYYZz3Qw7fa0RsZRQxHN11qqcoXKn
pskGGbcOyfqGrCQSjIosLo/IQtSqvyMQs9l6L02mnFuAkiB/Y33byGnP4iMIu3HqDSanPVqXUoz1
DZNh5InbDT33lsXFMaysdWnbmByQzMQwPAwpzBBrYQXUZbklHQ3r6cpv8yjDoyRHOXVg0U6zOuHQ
FhrlMwi5Q8O6szO49YGw++iF6Zh5VbP28QzmE7ZBZylOHhrFcWQAzQnuARqjhewgidx5gqJxievi
RjpuDzIHfWM2GcpiOR3KMz8dtTxvN/2SAWWyqAzQaTm+QwOLb6O7jxqr4mjETU2JFXKFxvB4OEv6
En0UqgVtO4RO7o9FPwpu0zCcQPU63C3zhx3bh/Pj48Zx7USHNpNdUNAzwDni3G3otoCMTtKYst8q
L6emt0VsaWUynxelLrAPEEI7WwK3v5lsJupFSFaQHU2tA8RroruFfa3sBomSy+tK1xxAKr7tWmAr
BEsMRq0BmOgVYO02wfIA217QksRI83KkIIGzP8LRDN0q++8+45i2fF2cyN1gCYrJRvT1AYm9Bpbw
1fWO7eAZAGL9ZrgpRFiLQzvj0wE14XMs/XexpO35895iCvKZhPNGpOSTmwZ6x/7yyajUiCrMLvaq
soo1cWDwpMBWCD7yQWP6GObb3uh+39rddLhYPmnEwQbyE4UxKaXwvwjnEVhxSg9AYCXHbO+T7XPw
70UzodsKhB9ahCAGS00y4hhmsScakCvUfT+r+M+VcTPiVKOxNmsUH18uhMLnFZULiAgTfDF+aTG6
HO1ndRKXZs7hNwM7jI8fBtBwSwVzaVMBgsMlTTlclZE00w6c/GIOJQlVF4UhsVs7J+wK9+vIYcID
Bg1icuGE0xWz6fL1obJ3c7FhIboVPu6drSgeu42XRKdRuGht7zqQnzFuObvxSmHTfMavmMEtz/t2
UQupPBWZ3fXk4+o0p1Ei64YjqjuKP3tlOFDFYu71p7ysWqFMlUQmh2tHcP7yQMIZOvHd32bA3rTU
k3R/JGKumLhTjxhl+ToGPr6H+zqnA1wyagk/7Cy4Ly+SvMH1Wk25XpBdC/OqnHhCd6zrfY42WxT7
GHMbM/+K/urwPMst470fefuO/FlJwOMr39BeihL2LIEowpeVnbHdivekMAPdGtXcw2CB3TOWHkz6
UL3qGH/f3KAvbVWaiC5ziC44YuEHKXMvA6keHk9ScECSHGuH9oyfXhmgwd3v5js8DAtIRwEs/YXx
RhVi4FUB8l4qYjYXrJ0kJ71pEUpiJ0ZcWfWn9Y18wYVrf5jQFOeAkYoQn/ytUqy2rLrZX3vw469R
qr4hL2KrnYhPsEmLI66CsYhRf/3kwMjKDg38jAoi9qvB8zdaXUUWLkFFlM64oYucibTXu1GSPq4X
T0RB60ckr72vawGlVRlGZSurGtYKmviUmGt8HD/IE9QFCXoJSXlwFNa3EDB7NN7Bb3HGhfqKfsiz
PsIxHYD0MMzYBoQ1oToEPdcMhYsKHiMHh+epFY51ZH8WE8FV61CR45sM2z6sXkJiGV7ChUaC4rT8
oR0FGpNsToitc2mAuROjOVoPxYYY3l2QSObwFjaRvPq1fdo+KPYvypz14UPb7zjQqfvBkrtdtf1A
xy9clwQ2ohXJTlwguDMo9YfKdxS7jDT/+zwtiPUi+AJ2LoS/MotqSn/jXBwYDY9Nai1n7Inl0cqx
a+5qgd9uHjebbucsklJEb6IfAbSpt89rsfUU/M4gUJV4ApyUc/k+0GQ74EK3APWJDV7GA7hm63jp
LUXBbOd2DRFzYEpelW7J2VhrZx1WS7lvf59wGb9qtPjkPwiWsrgama15cc5FoZ1DcXOtAnbRByTI
xJ70VdBYzJfY6K7BrAYA+0xkBXNy0acHK/BDx5X0CFBhhGZR3FbN5HvYRo1hpU2MU7q/zFSw7ok0
XcEUn49hah+QiseLTQ7jg3Ia8mV8qjuj5vhoMe0zcW+NJtltgVM4fkwwIXwT+OPUdPeSvBtQzO/j
9QSH33UxyPPQ8IdcXbU0lBIKJI626guSkPi83MHucjEHu0+GVgczrhMYdii6gMjVXnKi7OcAz0ZU
9+U6oYWf2hPRq7026Pxm5jCRnNFy54tgvqZJlTMfdQljaiVCMyj4M+4TnhsHfGgbZr2ltIeAtfcB
Xb09mhhuALhzoVi7Nu7D8bjXDs1BfCMnw87yb6ku/pX3505xAnk0/bgBv+MizcVcDfSe1taIlLmK
7DN6DcpDmoe4lwi7HlzvyPcDlRjYRSGyb3G5JTfodd6c3GeXuX49jZUqaRvm0ykq+Huzk0Z8U8M1
6KngUOVWOd6/MpbSZgdy8F57L/rEfyScbBV5arQMxeEFGn5dyalSD/2ITpDYnxZX/WbMNlB4RqY6
gLtQHUAGFv5ucxryLwVgU/J4bTqlA2PNjhhu2/qIQ9iRrLixNWQ+A54fAu5sQNpunS5qtLcTmgNb
00QYT4VUN1CrNSAYWMSGLNKOAA9hJ8Rd7qfTUwKb7hvIu5Wgsf5Tq10XFivKaOIjFX/PzcBNVW2G
zkK6TS9ulJycD9zNeWNvEWnX/8/Vn/f8a6xAmeZFxHYhrRailnKazGLjNdflb8VA0QIDoiBCln5C
rA2ZwtjoQwXqcXYrj/zwmRcnFQkex6Dmh7QnBlsbF+IJTcu+glJNIn5ImA98FM1r4VtAKxyHfaoU
0YAdYt2qE6VPm8K23Hdd3l0J01HiJA+yzCknyzhAKB9bYozzJjJyqwzFkwY3mT19lOEugqdSxy2d
A/kAK2eRq5lTf3pDoneJXKDpi7avsJ9Jdxs4Jc/R96mi/E9UHsCCab0deuc5EaktIU+E8us+6dSc
d3qgZvA7v+YFzPYWTWm2atqsOxd6jg8xaDBBa011CHQrxxU50kRqxPM51AFptGa/tEzEq+ANspXB
xGfvph2p9/vLcBEKaLy8bU4zprS+D68atLGwNdGCNc/Ydjz2dgIjzs6WV1EKkfeQ7dUpiDTb2m39
pCrcWw9uM5IeSakZam5pnrc4s8b8QUUouj+EwNFuoTvxR4K0t919PsZt6EAnwO5HRrxZCSTKeNuu
zg9aRVzwnz9ZNTEw0ZPVwVWCNIpR0W1nH5OuqtWsdLiFKhzJtXQ2LDgCpyMfCjGuP4fgTgdBJCQR
RvOuVgC0xWyX5j6pPMWHwZmUIH9BZp0Rkohqc0xAWFac7URiUlVP9F1M3/0WF5HHFbjKzD6c+qfL
g4rWZenBwWbBQSQUv9SaEgIBPG+fbdbfOPL09+qprIupJ48avgjSnCvzWpQCIOltMq/J1RlYcQh8
xwZWz+gnZM+NacfWpq0o1dtk6YIJ4RlXN6fCM9q5yXj8X3lKANREMJQVXHiKitBEIEN4hyYYrSPB
Fa68GoKpPbOQlFh/HSYHFPEGAkwD9MeMI6AWea/BFtr5YLZ+3kOev/5AweEm9dquZSE5SsWefMcg
hfd+97KcEWHdJ3m9MrfU56dRHj/5dMzHSeQOiOVMvmsi3o7Srw3l+qGkvxIAgtGEOgAj9cReoVF1
hbcrkViJp3RQ7DeIp177Nmods4X8AwUcWbI753rNB8akj9EZxOQjVqs69FKiFnEXSJnGQjw7tkzA
L4PxMVtFFBVHmibaCCKCIE/RyZFhRUD60goJUetKY1b6WZn6QkZz+kpbjB7PIrInNQJ1K2g/DeU9
F9bWi+O2lp93ADZQumxDe+ulMJXjD00MUy+vRynueUhlddwi7yEv8YC1I2AC88Vy8zzsu3+CK8cE
dAOOxAfcSHgRyjJ8yZsxc4vmQ4qjbekNeEYxwW1zFQ4WyurOcGi5cUsaVrPgHanlOXR43nQCqbH1
6SWhfg4pOwgMfEZ5Uq9eqRZSjtcCLf6uMfeqV24T2y/RMr/OULIPNy6oLM4h/Vjj/FVLS9lO7w37
TD23QslIfpXEW7gYnp+/RT0IkSbT6XtOZymzLrlsa2hffrW7pZkadGXni0dJ5FLzuIhwLAVIXRCd
6S2/p+sibYFdPxgO5jZciDvjNXfWwK9E+Tobsbny1RRqTdR5qfbtB8bCE1Ih4C7+UpsZvzLYD3Jx
tw/xSYPaFC3Asf470Sey/QkvSmn9ooi2NMwiuQBLSP5taKmx0X9sKgk5iRRDlkGkQbtidd/obomk
ugRh+gJeJoW+wYb0CfAitS1ySYSDRND5je4WJQ0tUfyFQAlFc4kIehaYSlDojNnfJkg0a5eMpgIJ
woyFxdXD3DcmEBcBT74Wxlu1cg4RB5z2sFhmrm3rhP5+R6hnUa9EatyArAO8i5PrbydUtRTghhp4
oTj6Fh0oJakRTTrJTr6HzRZFS+5eGSY61RQRAfRU3YySWZUXYVgxU1LDrGBFrbuFVgFMWHRXgFMX
JJRRdmMVMV17IDNBC3m/7TGO80mluMpPejIG/pJ1GkJfGuSw42ZgEuRIqRU7hKrzkIuq2p5q5w5a
r7Qc9Hm02yumLLsdzgGK83jtriLgqFRuCvRjKfFlBVbhgDggxEdA0k8zgopdWHagSCvSSARfgwBe
arS0QcrGeqMN6cE46ST6apzxO6P1pGvP+Okj5hIxFnwtX36u7n5vU5/gVFRxr9I8oT57WuNlfXO7
xsMWxVXGzY2nwxgimIHlKHNw1b6v42QbCuXFtO4GlFjtBFwLXVsy0NwVi+xJ1q3FSUJIX3a3njET
nXch0Krcd5HHLDZh7PZ8LeIC29ObfKTU8YKSB/nDQVT8XI0aOqTFio41ONxf7B+wVZAfLRqHJM7m
KiTNcyOSdA4n1mtJ3wv0SC+bzI0iFWIPgItgi62kExG1pLgwM8jj71nGh2KjfvNR5BdivYKDROS2
3iChq0b4y7uEDzIBCtmQ2daFzapePhs/KL/lq6WSqQJ8XiayxnNTGcXW5s12UlAtru8ZbSmmYmBv
px/zbo96gt4oyWwIqtCH56TCw2zX3Tx7X7Pcma/9ylLdlpqLeiMnaZrimvNTw+qmizllcLf+rb4F
Dje4q7ic7PV6DRWK1ORZ6imXA/AeNA/pqPI2M5MT6LJOEQLfszQJc0zHw3EZm0gnKrfGquF6BEeU
V7/rfxeKbydBCeAW20+40MiYu6dx+WYQG+SikbxoX5UWueG2mmtHf9Br8Ur1DKUsliGYBJSw/WrH
fJYff/kkcnYhzs1Lq3odVBrfyBawMkTDnX8iWbQuHtIjLQJml6/sxiIgkFRRilUrtyJ1EzoVYYVS
W4yPlHU5j9vHGezw5xsEac+79hxpfizbjjjrbIfNjgmNghYboKI5QQviQF29yZ089ZOnn8kkSsLs
Xfh8wX2qu8I/Y+Ft4jw9oKPztpD1f0x/oi1695P52q5aD9lE68oDZpOETku89EX1eXgxanfLKjXk
+j0jb1ov3g/stspLZd7NVt6N8Tb/vnA0MK0+KLCRWEXhjWnVMv2MkNSS0dsyJGcD+p7qZvY+eLRW
kR1mADo025fXtu3+UzaC0ZvXAD98NtTJZd9gImJm4dY1VUtoOP2v7rakL8qSaiB1uRnNPEoOjGHQ
7dVyPPLPIBcgNxtDvuqVJVvGGlGWHsVWMnPU7WSQpyW18zNZ99oxEM5qQZWL57ZyDkhF02vwcZZQ
WCx2MR2U2Eh91LYk0e0kIZXrlUYWJTxMiAjFaf7ga1Ax1s+YShFOkHqJZmbT+b2yktEqRjk8+fxK
li/mw+V5uiLfm1opUrt3zZHEU5BUDpa2n2bI81qP+T2L3JfkJRMDcFLZR93yC4tvjdAMIruhYlel
QjiPGEAOzUCurLfrIDYxs6PZjnAc0vO5AVIedDPQSRulq/ol1hhZH2GQc613Y8M7IB4iysn2wLvq
YkrJb8G+g+oq4vowPHAxW4/VnsTIUvXZxxH1dxQNoosAcT7cnMtO1IXDQ8B1rhuy4NsYpvOnxkHZ
d+c9dxgR2qYyvFLLIIaNcgGvqGs7lcI/Jl3TQf1cb9Xlj6kIscjmXIo2VIGUBeQWnIrJVHOfmUEx
tXBpLbhF17gS8/jH1ruiaAgj/8qEUgSR4znhzGtGoV0MyLRH/hjxRpMTtg5BoigBilQnEx8uk1gr
RsfMsNZyPQb710VscF264TQ4l6kOSa7Gysv6U16x+c/h05p1bOa99a6ZIEG/AoXlPa7DHDpdG7nU
Iceruj/Wu5YKC9NQyigXc6vR+KFTeGmEJLUjxqRDfeCVPjk3j+wrGFEDSCYdCe02RPjC71AcCTAe
WvzEtutRQ4C9/PwuXKcg4JXjhtgLQaq+2jN8Pei0TwZ921N3IWBZr+4EOhvJ3gCvwHdCiDH8Tdtl
BTVi+L7Spby4IoVm3vNXLb2pMCnD21yIi6YwLuceLY/G2W/YkUZNK3Maoh0uIOwyJcPFqCSLeWHp
hLTPoha8U6gURmKpsJVZied+8GE8+T+Tt64k9gJWVarf3xdOgZW3oIzYTzZL0onXOCdOGsvS+Fu/
ZcEkNmv2d80PejLXL5coI7mKyhNXxlvWrkbYuoAO9uXrPd7daLt+FxGdPTkdlSv1oIdz9oRRbsww
Sw/wbMTOMd7341PK81KiHj4CTvGW3kM3004kSmwn4duwb5PCw8+/92M0pOZS7thQ9wcX7aaETzBB
V5ptjw1birNF4sQeQUFpj+Ed1RRLWxXlL24SxfukD6U0WemFC94kO7IrmPGqKXlz1KVZ+ggcW0D6
AvZoP+nMNAoBRqbuQnqfMbPLfx8bch+X/NvqREah1tf/YmAE4py4VIFE88n8USCdFbjRtBH8Vxf4
OyK2a4E/+wLJJolhj/JeuH3p/hQmrDbpx8F9GY07wG7tI3K5dV+8Cvl8V6cP5bjIKqNR9o0HTD5k
/bHxLlHYa/rGm6lWCv+gDrSmKFBarnnmAHMUOSVrSEaAMYjg81+1fz37rZKoNzhMuqAl9rsgQz85
Jx557cxiuWiu3v9RCfzF/TwfTgcxdGiJdMhbeVGUgfcIZcVvQAJv9zvuoIcRiB8RXw2i3TCAklp/
xhGs5mKAh5qVaCQsz7ZLCwPN+n08H8VrNYYuirzArtQWVKiONYdkITXjQSnYnpMCdu9R3eO6bFkJ
Ejy4U92O8zyEmwmZwowwmySseSgOdNWgEQNFm7eAd8TjQZoBqihBzHH8H0NTTKE3VRUjYkp1Vsk6
bRfY3nO5C4KANweeePQg7BK6eWoumRfWt9DAHptYrLyl1Bmkag9tx3HHS2HDYmcb7UCAMox5xRB0
oK5+mEMxfyRerDjSxyL/iGHDLuKh1zVy28cSFEphBPSovD5bV9LTgy5riQh5L11Z3wCKdTXwktBC
qODuI0oPhuhN2wC+c8f1qY1sA35C0alHcZ6dJWc0gGeAo4BDewi/sBBVB9zMnfmrDA22uOKId01+
V/pZ06pQ2shc1N0dVqcfw9CFXnqqDAXn7EHrpe4MRwqU5Lk0hgIJIdO8L4Y2PqvIfJZu7MRusyKB
YJ3JZuKDCiYam9RqvoJyzFdHr5htqCklQXRNedFht5I8jSPaOuijg+z59ayzsaDDK1Eu97UuDfFf
bdp9nAV0ZE9xyuDOmh18QccxunrHOt1E3cdVHGqyrWm0tbsx+4dYbn0zWz5vmYzOf8SL3JHDF/Ky
aAt1RBjG+fDmzkbjOBjtu/FAFa5MMEb6JuNPVbhmxH8csosCLCfygLcS6MHyuM336kwPWMKQdrsk
hZ3MRTDxNKsf6XcESop2vrk3m8g5pEraGDLGu6IdDw6sSxulvf8RLZc7ZeIK2JLPrC0FFLYGQZuD
Lp9YTiYVi3fHp/XgtvUTVMgztNtPt6yq3D85WSjTeakpe9wuGmfhxrs5FTrxl4T9LKrFsnLZvSRT
Jx9lFtmSR9vM65r4V1pP2KEU/zKH/uxxFYURXE1n+L+vtCxpARtH3xtQmVcZ02DG55pOD/dbMnYa
kEoFMZdJoCoIgnUG6KdcYPymY3Npz1CDm9CdfIL5GmyT8eEBln4sd+JzkUKgLHrwk8ruHwcjbY4d
wrNj7P0DdCTL2H3Pc4HzKacU7cxQ4XzOw+Dr1O4DOpKnJXHbpzbdWJ4jdJteLCfZOVaxaHdPtUik
6AM5qhd9wu9PkjB0UJmT1Te2YN89p0RZwVK3Xu+GUFI1cuJd3Kp0hWFN4DSqWmHYXTeGqevgeCIV
5QuWdEQuix+BApCj/ekVCVb8dnm5L1gLWDk7vjoTHEKKgOODZPHJt/iekBAh+cyjvDiMh7b+HjGx
hJWswZdrc+PvvKHvm4zpatCRqDvBei56QYXmcxklFXNjwbzRJgcE0HvfwJtJdf6uCngsso0Btb2U
d7vsS3+iKDIDTwqzhzMJyF/pxZAbt74kpy0BFNskzsGXdgoC1/252Dx7O5oF+wKuisiGC7BYXnR6
Zv/s/uMpDBgraATyilI44/xrax9q/AZGfpEg1o6onFLTp5NA7t99uXA5Y0rES3x2OwBuLp5NKho5
Wtdmb6MlMjtZLS1/aVJdYA8QZYvArNQK+T+TfZaOn/RBlbnwjeQHQXqhAtqCVVSTP4NOxGDOF86x
BQ4So5Z7IHzVtOAO+BV7E9sxKU6ZzFkK1l5SQdXpVMY4cgg3oVArHtuMVMOX1qB/daCp9YGZlQvE
2BnvrVnao6rYD2VBRkm3rqQP/JyD754Nw8Ug1ETrEcZXsMsAt3NiOif+QzWvEYBwnhCtbLXSzDbS
iK9xvkedBveXK+s6+lsushbwiPtmffhIUZp9WFtydKtX8JjwXpY0dagcZ2YBxJ1lgbqUMx88Oths
5SX+swjSaexLKKjQdPRtIkRtLRVFxAeUFXdYi9h9PPVtTWyiirrseDH9BS+Dl1ich5Gs1/Nc4PzN
4aUZ4sFSDL46GCmAurJNOg6BugNEW/uIqK+vEcel6NCx0zgp4m5WqJqgjj7hIx05XN9C13fMDxDz
cBx6VKhopIOzHAYtdzBKsD/pXM9flIF6UAWKVB3L7zxwfAP6EgTytmGdtZamU93WGYOknjSEgu5f
nd3I8AylXFsi4tJz/6YrKIn9BYtlIp15qWWLOgevAsmqqJ+ODMYos0HxZ2MoC7HK6buIGevcvd//
4wbT68dyOc5tkJsPd6+7cZy4EuJq9ZrtAHFt+znkIVUV1N/bW7GFXhCKcJ45RUwpBBj9I/Z2Yjwg
Hrs40p6/Xg8qozH0/yg3vLIgXMJESMwq29DQBPc3LEtjuLe2DkBAqWUvy/FqZvU1x5kGTwx0m6Zy
+y1c/EeGLI2CnxUQmFCBNc780Rj33mPCcphOrbur42n+bKkn5FulBrdDKVjdMGnLb7bl5k0WFt5O
IO6zKW00Vy5tAAtHwrWSBFXalZPdKekfW7FHsSAoHtp9n57UkSxnaLUdVI2wKwTh9qyet9pQ6C+l
u2x86FVSGPjEUK1OaKFrou4ojAqplF0MxOYbMPIyg3agQ7N8Up5Y7gX8CPbYoYly535YdNk6fQsw
LtmkLe3lG+AeK8oUurwnf3HWOHFfo4wwJ1S7A3oqC69ZTlSsTmYNZLGA0S/vWHOePrGtaRFy5adY
CwD/cLcr9FUIv5s7ZHpzHhaFARCq8D1tW64IiH/uvCOVyzi/t4Y2hUvGD7l/1/lbBk0WAVnqcNpM
pA18gQEFGoyoHQ615eBcbxtFmRKdwziVOWGMlayziD+vRg61ynZO7GxZKOs8BFMVOYK+NwYMgl5u
4adjCHBGm7GUt6co5w6fzY/Dcva9xChZZhkH5YdPicbiVOO0uuLu7L6EjCFBJwOM/qNShQqB5gxZ
v9qirpyxZsFEE+BVlx5/12goNuBvulCsDJj2f6W2/+ZeAL0Ws6T4Wc9NVZJIPoOjo/oNBChUxS0O
KdbVa9gqnqDkpoKDnmcnvdSOmxcadEE8nUrc3F1nsF+SOE8CclrJMcwUBTXf10ZXEK5lMRZrXjjq
5+I6Zan+sNJNcMdesIJDoSHy6m4rIaQEphAr1nqWzHlFKMMJh7T86BLaJyPCoRcl4kSlwIFpgM7O
ZqPVZsj7tlDk5c3+gKftwwXPX7jYXf3hCwnAar86c6by5V04fl0t1V89wNEQLt4DCX9NJfDWH88S
XCckGQfQ/ND0C4wXRDT0WYvQUbERsm2PKvg1Jr7bkK0+CbRcbvaZHUCej1rz9h/KA9NG/m/TW5JB
glP9IXXFXzo0nYwp+c6s3jIsRJbFqd9Tx5XvBMliptVINRSi8aYyNxp1JPsyxwzyPImE5It8Mnuo
ssqzfNQPC6MdfHfVvDUlbW78bWHMHHO5ZNst0OVGAlW5PL4hOpv+VEBguRYhOUYEftWqSLWXEn4p
/7YWqj8PK7PALFzHT0FC1mH6rAy8VLDCWdENq5r1qm8Fxf4JhmSr2+k88zSk05TBI3EDcNzK1uEs
aqYsAMmu4TQcyhC+cO/la3QvQqrZ2bRvheEjNV4TcT+idK2McNRr6A5yYsfZJFhbPqFwBxKRpCys
vBeAbUZ63dh0LYiFRDZd2zYZT7PG0DR7HTuKpg1ipBEmDveCpQgxxwZXbxyYZh5YrgkQdovmy6wU
d0AwjmhaOszruT28dJoM8EJhGd+KDHNfTAQpMOx44IwIdehN40v6UGXZe4qX666Xn3Z5PkQAKZDk
qflKwTrj4z21XgDpylTJX3x6bCPZKQYNEJbYEZ9e2+DQTsGFFoMLnplsW96BheWkCndp6FJzWUri
HreLotNq+bkGgOYGQz/Bv9weSLXlHCogskY+EfFVtWbnnta5bnmLB5cCzz5k8ZhAYE5m9o2XrIol
niEbzHJrt5Rk9xkz4Ml9FuT7sl5RXqFbMsLuf9GgpWYTLe2j5qXYO9VyIi/QiTyHf5Rf3Mmg/4pH
E5lo2IKSBtzk/0+aS0GcJAQZRadZu8N+ogZXcq2V8k9X/Sx6j73jKMYop3UO6mYSqoQjAmU1o56z
2HabO5KFFrwkH/1twcMmiowEb/8lLBf762ATUSbZ2sMWKACQ/QhgpLrHG3TqN/E9hO0FoWuqvHuP
P6GgRr9HdTljW0vY65PSY62NvjH4Pb5bGqrYKVS20g4ALXU3P20vE8Y9OxqSxLOlVetFhF/N1G+r
mwVu2pTF6W2Olbw5noQuhFEiTsv5bSfkXrUuFCtNLeJmNSGP9IuA7o5vSYYcPK6ziDzlU3ZKLrUv
pnOZk0llY3yN0wreSbuuo1dx1xK8c50TLbCU0a4b4yiWtSw0Cg/dCw4a3UtFXTQ/FwVvrYf/6euX
tP7L8+D3INC40QiMyoX4c9mGTc80dkvH0bqI8bAqe2lEUcYMB6RmURhgvFpE+yDt87sKsqoy5mhJ
wwrCHAZnhf5YOuSqdi3dtZHekKSb54HckuDfjrJfU5md4zupsp9OWn9egdLAwJz9BrvaBNR6qfv9
sUe0wxc7vbjgLguoepjyqiJBT7nxz2yNhYp1yl5dcDO71a2ggH6eECWhIoV5VvnEeNpYRzetgele
PttjomcUvt6jl/fcws76hpzRBpTA+gCOdgEV+/MzR0Vls1P5HL+Spy9ztVLG/v4RGtB23NWTiRqJ
3hYNNfmoZ7zCFT3VtXAvHhD6aWWgXuQLQdDcp034FXqFICSxeSQ+gkcoExiDCQ/IrhTXcjC/HG9s
ZBqd/Gf77Z3GPnmJVl7NflWo52+y+siJW9+1PzmcAZFa4aNVznuJnrHuFfHDGyQEgigl7QQ6Q+QV
lbx5GZZNOLZj7OQb0Rg0zsSJHl6I8L9sYRaCT0+2jBNRYaxAI8pBuxfdXvDlVbfx7fsH9X/zEuHW
k4AmfzW/Nv+mxgI0E0UDVDMdM+k0fKSOUBBqCMamNTojIRHgpHIXd5IMww3DLmHrah7ozqkZQoau
fusy33rD2w/GHQ4ZAUA7Jfw8vfC8ZLCreqxzuHK1f3s26D1TIomQcwWNZug39hA2BeMFuYARFZow
1/QII7DqGE9xJ5wOaCpUuDocoaogDNcHa0vmMsOEGzcEVSYaWRzhk/Ulblr+lgp2Qj9AvKVansPC
SGemhM1/A3LYAkHSr+MUw0gffudYo5BUDUCnrKCKL68MXuXlfToQNEjnnAEZBnB8qDVv4Nu24sl8
bmoRqJwG6FkqFyEXxhKG/rBQyE3C74kgzfJ3iaCAtJpj694SLAQyVEUljSLFu6kUHVNekFUcaTEz
O9uDqwEFB5i8rK/iVxfIPasFttPLQ00M5IiQ04xyWzJBOPrxQubg/VNISXAwcB3JYQ0xRqUwZV4Z
XwfN7o1ktQ4fsb0ClHikqrqXbTNZLFirdfPaWgxMLtm1oExtNx5I/HORfNqEjRxfeTwzGJEUKDvp
YuIJbMwcdPuajV+3i2VurSs/t9l/Ln9xhJfAVhTe7cBdMDQWP76Gy/qmWhVfvLRoGFpTOgIIZsli
wYpb1fkPSxSUphfyyEOIpmRP3PP+kPyESkqFDqoXxNjtpiseWcYMKw0HLFYNX85sefiHatzpCjIb
p0HpL1fl4NZbGGKPfNmlEPYP9q2DpX2ANXqtCfR6WD/4/L3vW9qSVrv0l+14ckJdECuZxzs/hcUu
IAdl58fi4oFs1CnZ9Y6BFo9rjW0kpYxtnwLTEw4LwmPJpGE9FbHQsAVTDpCFfCokOf5D/hACJVmC
gitDzdbch9XN3KNrd7BqWOZ2flfyvETxgIoYKBJlfsiV25qLp0gHy5cJOwWsqfk/Yrk8y3D/5FHb
jz3IrFwqF0sUUFkTB0m8g2Q4vgUsWtqETlOKecggkBLzyJ6mtFRJuknl2rZ9I3SiU4rmE/bH6lQm
9Oro5LHNkzMoI2XxIp2Adc0pKSx4xUMmrs1jDCy5JAdM1HUTyIQ2VuMI/j/yjr8eZun3I/qb9UJM
QAuZLGNhnd+P7G6LvpdCiT+u0s7AYU8UOa0ZE2ogIILN8cd8etR6uxr+rb/JOTbYALeavL3/0z/Y
U2L/GbtzTvrpIZ/Zw72BlQan2vWxQd5+FA88kem++l/ILOo8EZdC55RX/a681QiRGSTbaLeSMe+l
txzCax/DN48mVpuIMjcsuLk0L8XDn5dTtNMzt8ZPu9ozgoLKsIniiyTLLhTOMjU5z3IAKV3/+S89
oYNW+nq2kenVvJVLjbz390ewWh6LHau9hUzGI79gJRRVU2tPxPMbb2r6RfJPkq5g0b8NawU84TSr
ZiIMXRLkivWM94x8a7ny0J5UdM9DzZUuN6idMk5NMzreDZXf+ZDSQFrYFnCr+6Ia45v6MOYH7Usd
qVAe+o1edMPSQClS9kkacpvBZZ5rgkT6GBb7Z96S2gnGPZwacw9nilnJNiml6F+AHDdisfj2QyKx
rlO2JhcmDRPs4ePP5ikCTuwo+HjO9yFydZjma5Vsqgz/HoagRGs4K8Sbrv+1TDhqNDbZXlmz1PMZ
6GAH++VsUSqoyqawGylfh7U5ZolBpyzwlpefwFTYzay8yGXMk+xDAx0lhQlj/W6dzONShZYcXpbu
PunIJgU87sdN31ndplh2rFrkzDtKEecCgfeGNYt0g9gEDiON9aNRYRbGuIefClZnF4Q12kH5enkC
4R+fMUpX1SYlOvQlrhU4bJ0K91/RXAZIYiO7GKitbrb92xRrHe0jURRLF/IOp6abIDx7KtdIYV3O
dfisFXaFa0B5QzZXcm+nhc4GyPlACzkEFZM2YP/KdylCjz10c0q9F/Qdjc1UNjwI/74muwp8QTlo
9Cb5NMLiOCWg8mUuvo4YVECeSw+b/qFM3uAuoQ+eTIMAVvZVJA+uDjFpsdVoLSLTD/QxP2qW7RxN
m4Z02ZHrTeW6knC93O83X7UNSa2ufC8mZoPaEtoXmbXmpwYsF3PxYGktsvD/Pu3/7Wr0YqyIq6mP
BwMgR+ZQjRl7Xzoff2y+SuT3ur2U9eoTKx5Ewfg9AeJMuHlLQEbiFtOna+ntdGvQbtoVQz4+I3PH
ApjYeHsSbhdF6y378TvVu5kgwTNY8OR508tQ4SKDUqRAgLLAEleJ3Xp3QsKGvfC1vsFwN59DYgHd
OI5UXmkyiS0Frw8fmb7PXAm9c4cFWWxz152MwkxaJObd5nkTvJjJ0Rb+r6YPndHHpIzZ4IHHK+9L
TPwRtANzHUJGtjeuMBUx0ljzW6RqCQiGfD1soueVCV3mT7UwKFmnqB2fOPzmFIkfVIVTG9EsdXdF
jQxMMPNuOCcDhdms09y8qlJKQANiCXUbMPj5WEWVq/8Rz4vnF7C77e/LNwtbMJYtmloxEAUtt+bn
OzfDDxMIMrC37fMyY4vAr0HTeu6khg1xesXdDc7TouqIf1sEoeCfiMjIAbZxJbFi1Q7PGOrPkFFp
IIyApLyfcRK1FMvd3QxcIvcTfiKhHswhkxGzHcD7xQ2fdkQrUPfZkdyI+vIrR7w3xxbDemOgiseT
vMedPiyfnsSn4Se1AoYVj3yVJepkr0WISfUE8J/x5kxSBxLYJXWw/piTBuatqHPKnT0Y9ioZ4Iet
UG/rbE9zGkjdFxZtd7xgWX12WSBF1AL0KK0gBJhDNAByqR5uuQ/RDt6PkpgMGK5KyKMnZaWPjtlI
nyNRe3dw1Oj16rcUdITqNPmtwoLJIDzq6235ve2hJ2wusa1KeUDtLlbsJbFc0AMri4RaNXagSK9T
u45jQCQtmsOO1DqpKci6gNlrXeHbTPAPvaakdAHRW6MM0ptIpFfmFigYDOHkGDmdaBrwuA+Xl5G/
hz11SCkg9w9LWEjaFIMfcVjLD0oa09DnTJhCpd2wWYg2iYxqRpICRHIAxnUc1P+V6RnaNrPQHnui
8oNs4Jg/nHrhF+W/bH7GZhP95U8tGSqDc8o6wCrztfT1Q4lULLBN/WuUgnp4fIMyCGMRnXzqukMc
dtFXy71BAzPnK2J2AELqMgWtG5TvIKtvU3jw1EC4lz5zhc2CpquU+fw12VCWGbT7t2zsbfDdFmgG
SNooaze/E7b49CqRaGrrxtgqvup7sgjywEP5mrUNSkoYnW6vyOIpJEqE+xBY7hMSJp1Pl4ErbYzP
UAwn3jEy4lysCFa0bvfHgHRwCCtGUmTEqbWgX+DHONBTJxNnHtUV4/1G3867BlDd84bKY21mrUF7
/iaCwmg5Wza2yZ+Ts3ZyvQd1MTdevN2pyTVwKX5LVH4aq5RQB8ECyB2ExzDKxQFJjfIeMJCYRWiD
K0UkWCnfnquu0ZJfS4W/d4qDPnG6TzA15ZyDJWjOxosk3RAN4KOPFc59C1Dz2QNUbikJsq9PhMxC
HlroHhonQNVxd0o5QygBb8KD7uvyY0TKWVEL6OM9CSchioC+WynnWhK1Uuh0EymsxAg8ZVV0T+Q2
Xm0oMJc6osZ1j8Z+j2pQaUMtWikDpL6Av3MnrXKhYH4uuy+OSXGvBdlLmWmh0+SWfiB3AOnYU9mE
b6ad6sqzMqf9IgVJ8TAT8TpZbhxXmLkk33xbPvGDF/9FMkcTXQYpNDARfSO1lrNcQScaWy1zwblD
Z+FFT77sWRhbneUwqj25PbSTdyBgN5hssdqg6h04RcF41f0eDx4c8FZNgZjQke3yGQrLHogMpav2
ltuLkTZZEthFVdaKleZ7RM4MVlZzndHOKp6anpekB7qMOmV5T0CxiixLQNZ5iB8fRcw/mrAdypv6
stdu5DXCPqVs/Skdb2LneyLINENHx+cUXLbaNSl6EzfKm8mOSIq6bzkwrEkwhFmZGQdFvBwsStU5
ddP1cYePXRrzhc0I/2BHDdvw746lliPW2vDy1HTnHqNILa4vn3ak8oKmB2cHmq2aNEawy3pcatf3
jAUKCsm8EnyRZAN1W1Vsd6vlb9P06rQU6DmiA0EgCLpF7aFa1TZkjmofcU3sPkYqNhSgHHI/0MCU
I7LNQ+9UnE7CY3WTGdcD8sn1foOw9Qav6aRtCkZTE4Rf7BDUYoCM79pC9aUO8R09YL84xcJQZPAA
2irhTDyHqEFGaluBwbkJF13jdjjk7gU058wGlRtbuimd2K2LJ2KAQM4eDsDQ5g1h/PedwInO8X6q
1eRhrxevsLnCDYyI3W/XqRvTK0DD3Oumzip2QBKFzkOekNfmLNldkcsV9/TxeFtowv7miI9YDfJT
A5OwVXCiSZ3OqyTFzK0Ua94urhaa0EqHCgIgkDOV3JrlUoJIMM15kzN/RdZ00rxXtZLm/LOVs0Rd
hwgmTBGoYvwv4rOdEdSMflu6Lm/KU4jw3pD6PR7n5PyDQTqgY5FIlZ4cQrapM9z0tYuSrBhg1nHm
gNFDmcRD8x9Y7BOcs6ryURzh9OiQpxzECUE9/WUNP+4gNCyb0p/hAewBglm/y5zlcLsFsPofSjct
xY1bWEp83FaCnlCVlfpuwbumc9KwEjInrE4pMdTvm/O9ufY3+iMBJ612F3ZxCEyjC7wmKZ92Rqxy
wvmI4tZDbsOXUP/ZEhNRMcJGh4b5VEa2s4V+ravvXJSO/r5WoaIaAiL47/7N5bC2uJCuLZCoKDDv
fjZlZR7PELrEzN4pPt6O9+Pw3EJ7FDDBfWAJYTQWyaT8XrMqXPRGkZeslTU2wX3kMeUs2COonlq+
MLgX8plpl/1pjKjsChbdHJruMpe61K4BH7fm8+TR1SXrokSuD+pNzGjiEjrkpThAo3tgKwvIa9LQ
P48L8sL6/6KGyjHDe1mrBm63GrVtAcFOOGoi2uuGKAonxThJSDKjIejZp/WbnSfpKMeWL+Kuh5oi
UYv6HF2lfyZgIZtiSAsDg3fTRDScAVnfv4LxFGQYl3e5wT1q0pb+OafV69SBuLNBcu3GHze+13qL
tBq/q+N1I8qU4nn60ICdzK3mf5ynlgdHnS5QE7HC0kdRqFvE1Kon6r2+dg38jgYHbNbxj/ivQxYM
D/Ue97N+q5bNdOB00lLQyStI3MA6o2NkQxwgheAsDi+B96HJXvC7B2sEB5ZAXwzLPVl+CCdE9lDQ
j3R+jv3SmFDtYKYGmasqrbLJ1wrkD51HTmWprLpaV7qRnsUnuyzzENeedo/lIR++vvC9YkKUNYo/
mFmUxfU9QuBB2RYwkxlP1Xx6N6y7TgHZXL30zEzP2lkb9leS3lC9Zi+vnK1IlQB0NXFlpxvEPF5V
6uwnAtMzTe4n0XxLqq8oNOTdBxV++q+JrLzNJevOW/VkJvP5/qU54aoGbEnWxn6V0A7btgapWH4m
XqhtGiRAobWRfoWTFZPVKIMAGcNEn9E/r+cacHOAZudVeLJh6od3PkNGZryPO5qtjUdJ755lWepN
sqvFyKVCPCKyYkYDioHwRXYn5Cs6Xxl0PXL2XZozIYH6p8WzgUavmzKbk7WmuUozqb/DnqzGtROt
nDIh3H+XPGKmYXDH+UW/cl1nqb94wQqTxGJ+dCQaFSwAr09VsYUn4ukOc27nUqZ9/S6vRKuG5Zy8
3bP66NKzkpytv+apwUlcof9fH6EfUNGkwQAQsGIx07EviZfV84w3RjnimGBhKvy/uyx9AoSoyFod
gMtVEtOHOvnWN7IHom3p6lqZMUqokq2l3FmAKFy1mwAuauSqH4jhTOlt7E17CROrnL6SsaVKlbPG
lvUnHVfwVpoB4Of4TV57441XBXNVRLXIOeLcdPcBUqvDJHGxN/bQBUWmQ2LXY5dGwy1ZofufTeAE
LAUX61JFJ96g1qUTVXehO/+O33L9x21PRtPpXp7g8N1sYWwq2M2/OHPe4MDwtETXyl3BUrIUHJFu
27p5Pnd9XHhsXBSURB6cEYJDRhAerrWew+FtgeWfRS9f1UeRfciH7hpZK2xOjEZjNdAEte6748iX
IxQBGlnU+3gUJGz/wSZNsmA5uwhHkOoDJ6Y85+7mJZiowSSUL0yOTlVvjHcUeF2+yy76hNc5nsrA
Y/x2BpimuiWLtFzCM3XbDulLUeUK71kc8gpaQ17RZPiKTA2taBPdrCd4M+hcZmUpS7P6kejLkeFb
z0Fjy6VEvfpP2Y6BM0JDEsg2iXolBKA/SsJeWm6It3d2AyQ4dquQnGheGGjwOk5KKbg9qQr6BXf1
uzLJsYMECv4Afwz1n8XqjRcSuvk7j473ux7JGglctIgSSqIPbxJ0iClfe3thY4md+CaRbo53vFbh
BQe5akeqio+E7cOeUCxMXcoZlm0f8LC+O9Nd9DaF8I/hQErIbLU1O3t5fPnU93J+iM/rBf96Cjy2
E3hIV+/N2tkO40LtdVFqYsCR2TV4LSAWb5EooxEtEkSAbKYftnvUN56h9h6fBGt3J2B8ifbLtKcc
oMmMsHAs/aCxsEI3T5ZwZViYenlwrchuXb4AMYmYvkJnw4eN3qzyW1YGrmAMyD641O5B1ct2Y0B6
EwRQRBQ4XQeutKXSEbSid/3m/J7wtRHwU3+9DmqneybQdSJ7AK3stCVDpaHKeobkTE7taE/+ZiTf
BcrHxM6fNhH/SlEdrpQ5ypjtMaMOCUTInoLV++6AUORIFHdzOJ3zf575pKLfu4qz4aMKCvZAoRSO
iuwOUK5DjdDHe6Tglkze95W1kLJyoXB6FrrEJLILVg2y9bSwW0k0LpxPiC6qwmqi8EgFChiunNHA
cHGsCmHrEmg9jZwDdzCe+3Jiv/hXWEYo+UIkL8x4nvbJL2oX/4mMFTWSdL6LpvjMfMbmO/SbTWVT
bJ91j4Az4XCmQwcmgpdGIovfx72sPHDc/MZzrPywiOmPnDyhH77+miBw2j+VDmpK2m+vW3ZdDxZS
C6cwCcLVsSPNG2Zakx9Zl/W1ROVN+9tBnOsYKFAasJd7vSLF/MMwgP38ERRNWzC7bCHKif12sCyN
kIPd3uyQHFzoE3/LOZvn4NpHn3eR9Z9b2USbxL4TcQM4dIYBG0EPmpG0oWGUYHY4V6Yl2pOLPZMY
u29/JrX7EVA/ytdDWc0FKCgBlAXQGrXUOLp+Y1lJD7iZITMLYoxR3lhqb4fr+3UwMWy+lBVxpyeI
qlUVJO9A8S5m0HOnulu3OVxJ6TEb+sJ6g5UXkNHdhgqJbyMaBHrbfRFnV0uaXphRuHrsLm+MY5dA
phJ5ersUDnTMZJCCS782kbVNecNW8yx34afuSctcFWcztIJVc50zyxJQEDtUsXc4KrmdE17ImFNO
hKXWcwq1lvb7VNmFYaYfazIWSUeVByXT09MrpNR3+glYOQkx6uwh5mc3gT1sUm99kMRh2PXxWbEG
+l/STc6vb1qNrctdpQPnY2kd7D+XJ0fz3y/23ReXtmWlCcqL7HeQff2/90re6M8KwmrHqrUa78di
/ErznWby9IzMJ7/Z6W9cp6DDXJun9h78vsadNu9QoNt6y6EKSGwNWWflgCvVjg5DIezZUAR6O14x
ZeWv9hz10EZ8breHUKDfNDBnynB61KelpS703Nu4Rgtl6cVyotKqdW1uxqkAhQI1u4RTSimsReD4
7mwH9Xw9DBdKX+52RXPksNjoV0+RFP4ZhHlh5YHt62UaiGvw916EKcoyGgZemENLrarrEveeson1
2vfkjIzrGcJSy2mpto/Rz/pwW8IlkrpHA3xH7TPnbkAVHo3lFK8GFMSnsuCvVDAKEWv2W5xQ7vAS
YuLIst6spj4RAFeWIxLtQFaCQ8i9NqXExqR0o5m/1dGxTuaftzbKpmBaN+u//vtfTkwrd+gYJHzd
lYHxqK+49CRSkJVNG/LEuBebEaFm+zLpVimsELARrhQ69XHcBRmFvT0Wxc55SJKzdhUpKVRIgHUk
eqimYfAXzN92Xu6vcKQn6r0/wdv8NpqSm4BPOBryG65ZdPV4I/TLNnDKzzzsabExCDCAqo6teEfC
xdUtP5x8jRPJ1knzRG/458mKAw5b71hAAGly/Rh/6WDE5LN8aBBnXpd6PFi7iAYeTWFMb/ojfEIf
+mJAvXivI6zMTqVKHUGbkYP/5cvMd9cMCuZeTwBvoxY7vp8+za/bTq8R97pH4Dp4gdcinNuBQJze
SZs0JbPl+RqXcotL/9x2OkhNX1PN+kiSjXx5I5DXm3Jdv2wqZyrpyFdAci8CixmXnnVLR82tWCMa
4gIOa5p8j4QTAaK97XApXLvhIoMAO55ahd6J1WnBkeKZoM3bkyfpinRX7JdsBpre/nQyKkOq4YxJ
vihCK9LMC6Mm7kH65RgpNZUGhG6jwU0SFB+TEg6Axk73EgU0tz9QhXvR7iQ5MXueeuUzq91kzWBY
UKYLDly9mopWEI+NwKU9KGKpftgPx6a68RWEQtPR9ZEobjbNm4dmljrr2prR/lCpiAsLvUJU2XDr
aNF6rit+cefXo9lTdM1wmk6bAUUy2cTJ09Q5mDPDR1H+mvC0XIyELR2PuNomWrE4E5SsCxWwAE1C
o/4MnNt5ZsUIw9UnP1UPWQ54c1TcYwVjlGzhIDnRu927Zr8R111L2yOiTOCuyBoRep4jxC4pKyXZ
WW9EIYjr8HEejtwjDdLnYW1Yt9ts//BxGZAb7Qfrt36ia844GZHixvpV3GNS9Fm5ETitK1ldO8rr
e9Yi56ZNnXpvn57pwc8kdjCepHyX6lj7+TOZzzzYpTzDz/l/K3AalONCuq/Mjuhg8DYrYkxiSHZT
RXf0Kj4muavEgPPk3GkTxm+QFt/BMS4EBc18Yi0vmEmLpDLxs+87PMv2BxooLBfPY2XLZmdjx7Pq
5jZi5qGKYzaeOWh+fZVb5zj5L8Sr7ckF3cpHv9gdmA3EtBq4W0u95GyziNOvQyIBxZSPFvVJhoWl
LdgC2jSSQtZh33KSrZQ8lvwW2oVZSnbf0mADXVxzIwqirba24tk9tiVDDJunAWwbS/9LRCRnMsDf
c0isHVfpWoZjTsZgacZcNeQPcm8d1oDGBUTG3+QhdEag1LXSvfdm/b4/h3gcwaUGwdDUtZR6qUCk
cj39dW9N8sY3yU9TQ8LlbBiQMnOZ3Dg1CI+zvwSoQvTJ8hZk2byLyvQq3wvFT0rc3myLmV7/HMYG
iRU/TG3VaG1Zdrw3V3XgFp+Lh6YYk1Z2DC97ef5l5ZcrzM+hUxXg6ZJA1L5UCaPO5OxzqYi9je3P
lqxoDAUD96e2Cr91kGimd0vi0BjLn8IDeIOkn79dPb59Vj9hiU+GEbxxOqKnGXgT7y41DSp2Fa9P
sEanIAv2v2XXbB3YBQH98jGPFdLyaFowEBq23j9YnY4EpGu+jI9EFmgJnnNKo7g0bPAaYNA2cTfG
9hq1I1gSblNBW1U0IJRb7wSB5EqqxepgW44U6qk0q07DoSbod2beb853/yN1iDi/rWP1QwWnIEP1
OOk8RO86Ofsd3ZU7HZd39Mz+EtaCiohzbTcDyTORpxxPkc3bOp8OYRv6nEeHiJjJMW8xikIYhieA
Lxt/Pu3SLR7pzZ8VjQxQqQQqRC1OUMmb+z2Zyp52ns9lioBadKehJ9qZgVQ1+VPXMDW4rsRuQK3V
hDr2l8gYoFutB/3H+9NtMK0lHZu1LdrY2gG2pa89y4uvSyXlBWgJrjXleMSizrM1wHgmQPZ/70Ut
Qtob3YlCOatgRykWLBEGkHoEVb8QNCBUuWYnHo8hWpTuQF8tJUNP379iFgYpdiK6IzXZGZV4Y/TW
Ru0+GelkSOILmSTUFORBOl6469MdPyNshkf4oSQRnU2Z5FGSXd/tV2tkZNSyGz0G/8WfbifQJAx/
igDCVcr6fKL2z+AAslLFIY9Sg89qN3nMPEEJd4+eAJFfmc6s9P2xMCu6wCH9TI7KRbGepRG9xOHf
4hDaqvbqZWwE5Di/d9+89Y+J6T5+vrPOwio2Wx2tWZKK15kzudAqYZ9PR284FNDEOHBjpLepbHLo
6M57uC/eB12tvizSrrCKOca4karMi+NnV6DyqAnzen8t8heFplDzCBX9pUENADYvLGeHLwqsMAqv
ai3GeaIW31f79typBjJ3bM4KAVKTYX2oSoETHhKdv52GTgwww8ggJ22cTHieNJepowbCkcorneGG
h/UHoVdgJBggpgOpC4GqxfD2MYOs/ff9gHNc9qDv3yTvTzGYTFRLt4Hdjm2qeKGOHOJEcLh6KnyJ
JR5M45P10qmLmseQd3VhJqwJa08uITqhEwhuWMboNZm6UQWCSPhTnhaGWzYU3qypaCXfkbE7tl/t
3ZdEIQVhc6rXmI6iYwmcPr3WVh0fq2MmujiKk+rKVMRAgseFGf1srDlm7fEtiEdCbAlCFb8mVsQd
UNl7Kd27u4Am50E5G8ESe1pBiUfsvqeDGBiHQAupg/xZ5R0UQNYbUevz0KW1fEe64rFfxrtlJjcM
NCfUh4UV60auBpOaKzP47+DfqmixqjFrC9W2GHjmAm02zs8rfsBRTqDlDK+zXDt4fJKwRHKsYkPf
leUPCRiv5pPozzzScZGXBZk+b5BUXu7x5JqcPXq1JUNXukMtK8iyY4rNnascXItnXbxCVgGDC2pF
L2WZxhZzcllc4v7M9AhF3qmkEhVnkPMxOGD5uHFMUpgqRHp2wSLvmEBuWwed0HVgT0kH8ZuFjWfB
M8+o4U83PrvVqPyr7ZV3FTlhcc/D/S0m9b8krf/4PRyUJ+MGBk557uzoXdwL9ijKnVNO7vn74HrS
nruKZHEY811ACBKZKqvlbdTUDPfmLHfz3bcH+97iP+qJ4aSR4gbjaBFxKTWPNs2yhFSMbrkgrRGw
cGtjASzRzRVCoGrNor4k09mOnB0flcjBAas5V1cUG8YVYySLjwU9zhZCiOs5C+WQA2ukSMCEaUMt
z8Uqd2I/ADS5daW9Mcpk5/H6NVN/QP7pgWBjLc/6Q7WQ46fzjPXVHgM1Ucgey5hRYaAW/jvK/c65
MEwsdqYI7MZXiwncHVMWd5CX94lUxKBV+BevGfF8Ts3oFXPkYFOTDkiu8vHVUn80KUuzxFyPImXZ
v6lC3yDYVB2x4V4cf9Z4ZMy2Lj/MyNJMWLI0LMoUhM2MfEOK/pAF6d6HEiw8Mjlv2lFFe8mIucDn
uyHU3W+o0J2LkqyZ1uONuFDYoGSIG8HFEn2BT1RTIP0q7y0XH07iPSE7tDedoi8tirS0XZXFRdwe
D4aS5V3FRAogQvoq1zu5ixvHDO8Fa5fsx2mYaMOs5zkrhYDusHydgxvJVzqd+f+iR9XantIDpxwO
L6JVs19GIBMOE4Z45mVqkrHWQBhmRTRQqTiW6Z1oiqtXVOibCSlbd0nx4C8/cEHm8jV773IfiB2N
L7URzUGae3ybg6hA+onQYltCVsw8NMzRECj6hztK1QELyUpopKLoTDtToZatHcMJlc4kbgzVHkP9
Bu865/YfYg/hjnTezBLvVTehNjc5F/HVn7cs6dNYDw59WWMwZqFIaXoHHhQbGE0uFNflIaqyqbSo
Zk3NKZP3OwjPxFM0SovbdPzcm0mw0WRqNaBmE0BKX8ftLY+qCgxBLIdAMpBwzfZlJA8AGYeZWoAJ
9Pv39iAxzERbARPLjfE6A2g9VJHRk46psi2Hm6QKjkdxDAi+1T0iDUysW+ac+ZA6qc/9+hrRNIQA
FpZcJAnkHk5IN/XhiXlxZQebU9MP3FHDXjexf1FhBydCLy8SwzD3vu7u/X+wabx0dxpeDTNytBVS
oRwaohjuqbWpX7b35Qukffhohn6EhNvsdzT4UHjuh0PAx/pz45ozRFTbEKjzOvu4JNVA468CwuXn
td/eAMmC5lhsNUZ/acwaS0OiyV+E9e6zEdcKC6aPXbtKjDW/43pocKfJP83tW9Iyi10EnFznr+Il
MdQQQwmQj2V4QtyFadz9rgE8Xb3ShMO4p+7kUUNvFkmxUPoG00GrjtEkUO/M09wHaiIs1aC31SOy
1WUzLah4dOjfJG84ncAH50fl/02ux0Tjv95ySthNNkBmM/HPMwJzZuU9P4GDnuMkiEy+aSTFix+0
5TxjAZzmQBxn+KCRGilvATY2hLMKuUT5gY9vKGeE6FEjLb5gwKDKWwAbnaQKceY1z2Fy8E4Y9TuV
hmREmUyxUKn1VmPNhLB0ie719pIV3Jkha2g20P12FJ342FX92aiBdVpMxOk1lZrb6UyWsaBuZoUK
LIx3usfZRP6eL+zWef4f6a5wOtt48VX9dPXtzv9WF17rOyQ9xNlphL7ufHe6J3OWavn5IIPgOYkv
HPEfcKONh7V76Fl2ALnuc1oMeyEFW7xnHScloNQ880Y0CWqDT3lSfrorgWCi1ZTIVjTZ7dH3ksKT
9fvdvTfzgzM6Dp67OFupebOQ3eLO+ncZAH9hdZeztTCSnXxoIgvBDP8Z1x3nqD3aFVw59+QnKH7B
tZ4njoiRiLCJAbHxjt5+RRY8Bd5qv1Y3HmN2hkufa2O2kFLQ09UfWU5lfL/DCTQ4va1WW4UUwNJi
xLYnWNd3kfeGZI9RU/IMGzNrMbUsihB2yPJ21K+LifWcxBbGidg2uQFmL5fxSJlPsytOHdJSqFTp
iQjdTfz5S/y6dlzGF0D4h1e5M36OxTb7BUDmRDAl0SX0UJwuzvjr/TPI+sxHtMALuaQcd0oQOxJ3
nivjRSsOHssWge+vyPmZJJA4SFg1xs8CJaacT3t3GNjGJPKjVz+s5TpTpKZsqNdlz0vb78AXAQK2
mOaQUmwQcjsdYpsVWpu/vyixLXXpfz0HWWVKJBQqY7OAxz702CTqZD/aFxTL7qjWbKUjaRTQpWXb
OMIaROmYwyXEtwJGGuHfU4xINqvS/HWZbbctQ4ADF0K4tPnQvpOOmav8LnHF6dD5v6+bn+vNUy04
B/Dd6Bc4vrU+iZotg/Tx4+JI+bivNJFH2MHFxqIdIVVRf0mQrueM1Kntj66BtimPXHwSpQuXma2i
cGcBkN71vln/ZUYVZuA7bM31A1WiHWyB/PBqZnW6H7VgQME8J+0M4yy8gnv/Ld87QN0qJtopeK56
+wbI5jPui1IcRlsKDGyco3yN9iQZC8LVkX2wAOeRQzBaxVJlbHx13gk97t+YARxOb0NSSdYPqnJN
FP6jFKZGNhcmH04hgRGyKlbqxYwLlrzHgz1wa/6JgRDYSgShos+PiqqWPbHmfKCkzWEZkd133Z+5
ONc5SzYgBGxk1cMlu38SDuF/bum0Q1KkuWLCFun2QXRpFGKZBNpc28ZW52epNPijccdsot4UQdlJ
XqYknu7HiEwQsafBonJvQGh3lHutw0r8vnLj0Tmb/QXougDh4Zp7q4l2UTf4xCQmFmPxMNmidW2n
OG1l0dcgtDRdEN8nZiNTRgT0hVmlfwKa6Iq7OWfb4iRkTF9dkHw8prOJMmwBEJhEfYsl3F4NHSEt
JWN81xGiEkJrHZR6yDYeoMHSvv1H1ZzOIdZpYlXBYF1Q4coRmiZLD5hbpO3byXYyuXDmg1lcJ2Ez
YoOQNBEq68448+c/TKbsopb5LwT9yIqA/9xnJePPDk/RrMT7YKZtoI+x2/cfOzrCNSGTUSO5YG9L
60VcryuBIr+ugFDjAP9KZhKnHWlBR1oqILkRtWbwX8p1WT7+LVRNow9GqxymjiK/f+7XYBNYePQ+
0F2NSeocZgqf23f1cX0pu0+wlQ/Nl7iuzypiVfqKcxqveyTY/C7xcNTHd0wvCl9PGl+61WR5PEF0
WUUYIKrhG02sqJlGGEL8L78Trze/5wulZRHx05RKj2Ep3wh5NVhOUpd6zxPHhuhem+M9T/iaw1kP
QJNUFfOMt7iV3+FVJfEvuaoAbA93p13ni5C7bo2IPPaqRQYMve90xBSOiSInjZkhECuUm8smI+hP
i9z+pQPsQLMZDIgeK0k1FwWtaKQUGCVYi95eViURhy6MS4CPwVglUm5JKPHR3xDPE/kfpcq2hmgu
SmmoyYQEkwyU+dnKmfpcvEFxuKFCfD1W3cjy5v7/M9USjmHaa7erSgk+HnqijfrfUcrhLiedrq5/
6HfExOVbd81P2lCRjMwnofJzlHpegs+RkZolCUO6PD5F1CdL82Hym7jN7iKHcu82j0pSxBgg82rv
MehclhFrlV/w/Rm9YyXD4jqZD0XX25yENXOG4zoiqd17MMCg/3KA7qjKMuNh35iszDbMHUoGYDso
Q3yZ7S5R0gsnwqKJUDjJIDqbojmEXjOPPdq22IwZy6E+RfyCemkWj5Saw1/DeElPzPiFA8+SB7Ux
yvLDWjcPzPMaXdC2dujeAW6NrtXgbupwb0SDpaojJn4Bb73PLxFvohyf0vAwJrXuTFBm7hB6ZTX9
HdXfdWbybs58UWj8NUuFPJsvsIkEbMcR6aOHzoVkLsp92esAYat7OY8kROQS7mD4nlr8/BdBRcqN
OUqVClZFLKDjs4gM0g2CnB5VH4yztesU0LExhKTWIA034EoObf7cs9+c0H55UneuuzkY+7akaadJ
ewvp44hXKLLRn8qbScStETTuqXbdxZ+mOTP3CcaREjnHQ4C+QeksCkzXvwQp4tsSQN15NM+ArQ5P
KRmJot1O//wWIlhq1BhDgRf+afzoLwVLua5cm9YPVVaf+LVrG73iy3bp6pK3D6y0FP2KQwjc/GYj
shw1ngqzrtfbvtmtpJTid95XmJTftbBhv8urp7k1M0bAVchuxe3TUkyDItm6bTvmMT3NOEepcL1T
oBnU2cUG95+cGJ/Mo3SJYbCChY1vXWZD2kO6h8cOuud7pMjEssQwE976ItQo+aCyJJtncZA4/mKI
LEjg5n4fJ51n4oGtE+i8JoixpVdWtyfQ32lSnkZAfA0ztU82usdFAPYblGcJtVtmNExcn6hqzigs
zCPky++T4HyLw8uC1AqoMnJmucXdQLhV87r4sjKDV1HfUV5PEBTq5fsvI28PEruMLLdkdzUg55Af
s9nPDNmR9/nmxoJpSYuhDAnJL2ON9pABPCHxabmBzbilqbB7JaeGR781b5fC8cIyRU6OaW0QJLa8
+jMBzfV4NOY55Cioqj3XrHC0d/TpdJpJ6gA388SSd+XlcnNc7SuD0/BQ2kh73pSqPgwmMMcKfu2H
V8UPGCBzGyBc0RSthYi+IAl4cLjo32n0illbOH/9qkYoFNbWv8C4HhALj0XwWObvjc2gidwqLQ4m
wMQXzb+ztgORj6FcBCoZPrEeGOIU64YyRxp0ro92PTTbWgP9PTjj2qSSgoewKUQZaH4B/9RzMKkY
y1dSE+h86Np7SzA9/9vaC+4juctoDuozBCFBP00qobNam6mimWPtqoWjq+JdIUgf5ESdh/bHl/ER
S4dqQ2lUIzD45muq7AWXzpOhw/VW9WutuKCOZbax+jHqP7REpw6rMCF4Q7SFNY8PnZXJWgR1IwPP
fZ+lRD1gQiLa0aYV3q8iPpMm2exLL78icE4hoKoLeVcSuV0EY73+5Ed4pb8w39iUHVCMu88YfBNs
PU7u1yTBgSY/zYqjZr/EacspHZG8yhJIiRc8cS1kEWOI3pEg6lLmmI1CQkLrjbHJamSEPO8IEi+U
UUygRw2j+Rw4WnyA7xAIYIQwtcydyZiFTUc51fdB7YZjelp9szXuZf+Fu4mTBhnoAK9Y6Umsa0m0
ZCRF0OoFQY21t0KvVRe06YZKMsSUBTqEtsbXQHuEzpU19d2ZvSLIwaBvr7byJSX1emRv0Zjhg5jm
ho5BRM4q1zHoX9RFt/SojQaIqElYcSXbNqwuVymJXuezXboGe6LXX2JtQkUvuM4ew8hq1LG9VZkG
v01wgQDEiWiTzTApNHBFDjayGaK5jVbd4PPfB6SGTceYZ2PDJfGnmkxB5u79A1nwWu/EfHPyJnRf
CLsEM7LriCmzgC/kiRPnh6k60K2mu2jIU5oe8qx+iPNna+J9mI35w/uzvJI9bPkGQB6URa2VL5v3
hPCAC64GGQIBmGLNj+IkrIO26Py5nSP+6i1atb2lYj4K8ik3rU+r2IzLz996iiWzS7gxTjgo1+SI
k2Lz27aTK41SR2kAKaxRSAGRw9DF28dwT6XPpyrjmQgcfAbLU4d2w2E/XV7A7mjlh6/5UWqvv3db
AcTwzDsM87LiPDIOgng+ab6SyAQ/KQHw1wHnTmEC3r93aVnD5KZ2Re0l2sNzyndF90No2yusAQ3p
etfbGSCe+qdzKZvn+a8T/brgW3itpp6GRkskoMCAQ2ED8vcvKB7RMUj0zEB8koCroq83ZR5iJ8c5
GVxhZ0u0quuNvTqY+K6DtZgDX3yI9cVCQbijwsdXIPuPI9GTYhMqH59Sk+r56Kgr9a/m2b3WgEhS
6dgPy8lnkP8d9TiuihYQTpcW5iKk+FNQVRFu9eTpwAy4KxkrfY2d7HMDOjLPme8kvRa8+HShI7ox
XUn+JTZTd0pbGb8VBkiav82uf51m9YXkusNCHtmEV3dh70N0U+cYrV0b3HU2yUieqiSYL9WYM6f9
lJDH7SJSIzPSycHxLusjW0uup7jbiiFMJ+fBHveFZ5qld30235z7ekgER2/4oON1mL+u884kxasn
8mkKXbqVZ/NE3EtGdou9LUMC01LlQ4uvZlnDAZtRbk8/w1ggS9kK3TIms3TF2e/paerdMTHK6Sjp
jovPtOuNy3BgloxLKAC58T1gQxbNuCn9uHRGMz9rvHOkzjSl869QiQ0i1E6sezyHzj4Bc1mEOgfy
jIpHi42UdpNx6BVR4e45GQMaktntaGso6nRP2lNem4ADMcQorSKwMtiu4FgH5E9md8n9UcoV6/X1
vKCEcPYO9/irAf0IhradNSGYgvmAiNwQXUSEZO0dF9wZ61hLwCbth3/rU+U6JQGyI5jfR3Frm8Sq
doC++8lW2nPx4TGU8Dj3t2t5j5r0PhjzMlAgsUju8AKhyHO8HHRdO7ddryG5hoCmrIFo+8h79osJ
OlNxnOpKZ+pGuDiUQoB/isi9zdOLWlkgaP0C5ygBSqtNuBDonBE+v+M3kSDgjnKJeWJYkaHdjoF/
G02Mw6xBbOWmMi+7EJjtFXavfQhDD3mrs/3mI8wrmWMaR8dwilT1OBYRyvNURdU49aC3hilyd2D6
Ikn6UbM7J3Ya5r8KrvUX1O5BOh8wXAxfUEwSKgbcwsD9BXt0UDAZQtYLxm2SIHG63WSKBFyiC1n4
7LI99LezZ8j+X2VdxbZaL6Tg74VKwsDBoqKJ1XwLxEsSec9hRFj7Tz/8V/Ez9RuVHosDslDIeU57
0Csetp70h6/Dm6GrphHAWUDYaXYCdKQCOUnULXEz8JqLqSAHg5ipoJ0schsGNcsJkcNgMzLi67kQ
bK3i/gqOsx6uGUMOFmlaqfHDRDghPYh5dSQIoXA9dciiN6QRD+1s1Iu9CsbCneVMjZp6B+MQ7KIv
a44hGYuwCQP108cekSmhUG4vxQoxaDuiawcZEChb10Z5xiBZOSRJeShZFHJleL55hUexJri4MIHq
bVhzSsye8E5JDtlFAGfz3lfwjmQO4NzIc+5b3W2rX6DbG0N7Jms8LntdHQSvPwq/9Jt22MTGiRuO
HgFY94Ep8EFwh7VAZQw+CKatZWQ35k7ULh2qUTxj6Moi739mx/1a171QEQkVXujl2opF7iQGQjhE
8IeQH9y5NikuzElUSLlAlw/3h69NRRB2QTOdx9k2BxfN/giMoekkZnfQO15LTW6KrBMBOevYAwH+
NJxCLmQKAtyAdS8F25c4p8D6XgwK5XeStbhA0kIzVclAuq2sX1/cxSRAl95ai2XFskNLrwVoWwOs
PK6PJrXkid1XErmj+6GuiKUjrs6JF6dLjpu4SxgPrGg2b/+SVvilKwTB9duxIMvXHd9TCJlBBdKV
Hk2uuvypH+IrUGnUtjtK5jwLpClsUhMIRc1nSKgTjnlbbAcI2FPGmC/jqpjiI11s7WE2qo16fisW
xTAIlxLLZiO/O+ERpobfXDeWo4olq4nMbwqJQj/RFwHmcoe7lzRnrIJC4Y9H2dzbJFSuaMRAHMef
vxeRqEiBeNUoIbk0gfsHgIdQTH6Z1C5EgXNvYmN3V+dODWKYMSKJsc0b58nRtuHwV5g53e31ZbWp
nHdQiLh/aPps4j22cgZo7BP7e1FR2C1DsCzgfVdyCgq0vx+4KpaVpYW3lOn2amFX6yAZ7hV2QkGa
V2+xA9/Onk4y/Ry95F1Op1mh1qr3SeNJtT1/XS4ez915U6qkeIL8pru+L7m4itrKyShxIDxP/Qta
FDyDvGUmEBwnX7YUASqNfbYBY4l9zi0osic+1lsInUfWd6EJ1sYb/hFL6Ft2MKBoBVxjrAyMJ8qo
zkbtwvE3Kfcdwrwphs61a9G2TWqInxJphvXLx8qr7eD5BXXj/HK7hHUSvT1TUCPpXgxJLklU7Kr2
dPSYx9VnaJ6q0nPDN++nfax4B63FZrJVKPUygUEgYI2U74jFiyw0EkcniZ6s8yiNfmMc3FB7fVCK
dBo6fi6LETGyGZ4bmPBmRnB5QkpHrqUinlymoG1hvHYiNbPx4sAazCM5vM3fRkPQ/95FvKq/RKch
KEh/RvPlUpb3drGjSUt3d5qsmK+H7/Pke3RwyGmy1PhI2PZBFFpd/ypmV74F09q3So5HatNuys0/
48v++I2+Ha/xNT6Qm7olKk9R2F0TbxdwYKnyUzQWRbgEhCAlTOrNgO30K/p9MFOjKNHbvmw855ol
QVcm1pEzi2Rg2Ce/wmNSIRJ03EZAEEE1hzFNNmwrN4Lh++NVcVVCbS2jIgM6BfV/V9FqaKQkZmSj
2ddnqNIgaFiSiWHHOrb2gy1v5H3OpRJ4nOR4P9AT7vqM797buZ8ArhdfAW7TRFc0H1QEd9tIgOqS
cqU0E9qtGF/zvXS+J3RS4IcVh3fsBI1sT/Bkm28tkCAHOOBf8U8sSvJC9cbjPlDK2YJXvYd+hmxB
PJxmpJl6SFugJ5qcBzVYKEkfGO+l0Yq5D+2+eyusLLXl0tEACtZrgbiP+XhU05YpN0S0gxV2ifOT
lZoPbF1ev6c+Y2DDwOQyjKFqxlpJUdZO27w1wzNHlmkHQsEwADmParw8M0uonE7QjiXxBBoykiZq
icYF9js3TonkbDOw+GvhbjJ7ypyTQ/xv+dgQYkzDREgwWXBWUQit7g6iF/rTkj3hpYXsYcA83G2j
Qo6uEJcVFjUEngdSSc+spGxN/L1o6UqpOVgJ+9ZThQ5xURIp0cBb+8grOaGfEcykUxObNsocW7Nt
INTzsbQStHxrB3K2z8bafza2DobaL+xerG48PbP8SnpBVxOG3CoEnlQr+3nntZuMyTkbUJoykdZw
pPq723/QLglcVg7NwhF/HTEl10gfjOi7Z04x3Pg7LzjCoDxbVRDhE9TX+AAKvPzNaNwfy1iJqC1e
uuazKxlzBCFoyE6So1vxReOhszNdHWD42h1qWoKa7Srol36Enm8WzTs1nEF97DCVt2oxWp9g3mmb
omEo3c04artfJH+tuVb2ZtSrlvsl/DuWWB4YvcG/K6nUCA4esY7ren8vSw08kp2odXllp85n9NzH
a37fRabdF9UpixAWAOSGc547sAZ88Snmd3SDQBw3k2RrZbMIiCT1KAVp+LEVyyk0Q0qRxwMzvem+
mZ+cV2hjKAqi72I0s8fXAof+y1OKyrlTIz2ysd1xXYMEwSlu1apuFDmd0QdxvZSyJI3I2yra7hwd
ko+hd9JGwegAC1q4ATG9s8rYTrOzufA2xkqZB+aJpYlnX2CoMGw9i8980dscQhBOe+5LF6VXfSgs
Iwz/LblWf/Ove6JnYkjdxzK6It0b1nBMeRZy5j+c959xJIvi6Y6WxYgBUsAx7ED9c8PkSgMnDtWs
dCRygkvvb2t5wgHMM+mzajASm7ihvKXv4wcN5xnV4hK+Lxw7KAne0mXKZ0qvNlKQPQPDVzxfXadn
+d+eGpcy4AcV7G2vrXpettNHtg5hQxsHCOohjIFd2W6GE1iyyIqola/AHFrR3rrKEMbFqTrP2HYq
HPK3fKI617T++d1uEZgHFj/4x9yOqK81SFe3JMcl2tWs08jA3Y7NkatXZd0QGzyiumTd+7b6ur7k
LWkALP+3OiKMNRgRaLsn2OBOMnvi/RaT3UC9Qs/AqvcyR3YEOVLvWKOIq4FQXEvvTekZhZ1DSSvT
KuSGxtBzTFqmQpNXK2D/TUjqnWbcs1Un7ToTHsT47OMxaH5sCjMXvNIIEccV4uf3xLcRbQwhUJhB
viBhEv3zRBmKfaPW8L9PqvNPq6JssOLq5o2aeiXqpG2F7SGanI4Ic4R/pbjRUrwAs5Jnh7jVe9rS
cA5Z/nYy17JLuh1QQkmuB6nu9IM8Xcwa4T5YeHwqkzk6p+a3NSFCkBmnN9jgeaicVgIwYLQs3RLv
RuYFHyAXNNfzFJG/NhzdS6sjNfW7Q+t5xYTO0jwYkHYbxBkG47nBbRvaISBec1ySVvec7cZMLJFT
QTReVNdEEWsZ9Vgtdx2zAACRCEXO+iWixwQywfCgfenBbRZJJ6CjsqJ3EpbEAUjMnXOQ6IpB/7EM
bB/pElKp2Lw+GZK6+9V1YRQ9XmIH4ILpyNWDf8jXqwPjr4B5TYQ3MsaJXuNGglx1TFse7dZpd8Ju
z6VtChbKLqzsIEsxpk01ky/zav1EABp6v8kWj9phxm2dBNYmZ0nrdYWWOmOXdhLuXnohH66iMz56
lK8deA1Vh+tfhQz819STyton4qszPuFP64ejGt8Zf8uzfL/Uub9Qtnly0pX9JiMTKNooOewqywM0
V/kQNohrX49EKuEzxpcppzZ6MDal0eFEwPCJC0ETOIZr0SaeKX3M9QSRJGC7tHDekcSLms1LszbP
lTg6whzL5OqJ8m5EFlzhwMHwyxhUOwvgTB5m9Q+Io3lAAlBKpxefESv5fjE8tSLmmDX8mRMVqfqm
CJSWQeDdmK+5cWTGfsxH/3EuJ1SuXksDem+3BDXCLjUlt3oMZ1oMSV3HEoIkSlxsL5o6Hk/w3juD
85mWgLoGchjUEpf7vGB9Vx8Wsy1ZfWrMfW/g+G2zmhlCKuV+OeSnCsTJqi4649gCjEXKdzn6Y8jr
AtDoCYswpBbgrDA3pTLZTEG8CEigEnwd+Y+HOXKPAhD1k2Gay27rwUrDQ2kqF55OhdKx1V/Sedlc
U9SnjgzLcfbUuH9mn4jz8DJc/eSHdUgr7+0is9Kp27BxzNIBQJlMX14kJdjQOABjNW+XYmtpbPOb
TV65/i7ZTRf34Ua+WJ2Ra3WqQq8zNjVVCr/jTx9nY1WyalDa3oGruykVBz6CLfsFK0Dr6tTJzroZ
WcQ7p6rAdZbrDzlfJBn952yLVJjHhhcCniMb1ytU31HElf9n86c+F1ZNt4G3zItkwKJMk5G20WVF
p854+54ynOM88nQbWRrCVGEJavecd9vLjkNfiPYY6jXRWh9Lb0XZeusFQSX9uXu3DCzhrl4kgQMf
bVCXnTihw2OwC5LOCecQYIXyRur6bju14+dHi7Ifb8ewyx9k2bKvbxoGjZ4jd919yWMe0Fwe2o5K
70dgHvAJHMj+F4W40wnK70ytYKZwsZjAnGB0TZ04b5bx2LJCGolXSnNTFLS0sRD/UG92eHj1c70O
4eTQv1OF/G9Q1ZMO3csYbxgjoZfUorIPieaAhaX0z8sxY+lPnIezS+g5wQCNq+SYkmwSEB4xWibR
Y3s3ozcL3rYLT3RC2Z5jPHx4iek+KY8/kUhOSwpW8tg+iGTLiaJWyG4rX4ssnb5gyf7nf6fhG21P
0rYYiVnyeA1zuqV5/g/+pbbV859T5faTPfzgjLZW5CcDOwzb1icisEDRG13qBXwpev8Hd5XsL/db
YvABfvAJ3EwSxs2TGqGIaQGpI5kl0YcgM6VbJUFzOiRGEGhrneqi1F14ic64sb9f+WSmZi5mCHSM
f6Bqd3x8uTLzEavIGhSHtPtpcEfiiQaLwccKXWt13sK0axYY/Di0iFTzl4jo31uCRgMB650WnFbo
UzMnBe46jNrzwSrfqagV1HvWJNbFYes3EKFDc9JmvEyEUgGeBiagqwT6JUmLbXWDE0SMhsWPdB1t
5ZT8XXErRRBitwmz+wF1XP52zmqiQJvE9qsxYWFr+dgniJJl+U7elZsa45QqVO7dRE9v4SSHwUtT
5376t+kCi6ax3kcwXvc6mGcmJ7OLteZw0HqHILQtY1QwWWD8RlhWjJZScbSQUfIhlUkda3fZGE0+
zoh2h/48i/fePFCuuIyfQb/pDm7s4l8jiIX9oXmrx+KXV0oZf1moB1io1NFGBN2/moFVu6RqaR7w
3YFlfgl7YoIUgTGwcOod9Wgc6HDunIkf31yos9qIOQsBLzRI/OQsDChxpEbx22iATiFmV1wDKxLr
rpL0yl5CWVsq1O88lxHoDQPECUZuvGctQ/nmeZT/LGL1BSpizYR/YTcWF7RS8bPyW575ya+EwwAc
G9u2q29ZHJl7breZPahtUiMOs9VfSBzNxvOzCM8tJTx2NNoFml2fNlk/bHw9iPlh4L82LQPVSrCX
D1PLAMYLUAJVWWi4mMmT4Kc2Nxejsp0XFv2K4tpXi0FsJaUxOqwVOkTwl3AJVwaVZtrpxmC0yXqp
YStNBZ+NIydWJbr2McWIFC0MKtbx9Gn27gWHJePdjeo+T7RrHv/A1m1INQdXu7BRBZLpYu9hTcu3
rKxOuQCp81z/gezyS3DZKcOQojBpxqqIyl0Eo7c6rYj7sWCLmujMHo2OiUYbv3njwxdSLgK0StPe
vJqSevkEB/LxwKGsWyy50zNP0+lrlqVtRUzV18lsa7SfpxXJU9j+9D6ZDIHKZRKAeTbk2cicUjro
SUq1Wc5RWAOfIh/CKUEjhs+5+sPA85mX/p6gKJ1VI2nHgDn/VXdpd5MPnhDz64MNQ4nrhf8DgGJJ
jDlzhPmskkr6q7LNXrru5wVC9fmApnR7JLlYoaPcPPOUQNbz4u6mvmv01YLExQYJEk+ZAvz+hfA7
dsIsxCV0WkbbLD9WgCpl6j5TrTneAl2l39KQkCg8PbCjCUJEDup8wuzKVoSARdEiXCt6Lj1R597s
puB85Mk+CrrLSpWitf8Vcbjd8LjOmoFy1QzpKCMsksl9jAkQ3jOamCKSVn5dbaUs0WYJADJ+J/zJ
/TtEZu88+TGDVxG7FxvDyxFL/nB46PfPgOTgFN4QRW8XjAz+COENWjZPnWSHDFzvEPE7YTrC8eYR
anqhWXYdYB+0Qz19S0q1eUjAgdpcj2IoOtM9STSYFqinF+vkOZ9zH9+hD3rRkDUbXF22NDonTofP
6C79+6GW+cb5qt+rrmxXLvcNxC+Ex1vCPhj4Y1+B268vYX5a82HOL/an7Pa1rcJQS1GJP6kC0TuO
I+vappzIML2w0hmvr48CiRGze58Xe6iXldxAKyLL5SniLemE2nQIjFBk6iyxNtaYknoQZpwvgM+1
OjWSwfWtgbrvkgxD0mDvr2UiHKr1v0JHRyKaLma2BgXeMA5SHJ8gJHErjIBjA9q1Yeb/zeI7Wsrg
0hLXz2uCb/UtAqmOX+ArZVVpndvrKLeGxxkoW/IaJCs8GVsru3nXWlAIx4VvKoACJYUqFnG3VQ09
JZrCCoYCWLYJErzQmZ2kdLzQ616kxfYi3oYVQf9eCxf276hxrF7pUBa7WEG75BtB40bRlShVcC/M
hQM/JQkXP9yf+Kg9MTXJ5HH5gdlhfp5FprjAenLK/eteNA2J7tqS9Byg/CkWTANojBsF1iQfsfFB
fL6WydRLGyUQIcxA5JBeFtOsDuXxKXSJ2OnTfT97QDY8rZoDdMn+HDYRkNn5EcezTodGSvyuGyk+
PAP/Ezn/atYKGiXksnDoF4SrvV95VyN3sZIvOtQDeWVTyIiIjUCpoCHjKd8cx/m7DffzQ1P046rL
5rN0e5gEypmzPD6rzLCLq7tNKRcvmzXcMNJlO3cPG+XTzU7RXo6JiKVuptD7xW+NqTAk4gPmxWqa
rVQqSC4NgkN7L9GQYwSkntdvx7KDexgVS4yE680Ky+sdKyYnLckN7LjgpfpxQisVs2xFlb3qeAd5
sVIlFnaZytu8Z4iqsdomIlAbdbsUUrIK9flVddGKa7GFy5FUQxyuXFAl0ZXMkVDHcAYqMtHG6nwr
uuDuxoFlJtckftsqAvbiipVqOoTpFpYRv+vur2hyaZ7sXinO/3qLTgNVmXgdVrTPHhFq9Yc9gDfZ
HKU7PiYu9FU2DTyo2FBKl+cC35VrU62j55D5SyBhHJ5AjQK9uPDY6mneukc8rZCtWTzLVAgH4Y9a
ADF0v5ckBko1RoCtx+S2gR0T3D46VzVZGrY6zi83x5bBNYhPwXAAHudEyuWmhQe19d9w6rlIUsap
tiXiO2g1dayh7z6zZ/tiQbAJdWzqLCgOmRcyFQec7KOuJXNsONb8lKrzxpWbyPH+a1Bc5sEY0s/8
c+CIZC4mXUVfzIHYi5HjYF75lw5M1eGLura0shUw8mgrQwRkja98vt3VoquWz4rwsTxaos0Rd0KS
cWZR3UpysTULJBCoyJCbEby7r0xh1ZQvVnUhvcHJhM0RQnG7ludU6c1hrZK+9u8+71PoefvQPKez
VnqMuieIqsa77K47+YQP+i/WI9yia57LXd44EiESa3ogQk4HYwdLLad6vNKgVWi2CAT9eVVTObtK
jej/hrmuNW6MBR8Ry4kwqyRZmprq1kUiOv5ucJ8snDPdNCR3kQRCAPSfuQlJd5A1RpUZwVeNfuTl
ChmhISwe8eNkIQInKX62aU0lj+SXHeI9KQsCwkez0NFSLXh9Hs0K913xJIzJBrIAlvQzRNgL/aIP
QiGXUAebmMaQeLJw3ABEw4m5pUgIFY/4cCJzZc+3gJQ78fRgCM3IqjppQrIMS45O78/YvqHYCiOa
pEaicdhFyGpCdFjA3IzdRg3EZxqo9WfpF5OEHiZPjZysAM6u6a/3JnnDjXnY5GpwKFsHNkaHxIUT
PqseuqgsjgUm2jltYqR1O37mtDfSevXiRqKWvfl7nqvHcq8lwRRkocnKEQvcEwPCMA8KOdhOf/19
oYGReqJHEKzadEGGwP2geg7rFL1LImDAituRyWcJ/SMXUqNfz+Vv1jGlPcD23kd1Khy16OkgXaTX
neoR9HsJm5jm23SCg7hKIXSv7KekeD9O61O8OQ1RGGfXaXEF6wA+xI8JzNNf/3VmeTkNKc8HN1G4
hv5QqcG9e5Bz6W2MNg51hSlpn7+8iEwFWNq3fmKviwTg4UfRKwwUe4vPyIpUqXq9uxlD+vEts3jc
8I21pxyY1SejoWBq3bs4muyiEOMLQ/2XD0HOHUsVGUrTwd0bbGTq5Yx6zqONmIHyH4NrAKX4L877
Ep0PUs1FokbV1Y46UW3JQ97++KSllLig72fjGIYobgllcp+Hw4c2ufAnsMdnNNWcgOMFseayfovZ
XU0s1hDj5PFSj4b0L1IV5MEiNYkrF/3hs5okWnB1CUAs8LvWH9a4MygCvOpwei6P7s8rgTubaxgK
xGukcQfXwTU6sMBJWetVX4C6ilBoN2Wt6K7+QAUoojGcGQCHCtW8Htl+DPImkZM6gaxA2OOxVaba
9+HIk/8y7U4MxB39aZtI9kGGQTkp95qfjijEyqE0q9O9i3uBldjRHEHB7+7YM55lDrcTSmK2QaaF
Ns4NtwlqP1CS08TexATExVZ8ESX9kPjOWaCgKhR0u1qEi3xScKyUxOOQuhUWhgMHDQtONm4VlFzs
5gWa8puWGe22MH8zbEWd9Uw/oWJPyMcHcjsargK91839A2+5r337TenpEI7UBoCfZg0TOavCJ7dr
xuGxB+t1D0CyEW0FC660QN0A0L7QP/MBzj88W8PPM2eheB9Exz7KnbrRXAJ1ROGGmrRKIqaiN/Mb
ELh+SxQzQ3bVhAXcxvG0Rs/Fl28kDt/yjslgC1uUbYVNE2JtANOwWGMHFqc+NK6HKqpiQeyLuurc
9RfQ6TvDvsMciQLS94diuU/NbfXNfU4tGkcgn+oaj/bmJ1kccqblJ/nGyKFVrRqpGkv135WHNzbL
A/lv50kzqa2zFl2wmDXnEmjUzCD0IQLv6FsXBSr/0n+6xfBvSsLyEGbmLz8hLjc8eIeWbZk8Xnvi
NWFzMzwE4b9DVdBix9FX/saPwRUyVoWT4zzmBHsdcpccO1zOO1d39lLJQuE8mzG1d64zyvhUqZPT
XXBqXN2D0HsPnqIefwlo6R/vy4oinwM0wFHW5jocH1+hjLl4ueh8qZvEyYiOusSFnV5XUnVU5ZSc
j4k5V7ZRQcZQlt/TZjB5xK24XeEw4QQ9CsjsmglSP9GOlIoikCJSgaYJeWR/sXbAbI/sbD9umB6l
FtXlgzroLWYG8WxM7mQntlgPd5TAOYPsgP+y1NHlBoBNYgsEfybHjyxBIBaq5Yo/rI1g+PjRVwto
WxsXr32khVQdx88SYRTFDVKunOu5pLghCGYnv6eTRiuElNj4cbxNXV+PFQx/qXYjtxp0pk0Gk4fJ
vSzGNDPgfupBJ22XPUJnr4Arhww01+cE5uiNrQbQ/5ianra82f/CVPTVeifhrG/722ByA4dNoU+W
0vHhjjlGAAGtAtNWH4EkVeSqyEnIjHpTA4vKntXnlyq8jV8kJKn0A+P3WA6+NgGhPkzu1/z8JycN
m0BZs70bflXaZm6s8bTL9TmTtgZJZtho5nitSXAeUdirX9xMDRMG1GwvJs6BqaAVIkxkGXdXt84j
2ty67zNHF137GZtitGlu8zkDC8IaxIFzNg+P7ekzJG7/J0xDkRoHTbkzOEKj2p9IEmYbAfpLo/9A
ZH+dm/7saP7A2U0CpgAzVwjmcc4iZEu2kEavHWARffmosJeFohT/08GOzlM2t9H7ErxopRuGEzZo
DQea06oS/tikZdcwL1t7pfM0z1n4advdWwq4u/U5xWmnUTrSJKjJZ8sdS5ZYwN+B2VDA3sBYjmos
VRwgLgAFsLAx5kt44UBcRqz7T5WxA5ezcSqakMs5/JdUi2ZfmSYrln4UZrEeDgUJ46C7tB9FjdP1
D0yOpY20CPhJ3CNAQ0FGarUrvrC2az2+knwSxx1/RUFRIRP/z0PIgu3+ADi1VbiPpBhcIzuu4uFH
9ssJW1akZ4zVFUjjqGoAY2laC8JyBPJpTBEVTJmQwOgHOUoWoVYi5lhTJmdKYkU9ns0GrOPkajje
JmdK2bj4yzZNwyRIgyG1RLBTaDxDx2FYXCrV6p7c/vFSM8VVHPPUEP4AP/wtiIpvV/LCUPkOnL5P
362OVwYFLbhcenQh83kAl2jWDm8xU4U592nDS+psSnKWf1jbQCpddQNR3dXdaPJ7T+Guhr4HyMz/
pED9XataOw14WB3nOvfLFLJD6kBs8zXxLQL81Na7rqLzxP5/CyDNOi7t39IuljGHOCPVWnQnsLNH
Btk6we6UCrMj/wVuBH8cQyAuToX1OlzEvcUhN6vpGR9ltDgcZACsGaD6yH2olu/zOrOwAtrUYel1
yK/gz67BCRivPD01baKbj+rIqgFHK/0SK/9BMQSjZrxJ5LbGH7nwgi2lC1ZkEbfK2EeDclDBHsvw
vl5L3R/gLkMSWlJoCZ0t4iPqCiQpwRn9cdGfJtOZCLr/RKdWo6D1zCp8PsO6sg6Mu1hQAySvUQss
t8JBnUodzMLybNODz0xAZrebqLRFnCEbjCTAMWGr09FQl6sIeA098xX37/ahrtnkJtrqmbOYKb6q
EuJfuGhSB04n175d+oC/dCu0MKCMWTupJ+x81/SYgZDOMrdnpmUUCoFEoHGg7p9cEXO/eFBjvM7T
yk/AHaQoicjb5kiCYBr+QFWY31D1X3b60mwH8pr9MhvedXdU2jSyMgSHOjvI6qfNUL3wE9xE1dua
DK+IJt/ZnNAiWo5A1xX7TCS9BpPJ7xPLigV8mpshETYFklqEswTSyvzHxB6sec2UYSxTBFC5B5bP
GHhFW3GJ5/lL9zgI8pzUes22VCqTSYQOP6G3mYzidKhzPDQq0BbJQM0/TIHenz+iwy8FsR0wlB+C
9bPSXPRMDXljtnIzvt/63K5Y/Zj9PUkRLXC8pGRtoRWaJU8f2Q1/iziqKMPFHZiSRwi+S7c5Y/OK
J8cTCCQ8FhQXdJHsrbZCnerktVXJ+oQleF9++oWXjFoUeVbXCqvVgbw65JYp0K8SjDZ8ysD3Pr8c
RSi5Z5Jpcj3Fr6fqN5wNkFirNKSpjDN+ZI+J2tQk8NmSsyplXDcZMY7Vc2gT6GmB+CCdyOxRDSuZ
PXs9huQJy1NkMnQ4c16zCAxbWVQkMuSz6nFwJDzFmqTazjhJ7JzPsNEMMR4mn1PSn/b1iPkVr4wY
WFaEUBrqtYrXB3bHjwt/XonmP5pP3PB14zZUOCNIXSWUa5/2cFafKxK1VwPTsygykI09fYC/zA28
O0NxxVdtDPFYqE+yXr7LX6tVIaMk8R4v8o2WTX4rpYrNNJ78AbQJ4JpJ6cLEWl0zTjFxeG838rUK
eIdIXMpAIGx7ALtxsS67URTTVFB0DmY/XW6sznZRsO5l/pIOafr/C/qrf+/5ie7oxvsqV6z1Vt3F
IDBkHOW5saLPdnHac9GoT51eTN4+GGzn5QANkaNOeDOsWo3u66MyPNKWoOknFaR6bXP2sj9B2myr
PDznwx7AHQobs/+5MS4RsObHco3BNId8YL4N1MIqw75R81GerciGkmuS3zhEUacKKDtbyiPlVWmx
vbAn/PPJ+k2Akb39U15+debIi+Pht4o3WeLLsO37rrmNggM9zaeS05CfgDAoZ02rRzxpOpNjhCGO
026Eyd7iZlmX+VG1Has7jd+XqXRF1EPpUQs9sNzrMXNLdaR9sg4p4iO+W+MU371+XeFLYDpUocEw
T9l5n/kDpHfhDk+YsgfU5KllckXu8sQtz1g4tuyuUrthcXtWJSDoCgHJ3e7ISJEP8Gn8D7W0KozW
Wftj+APUaV4r3WjvWIe5SYrpc721j5niEK/UeuFSZxSVHGdbyVORDeq3od2aqBYbs5mmNAL6CYpL
CgRO1DTNph6J2I7pns7PMoWbDaO6AW+E4NtKieuaKOfrReG7AMtX8KfPnrrMbc+kJFcVCjkPaWx/
3Nn2sxOOVlF9dUEBFJ0NVZrUO2HWNArfI5q4Zqf+rWY3QdWcKVWaFU1fWNip2jsfXvusxGpfopWZ
iUw4mOFP5icUZD85H+XgvUgej0Gb13Zo+4oVaxTTz9XJbxvY7yv6OZ0k/vCluPMLbFO38Dg2wkz8
QM0UPGu+f02nncCttMdGgRmg+jVjdKBCnN3A/XKnAioFlnAheo3Jo4+m2ih0iNdcTshWXJpHwdbg
2An5W46cQpkPLY5/D/WwxrxKncLS7ZtXTs08JSoVdiEE5P9SQzBmulEdDl1On41ORCdN+RIdxtrB
LedrNg5VdsoqKTz5L4e8RijXiLzgps8jsIAU5HMP4jpf8g7RwqpBuJpUO3PMZkat+VVJuyAoSSrR
pM0mD56NH+yX6hnJkq667lNlDwR7fTpop+pIZcairn611sLbisyQQH1T0aYDFRg1EPD14t3rLE5f
FBaNPXTU12YLPqPo4P0TS0SQxE54Id19Xf0HoaCPIez0c0y15J23S5f7F62/+fnxJeY77XIi3baB
4chSMlZ3WpUssmXHrKuV9MP4Vd/HfgCz/10tmvZo6BhK1GWVnaBNZ8WjxURnopRlHNd/ht++bcOy
0/BfO6bfOMlU9kLxhkso5Zjsi3rO9FI4GQlnGedHW24W8AoEI0AaZTLGH3HlhiDD/4T+1/m/+cTz
wT+KV9/NQwQYrxmCtmBzkh3ZZvrA1SewhCqafJJSMzydxj2uCCZGLHKhe0ju3AWHUQGu9PBVDoq/
/IqQQ8iE4wtAB3/37kDSmohDhrc1BI2rSCWw5TZzyQjOem2HJPSxBUW4I0eTcYuAGjBWjEEwWeR0
fNsadNrZKDqC9Xbz86fMwfjlG7f9Mm9wTDWwCgA8l9a0v8ldKtAN+In3p/IW2Pu72LqnTODuIhS7
YZlKmq3jwmS52YjlCe9gTwKVYMIlHhkDGD66dMAJt8XAjwGUfkE1f0644NINipy0CbScJUAIwqm8
UnH7gXdTfGl2cBXrizOS111NIp1UYkWpa2nfM/YhT5R+fnghoyYJMGW3EwNrEh6TlgVddBXJq2GK
L1CJRrd+86d2FJNxgvKvC5CtTNWRjIqcSzj774lZ7kcqlxrPYYKGbKTI2wPaxALU+1L9B3bpUpua
C7YINUmVmUfzSuiL1ZQy3T7Pyb8XUqSbl2lQjb/mECA7L1g8u/4LNX2dgaR7kTGfPDCSyVqT/NMt
hZ/sI3t0tzEpcCfdfcvdWYcQ1wWEjb+F/EB1uu8y8BIRv//LfWbJXjmXUlf9xF4tvOBsckOOXSgX
Cbd+EuoAgsjgSy8lo9mHpyZrizkeHlyrt7g+pmOehewvyvrz8qS11kyv9AOerSckCYVAS0lZ7FSn
2aPbjDv4l8xv/mdLrXNKcK/xCXYgmKHWZHHLCinEOoRHwo1Xih7RV6xfKsDPvV+u/e8MmApjm09q
PnnLIkCF/6Q9LB10oLfdE1Zjl/GA6g2o+dl6WDxrhT+FNnv3L8pZiyJI6EXongSk6XaihzJosNnL
jieJdVjBRErTqmqOAwDxADlr7M7fOlL5v4VXTt2nyD82aaj4mpXgp27ZNf3teE8kMJ8j3uZYflOW
HB9dk1iAJI5Nepo73yqbrcKKcqv0L4+HEnU+UWb+ISlQ8P1zfSgU6VMjHqLEsqF+qtJE8TzRoIyi
YyG8hzSdzi1crsMGbJbRTYOBAdHJ+jX9pNgOUqKZbvuNh9XH4r3SS+CidKAkHOx+YeMwSDt0G1JE
mi4k+boDOlPpPar6uR3pybmQ0wibRlJKHz612mtzx4tXqc+eNcxAw80lWdpq0HLyZXqHrBS1DpWF
QRWisW2mwV6UNcFersWItXgECLToTHM3waSpCvRI5uIAA80eobFM6CiWpMDiDpw+xMgR2XQOMdZ1
mFTAAdJoGODGjXx6O9ZZnWMWwseFwHEwHRDu99D2nU5NO4oky/B85vOXagQvRt6R50qYHEO00wk+
iQJ3NRe0vJDgCS37u/hWnbzwFzmGn+ZI7gYidjuKo9Fa5ftG1B5jo6Qs4M6e1pSBOQ6fMI5nJVhn
gkbyAiHvkkyiudu1dqCV96rkhTdZbbjLvith6XumoQQk+i4jQUZMz18d7m+B9cAtDgoJ8ueXe1du
c7C1u4i1PBXbJaljzsHjO8Ozz8EeLK2x0vspjPOHQlRFmIanJu6Dk0Gs7vgsjzAKQeDa9lCgmLF/
4eOLkY277x3fgF9i8igBiLWLlCHxvGlOtpp9ys5Ev9jnvLXNDXCl5oue95/6o4PlttWyC0NbUrwJ
PT69Y5ea+TslV3AZbeF3S58CkTGWndwyOzifRzhuK/E9cKmEQQPGA3R9Y/NnIST+bvI5inNyppA1
PWXx3cleqNTLnTa9iIiYo2yCN2lXjiEwGWQ+ip8YoR6Kx8sn6hR71RNOJTcJQ6e4uNVmSKrFn2xe
2RzYTtT+H6cOhNnQlkENIoTIThuOcEzd3I7/xdEIPVFuwjKLr/pOgBSm+LOBtaeXd/slVlJr7Iw4
iTGVV/vR7Tp+R0D3comscC7lPLqbeYg1okJ+JuTf/2xZi2TvBR+Ku7q0XMJjvJqK1JWu5X/qICfM
5LjssBfE5xvz9loKzgeaLvxq2z+Fp+SG+flBD9rCeQyucZlH/rZ9PzeluUACiXX3S8A4SB5S6Y2B
AIicJk1bFTt2IxgzsU72idpU8vUTSU6EP82HgHBDOm8NxEtq5/0e058RVhEwyyG4/cefHqzEGpTD
bUJ9eW2pQDub52JCySo+SR1evebdck4IzrX0OzgPwtjoa2m0vzhLTnTu5Hqe/nt74TbG6L4Y0CTY
aSN7fHIuzXlg/AVJUdk8xXkfoqfxOErXl2M6Rw+QAyLNFWWtgAv6vhqKZ6BJR3PbaVfXxabDkKwd
3HMFMv/UbhCO/PD1fDnQfe7rlqIg5bc2JtJQDt6Fo6AKMLRv7VcN+OYcsmqa5GVL3mCH+WsXjEi7
4U8aE1Njs3Jkk2dvcVO8vj43ulcGT1Zmc6aBNtsockNH4A2Q4xVnTFhUh+z2l1WrytIOeNSrXi1p
3Z6NBqCSeaFQH2+FXqzY9KgsBgQ+fm/Bv9iGu+Q3IxSl/+GNo7zUKLoY6wRP6nYbBpqgZaEVDBYK
KDK0d1t5HcW4PxuzM1+mGW8jzYnpKmPmXhszS6v38X24wJ7AHw+4TXgH4eBqPVO8Q5r/IAGenAEM
la/gy3ZFwEGAkXqYwPskc1TlhlqLAjHZFo1NR8Yt/wjaQ9r2wYpVtOXN8m68jGX8d6ehWkrEWQ9d
XcSm/8yQbN8tZoRE5TqHclbdmMdcyQO5mRbGWOcTfFDjWIAyQ67snHXaGPABtiDUZFcIaX3UV0SC
GyRG26JLqXSYUcW5CQJ8vH/gpzGK86S/Us6B2ETRdLBeQ4sP5Ur7lkU69iTHhE6Qq5whEAXsFOZh
/IPrj2mkxJdjTxAQgMX2Eemvr16lrTmSckRQb7Nn62jDbqjiGLxOsGmsIzUKOnOe79OoGBkPe48c
ePOw8jhG/soW5biuqjVAIg2XwIP6viLsh4UDbLiiEU/a+q1bkk6ao+JEmXQzWLh2+4xbn19TURik
UUey/HZDqPyxVEux44okEIfpHT5SNUB+qTCp8+OZLZ/Jmmy5T4X/HmDQ4M9moEk2SFqV2iuABji7
Nji/zPQksH6LZ0I6xnNgD5z5asBt44B++nPCCWS/myZRnSFrof6fWeRel23FYwWBRHkhhIZ5LHdG
ufBKwbPjLpyXFXGMVAq0gz+ZHS7NMt3iVcO6Ctkdjzpy2BkLfWy5PhERSE7MNSodeC8h8MF8lMvH
VjwxXvASvxBuTEhog0Hq78bqBP5wGmZGJ0rnVhD7dIXfx1LdE3fNnIy8iFnskBXwYFuoHzhB2YQy
CgloFrNktx89GhOjR6tjEtE2l1PxfCBH2ByJnrGjblK/Xv1n5prD5Q0NXsXfXuiTkZ03Py0CiBa/
MJDR0DXS69jZgY+XcoZLWGz8idVwvpoklGOKoZTSOEr33/xMXtEO5FiX/JNMxp4dv9AhzHHGOrAG
gImm5HGcIVd3s7wm9MH2ZZOydm66SbE1/kJMRBAaN1L71Vf5JwsuuEhe4OKzPqcTckuuawpiwbiQ
kT84e4/WiRZ+mNlcOhIE2kLRF2lu7o23o4Xa6YF6FmsmhatzQraKobHg3zgyCqCQBL1qAkpozF0k
aeiyspuz2kwWTvGjZ59yJ4V1K6PbbHm3Lu6I1p/MUezoRRtA2AHYmaPCqs2uzH65A1vZY4ozEkNP
Jz4IY18ObRE6tL1I8anBWRWyMeOvpIHd2pcN5JPoytdQOuSaImGPwmprf1Clh1YrZw1vIo7MNDLI
LGmTvfYslDbE9wyndBAlnakbatcLLwtPwqPoC77Pw0N6Rh0IYNyhSwPZy5L5vaWbIbnhc+lkhVz7
OsUOkmOVrFD5kll/CcFq8/En7PRdcuXz/TSRDs+X98k5pJyxrXwTPQwR0wQ6eALREHq3+FYy4i57
oNSwKCIvOOf/YyPp3wEHJ9G+Pq/eAPjdp8lWPFLnr1Q8spLStEvYhNp/z1hqV+gwger2pUWS57XV
ylZi8fdPYcZprWGb8jLxj4twz/EgH8fpCWN0A8l5MPABYAxCibko1520GNJ8zsqmZIx0GhrYzWee
jF+n0EI2j3NQL5vToqbIQJIQU+Hdn18JqZOgO2UOLKZnEyqT4pvpvNHBfliiNnJxxZZDbbUwECR9
E4n+UNn5szZPdsIxFWjODeX4uimQue37ta+5JZ2bwKqJm/I8vIxIvTu6aXWp0QqMpgE5bsBPzZJu
i/kOgDKDWifp3x8XwG98YIeK4ijn3kN0N8FL3MZo1p+6Z9n8WcTH/fedv/Q22CTbNn8UaazpH28+
IHKcnLOBToqava05KZAbPnK45v2tKD9vpDSilQB5Xg1uqdhF0wGWOHVTcMZdhAPS4sR9727YeNpn
H9HH2cIUMrZvUtFDjApO1nnOhrfeCCUPjLGHtjh57WpNWLdbzjYqd333jRSuI4U/+BBgCkeiCGVD
0ynMsTw44RC8uDUJe3uapGu2ml9vRA0nZ7iIAnLmfl1ESAVDJpVmeUjsHspH4vp16hjI2VLwaqW/
j4k00QCQICj+/eaqzJmpic9A/b7bs0yLCqa3l8c9Ngll0N1bRXc5LGk1FsGvg8PP84STMDpyqDWE
jnUM1U32Hd0AIalgrhu2H5wQhMXpzMwrSvIiW29sNBNfcYjm2/o8sjgrF9r8bxzKE5EDqdMHd8Yf
w/PU9xmpKOGW4EvjUlLRBxr8mIzm5Pqi++1zeBNxNuOeuHafpM4YXAXnzvoveLpQnGkKsMv4ZQ9Y
UKKYxV7C/XrIj47KimCxFG1Lm6vB9OPcuIG14RBhqUyQz7DctaAAr22PeK0WHaClfGG4XzJnwDo/
j+WMsuOy+AgcPDh7+ZQe3RSoL1cHX+geGCjY6rFcZ3c6E7bRRewzjFdY1MQkzEI/XCCeP/bDQZjc
Ij4/y2wXzGk2mI6qDvztA94vdilnEKUvmhSk8cEsZOf4lH2gYgw/p6T2KbO+87uHBAgE0WyqjLIU
73zAMvVdrVEhuByjrmT0k7wSdjhTPp3eZjJqj9ZsxzncYtvug5xB1E6hN6nPt6e9rdmqdL+mrp2z
4QHthutwjkFIOnANLrJ1X5oHYT9wqxpjCBNOXTBmBHvFNBJMaEvIHHKw1TyJdrnxuPUrsFmrZV4g
ieIEbMuC4uC47WUqULNqU9H0uaWZKToNm59CwtOa4QpGTI8T6IoEnUUQcj8khtWATJQArOJrpJkw
qrniu5KEEkj92eP1E2diRYFCskMyj4cqkx3e8GeFV3q78OPgbCvTbfpnE20vKLcSS+cUWhe0eQ3w
kTo/ylF6QtxtjDvPiv1WdoJLWPOe6ELV78N90z3QxkkfIgHDuOJE99chLLllcIx2P5flf3E/ncxT
HHi4sYJ+qt/n+ZReyGNF40BqnbueDz/QZhuzN91v2jmdfxiJi9mH6va7NwfjsiaqUBwUStfXTL3Q
rXvzC8lJf9oNbi1a/wvzjgT6RlxG+R335hKGAmdxAS8uqqiWsjZOHbDS/ZPRAOcP+IMQkkyuMdWO
TbpXTsCe0kC6PkedkBp1IDfXLjCLIrENFPcczLZNcvBggsAt8vIGED6q4wivPjB+2x6wYrBtkB8Z
bdvTbgfRsV9B0gHbmDmLuvUQVz6PpDWQN1nAxD/0BLoylAx5G0ELR/oaVAA8t1/g5NDvHBcIgzK4
8QGFWfcuGfH48LcIyb8smWy4wrOjBjChoRnEzUw//+1uqW7SGmSl//7TcgxCeMhj/B5Y551m1Jm1
kC0NVZPiiDBHMBbFotoYwTY1I/XgJ81SJZEJWNbTm7O5FaiG5+rrpocMx2Qt9auiL53zz5NPx6X/
nuReSdu1ILiMoq8OM6LsSBlSolAYz9RdwF6LvF0GZNrID7CO766CHktB4WiOrWVb8VI06tk7d05A
FmwzcV25iVeG6TLjoUYm8bbaEm8BD3XMih7A8dDUzdvVLqaslLfl3xmdtIKjBZ3RpmxJNMkm3b1N
uM+3KNbOqNFPNMlVNpUva8OjO5gyOLoHExJVAd+PV8DwPmHka0eWbn0hNphcuQkV80Sfi5mXwZFf
75Pb7Q/zdBzity9JFphvcSZNBTCWKV1bdNUCvt45rH6mwMgLR5NysQfeIvOgt8EoE359kV6tUFrq
axdf0/miIn+xvQXAF2OnxAfQ+YDkHs8yi1adGOe4RdGeGnsnuv45k6tg0hN0e3JLBpap5QfUTbtK
3lssxXom4bA05wAkr5hzYC015SukD7T6BRvxskSoZW8aR5qBnldbqLyf92bMEkppRpsWtmFo/pvc
dUczuUfjvwj1lErkG29KWNu/b1hHRCsQ/YckFnCl/Z4mFQdJ6iIQkTkZKGK13ka9bcoSE84pF9cF
BFeRK8wILx+uCH2Gu5BZLH5CK3q7XgR6+CC7qIUr+Y4iDASFQCc9GD3xkCZKivye/Aw//V0Z0L57
jc8Q+fzlZWclKy/gl1+k0xSDeJzh/+y4CwKi6c6DpSM1XYtkHoPoeBir/wqfRCjr+oESTfax1COb
zjR7aJGlcICplTago/xwHRscFrpxXjIu3XGDYL4f67FaD6FNdvmBh8gQDEtbvxHwRwfMcJYpQ8ZY
mkUO0kZsheR5lhyrz+2ipS+//ZXN+Dwbe14H24vIWJ9lC/U4/qmWSFXZlGCp6if0L5a3wzumKDfD
Mc7G/IZxllMPHN8bjIeOhGYzyuL05uo0gl7ZcDz+yKDlyTVPECxt+tk+rYo5SguxEQYftjMwa9Bd
jIHb0oZuLizQkFu6HVurfJ3DfF8B47Yril2pzDs35shSFOMglQv119HD258Xym0kGfNMVIKlzY/j
uib9jyO57UHsO6LSRuXRTarKlCBPRB5dKwd7kR2LtmglbBox/5EYRM5VP26ifslf/LMEKOsPupVe
XmThNdSpqA8MeBpYowH45kj9FGOB4Jgmcshk3oUsvXblgd1PkByYSDxHN9F4VmwdhPQXXgJcXht6
XJnspH/Y0d5hLRZbLtaHRzYihwHectw+FW2ZggYv1B9l2pi5dYYLxo5t+nxelm1Svvgqy8dAe0dN
hpsE3J8KcfjYI1AufQnwjeBoudst72o5nZXP10Omw/bYYOuqpxDyEGOmAW8CQ5EttyUrpP7R/4sO
ood/auZTCeStR6IB0E8mpk1gKkBcbP6iTN+He9UeO7AV8piOfdujJXqhQzwQji2mcZ2WDkgxpwA2
oH91vE/gT38S5+pqnwde4vKFh3OWnaQJH/ibG7cyE20BsTRNsLpODz2EjqmOqy2HqqHEG0SIGn/B
ci7KyGw8eA7UC8yR1Nc6VnRd0H4X4h34FwaSJseuPW5CJ+pYftqftoCq7ytFVRVuPguFzsKXCauj
X08967j7CVTns26aDWoeM4U/+smlH1/liS29/mEAHISSr6BiJ31H0Fu/1+mpS/ekjsgNUpVYyKoQ
8cau/ofeb7RLUk5isD90p4mQhEYlQakmBPSDcVEUVcdMMgn/3UJkShCn1cn5bkk7/Z+Y6ozjWE+y
/sbm0baHzlDf8HOtwVewVkyczGAVV/QAWH8l1Ir0zPC6QZ0HMyoql69v7kE+aJwfaTmtZtlreWU0
UpHFj2Sm4t7dOVG3jITT1TS71nCQH/oYy/JJGNubtX7u+oVwkzfdm5PJry1G1nEhHcIrA7lCQPZg
vgAiysp3XOXrWhyTDpxynTye7r7e3hRSWOYbJqxPEtFN0FQsWbVJ80jOK28xyqYC4zuQlW/MqJIz
3oCOgxQdGts7aCVSh24/lgXShKvRNsAA7xBS5wbcPUQL8rTdbXIUWU4CXZzofa8vBTf+rLa4ufwU
eoznYNKJQ7gDoAJQdiD2uNzJmKaiIEugA8o6nHt85FlgrOR3+NuIuGqeEbRqzHueYgZBX2PJfsH+
ycgjsjV9Y9a2FCA0pbzQMNcQEGztllF/RFKgbPuypwcFZvy2JppLb4Ss2Y9EJ9UefAiKv8Hk4JK3
QGEkgR4PrIuxdWD8yI964vLSiBnV83HplQrmFWUtR9LuE+mRwIpLuERICyweq0pU70BnoEw8Pftq
wgF/6HBt/Sv4sqgc9WuBJQgMnxgYlOPh6ibgFqbwoAGko5ykZYA1V1NpQrog5jHrsjSx93AZft0Z
TIRVAiC6jQG0ow26tIddCwr7262sy9w1Jd7O3JxFvn8cJ38nPZkus84uU2UBUKAq1xsv5jAs0iak
+jUuZWVdzixamGH8Y3EzS5tK8mJ9enh0IuS41SJ4ff3AmA3+5K9SZFwDz/l8RzAokUFzn40Y32HE
Zi1pTLSzg4RTfyMdDh1V4b99wR6wWHbDygPIYR9OqwtEPVmhCorsrMAhPST+2xPxzNC6T8Qu+Fa6
DW1e4WeeweCi/iPYlECzK6Z4iVGFHReJOEbueIlwsT2BmQfx0S1+TfLmjqCXXQcMZ9zg1Md0/gMS
VQ4TUIYW3plhYj0IMQ4TPUVm8QvOE7nxORGyw9HC2dYpmkGmkssHWX9hXnFiDIneWsFyXJNCL5KU
WClbRrrT8YK7VAoKB8W3lnEk7zTuOePY2wEgU1zUcplooZKf3HGiVc66gNzST8Tw/dZgY78kWLxl
AOujzcLOt29VpDJdl0aGCb2SHcTP8wG+BDa4lIkKYuGwjH746eHPktbsIryMGS7+e+Jcl6lag1sc
Vfulg0M7Ifear074hvwemknVgBVWHYFBc9WHaYeWilFCBXc9xz8H1f3Knac9JTCFkise178zlpf2
CQyLY53d2jch27g8SRUwz/f0QV7P+9VQo6kvTyUeon9g6Ms0Qd2p9bxP/gmwrfmnITI0hpAxwA1E
4Wa7YM3FYA5uw/R+25y4tUs3zkHLVLHW9NVzHMViPR1VCPYnN7TWjiH9HL/8fqD3ZvX4DR3TYHLC
wnX89Oft7wB1U7zg9I4vxzJlHIeBl7HZhPGErgI+iOYYNOsvRf+zM8r1qmldJNt0fH7GiEyk4wmS
ap2r0iubH8Ad/jFXwcp8+A8hxxZrzCBFPFt7tUbpaaeLA76ZSrq1rCdWSjkaPtUMQuZ1leskGWhN
SFWCQilxR8Ut9wyUcgajbD0bYmmmpmATohB1lg5uO98hi1uWMmx+pyHyMHPeqUA5hyH94qZRKFfv
AldC/mbwCyScO2IUXGNOHBBg/1dsoLszANkDIzZvWUn8kk4YrcS8/xaTDQmP/DMcp8HEl68PrRZs
026gTrEHQfBM50KfFA9pivf+e5TjhQr+05JcZONXMt84uvfLWGgPSlsES3A30ONrpGhSyVF6P4nP
Jpzix6I6O1WMWFZPNT/hCbhxuooqSTT5V31pXLxZbCWuxOXio6XH/FGuvJslJaqNovbvgvotA7uW
dJIdFcqq5Xzz2+o6XvsEUmWpVlX07IKL5Sr+tiU5JvxvQEHLynL6aLGT5jobMJV3EPbfZ5e1P/j7
z7Ikd20y0KiyQu6tQ6gBlI9X7ZpIuneDUUz8swEhIGt+u/8eWRt6o8Y5mq9kn09vWy+Uhm5DJ6/h
XBa/rQJGjip2rVcRDkUc+pfu1jjKmHB+AOwQmZhfR+ebZ1i2f29c+MqqS4aXV4n6BUplFCMIcKXc
8ZtRU839sAPdK4H3LjULYJKp7fOKHAU6CD6LnRy7yjNMqOt/KfffrRkZ36w0GmYshXZeSVaN2bCT
miEB0QYIqeCd61dKQ2DsPOSsLi98EKbxKrCQopemzP9vDbvErtb5x2sSY91iE9YCxcfULxLA+OdO
kCNtD/ebRE+ozy73UHDC6H9V/Wdl9DfaPt+PR0r1T5t+s0NzqwTYPeDSpPXXlfJ4l1VPQNh3O2pe
iNdiBv/yW06JkctO6Dk/nIcHxrNSgWyVDYFOqdS5Lymd0/QAnvr3rvWIEvWldwbPMTc3Q3RzL2gg
UXbsgF5N8jRTemjgb6lGmwVnteLh+Dhd7AeUD9e2AQ2GcPuXp/fKvrqfetvxFJhQ9EQt686dPt4x
qDHKuv7cwFHmNCO3RGcT7kRtRsPaM8VZcmx31T6pyQarlgw7hu/vpY8L+ibIzummzwnVYzDpWxbq
EaRipcVVk2npipVt/D01l18dTG5pMpYcXfeqlOWG5fiDTnyYg6WQp8qe2YMxuUPrxcTpzp4JuJvc
AS76e+4XmyrKXhWWFqs40nasQbdjrPflXRFpLnlwii+TaIL6qBqNETxjRF/MN1Oj0LNqxlO7LrTA
+dBETmVd2jJ3mcL3xnKjK7CsbMa2dgU5FKsRslZJlrs9JcXqPkpn9Bha7Ew25bUiMJKQzKRv1RKN
yeesK5DJYBfJ5evCD8Y28rpLKv85fUbukBck1Kc7tHV2Wgo+n1UE/IKkJ08+Z3XGbQ0aPyMz1em1
okmHrIcsKOJiwDfjh3edHSAfDRnVbyCVxCuIQcQamDdVuNLjXOygFQ1YOqPOcvcH8L6DKaOu8cHm
N/wFKGDhLdRuqKUEWgBMUP+pE6SFngTU8T3DtOFQQp7iSEN/OGhT6XjQ8SQjWAbYjRd9MI90jGUI
YAHDBfuQY/LVegP6nMAQ9g1zG4GrpT1ldacE530QV8Nam8mtzCTw8aX9IMa0iqOaIdUFqGVTIxUl
0lNxBiHAY8+6qm0Meu4muPCzFTZyxVvaG1I2l3LQEQuGu32OUcGfaYpspOrtOmr2jomKB3+Ymu4T
XahzkedEwz/iu145wNmdKSCXdDDpvdCofylPUfHtNPWayaA7pAYPLMINb19NWzrAWM8wi6Oa2JJb
oDjxnFHy7WZO5TLmPQHa6SVL7dhtcxUpcD7aLhc/kF5X9u3+c4H0b6zfSHDjkbUuP5G1UD19mOg5
hdrYZSzFg/t7USug708+hD9WweKd8UQcBrp4IvADhbsEk6up2vB+3r9F76LX6eILQD8pYTaJoUyi
7pca/RXx63bAlocLxqFQNZAlZZsJX6xGnpL5Taj6CQO4jbC9H2vkhvoXiX4LXFZqbEv7ab+Ec/PN
Ka2IhxI29j60E/RsoN6Yt1UZ6LhkjxKp3Gdbt40r0bYiR9GYTcByT5b6wVStz6skhV1NCTGbGeqL
SQJ1SotAjPoVzsoQam2DH2dNPzs4xfGLob22GQZtHjQhQUjWIiXUWCHgQogBv1B9xu/ZitaNUspE
RnN2HtMJj6hY5VxYyq51fs60Da4AwsRvpwTq01sBd6ZljQ6JUE/d3BK/hX6N48rkE2seT+1ocn3d
lHHHnN4T51hZ8T1v9HA8VwxEMiEnBwzV80l3s5gCzVVSk9QvS11iF8R5X4aOsJeQYfy/XsHX4m4y
wY4oj6ae+Etntz0NGYQzd2Wi/+GHO6ugliYIYkiveeRqeGrX028Jbd5LBWg8ou8FkKAjsUWh80BO
bdTEEPpvOdFch/XTP4N+AKO9eWSIar0RHEMihgcMrNjrMcW9uchu+dj5u1SMr9VSTzl5WLEYKyyd
sMm0ANpMiAmBtPoY/EOiSTAuxVKWBf2zwdCW0hTQbqY4yf45a6ZkPZEGWnD6C2WAwnGoYFxZHYON
VXiX+H0ixSkp1GHt+yAZoRMDicgZmkaAnV2mIknZ8pmGmuDsHK9y/6rDoK8lwjYkPIR76eX5Tt06
oQqKBheFyxETTfy5EebDxmObj7A9BcqWzqzv2PRr95CHiYBKv1EXpigAyxX4DU7x1HlDxfKSxZjP
zX5pJIPK98iinULwEJ8jkGrtC2Qg1ahQ46pB7GRluNwr1XC5JOSS7UAEhCFC9rw6RAk01WO5500z
W+zafdyPnay629OZ/wM2UZ80tuuuWMuVZuHvYH2IhVVjH+Aim90ZO3swx0w5q10Co7mRNDrMBio4
CONBlr3/9QMwNYvqW6utTL+S/WwPKbjawSIOGQxEvQfp3wSKdFVj7rdYaPcGgiNFHqpBFy4CuIpN
fxeEOh5gBy3C3qukRa3tGDk0bFcebhCrvDRiYguFc1xQ3UgjrA8hNQVF5XNSoBhpC2vNgdh6crOf
s1RmafJWWmM36Afm4SasxbGij6gYwtO5paVIXm5sutfirouobk8EzOivRDP6xjvetTyWBem8tusQ
VuC25QVhL5OJSTqZxU2mukZRgEtxmlBQZg+9zds1xdEvDT+VUEhjIMlR9hZWfNcqX67bcCquxouv
sw/a7Obl/wsp/IO65zjIRMNVt6cVc1iIP1ECHtGXe8k6pMJwnfxlJMmgFd38njG0wsXlbvH9y8dZ
tB4DZ1nOodE+Y/f3hfXTlU3YTt2au8nCaITs+UPj4PbSFbuUDkk2buQa0UJ4ik+SVUQyZhSWoxMh
1MnrUZnvufvdsEj9k3Mx1UTgzN5smvaRZ6XsMJn5PJ4+XRb7PBbh2/nBha8bWjT2NCgKVJuB3Alh
5DXjcmz6Ti59/CEMuAWElHDQm3lk3O2pA5Taxqh+QhyJx7TjGgVmvXQ8V2+kjrF8FECFDMM3hrj6
/kh0Yj2v9fFCuHxKMnzmhwTfVAarxfx7fiisWu2vaE+gQ505ThIaXVYIuvezJwCSExrk8J3YpUZB
KUp5Iu6znUAzq5qSTn+/vuYDrvOXJK9LAHQdJiMpHzqtoJMwmJosjWQFfyPSY3/IdK/gI4HoWVfK
O4H6MCTy++J70/uFczGy97NVtETFcMOJrcrKHF7M0GPq8E5eFTc4PEJsTlQXlkRyMg9ovmQpOtdU
+2HBoZHbqKLBkzomtMqZ/e6GfQC6CVgsjJtz8fQXKX5PaZ1MW4hOtU9MHSIRIxAtzyitsIbIY+Ng
BSyqT72UF8oMOFBrPFFkLEWL0L750/Zg1cyvA7eloU+R4wxrZqJLNX7Zf8NmyVTmTaQ13eBPI4kg
jXKqIYd/AWFDBNlnaD0gKAl1pEx+7TpAhN/SSXTnvXkQ8MwobQaKG8Drkbv8bubU62ZfXx+iaz90
DN+u3QGA8KKp8/KatNqIQcQxS6H1HyFJPOuZg2ttdJlaeZmNWGUpi5ZgxmNFO4B3TQNnF5i7kjxb
3R2Bq7rZiGl6ySOA+AtxFPm1Uzs6WQ7DgBRErp6bJIXiDjUF0UwXjZc9Z/7NAxxdoxieiV3JD0RQ
Z00S6qOenfVzCG/Yr3qb4aNaFnNhjW+irLsj9c38ChGkKJDO8//AgO0grO2HcaLSHkitV/8QAhLU
wAPv3p8mUgkAoN4Hh/imZK7KMELwRk2d4U7i61tklRPh5H7bNCc6/Y32i+O3/SJNPuvBtO3KAXfU
MZuRb2ORMhcQG9+1bajscKhkgFXMTkPSeniRyIqIQOk91ZqUFovRVk8fNELO1gD1IdRJUUgGQiTC
rpcF3pwRmZsG2YxBDbmbF1kvbT43n++XwYKMsOz/QQ/bR4SKib8VyVBkUfSTCJ8pdmL1VVXETAfc
N+Jbg6vNtVEUsMdkuW5c/zuo2p52RR7FJfbDL3HfZ62ZfAo5wKuDD4oYR7rxb6go7D4XYz1P2od1
o4XamOvaGQ6Za44WSBW12lF4xWnJCCNWHxOhXEwYzGGJz3K3JhgNcVZtUI/zlXQwOKTVzECf0cDY
ZiNzqdzoHAi84sBm4DlLT0O36s69ztGviLnkWr65eP8Fs7kaeChVicQ3SYX5Se1VKSTCfq95VmGV
rlwDvfIDa/87JuA5tnxs7uhwrM+KzJ4/v70aTx2gSjiP2Q24+nyW82dPQ8Tnw6SMhacqNs2nqa3P
xVDOYCTncp+JcV2Kfmu845DME1zrS2c0uC3UOlQ4yWeTSlYVFq5oi09Kac/EiLrJqdQkf96ybMLa
4xsGdf36L8sOaHnIZzwKG7BZbUG02rcU/nx6nHrPXoLpFvGaxEnHDKcljXk+jk5VDDx0tPNtGyKn
+vbNLcWUH70u+xh/QmyqcWHAXsuOnUdLf0fc+7ZGyNEXhgLhoxWaV+1YFwhDRCNAMMMkD/V8Fdwp
u3mm1io1+tQJRJWW7WMolhMO4TAoNIVJvSh3Wk7FIZr1+1q7K2res4eewnJbuQXtkm3QEQciNsDG
NQJ4WfTn6j4aVqlxmdpNgjp7YcYTIyEbm1KIxngrd28orGzqCOKIeAF6lGDmff2vUcoLB4aB5PAz
UyTOyxaniYEB5WnTNtekfQd+laT2QfEczM1M+DM4XH6unC863Oo6XLHuzVkZrKq4loa6PhG/ZJk/
6ARuJv7Y65m7yJOOJtDevScjl/0cSj9TCwxWR5npIIjC7XqM00UFlL2wusmziJTFpq5Ai8kMslmG
7duZzxY+rV7d/Bd9Ltl7jVb9QmUYj7wrMr+1ICyH9V2JVBmbXVRTnF0K42qr4b55EwiaPvh47uXL
E4/28AYT2eTgTvnrZwuRRVl0t770jcKQNQQYdFdlDgl+joiiIgAEViFaMfIHuVusSip7mf7j1OyY
qFAZP/XSs2jRiGoNJDVUyqxiuuJv2w7jLkqh06uW8s6a0f+uHKJPplLkq+N8McL/5aXaXzXpiXbN
e/PO1cBFnvMkWCKAPXvSby261H0qyNbPKKFigFAs+KrVy0vs/FQmOE6/Mn2mbsvnXzAzc4ziaSs1
SxNdJGzMzjYduMtMGRSvBaVAEUq6gAcMLVJ3/Xk+vFrYPjmVlzq2i15kXw97/sSu+uvw2wB8wP5c
TJ3WzNjoWhGr6CZdswBqEr8WdoPtTRKYgA1gWV9zL1wMv56181ux8LF+CAUzi4Dav6zQ8+8oqjyH
P3Mha5re0uI0JyJBhUhWHrpWq2POVL+vJJr+mTb+rTQxUbCo2VrXaGx5YHN8asAketHQ04YXqcWq
z+9jefvQkVva69Udah2m1GNlWZXMaBG6vnkHNUBcD28kV3DxKVVCBll/ZKelw4SK32iUZ0itPXxF
a1j8RXbjTvAE8692LEL1GNxL8PCugIwBmk2aiL1keDxWWmD/Rt7AMUA5P6FB3ikXe8oMMdHebqLf
dsT81G+2HvRDAV64lVdjj7zDVtRbbzuNu/CzZ/5w4SzThJcDyoYLD3/KtCVt+G5l0urHeXxHBOA3
xSVtHo7NPIOCeA/8elMqdQAY5AX/pBDUY+1hItotsjzbpPNmqfbGpbZ64+WGSxSmcmqe7UmI3VAL
iDTVU/5u5ojax11ppK2KyXhLSBbQTWyM9pTz/EE+3em/9NnB8RJnAMnSdmH+1H6pWc5uiTOtzt3N
yOomQgDtd4rq5qxeDK5GfhQRbLJjVUUZcNppL/J4tqqtSQ38ux7RT/qLuv3YH77Ih0+S5PIYGdIb
qHGDa7dQG3PSjXkaeQC/2beHE0EDaxyM1npy/xbcCJ2xQ5w74dnosTNLMXz0OM6sDuQIASIPLKo2
rZ8QTVrbMMSH81N6XK5enntS1ya56yv/X5lYLZsf7DrEA6xp4ejdzJRyosElXtwiuUbgtN2x/qK3
P50Jn7yt8jqQVpL8MfbkYOmBcg2Tl3vsJX1HYr2katCZ8ToeSTUV7DJbhChaAIDNyXGYLVtCl/+d
lOE6jrX3g0wEjDmOlfzeRHr12Gd4yKt09eI1R6deHHQLlwR0p1HAFFDJXOZyGwJuA2KDQMag5mJN
diNaDt5DyEdR5/CmHdnKhQCrLdC97neIslQN49cC42S5lDpcdt1MZGYVesaJ8WcFTLLNZSNcvtJM
9MvfgTsrt4O7cJPGiOLBRrS3OrWHfbExrjOw5XSsEq93QbNNmeiKi7qcrlEMpkHJTujEJl6wNFKb
nlRSUyit5vGkBfgweriVJWTrBttkr+dteAMAIXO6qcAKAjMGTdbgcaL+stgt/Rzw1fDFfyMQaPZm
cJ1LeCCWxhQspytvEEefa3dsjpKfp8m6C5ZG4KNxb1o6r5Mz+UTDgTkSmT7HEKzHEzGOhIP/JFis
pIWu+RPGPwq+BYQuHhV+KOdL2nvn3f0PCmSE5ZgNlTG91KnK0UIsgxxDP6uu/uJ26CsME6QguuGM
OpMqcZshVUkE1QVkRZ2jy3VpU9XI5s9ToRSgw2S0HGadYnNpcS0eOTNsnr5sDE/KYHIKIWfLXX6T
QOoz7Jzlz4T75YPHJsD9qmnpxjJY2Qu7Tsa/FhexAgPYN6nZKYLKWlvrq6S4wa0+5GhA86XaVJKt
iMG92pnEZ2Lh5/4l5bQOW/l/aEL5GaIOr1au4bRmzH/bS9Fqdg5a8R/6E1u2/F7a9l1YiozRLaHX
KJy6wZMABdDNOZ0QZuwaB6PtKz2+f4chLGqp7O6I0zNY1Cc565j3nGTdQzPt75WOgTNhRSlf5swa
BFyLvdM1mgZDy8N6Cs2WrmGS+D+o4hIc/DQ5upHLVJeu1jnrmksIFkDDIW/NknXCcOUmlaQxn6bT
SzJF2dLw71mEvpqA3fKWp7v7FDPpyKOUNG5JF+qkpQMBIEl0Xvf3LZTY+AwGAoIxR5O19VwYBtuJ
QBEUaEBdIn/vCnZTip5K3JaNS3DeK9Y2nglrG+GLFlNQ8s/PWyCJsTdZI/o++Bq7TF2ZIDND6JnU
I/5lawPNX7o6hxaIgyAaRFlNMJRRII1QnhLej3ZTBN1rezhGkz1jFKMeMyrvVNUSRJBv8l7RwP97
F1fxt488byx2ThkR/EIJIgViRSkNR31Ry515KmSyNz1L6TO7tDhNv8U/cFNAA4wcu0ic/SKX26Jo
CaQciZe+bDwWJOcPvP0XNJPwGdnFqua/srw4HMtTrZcLEymAPBz1oCyAmOcIcKOkz1XhWDJRBhp2
vrqS8oUg1guy0LfwO3vK9fHlvwKFPjFaGsby10rz0Qi+8wwdk0sTkuQpV5P3Mit0JMzEU1f6JtNb
B2dn2GieWGyD4bX5GZ+A4Lcqfu53uXdYOHoTb75z3kGn2uhAaaL+9EQfeEa5swF93QAk/bJtVikr
CBCBd7aOPjWGJUyQXRjnveCGgVeWcq+O2Y3twK4O2aFz0RjzIBYNNZibQwrNrVoaJNX2OurYcmFU
E0degu4uGRwl2lQzZfTn1DUu8hqaLH6m85A1mEQP+c7RG10khtgGc4WEH45cM/CK38m6Qmu/oc+g
wG5LBo/V7cAZn/69frfrrSmGiZnuF16kCb8xuhDRDlvGeVZtc7n/JLi3fEiKLFQZ9NNO7PMhAyJ/
nmYjR8ZXvv9GkRrLDY6oXwPeHjPwTHG/+Rsw2ymGMHGbmy23f+zCPdJq9jDOGcOW7xa87SX3hUSB
p7ZDMHAJ1Mu2wm/yrVsgjZY8FfbgZNm3Jc1QmjePAbzzAJb1U5ZTMB9HVkcBwNMHVHnXvV7iuxXX
ITN7QyXlnwNo1XGpZADIEbjFN4BJzsHDX52zePH3pWPEia3udXp4sb9dlGfJCaqCMI6+dBHz+qU+
ByulgdhfkjVpTSWG0Uw5y5SdL4W4oqfckvehgn/xuD3yC/ASEFxxTdw7eVzZTRvgQa8vF3rD/o+s
lWAa9zf1q8C4T6EciwZTCtffoLNEJc9Yauu6KgfO2kLnU+TkNnAGi7xCqBOtrLtl/+LHUZYvmdBK
TC/+n3JwdWMv91WfSZodW8JHuV0VNvoa3AnC1nfAJG4ZUnCSfc8yxstghIkrr+dqsk8DgwuqaJow
v9RHJHLN198MCJQTitoBqgrgC6lgqFKKl4pNa9bONPhDMIgTJjN6kTV+dTVWmj8dptXJq36pp/8e
cVWMA8HSLKDshNIM/kNGORs2IOji0LgvQRypdHmRo5STNDhIH0beXUMZUjAw10/Ksw6Fo1iyxhXI
Ib4tXsytriV8LJJhOgVN9m1TcopN0hKTWgXz25URfc7B8DR7a4Xj+2HkTJoKyAE+urgSvnXY0VjV
d8Wwmg4fmEbk7A5eS7GgQ5jPUfXUScDnXFmM5mGKzUAn14jLS1gdeXeeRKJtR+6pwZP4iY8nW53r
iZQon0Ul3tFCpePJPXvZavSBjr00FQpLaH+aSwnZJECpCfQhMus0EwFB3znY2R7LPC90HDa49vvA
0vLlsRVolS8A6lO6pR50E4MYjpF9vkw0aZOSG8dQjb8E/UY3e6u4RO44HCMhH7tn0TUWJDirlG7V
impBzrOEhi6h6Xg+YJg9oaLuWaV7tIIfeXnEfbgXAG+BOA8syL1vl2L1V4MwjSyCZ2+oWZFumCum
StD/Scrpjbgl0/L/sMHTYS6fzgoF5Pr/7etMWvPKxu2UHUiJ0lm+7mVyZDIrCuY+U8X/1YCuroqS
3+dXJxT5KUg9XmDlY/2ZSUKBeXWV3bGrnVeZ56g+OLT14D2qZye7f0QScMc059/mefmXCWxD5y01
+KA/zz4GdAqlWh3HAdFCwlYzTG/xoKM3EixjSTggygYKRwsnlaMST90hIQR6hqv2Pbu6IYaf7/Mb
/UwU0KShOi+BcQ+ZL5pwYdN83MV4cjN8f1us3+ZRnG6r8FJJJnBiUD0FOgLKHFbaz885Q/mHYmXW
xUrikiltmb7wDHn8AFtI1GEb9JqaP96ejN28XJlJ7bevljjRLaJhC6VCd4UWvAuMuXmYVoCZm9x1
qvUkMP8ZEVmCRcioTSZe+/ccYn+tu2UgomEvbt50ZHC7KnB8f/gxOU82nsQp4VCKc/Y/QhITnpak
pRwpQMeMhrukTN6LoeOlZsbLPgX6L4WWdLfB5hLaroTR85Oa/jbtw0/K5wyceMQTPSjSsC7pH+2I
dApgfTeuwnetoNCo/fHb98Ukwf6irkZ1HmgSTMuH5ChNP0CJUd2VuwrEowW1PFSSChmOqSKkS4nY
PJSqU4mPz27E/xpgFHsQRwZyDGCJ75fs4xY/R3XNWoTjTB6LkKmJ3jYQ4M7bUxJHOR4pU7Ehwfpn
3CTC/y3WFvmd+2MccMw5t6znNeE7l95B308T/46uU6dFsKebIyWxqA9653Wa7hYYcVdFLywc5ZQ5
4AUX6FTl7G7rBy4LA8/H65rnzfaIoBUK2fBuggh4wLTXK4jAqR3BOke/4dD/Eqf34pBT9SagzWTS
n8VOFkposWDdVHZ5PySMibk2QafJ4t3yN3idWTKIjzMbiAByywQc2vd0fvMgFG3EXjjW80d2AQ47
THWDlA9if2N6u561kMh1ADBQVRBb76BjVN8TlMKadsi4iwvCZp6MjnF5NK/wLjYRkoS3zVK/kNhk
qkMbOf5+/9yqvTRW7H/p4dJhUMCvSkL4UxAiDZ6Kx/SZ+uAxbKSyfARR65veX6pr9xhP3UKIg7yB
BLz4RkIzMuFTE5wFTanx8Is/IJc77JlODXdliPRfhdt56NAe3/G2m53wZIW2EwDqbdVwQzk31B+0
jHyTHuTDGogJ0PiAnCNxpv5RVI7bvZkw5fFpHSvT7f9ggInLz23K308NuMnv+avAOjqqLqCDTkQ6
QmDQNl3adVwElfrOkiOEz7fNvudTHvec5iw9n6J+ny82fXtX4u4f7CuAu61dXRLdfRAu4TJ/jFYe
W4un1Fgr0HXAigxHrtsKNQh8zojAFdkIjEUjZiaa+y2f3KVPkUNa7T/McVCn6c4tvmwjjexwalf5
1kmfkOZI+WNOAidFGxQWERSjFJDxO0/8INv0dTDiZBOgemupFYbfYXKdRuhSYu4PB/4qvarzSiF+
6gN6LN0nbBYwAMM+jj6BTlh1wF3DmZPz4kX/tYYs7RGGBweFJj0+HldFRtJvdV5/gUFh51XRPFA2
zkeugCXHQW6UbuUu5ZQscFu7qJDkgS6Nii7qdojtbU0g5BX26ytNRS64p8HbC1UJ9OOM9k6Q6doO
qyfigEEpMr7sfLROy0Ui8IMfWn30YOgYuP2eXW9oExaAfxcGqcehENioaZ5AZgqrquxEEgtll0Jm
5KtEU1G2XylBEIICEskHVxs0Ghyd2SW88VGTdi7wpSsLapg3MDksfKGViTbvNRjPovqSfRHoECCu
v5T3rMKlV9QKGXH41vgGIaprWxuFYWE6P38mKxH4scwWLwEGAPVJlSVQqqtAdooAUhtxLpB61WaN
ch9hvT0oZ25DdoYrIShoNNCf9O+ZcfJE1wHJoG4pUsBK0d4F0Q+p9OJxXEt5XUfY5WVYTzm+U9dT
MAWMwAan2yLIxEsqSHWNUR1puR7WraFTMZJ67b+nM3j358LrBXn6ZgF9scpFMLc0PFxhVr6co5vV
ygPkyA9gnfHwoXIFs8NeqETQQM1ZVk1kwkrsjw74M17/UaAVx8DWNz6QOwcX+/TMZAf99szbXHUK
1FjjV5udDwLuDV9zQxYPjiHcJYtulpNSNYXNYHnEv745QsbAFcaiLdiCmWjQsMEQ9nw+toZJulsD
CqAQHiliqoN7FMNOjv69Eghb0Xycp+uXC1V4ExrbdFgMlRpF3zG1IPZ98Cd1Pyyxb19WcN3mm7t/
0KVAc5idQ/SJjtszXN0sGPswdRBuo2tHb5Fg0f4WoGDDFTRQxcfBOCYTyYzMjuHrePuDNr+gAJe1
6jqD8LwxGc9/68jqzBCIWkAkI2gmh4h7Fj6SeXGbdTIyRraL8J2b5cK2p8TMgbs5vqG7Z1/gKp2X
MpeWZlR85iLKKjTNdGAsvsPmTiDTTX0jVkgVx9OcAcOw/kz/CS3Lk8U0ao99TtGVsX2Tlewv9pAC
L2xWvCtfAvkziTcT3UghhHpDxNiVXUDEYWLziQh4UxbMOPiwZ2BRRXoJTUqtVlgqjMtIjQqIicsa
FYqhm1dwf0oIvkDG4tJkEvfYUR7kA8CT4YaScDWdUCNeTVL8DB6qHUvLqZ4Y84Nt896yNUoQAUt2
uUye7kVEuoWB+nlA1UPd1ogViwLUJz+SXQwwixyGkUhbspuTBiMJJbDmw6bqIHNobskCIKGFBq2f
SKajdUN1CIRz8C2pYBPV4gG5P05xI5AQxS5xndKqVK241ao9wH65J5r8qcth1VbEmZHCTv7IN0LU
QebtbfV8qcCcwagYuVC9OuZiVNZ/KndF6fHgR7t0zRenL1EoNX6E7CLIqMXY5Rt7aXuL62z81lvR
6Hmls2dZ7lLm2SGJJRUaElC80RdlBwzN2ZeffSom1mYK8u6imhwkwbf8ZkYMUZClUBEEezHguGb4
rwG/Fawg+BjAz/4gvZUh0+TKDeFTXHCjONFSpipwoiSs1K4o7FgJkfXhqesi7G8cGpZa7Dl40v8e
KR0lZSmdBuJ4p6E8BEbdpDi9h/+4orJEz+oGzf9NtIszOWLUGdw6+/OZiZekPMi1QKfyvO9BQNG6
KOiCrQuxm04IioDOLsSb3CKlsh9cQk3Sdp/cVzqEandFt6xJYTUyI2VOweoydI7+rLjymE/+0cm+
p5D6IVXaONj/ZXMbL68NHsPWevLytzoi4s9A6M4OllkR9pInGxNCiJDR3Qxb0jms0S566WrRIRtB
t3Okt0JO4GorrRxFggnquMfLogs7nt7wd8m8uYkbZ+5+G5dvU4Sk44SSAwwVHq+WAzILCTyQH/5e
5/7xB6EqgTwDNzy1WE8z8OmK1g6618fmT2ISVBFsLpm2Uf0CyLgImp5KeU7Qee1yQwJEy6IEr81i
SoJcuMUkN1Ceb8emXZhvVZeek+VJ/kjce1yU6kK8m7pooIFZ8Ow/X5VkWTKn7GQcM4I8tz19taRA
eVjF5rY3u/gnQpQDoqe1ejcHB6r8EK1IifsynnFEdjhRlXTm8bvCpUERfrMJ8D7ESBXJhxEkSfkT
kR7Z4/FDicWjTmbChUiIfIyMlexXv0SfWGjEpViyd4/Ug+83Pjzj6AARlx8p6wiAFbbEj+lH2Png
NYwqsfVccn/ZycElrsJgSIhVtJvq5zMyY3oDfHTQWX8MoznChqldgiw0Ofas9SMghqKBcXgHeJYF
mwI2ja1nB0O+Dy4pAVFCQn2YYcM/WCUZsefII2/MOPhkLlSii83/IP/kLcHaLM0zX2BTMLUcYV0r
HvWDaxSO0k5qYdxFM8S+NpNzixdFkv0vonCp/Yep6XH9zbuoz5p9F5uHumaaMU7bz2c3yPLnxZHD
7+G8FaK66vY1Ohml0L3JfIwq4b0ST/2FC0WgxZIO/dhvRfmC5fHtO6k5cYQqU2d45Q3EstG/tJx7
Yuzba2OCaMmesL9ai8+VWq97UjVhslY1VIhrjLdeuOP6SJEbRu9WMzTKs0OwdhTWAFQjsSF51l2f
GDWYrjeaHKK1RHjNKNSLF9kFE4JocU3vUcJJqVUQ7ln9lO3tLj1GDTCxWTj4076AEaW4D/of9UDH
EM9eJv7yyzTRF4WTkNa04ppadAFub2EFVFQnIVweU/8k9X9LWa0QoVKZcurAH/40Ur4llM4Xvylo
v8YwGZyWeeR17DojhOv0lNhQR7uIMNKtcKUOj0Y5ugGbP+SWasLgplXmYf/JdpbBmmO5C8MX2jl/
v1MGSpBfaIrbL38HCn7YJOYSq/Y7lU4Ak6Yaj6EH9MdcHutEUKbsmzWFF5teDixNEAam/mjnVJ+M
RFHsbf1feUfCfr2ZiOSshCx56iqxVQOWlsHz+TLR6augW2cdO2dNdFFxRPLxDCmqUT/gMgY8UVjB
N9h1xztil/U3JUA+R7/scE7RErGWiIhLS9ER/pKwUl+ZCFutrsCQ/NEb8clY1KOzovxhJdJQ9zE1
ZB2G499cNQd5RlZabXmHpHnNiIJDym+gtuab8Wr8tp7/PQacd7XPNof73SRVtpiE4TgLl4jMfJ88
xIamDogaJgK9l+aFsaZPhAHv3K+Neov3YHzau3zRgd58+gyphwoJcxgAbAx95xzOsXydqBj/ro0R
hKbgEQL/oislWsT9ZdU5u3r5SbANWmfSmDXvUvx95zOUmnV4pgVWFocX8NtClBQTv5JRwMrZJzwv
Pt6KI7+DrKnN9hb4XyYVAQZMSBLMSemNN6tYfnIBmg2FP05ewLkgqFlHuq+WZYtOnGVRRc+8PTDN
CG0JthQEIazwb9ESJ9yoq7yMUlyt1hd52HeoHffe/Hw/kmrkp3RjUblE3/Cgwp4yO35F19YGdxDC
iUamKfp/CxD9eGl6NtPZTewbsGUonT5YrkSsRZnW7+B0fB89u3zQJ8ZhD3ZNLpYdd03yd7kOlumG
qpMUwL4hV1jLCOvspc6n8zSc0g5LY7imnhpuPVsuFqGTrkbPe1IlJ2yaLjJBmdrsHWdxjgMNbUhH
F2sk9GOPwMlBH2CmALJB8Dt7NRIJ++joxg+AxFx9ZoF5PFC1Ntp8WjPMWEtLSxTD6/dZFwA9NzB6
U0pmeuiY3qFK6pD7n2rUCRzHevBN0U83P9bnjt/irwRpB5doBjjZgPBFcsKcBqzxpXiCB8NOUbGx
EiBTdY64qpZ1UsMNef3q8vO0g75+9rIT91zSTQGLQX7PPHfqnTcTCkuZjynY6Bt3i6sJSchSw58q
p/5LvPbukp5JuWSfIATeWZgWk/4bbT+m7L05l/UzqjhgpkyxyPmWCuMBX2csipC6NGRnA3BSt6cj
YZ+IfT0BBSYjj/DX8rpv1xh9BD7J/Sy/8vE3GiDuZBgDGLSg8dVrh83V2Bf3yRf92OKuW0IWME1t
+7s4DowAdF5NnRIhu3IfE4I/ffE/MSweXDj76OYm8MLFYmNPieDVhZ5YqKwxqRxBSMD5cFHyXbJD
8Q+KjDNJxi4A903FjVsGEUboUmG7i9j8S56UUeIwGaX8W6LDyVN+hXU7iKOPIhp8J2Ye1kCqwROr
OIVBlmfRjWfzWknDr/+QWkt3NkMFRwd1rs3LpQXGI9vngLmmsEK0zI5nJFRj+Wxq3BpxNa30Qkra
O2pMSIxAVrkPkv7rZQiD+RkGZblSdCPUS8ZcbE1PKIMn5qMe05G/4ooNNoXPJuQs2s0OeUbU9C5Y
1F8Xq9w7YihN9IQVOmOo1pO0tHlaxCRbiW8hPKi3YxSx/p540DRk1sOuiEoxVxLAZsR97JL4Wsgj
kym9IHhV00pN3uKPasKwXrHUF5I4Aue78qRwc8LO9mlEPcF2lVX3dhtifur/jhKY0qHh2YYR6xXq
FMrSgb3q2lh6M+kIIbDDVBSSep8KetieEouReN/11NFT3Hc+jDUyLBj0Rrt6oxTTl2zZ77QtSGGJ
h1twahhYjgEYXePecyaVfRdTuj0+EQ4oo6BbuVbhLdk7thL3dZ23bK2cY5YIya3w05ufqOpqKNkE
bUbj9YaDSlMxDpUFL6OYuMTFRWdyyieEv74oS2J7gAMpVoQaXR8zFjq2qHg3SnuXXJD+I9cgq3xu
OH5PgL3QdImCARBzQcQR9X7YQgHFvDnOr7gRxe678I80e1Cm/3+aPuRUITbzfHHhNaW2QS+v/SEH
8YeubEgyWTwuuMmRHoWAzuxS3e1aud1OA6suhMWsXwyvWNRlVJEAu1i0+RvvR2FiFQ+Wc3wcpV3F
3ElcQZ52ZAlfVUg77OlPwVETZCmsJOHtif6cHtU2Kyf8WA1v4aunIJxDFZB1A9Fj2SgCPPx6HC8g
98A+dq2+SB9e284ie0g8Lwpvko+GufC1Sj8dGrAKok1+tp/qhwFfpGTx87EjwojYt+CiycsoxdTM
1mt3jyeOpvhLpPKkAyS+b/xyvlbA9IY8W6O9Crm1p+WAvK/tqGhI9EhvdmLgEBj5+OI/dP24Z9Ie
7rvm5ESB4ncZgxrc0Uhm73+BE5rbXtsyXbRJSwFSwEnxpu8sClHeeNyKNcqLyx5BUQt9fhqFm0zA
UhkKj/ht6s4DbDWcOWS5+dR5F6gEQnuJcan0hwQWMCt6ehBKJ0a9cpJ/Luju5DHUm1o07XvcG8EV
AvNHWoj8S4plEVCb+tqqBfzFTsLp5J3angCYyc8tDWl+PFEx9q6ZIUoPVGzkPaV7CUX0sdlCOO9J
6BkSTfN+IdR/8lPJ96MzM6jDTUd9MUuzubXbk0s6vau4GL0QE5tSDXxMvROju42p1IpY+6e4DER/
5Sm87fQkUcTx3K0V9b0m2cN/jo2GAsWot/jx5ncnXRT6WPPgqv5wcwJ0/ys8FxsNrPwbO4NbcQ82
HBGsYAFgfdCxnqgZfMHK2LFi1kjNk4awoSexcxdqUr1zChNgUUixWOL2uZnzM9ViT1NXGjdFLeK3
kSAAVoRKXyaQHCVjgFgPIby8h4XqUDFNYifiXPQ3dpoAWG8b3UnEtiH3E7PMAm9zMm/JW7bkoXJn
02e3E/57+VbO+39p+jxTRs5d+fhQOS3cIuH8llKyl9hLxpVUIp7j/OjoNTz1QLuM1luEzgfsBaXS
T0FUnMDdiKvG7vGg8tAYIZinAp9O5+2WzExYGTupIRaZHgz6ec1l9lfnNXRdV77u1qi+kMcPzPfZ
+Tc0hMgPjjEnh+xpEgPeNg+uauRLv3dad90ddrdzYkJe+l9zbp8edoO6hQ3H/LjVPjGWFiVuF932
4m+GxotIE6U8/WgqVj0VUpV2x1E2YFgpCVtebPxsOCjIy51VtqA354Mz7mI0Se6+g9DRbvDjsb5E
DZsr/3PUTfui33/s3WpIkte/LUR1bAx01/TXCjd4L5Dz5ECFApxJujzq3ZRXtKQwUWFwgHXr4N/n
IhtRAIpd8JqBH5f+z1rlmPv5k+kcyqsBdGP30gKDYgbo4i2EbcQIkjWH1ySgpTUWvO+qkVCtQ+7Y
CaLCrWZ4+kpCD2M63WjE1297F8DgfLgyHMtRy2fEB7+fyCYojoZWaoczMC0uItV0fBAQbCrt4SwA
TDcoBNpz6pK4HlWy7xI7yK7UgJk0Vml710/uB9P+BljbK6vJJJqW+pXH424syeWUwRRNL8b6I3qk
s0CsE8gzkTTqOm16DWRpYD43d5wbUWmAyKh34wXHjBLypjFrFZrRXyC1AJrcMt8nGAjRUGmOsbMh
+dY1EOpbBouFnCuIEHC0+xGrV73pYFV5vwMl7eEL2jegLaK3YUFv/NCS5Crjdy1mxQachb2pKM9B
3e7n46ADjklCsHiY3WbVeTLSj/hOMYK2PlynUX3EFyX/xR+5+rDVeicPKh3ghHyaRpZNe/DWRIx5
eD/9B78b1d9RlZ+mbvJitx/35BbJW8VCm8AJfw7dffYRmwljtT7cTkkR/7mvn8MnP7MguB+61Mf8
raDpK+2abAUOlJSbbTosfSCRwWTYFLMDGzv3s5/3ZozvZGovGt9NZK749/y2qngJvqG+vdRWDiCs
cuMR2kNr24FppC8FNgFNwbXsfM0F09qj98bqcvn9tdgbbEiTgxMqTKGEzObWIsU9oYkcqhV0MxSO
HOpiauxuf7fLbHEy5YGLCPzIubaPts/6nHvfQ+R7J0vXNvWmX1Yucqc2IO+cxEhKR6IaPkse0xZF
p9b69TT+bW4uk3KMX+T5dIC2E5bYdJutnK3DVN8mn79hynU0Z0q/zxdaauNb9XoXD4oiZ0sWcYrR
FNnHuB5Q60bmOtx/dgelO2CaKtCRG8YaZ1SWry2EuYnOq/OR3t002c+H74EfCxciMwNgdjH+KGiJ
fCQvyPgIJ03UVZ1WSG+Y/Q+uD1GWjmC4iqTfEEJSCDZ7C4kvXScRuGzkrSjOTjUyG/k1RAXOfHdw
sxu+YxumaZu2tQ8dDqyPdHLsPewqJNz1snga/EoOC+gRn96SoevnBpn3cTOXR5s0sQX4pOBx+boJ
FqCfWGBOgq/ypje+/Zlfzyvz2Z6reMSIyG4PtNtJ+i1udC1T1czRT8dQdfTXDbZj79zCLXElcrDT
Qh1hxz9RIIzuE1ioHHAtr+Snxjuw4TjlBu3CYMMLGch/1TttgxTe/MKDKHQIXAnNjQEY1y0HMkdY
oYfqWKIoh7OvkkBFUWGg3g+R0qmSQNiCxLyU9m4AMnz1mts4lX/aNYD8+sDdafNAq89OFSr1A8I8
HCsfKlbT8xUGdrla79lhKAq6U1dSgFWLsdbkobNb/avp712xN/Duev23X5dIyK0w71E3hW33WD6s
3eE1sTxZ/OZPMCu4nC+k93yHAY74HztocSKtJTao1Q3qx1aBGDMGJzDTRnuL0hcQuWHpHphgW/5E
M7A32vKySjV912hzKBedck98YDo6WT77gyrcI3qnpV1NCrG5q1j73GZg8zYOm45GlgRg8joaU1AY
+ZBzUCxboV9HEq8hiPMuw/SYMmTiBj9CweJ328frVfN6km+AjKvD7ScedGXIKfFoQrfTUsL/A/1w
Nj3YxvTTewhrOa1fsCEmPxK8UjcBFl97MCBHwbNgi89QWW0iC+4RZ0gPUbNW4+7BY9PFOKt4TJyV
xyrCXGCcGoAlFKFCjK8PndXiG7sDant++VDRqUTyD4vXnhRJSuGvjM+AZ7usfnO5Q3R1x35h13un
0V4Ac6kIsX6TmEb0iLNBOfwG68r+e3TAVJhbqNN4Krhp5abDn0lqIYCDbLCqgYz7EUIb8tQyMvwj
Qzag0byOf3GqcMpaRIzU6LIj7jxT9+ZwlAha4QH7XBIIm9jvqmVGBi3d1U4osh/tR4W0inotPlQe
kcGY7ti8NIbMfhOvTy4RaSIoRhaQ3yCcIg+7ahJ0vlR7IKVSZm2Vs9NPZOkFqBvvZXKZg4k0+77J
JjBXkr6NO6Kn3qZMCaJesxJtCNqE8py138SyvBqd4AfiAXL/TDRDvQUm+9MtRQeWTUZnSBlGNaX3
QrGKbygfe1kR5WyEnKw/xodjUikBY7z0V+ra0U9n7VtSdKWJb4/YwKNwzjMj1Iw1Y9mmKEqVRtRM
DDf4c5HQt+0hMAQjc5MHRIAjuhSP+fPnCSJNwRCtGaeAN9vFBo2bg2PKTqWQNQc540zbL+3F7Pf/
i8SiRCOcsfQCDJuQMlm2qilQLoNt73m6sof3RkkrFgm3GNzqYuE0bbVovsyKYcTooPSv6s+4bk6V
f+3hWvFWegYaf35wWsvRsZd2RsFYH2NVtgUYwx/Qpa3+Fhg1QFtgJLwv5NqnHuCSKl5KVScn9EV8
UHzlZoTJ/LXjps7EA9ZnSwmjhtZ+UCryV3+ZQmXW8f2ROzaEWGGoUVJV/u//kan1LG3b9Rrn7vUt
j1delbA7lnCY8hJgEZgdkrQaRACiHFP9J7L62H+Zd0t0UC/ynsZ+vAMR8Z3eh+whPa+R3i+2CDgD
Xv2uvKZAZ3uwEC1Y1v+vOc/J6UwJsHN2k4d8PMVSwhc/zn7RiFRsRszBxfHCVWcjvv291IiczAAw
4qaS2BgoaijEXne1en7J8UqjHXrRGumOYuEaS3Hn0RM1sFAIlvySjct5XUOsHamrSQWwfvDfD2Bq
e+qjIs0lVem6P7D7DYFmCzMlXZKMoai+8oZnk93t5IbN2yb8ljNJEokBYPYC/HXOJRImdgzdv2rC
AdCKKvd3hEdM19cBKxyKy6e1nppItMLTG9lq9YwFEqS5eDXRx0n4tcI+pUK1p8wfGraz2CjH5b4X
nspWLyaNnF5+ZqB0npmRjfcMxTY/cciZfV2Vqz5/2rFRZuD2ZeVA+VxTkkhK6mweVfBmziYJkjo2
4jly1BFCav7zAlhJrvJOF7odF2B09hD8o3CoTWzu+1yIGv8sNYvAv0Uf1koLOW/mxIWKPf/0NBtT
qtN9qq+qqrkxGOtxOgGn8OmM3oKfeXuxKZNqguIWWXfbqQalAxTYikOsyTQyQzNdbVEvpXl2flE4
ZTvhrKORVfm3ceZqvhPuuXdaqyo6Qn+bl8kPheYyJHU0Q6OtfBfYlub9YcUkvEiYNO0hBBJheKTY
O7v5fb0uXbhqNbQmCKVH28goz0jRtIZm/bAev3PnDsREjxSoodZaSQoWUBvJryNQ9xVLCgFVz53Q
Hco/5mjr95gZOKCViwvlbJmEbKGorWjsuvrcVqq/5ZEspdM2LLu9l+3AOq348otDYk28rn87kUmr
6kQQWiUoKYRHujWLOonVQ4X6AYHi0inzxdUaWPtL1tBsaVyr2HfFr8fEfVbeNhN8tXR5/GbEdI5b
421Nlc8E2ppRfcj17WVHO77Ahf0j6zQMCAI3YZldPV+uYgJFfCjpDx7dX73NDs1BfiL/7RRjmRb7
iC6MEaW6VabxPMbbsl/AmNWe+F9ip5Ayxs12P6VVeDNnnOvWhU6WdlrniwtJW1V8t+x0Oxphgf/8
+dmKmfE2tSszNi9S8wuFbg7ppcYcu4O7CE7VuKlDzVI6zYTViaaianIXn3N/Wr+TMyR/6dYmOpyv
LY0OTOnw/GAxW6pD84H5KmvGIZY2y1ta/CYT7NjSNAvB/RVX95SVBEDSjNBsYeHZs8+cYS7dj4lL
WKXJPc6uPAhCgs3Bcz8F1gN5MjMr55+HV/mTH7XmSC1d5rHZK6n+vljJGHbGzbOedUp3qva7naVq
EUUqjIYvir8j/S09mE6e3pqJ4ZDPGeRrtZMMORyP/aMXJjODYcdi3TWLZnFHeVTDFsRv2akMrEXJ
HoReus0Q5Vy3SfwP5yfZ/1VMrNey5SVzJyP+NWnwsg95x4y5M2fJFTBf7dHW1rdmU+0HWead0xoo
b3AoDp9BmfV26OIXHDFX1i0n2UeXv4PZDx8qPLG7Bdxc7ReLENrTrjVAQSl8gv12Yp3yUc2o6aRY
3nfAeUP4/x/RBdD16HOQHj9dt2KC+ecBIWCDvMh5HjMjY0k1OuczAIggt5jLfQkDgyL8fo+gdIyf
ioe1cDd2q6ayG/574/srQ1+lWpx0BSfkltTEEiW0Zrs6UE9yDqSNrwPQewIW3gIm3yQkEFjyNdZU
CnZIYUZZ4yG++uLri6jYhdUyGFJxto8bRtGqQERGOoIFwGPyucZha6z6ERD68/mFLL8yKPwhCRKr
hh0y9O5EDOJOkJnW9RiT+HTeySAGsbcXlDBxAt25o12aoF7JhIcK4tT+fwEksK33Nf2uaCnUkD5Q
ivYSQhWu7+TdCyzBP5l5gILjxRfuulWwldXThVLkMdfq+VbMdkIIvlNw8VhgkF/pWZSDrF6jkuXa
mi1B9rH4ILGI4tGjaSa0HBoGOLZx/XUJ3CYp6t8KuDWnzSwNkIuv2UYf/ezFdichBQkXX6oIS4Mx
tVHUjodQYbOl4imi3Ire0+uDSb4uzGvZvxQDpWvxd8Vs5hv95wC00Mj7HmyQX4ZBgp/awIMxxGWX
x0nO3cuStEBi2EgvaZNwjbDroNF/fBfAGaA4wRqesrT+Ygj19Lez8yWHjX/VKgFsFqT0JxCd4HLa
Yq5t7GciRT+2v2vrMabOm+aiU+Xwour8o2R3cGmuItqpW/IoAvlSTAQv7AlfofN1vh5zdSnyh6lD
i5UL9YNi94XVJBHhf+czYINv0t0bDAnKZ3ruq/19XoskBGWVelEGyMjlkAGaxcPMyE84t64GKo0i
n/gsB5La47+6Uym1T/lBRawRORY0BgXof1RqD1ttRr502oODrbbZEF7fAL4AjYMmImTdjCInvluV
ag3yC9im6cQD7hpQ8FYKuEZu7kZNITu50auEe7z8CZe5n+5+R0s95p5IKeKByZbBrAt7nUeFYdxJ
4Pcex2gqwylb/FcIoKt1O0gR7GGDa0j5DoWVFWPwhADdUh5hcEvtTPG8ngrVXbYAVbdGCt7oa7bV
/vTpAS2oWiRn96jVN38cPz/li2FWVfWn8ZquPLExLs7iKxTgGtoov31GEyce4xKz/7Jjg4QZemXk
55tXv1WO/8rlqNJHDFsbZNfWfS2fOzoDjzyqnEWwCiZvJAtcBBvKxovHt2w4K43uAYFheg7nEXor
fK9TF+A3D1pZxh9EY++SfVmlpFW+Y3pUMWUlQg9iDApbLGw2aVM7ugUoFcuvTpBc43z9vvRLiEL1
OK/McNOLl7JIcAV+UfRq3m6hzXQCgRJKH1hwEftWvcNatHnS9f7t/uVtZGkMeA8Oo/AZQ/ok7z6q
sxmEetBp3AMQPGDIr7U2iFSH/yicuoOYniPzJUp5yav95wJAgj3ZUo2L2yc1FRpii+sv97TIg7J8
4mYcJ0xdLv1YPj3+e4IbvI68PkAEknDE/7bbqMNNS3xvAHsgPIX+QetUXFE1Z8rqpjFb5BSauAMz
P8me2kmUzru6eHf5zQk09j/rNsHpYTtSP+vDYy59/gWsYB6FsXWruNb9EBoXkOOLmskPLxYaxKhj
l+D/C5iJ+UgXMSpwEpcJ71TT5hWqs/a7xC2k5IFn/2Ww71hSxAJOLJYgm9cgODJDL4WXHMY9/9S8
j2rTIT7c+SifSFgKgdN91f10kvvXBmAChqmOiRFEqaxxO7phnc+o0VNcwN/frSiyaopaJySwEJAW
SxVStUucdLC7Pw39cOmswHfjk3MSH5snxxD1P35NTrNmZnmUwALtkVnGpBo/6+LGkrq7lGazJj1Z
ecKb3XAAIYS7xY2IuL/F8wD4+mLIW/BYUXJ2sLKaLVvlxvFN1Lmw157MirMLKLKwZxy4kHExcg9f
TAPk0csEbn7h+GGaLzlnQi3aQ0iaq19VlVT6oX1er4Uy5cijm1iRIJY7frsd+dRT9NvOnFpKZt2u
+ku1XslcG8FX+VJJHs5X4B+ZnNFaVsuiC30ESJhowUu9bdyoHV6CSoXa0CGV+nsC4AnhqeOeP7jz
OVVE/qyUBpujekmC+0bO/ij2Azey2bTQwjHH9zdGvtoZXAJe8xOPh8m2oLDS1PhzoYj2KY32/dCj
jUVakd6hLC680MiH6xnuDklVobK2ykMDzfOcuVkcjpnxskPTmfkca3Mqa/+keXVhX6Aug4at5TEz
HVime9rEE9th/E2RLuSZjCpQim4r4LuxAjSatL8aaXpmajp/WwgssdH+/HI0vhsezIMhvlNrJFUE
tjI0v78bg63JoswjQrT8XcDd68XFrp12St+HB9Gt8cF4cVcrCTFLvnj2br29sRFHT8vQkqePIwQG
cy5h3P5Nq9z1kV3str2QhtS0OddNWlbEx1VrIp4YNB6oVrvI9xKiY/fmQ/pl/6nPjyHjdW/SSKRa
nydi+hPTu+fJBYZ4E9Y9SEZyGFJCh4LjRB86/a3XFjp1CYl3zyMFFWpJyNqhQzCyZOomnlFKbF1Y
YrMm1dnjyL0m6inuJO42cknGRIb8O3dADy/BkQjybzTOq5bRpPX+Mc51zKT+5g9MaD10eqrNG3aX
Un5z1v6P40qXA0awdNRauiZW6OxKqcsMy069TcZGc0Da+F3ahrrbZPHpER20+JLJDtMLm5R1gzuw
ScPool+1SjtdUafUQNq7WSvau8xNFMQVaiQGA/efK9niTy6VPP3OJEImZA08nLITDSNcXFZk7OnP
8dIMGHiXv0zETCqCecagd+V04ny1+8DCZ6Js5YWwRqZrXDKhTBIf025hTW1tDSLK6/PPTqxcHTvz
wSgFMojxNEd0NfamAUKs34WJps9ewAQxun/e1gt6D6aXXrx6GtBu+JF6XMU872gMZtSEM+ZtOa+o
DfbBrXlZSz4ifzH5MQ+J7Z5A5fTMITXAbYaxJ1q7Tu7+szOQ76EKnS1wk7dGjGt2pZDj8x83Pjcc
iHA2VJAVGgVYf1Zs8KWRJjc9cICH/xy7+HBil42lAbIYgoPKScB2B97jCFIsd3mQ6gaf5xAw+Afe
n/erct61EixltGWG5TAVdtIf1r8HIDzDfhgX4/+qAHLoC6FA6VpYG3JLrqo+gOJcdRB/VUSVRCMl
954xQB6dJqEGyjBGUhz/uF6vLaFctyMUbFBf2jGeloFeHQ2Kg7ZAl0MK6vvm97o3XqNh7WY9cqDY
jOwNOQ3O7VTAgPwuVAWNwC0lhL0F8ZikfaScux5aLnFUQA217o0vXHrZDT4DI+kU9KQs+v9rr4q6
UvXOdPrHNVbZtvScK84UJrnYErxqqxHAdZxGOlW56X75DhpzEJDFocjB6WtUo5WiAJdt5ggJFfCo
rUbSnmh5mux+9NHOhK4XjChVby2UvyQTV100zS8i4Dsfq3OyqtuVD4HM+UiBevKlOI75ntS2SmL+
VkNa1Y7PFx24dIihgzqoD1t5aYcpun6hWuAoIb9apgfiY7bEwJw5qM1VGsTTaeBVwkGjSuox5ke7
MUWD41i2qLCSlQLz6XoOaEbBPztD9m1wuYg38gGVEoj6Y4Wd3drgn8M1TA4w+pyequ5mharFRiD1
y9LLOBi6C9R6mRIOBcklwirDRKNG1TYQvFuKX/+KiX6CE5RFu6hL6vea3SHlP1B54SGFzGYWBasq
xY+o7C4iSXbHKPYN/A9Ry3vXs0f96DKd9uBwUp1pFOt12YXLsoljcet2zxyXkPOs/t+ChT/4bSg+
Lljx+16DbJ5yXXkH+bOymH7W+IlmTsjY0jzsdykfU/CWgNjKzsaApvzzUWlzH5V4WxyZHqvAfhF7
k3ogL6XFe+FYMhe0Ru7598ZcZjuW4Viz7ylwyVRj2cfqUZE3m8Em0copz5aJ8JY0hHLCyAXGN4Yk
6jC9j0eKwFMeukT9vGHk7Kc5Z3Z8Y00xf94TVmUUpgbx5SfBhIYbPbvnIZUcddL1ge9T34G9z+us
kxlu5lZCKAv5w4eaiJzV58q4b03fkml9RQsqRxWK+J4pARHqUj8CLe6274g1vUouso0Y/IeBU3nd
UHOpTHIegyU5ARZWiPPI0H0azALbZJs8hkPzWQonbuRnU8l5xChugbdm81Bmju/PUq9y2QMGRa3q
4BdTA+DA4/Mh7NwnfDBsBkvrPXFt6xsc5TjI65ym7MQwYVp4o+O3jy4T7ScW2YGHdTquJzX4LNX5
RIiC8x9/tOU/XjZgLzCEtXg6crxse+5jaVxUdm25eLUuaHwZf/nq6a5Y/mYIgjM+qJES8KmeEEh+
ZxgS/C+YX6cHqn3q6UuMq5WhQiS7EnGwBmdU/6Or7XUp0WEylN2+b9LKeOy9CaO5nO96NU2X1/xv
ki4SkRLdytISu1ym+mLTFkpkny4/7oArqLR/UrptJA0bJls/j7/BO5sPOZfZTuIc62L1wGtTfUv1
T0SGq9min1U7/0hnahcHtFijbQ8JZfS5QgsMuFlSYWBletdq2YBpYHUPH0hAUi5FlAAseo6ywlRn
qk+8OsaKi7kLAh+c3jFFsbaddrwu/sYLAuU/hBwNGe5MToyxvTf+zbIzftdpC7DDbthwqwF7ljV4
J07pH1iLnuQ2poe/SYgd8S3iKwhqZQjrWXY53oVHVVoyyey/6BdZyKOqPmkHH4AHcxHMs2sIp0Oz
Mpq9vq0EXJ7q4yKrM8Es6PtF1xKCq3YOJRwUINd094clWnmUefGpk4T9bvLBNdm7oF+28nbAH4y6
dhfT5NW/xF4L+lCDaqkmG7cl5tMp0B6cmkHhJFIaWizOuKkdrksHKejZQol0If3xSbBXK8sKZg8X
olWTwK2Lp3u5jKQeQ/XFht4RXfLB61U7mZLCFWHu0VdnZMt48O7EAKWboiDeeipwoDd6KRjduysl
Thgcr/mq48xVvGLgDRF8s3ghzi6DJpphbY5IuZo7EiP4nTrTsHSSoPSrUMaAZwAY49KPNvTDzOF/
95uGv77R0wpCpqdBihprrqsUcHvBH7ZkFaiiEXOSC8Ajob4m8T8ERFq5xxE6WytUsSFMfoq6osr0
ZYKm4hVZvl3DPAqZuNZfuc0B7seKVQUHm0wTWfvw5HegajZl3TcD3JwYUwqXRM+4VZhvO1zzBnnn
inSt97OjZ8nri1usil7ydZBV5k5rIJtsBoFkMoxejdiuV/grct2fZIE9Xud11/cUoslbdzZzwwnq
FY+98avnQM2qs9/kvtjX7zi74BvltLq8o6LqJobVDak4uqkU2bq4oczxkxrGTB9b8ulU1X5TdvZS
CaMoKpZHvvRcH/iCqtcTkUqK4TM8VQdNhAtMFEdE26mOA0WLEWdXYikqLY7ScAthwqTYLun9VUS3
EQxWrExJluTvLn17OE6ndsJCthU9yAf5qsEke/u8Gno5FqZZBWf0NughANAY5pKzshC1GvOkxylg
Xn375mBLwLRwQTpwc+XXd/pUkwioNnquX3eN8HUz3CPV80o1V5Z0Hup58dUhGCa7453OjTKJFLOu
aq5whMKqqmgY5ftLUOu/MkJz+KFSHB7OScharSKBzAm3hHs3vSPGIJxZNkrmIe0OFbuaRvDlmhfi
zOVaPSQmjnEVxB5Bu4ZjQN66a4iqEa6TqFH2z+mw7qeQ6a+PZi1gspeNzD4YWbM07eXi4VNVJdGD
frPHi1HHlc0S+2VzWyRjzsiCJIlqt4iLahaDxaBkhhuPdj8zSZHz6snnyL3VQRM+GJrP3Cl0HgNr
8+M8B0E6/aXoMaFdoH7Llu9N2/XmYQkqqTw8U0pXF2+SHfVMk23FiJevjA6TMKUlcnsM6O/Nw4dG
ngMdZk3jRww7CLuQSdowhRCgfs4CXYksB0Mq5+DGeWkH2a86pkmeY7W6XEgKmqhCN9tTMIaC1Lwd
H7k/sOvFDcLFFsbR2sXsuRMAe1MNsdJqpfDhbR5musP+AEceo7AtV0vlyqqJRKoWqe9TCb+lyhAD
HMISOc/TlsvyykX2Drsx1bnk9D73yJVddNjuPqAgksZIRmF8MwYELqN3ZFZj/ssfRYXvbVIXPg05
jD4D9zcg4S7etIvQGTz7xzwpmokIb48iayLjtAw5/O7I734nDlm+2VjHre2uAvoXfd38cx/7LxGb
gmZuSct6KiiAa8nHViWm2yNJGj36QVnVGs3oEWBUue+UN/TEJRTrzRUxzueP7fhivqD4Bz+RulFY
/IC7AwvsAyb6qo0E4wfDoB0Yn1zWpqTRgXdgj3tAq1d84VQR5YjkHvYO2xS8yELr/KWExNs/bCCJ
K8aBJPWr6XGh1sZzW/qQHG73F+utUN1GVn5DPnwZyvYk/3Oo+EM6jqg9jX+0MRcg5wwT2xMi0dW7
BJ8BtY55bCMTqHEnZbg89QXEIh77yDsL/nNtc/czKlZG9OzZODwCPmLCzPTPCVytvkwhrWwuEGY7
KIZ8hCVPIbVMoNDyLZ0Jx1ly2A4MdIuXVPZalbgwLq+rkLucKTd/foJv6k0qB9OWFdJgt2oQIWiE
MPW42cF6/QCbvQ1L5aNh6JuX9835klUObRqTFiMvsd/fpQVC/4Cwr0p8GnCj0mf2vXrDGE8fyLYP
ZuWUB0JDrRxcG9H0FUBlEEq3+KM9Bd33R/DuQqknLbu2dD5KZ2GUPh44MEyYd4bIUMeColJ3S1Ep
L6d1H4TalTjc8BHKeaOJhFxlDVVZCP995YFLkpnDv+VkILVDin9ZsrErMJYEBfX060Vk6lKvMvar
/eXA5Uynhsn+dd+0bDAiyZ5asJMQziLB8cHHl36V8A2JN8khp19NFCbum1LdNTS3+EyOwGFLmzRC
PIE5qYkrQ33s6JPAiFwj99U9prNm+vH8m/+w6+sPfLz6NqkBuSLx+JymueBUXYS8FwlVS8EobkXf
FplHm0UlMPWUsAHAGrkbKxfXpJRO5d0HTkI7lY/0A8uaq1v7wSa2OKAji2MlgdvBIuIQGTBTL2pB
Ia2Q+t75k4thlohcIRx1gHRqKWkGM4fCSFO/idxcY23SI57OJcjaF2i1sRPD/7ARTDWwhdxlxjeD
35lm9EvJDS1yJIqYoR2xgz58wOB4SejsUsFCDjlHBkRC787qPaZbxt49i3EK6IisACOz1z7gGsZ7
OR+KTqBo54K4tQJngpXV9T21PkUdfkyIP3gt70YYWWHtFlnPgo/29b3K9g5b11Wt0gx03gYqp6Rx
3i34elPJM1Ww35iabv8xkVye/u22oDei9G1yQ6qV46kClcH7A7ARZFC027dxj3Fd83DffUh8yXHr
6gtZ5TnKMqExLHOEOeY2bg9kkI4NPn0ZDR+8SAM3jMdGCtRVx0Dy0a21TL9pm8gW6Va65F0nWuo/
wbt6A0RbA2HAi5wXTVd+TAFNS164c2RFDwpqXlOmqOYqzPG2JLxPa5E6QHdrV4jEPpG4bLElCrNx
Wip1Q9Qpv4gYP+cH/j6Bv90mod5ZJ85MKWNFR4sY8Czqd2NfRjyI6Z+e4VomFrBzMaw5XVDz+lBy
OUOMrd8ovDvj7un1WDN0pY25S94d3qj9U8rKz5babVfDRrMlKngu47yiz6uUaHH3TL+/faDAx+qM
xHOPbHYupVQRnvJ4zSFPWXKoKZKlNnXgVFDwox5gn/d/ozgKrEd2W37z0K+wTSQ8CXwhRY8xQbYB
KBEolXew5j7C4XUeo5hDGgMyjPSheHLsb1gcJWIHpKrzy2/Ju4Y3qt5gJFSnSrBZ5cjhZNDW6y2k
dIonLsIFqo0tiBPoSbxIOqdQeDWZgf/FZzviGlJ3zDXV99yWN0Lccn8H8WTyHLgqBFpCPGy7fcR8
dfUK7aIASaAoDDwqtEMKrrLL8ztl1+Xkh77KPGIAShi9frHqmHSHLPwz1++dLLVeK65Z2ow8sHtx
u4ODw8bA0S/Mr5XM1Z9fO/dsvjEsf/uDfS43F3Vzj/9Ua8EZ9U2QdPMryYUiDsgj3hsHEWbsZECz
Owe4nV/xqiB/ATPmyDZfyHo3eYszekFrM68PgrujAkF428iJeztJ/7JoipNTNdYS/jCJrcvDUXQ/
GtzEomxqFROzsASDFrwEJRDSaYOFphKMq/XGrOGo/JP19uUdyCBzTd6c+BhZc2n9qlw1MpUmMRUp
Oq/bHDrVNi7xfoaPcFc4G8rsDfRYrWgg8BFWEHkHyGTeJTRhWtMS4kt0I6JwGqd2dVlZu9ClcthO
7vBKyVJPO9KE8EIC3vLS9Hq+thkhJKEf9KKa0C6wGgy/dvvTYcNFhO5ovvtfEevTkuAeMIbs6RCp
QUvNnwwHU++RdSdXf+EJ91ysytk6El/WrzZ9x4inxIEmpid5kFjPJl0rTK6ooXnq/9gTR4/r9aWQ
mzcWGM4OjNCtCBE9px6ewF5sPMBDv0qUF1FhvVKvu8a70fig/sL43a1oKSWwVFy4jPtFIv0q+tb6
rku3H/Yvvsk+o/iDLePPooSAWhQGelMHwHC00jDc1fDD8F/Ztjdo+ROHqmStRtqMstRvAp29hjng
+Km58HIcaWijrYEk7ommJH50XEyaMzfdbdElyWsuUSwMn4S06d/S77LZjD/lDkSpUgjWGGUsOLWK
rAoLezA4HJjCrpDVKL7QMiIGnS3+q18alKHGntDDmCMWZeNR/iZyzJvxqG0WgIK1xqAPevyxWrnS
eWDikH1bl1nfPRYB8wmS695ZC0zcQHpU2VH0Hp0hnYmB9XNJuM2NgzYmOiFmX/wlIVZvg3A5celu
F6I779OXi8p2+NRbrjF8n1r1ltyxtPPRm59P7yaY+gndMQmpQAI1C0dga7JNdPqfL9RRvt/lZ9gF
+uTyjcYMn2EhwD7sy2Huhc5rAWoPWnaYO3y8/zISRpnG5CITXNQfZJpc6nIyNUFkdi5wBxXA+dRh
zXe1GSoA15oTGDWLzutf7tBvIAdp9Zxysmt4/7uC8re74SkOLoEa1oAMSaYp+nzMSBOoCAKYJ0Yf
1KKDDB5yBNL5C0KyvP4KVGwqwBsXBx9Fllop0+sZQzrioMWroWGr1pYgmehrWxA5ZOMLTb2Tg4vl
zw7hwxCltYpyiM8s9EFZ4dHM+6gdYnC/rzByRL+R8Riu6/68q/YjwScniBp8x5EsFA5kf/PHYx+g
IxFUx4AtD3z5HWrmVQwZBXhE2LwG1jhSazPd8byohZHue/AF2jC8jmOgLkZGAq9NFKkeaLzTg2VX
tLhW6vqz513RX306n77ceCkPs6x3uWfl++NTBCQd2nhsnOBp6BNEIUbvVV4IkQRAeDx4I5q9GUt7
VHJ+Gi92THE/7G6/cg6iYyBU8kraCZmUjdw3RxuAPiq5Z9cr23aU5G+Df9qqkloGepwJJ7xaD/WO
vQTqeIEeSoCcXzarHxXQFaLuJy7LIkjAp2unLl4OGTREvRD7J+PmIVWoX8PqmdOjMopy8FYboA/o
eD52y308a/uB2OrLQheoNJ0dmmLnD2onbSzUA+vipJiIthffXTChr1+8NXQInzWu7VWJvZiFtXVr
sJciSah1uZJteAmvgHqSO1I+lMlXfIxlhRiZos1lHCVlLGILW4xGjvf372Y/cn3zDv2fphbQ6Qha
f1MOOMoQxVmrmfjTzp0kHz/7TPm1cDIerk/dzz8uA2v6O3B5GTE2aZ5zLu77JeDvC72Ye53JfJ7K
u8UFp4Uig+qsvOwSF5QDcEI7x9Nyqg2XGBSe3tV6VPQeHjPHuvRLs7s7CQtQpXZda1uU9kfvHrCP
mMqGR609t8RZJFdXThVCNAmDzeDKX4lz7wni+3tIvDMVW5anO//dqG7MJKZjVg9ZdfoK8NnTTRWR
k2MfpiRGo1Vq1etUXd5Y1IiJa6DbhwZkNPYwAAfUWhgNAfLcddrl/ud3WpmOEyoUMSqLF9dKxOXV
ejUVjzQx+iV9WxhsjLQ0S8W9lpuLCKydAd8MD0498E6Ji1WHpsiL/1zxgmOkpY+VQYWrEjro78bq
rTEnkX/Hw7TsFZxA0/xRrImUre0U5WsLyvFzjqRhXPH9mKlgz+wfMNE1mrQtsct+mRZ5LI3L8MEh
57CdwLo6DDfO4JndTpNYQlBPwMMnM+XZmGlGt8fzqeiRl7yHWjn217az7r78TMaeX9KrZ10njSfS
4HLISVqUdvbnH6Rk1CqMt4lEvlP+r6EQkI8jJmEFVmXZeuOGUhV3AENE4Sqp4Ou3fm22LSvS6Psn
1JDKy4dYuVQvgLnQH+IQNCt/BqIRewc6afPs80puuDizm2P90PGqZJfH8CSc+cFAFqA394CGT1Lx
UOdVDPs3AyDjO+pMmsW2vQbKP6k08jz4YzJvcfP/0F74NIhT1NerV+7uxNQVBcCNkYoKsoSb14Xy
eDa29CZTbG/z2dbfrrLKtlUPtbXuKHUyl1jzlV+M4D+HdsHuj6nn/WAUAHVjvAaRB+Eo2h0r+aQD
4Lz41wFy4lzIflD+6zZWwLIt/Ucu3MNu6RKZtApzTatBD/EiZ/noDAUI4y7bsWQZw4TjNlPYiJ9j
gwewl+J9DsH3WXjV4Z97So1DZJjAhWr4ZVuegNj9pgzacQFpfeG0pS9Nisuqpevep5AK6auwcYzR
+t3e8a8jyQmf7R4j0NiFvEOlVDoJBJLQcryrOrJn58DyuRFZjbRCiD27eLs1wIiwtAAJNTvr5udo
7vpZytWekdmElPsheH5yl69si2y76zcLGbNNWtgh1Tu9k83tsDVj1F2Nr+xYH9MJ5CTEo0z67oN2
rNrRHQI61gSaS+i1kFbF3zdVi0fE0gWmzS7iwWEaconbxfcivmhzEi+RzfYRW/A1/NVZF86cfPLy
S8Lc/gHbNxV/8exiz6jQYKPYpusH9y3fANJtZ3ykzERDR18T56exPv67qpwODBsB7OlXYl0gnhZn
cgEtcxx7GP91NOteJLRzRFmRYAxUgvPiIf84zh4cmMn/OhciQxH7Hp8dh+j9rnJZDsFdiGgmpZHQ
kI80ypV0gjXwJY6f+4tFhs+3HmMXCynEvkDiwelZBCQHTrIaLuDvusgfCQdG8USpT+M5DnFHU6ay
aWxxccr9dkzvNhvffF+f5HMq3okrCGYSUHZAfho+wMCYLeOBzathXwYAIGwkZqXB8QgbsYqz0g75
PUP3CNkY0yjf7eWQVd9E4fRYBKwdB03HspRxy3zBzvVwrZuvN94kpQA4SPIHqUq2mgANrqobdURV
Jv7dJtueFycirTkICyT6o65azWDy6xGIAcVMGWNzz6Mf5rqYbqFzNvBq9D2pxI8jZXKTH4kaXnvz
wFCWZWTpi1xDNDnSXPN/HrdMf+T9WzqyQk5DuYYJmn3g6KepxJqSlCBTBSTrKMl7vECSwDGg3+zb
p01mrx6ZPPtk+nX1wFIJpYp7POrEqkJF39HPVLeCkXUWvkSnvyFeAP/z5DgdYDcPiBmtnVKJhYA9
EeMMFMbRyxIek0GgtBb9oRzEzTAUlqHTR8VtqymhVdG9JaCRCYRM7yyZJMS8Yz42NI0uSahL8Rvf
NJyAgyVDZoz1T2WL1QjVngtlLIl2r8qd/V0JWE+RWfNZLMOkmlWkACgY6o6gS1zRMJ7nF4/NGz25
sMx0v9DR1B10oMpylQ3UbY+nwXCSS4pe0w9pnEG1GAy+dE2DUL0tSer7jjfDdM9iztYu3By1hf+J
L+nKbitncH59kZ+HcFVgSS1kadODSjER4TCqyFYFu3FRj4YvqxocKHLczdZAKkL8Hg1ZjPkc5vnK
RqK+34QshMjwmTaZLRLbDwQusBHDAliDuEAeVo71uUl2cAQwDL0Wr2kBWwITUcJM2oq9qvDXk5S/
A77gWL2TVpo1wA1EDlJPkvR32jLcw/SKFQvaduOwVfhJjrrVf1TtZtCR9ghMjNonJKalmfCsNCdr
cwyBYhW6WQSFYZdohpkBxldAisJUjfqTSZxFwo1Pse+AOcAOtOZZztgvVAs1m8RcVbezeCSIZnda
gZm3qezH+m8JGS16aGEcigrtSJgKrghbjLn0YITtOa+c9UcfBVH++SKVQZNfoUQpykZnnA3iOjwm
LZH25JH1zySwMeuJVeK3WDg1zB2oQq7exyaAfTTIpHWfQ95xHvoqygC23JVWchQSbMzM4BaA0zZh
rDAGni1ezmpvEF7zlkoNtZJMimjWtSqX9rLSedBBgxBYTLKPU4gAA+VNyhXGO/Xp/urSZLpwaEXf
T88iujBgfvHCGbx/gRXZJtsq5Jgz+kID9nOxjIAJgtq0oVBfNWhML4RwkLnjRmzd0kww1+ZDFwPi
IBr0EP8KZ3xys5XnbTuraHhRfNSva2ynQGBHp8NaK4txcQhsElAVlFBtdOIBhhLO4gNLxtcjW4oG
J3iS4EQcKszePnSalskEbBQW6MqY9ii+tYy7m7ZYZTsRZEI3fpwIY4SSZi2c/WeD6yWoVjGuZtH7
HvPJYVsPDCwXQ4l1FIP+S/u5L+GC77y18WEDatabxQDFk0XCMsp5ZMCDUnYIHUzpulvjzJMernYc
70vrmpheKoQLES6VGIZ7Rf49TS8caAJ5VAzrCNMNo7CZ0jJg/+f+3SEFPVMLnYChBOwR6Phsb1C+
dHi9m38fkF+KSD0jECSHE/GYT5EHTs/wZ6vx+lwDO+WztaOd/R9x/c6vQ3mBin/grS0aoSy8mWGd
EQ1RNe42L73s+Ba4v9mnIhtfjZ2nzWTffKXGNB9VcqDFH46R+M0enJUvgwDHJa7f2AiAxps5WqJY
7lNIjLSpkf0TgX8Pbk9Sdq+VC681bfdGwnsgM5cBlSyYXDGukyjjjG2G/XRCspet3v+Cxz/dP0jH
a+oZ8vvW+I4DSP/lS+p3yqVI9J2jzrhoCgKaK/OOokwaDLqTw8yJqYp62lwPoHZb3yZnux67Lerw
fiUl8MpyQBDrO7GzrpNNZhVoyZT+ICLIFDYerCmcMLpRsx7G09qUdoN9K90QmxF6aPGjSQhH1FI0
24IU30+eRg0L21GutyB++e0LETrEThlxJvSSlUh3IVTPSlViyZ0W4ZA+xfklIQQjvIaFvH1vt5dJ
+zpUDEqZCmkliybsCIKMpVfSQtIz3rgDlaZJ6g1xY1znd6kA8Uj5Kfws8MZQbkQ7ZEpkoZlzfji7
sDUwMOr4Avif3sX3IAKwK3VIGHMCcEXIm+s6bjLZ1fAnMuMO5abWXxsGVa/L7HDAwCIO/8Xxtbpf
eXdAJlY0sstt72A3Rgi2i3G2R4UD8+Q4Y+L5KuHNZEq8jHOLGBkW2tmhNAb+7tQ/eFccc2LtU7nC
aPbNEz4bLL7OSwclt4KBJaVKEBWuuLt4AXL5gPZGyRBqfalVEg0ie5eLLmW6vZzg0VwOjS04KMEq
h64wHx1dVVZKmwSWTjz/uhZSRG5xyLaQJwGhkg7CE/liwiQ5d1dWdgdfV+hws9tZSZ4ntOF7FD8Z
cjAVCKRfnAesk3E3MCYy8hOfeSggJ08aC6BKuvmAvVWhUrZMJ/YOXQeFVwjoD2jUIEbYEUnh6rvh
nYk7a4H31qi2KaoevwOEEGiWXdwb1kaRxjM6NhFueMX2uMBR67iq+thi6g4hvnyEsNXnLPOQ43Ja
7U5vfGV1ZomuNR3XgUMBA23wVoOlh4U7Rm+AesNYNevstOzuwEjd62xeCN/LmkJjkZa9f1A2QxUv
GnMWekDoaKegfkOYhVOS87IsmXWx1VLuFyrf1hzOpwnsvYO4AbSMsYOt8Mqv5KZFn7qihvMou+Dl
oV3WtTFZYxKlrYN3KEh+ge/Zuk62og3ti8KAdKKHAQcw0Z0tRMKBxf2LXngkLzuQcvnlcuQZGUVe
dLk8+b+Bu5B27epcmJT8wS9xT/kbU91H6BT6iKMZIqtwCoX8urAU+aArZnSRevVcoWREfPsQExib
zoRxY8s1c8SLJQyKlaGpafx7B9HMzFxpsvNC5WYlH0LzGZtIUg8TSqeKl0fWAPAv28jZ2yQZihEN
cdsXhDBTBQA3jfT2LgTp2FDPmHgFhyGCcfvikeyGnrrE8ud4DxcDpAJrPqELkpyDqEy8DBmMSF6K
HGhYGu2sdh2o3s3cskigjaIXI/KUJCqz2IZ4zVBlsTJj5AhM2jA9J72xci3NALcICTKb918VUl2s
37JHCD3dDcDKDd5RCuIxPRGks5L5PY7DQrazvytqAIXXjRLcstH/rsQFaGW0fhQ5HteptS6BIHGZ
148robnAsrE2SB+RCVxG+i668LQK/Fh4sqNmEi4BambqzCD2PY0FYRvQN09dApOo6uk2eJmE4xN1
3WIeAQNHMioU5kbLae8Y5meDsbo8YEYzIUVQaWM66EypWmBCsbwRCrWN2MbMkOu89kVFTJNAN4Ms
bQoeVQBbjI3XKxlVOmkLBTdPMfYxi7JRgIt/Oe27VTBpXr+ER0TfsUrIF5CPM2JwHzGx6wjMyG//
fPjYXMcUsZfMBunRWq/+y8I+1ZhuryKbrL7AkDY5XrzRkkZMHc5ZrRM+DupxIuk6i/e4BaAQ2Ry2
ohy9gmSAoZBSgDYaHMfpTwYAdObdl9TB01WCj12BMJuPt5QRnPpVkRsLBu1LcmbV3INyD/ATWHLm
pEcF3IVNjfQFl3pOj9QifF4piFefMK7U3Vto3Hhkd5+z86fZZ3SajSIBEg1y/T8zVjm2y9qe1lcZ
2W+RtR2atIOrq+AarndF6sAYBIsI/O+0dVJ1oPQXzxWBjqqkilpGm+mjZ3+0kBeyjBkashC4nJRX
qDzahDsPXRoxidermDmI7Yd2L+wsPCsJm85PJEWzWgMhuspJeLl6lQhqmFK346ynRHj2kHigsZJD
+xCuUHNFI6eD1i2XEiNX/tbf9uBha9LidW5okxAX+7sw5YFjoaWkYytddcae6LRITfKathgkVmPh
VJCWrE1uuQUk60QXxGMwD+5nE7kJmgp/O6wuJJ1c3CsA96/ISvCO4ruQrGY2+v54hnLdjVk4npYQ
OhD8sFs01z3ix/fMQrW7xhtBNRTZEbMbO23mSewOzyiS5py6kxji3ap3fMmRdrwzYeCVtgwh/kJ8
ZcKLI0hu2hVDx+tOn4Xr1Q0smDVYwDhO1tornOEQqbqMP4NAK62FjKdVOuUy6iDnbSNHdD0381qt
HR91Y11cZ2Lp6jmCQFj3/vlRfSd7q5JSFcQLVwGFbDEDhHEExyi5N8Qg38cdGmE6GfYCipkA7Grd
OTXtZT6mZi2NRJsO+bPaBITnZgiwZYRa6PwRchoWy3NQaF/RTFgJXpVfn9nwuu+P5Mn6s2G59J3y
D/bX+jvd1ZZ/gtni/g8PSqY7v+I4g2D8sGJj2kYRPQspY/6CdQc7XTDe+defpURrlVWscmM8YwAM
wW/fArPL0krmj/hCBUzulm/yxOEBMRSQSbeSOu3LamluYzxtxislhmxEsQuzLgjYtA9aHsXtNybU
sxqhz+BUz16wsvaltcf7964AMvMglFQJWWfxthJJ6cT5eI/u9dz/jxuHXhAvUPDgAjaBnkMpAu/P
Bc505MLZeF8lb3GC0/tyAeN3bIBdlpOTOQWRn7zVr+7p+TsCmIYHm+vF/bENXXmtsmLSl9nIMAUg
h9Q+hogqptOoaI8vv3pzHOwhAAwsquNcJ+vyYHfHpJtSiD9l2+/pmz1ccLhxbKL5uGBuxEEmkeqW
JCPSDxnUZJDy1dBcNbW0M1kZckwJCW8HuM+kWn5NKyUTqDYau2ZuPf49tQxBHMsd3PynKLkUsttO
HTi1IlXV/zWwSLKadoROt3sY/EFNdkFP4ZJAct5JB0JMBAUYTYjcA7b1jKfkokM93bw1urAaPk8q
nOo9tK/wVKvXjraMcjpKnP9KaGk+l5RKcwVmaJceUFj8TuL0SCkEBg/SG2nepX0bf18OfQeDaCbj
AecLFTq+7953QJ4AkpL2nRjy1P3CD3iQTrOav6mE0V0qGi3OLRtyq+OYyP37JbBJ+lCRLgSs34Zv
6x7jk7j3xU+UYzh1iESsJiaXcDmfxkZjn3wVGmDGe9bNif8qU4upnVKpNTf/FXo7guJn2QJmEKNC
Bvp3JmLPnKbEFrLwSEgDGaqem3VKmPO48VhROf6JPj57o9e4FRV2VejnRleZebmH87ZZ98BlnVbn
x1nyy315menewq3lAHvBv0aimODs/SqA8XMzqbWniRCie6AkAKmvEI/IWl8IGiXtKeTaz6Acf9zh
z33UFlbbnJsjW3+HNqY73M46MCP8AfYJO9wCARNXbqFH5nemjPco79nKktXJizHDnEV2RK8KTF86
Re0yfQKehwCp09G0QU9nxZVwSZwkxf9wknSNS6Y2Jd0WSXfAQMOqeNFwIFuYwYdps6vpKSQzUTCg
r62UHFpq80p/fMAe2lv14YgBDnfsEy03J0hglKngw3x2WSjl7g6ZUNBAb0fRQ7qZIhvzfSqMUW/k
6Gk2mLPeF9JITgOMyAGzXd6nIhfanZuEKmf5NTFRel9UYs/MjkSSmeHaEJ4thotggnxMu+lPXtp1
SIGYOqUMY7SXCKACrxLuXzZxEefV9SvOmdIwQCEjd8jtfkVLkLRnzpYN6elMMLVss3HrzN1lGTxj
MQL5WkF1HhmGXpD/wJYMB5GCpfYdkseQA7UXn1MLwN35OrRczZLDqaOWINcq2n+yoPW9jPmhU4bi
dpIZYeSqoqwG7pT9mWtQHMVZPgoT/gfKj1d5HlmUsZcOJ7SUJds3MnB8kta+1G9wVmtC11NLta5+
ODF1xpL3oGNES7+/FUR49v50IuDFnOAwHORBHQVjMCDQgo6VlEUCw6DAcVlU0NkwQWPQiDtzEl20
LGi+6i2oC15GqEJdEJHYf5DKfOzbU0zswipYymfecFTyWdAFk09+ZnsgEkrBhOiR3R8niKUDYYPw
VoKvwzPOOaT5wWd0cw8UCOaYOzlPTsBmiVtJQFJw+vDI8qE9MA84PoZ6OwU4VWNNmFIv4GIrvmON
eKpMuEmktd9PICzRbUeQ2qhfb4/FLmxsnI43Repm4ROnto0R3blHaePHbnKZNYyLqErPkvWprKy0
EjmT7j574NUu6zObj8UzUYWDxBg601SoqPd1Xrzc2aZneuYMRq3X4k+8MOSWA3gzXidt/tRRweRv
hnZw51819BRrgXI8/n37ovAOvB7y9Ta3+w3RPZJ6JjoVWCOMyJce5FLnQrQF1/d3SfWK1ayMlgk9
vyKySiReWjmFyM4kEmzllXxv/7+VNpclv1wIBbN+rX6jVOuJovqCQao6S5s/gbAxZukitXIuuo7w
pNKR6XDLEyISRQO22GdfvwVh3wC27Uc8t2t2YceP36Q2sII4o7UWAw9kx9A0zEzGXZ0pO8bnNWl3
PN5hob/NZkrXjqBJ0mrln4gA1HdkCQ7xzx267DQi0vvmZBEnLTFyE/SvZl3VAgq94uikwYsfDqz9
jWgJeMOlu6euQq1xmWWUO1lqvSWeWMgObKfGPpyX9zoFKNXg3eMxNQ940b04nYs0HfR77p2NSWuU
+Hy9/I7s2Os3QCzrzNgRVF/aoHRXKT5ysPyCCDFZGiC4C8gPJIgnd5SNXyWxSMEO4qEd+IfTLOFk
U3beCRHnG6VokpoPO47DxpxAKGbzvNSNbrQbC0ytq0Bsrr2KDhII3Tyxm6PTwWUAj6VJIDnqCMpe
kQmw6cXXAmeAKxaPNSm2KJAHXFmunNYllsFNWIcxxHeG6P1MZf+GkidxHC9qte2r72yaA+wZPnZ7
dHHHvBPhDvF+xHMUTL1FYH/+E2IhBAxkVTQaaBox03V0VYG63aY85wHHZJez9cimKbkWaqHg+JRV
duntgxVchJ/k7knTgLLNduibLClHpFkGpVLocepDG90U6S1k9i6VM7+HN2THdGuBNvuch3+41rYf
aJ/HNLICNuLZxSvnoLVnaYl2591QgBkw9FGm9FU2tL5ZAj78CKIYbxCDEetO52JvZjfGpukQHOaz
nXOFugyfInvMvSKtYKGEFggNQ6kIku3edCdpWNvTDugn1pm3Q0qiOk+SFaFgJYTmUHsK6k0Ej8UZ
UKiXdFTxvqeU6CEs8ZEpGKcmqhk4RdWqx2sY6eVFHa6IALNyKPNlfnrZwkZzQH1pzrlXAvAMBeLw
AWbDjZ/+w13EmGEY4dEID/G27/gZq0NFrlz4D+bzWy0NssKJcnm06gIT29SB3oMJ0qBKgMTHxY5Z
YOzOVHgrC1+1QnaDZUJQvuErhCg3izTKKOC3NZIrZAS5+YjTDU9kmqAemXpvRm/tcACTgZSTfuT5
2z5+5iqDWogaO5oYBmoj5xNledYyzGlV8Qs77kRNT+iKzCoSNBC5QWxcOi4QXEcnJxLi0WRoXpKb
7FdvqjXR85zrOyM00un6tzdOzXuc7S0SnuzEShpEM9DQolx61gUwQyZaUUCtixH+DBg02hiIaStn
mG/JOfph64nbADm4bPU8pPg9otDi2svHS1ZmNOC2Cf1zWqwSGidgSDqY9/rGLRUhWb2R1ww4fKEH
WUb0nEXcDOaB+PQiPewKX5M+LJGbQ24Vo4vpt2cCxhafRuRV45KlWQO7A+4mWKj0+NABBI7gTFom
W0Hxp05w9ft/ypOZTjJaXa4S6GNXppAyPiZy0rpecYCveV/Fxvhf9Q0SIAC82NR5M4BF3DF1VmXM
49xhvcfDw9DhyYlLJ4bJTNqqhhuA8c/Jn1FtqwYD/yqnwSbpQVizjTD06mP4vwnUH2pvrbvlZ4Fi
B0Gj5ZDcjfeQ9TGNm6AnJqyiCMe1sLFCrgW9TOL2JFHPlc4acqxXsEcUlUuxNTARSDEP+RUBcbuV
h8C7V7HMtdJOh42zwgjiiUtsa5HhzNkrJRiVJUJ8GvVnQypadEX35Mbt84XbhGYc0Qrg4LMoQaAy
Zec5IF+IzhZnW8vGint1HP7Qu7xeR1W/SgMGEzjssaAHrVhvplWgmcgk7r/sfMlnghtBYLGtdsmX
c9twJmGyuLidMcdaCPV/BmcQYPqvTYkrYexygFcWAosIboONleAPi+NWeDZhvpn+GGU60VLg+jk8
siZtY1FRyGG7tGcvV1JfDsheXMWkopv7jyHwsm/Zzw2PzjMC1MZeDx7xpukweZXtDfNxlH12xoN2
f3bYvTdIlhv78+X1Jid3EpgG78dN4RD/h+OobIFOHpOf8u4SAUR9/FneKlpVlaF28k2Wd3326L+r
fUOB4HeGbvQyWdxDeLsF+NmfbZ4QjEEAjUS6c86iIKWl2s/G9fZ2c9+5Ud1GU2BFpHpsqmNHH0M5
ZenMvXZg483xA1bC5mcCs7t4wfq9X5DfGEAloxJisEbi+O4FMrK6CQEnAoEfZS0by5QUKNKgNOHC
fDreYO5skOllrdVxR/4qMsUshIWWJlSSQQg5W0OLHJZB2wFAczSpXAom2EUqq/BFOMFmMo8lZxEV
zqVCZplc7GApMG9d3hRsHbmujR9j3S6MQGk1AVPIcKIj2OJL9BxGc6nPW8NI5ZsXUNMOEnwgW8N7
0Tq/gApM6IAEQAhB1/IUFQ2uZr3X7QMMAfuMyatd8jNMPp/pkeqrSygybr4N89o3iEaENYt2ROz+
9E7MmBFA2cSeploxEWxqsHE1lXGwKQEoEp8hK7XAF8NWxtfKSauUsUhfGBaHjkVpJEknVf95ILGm
HIrZYylcAb/FZBV5oAG0HMEaHV58ce3qczgDF5zKHgETDExiCRbD2fn2WFhcafqzj+W2YfcIxC5+
WwwbIdEXsZDXoYD5cpLPKGKDIH6EWIUuXHL04Zlf3WxGNH3ozqKyayyt8cLiV8Z0Yk8RUNiGHhXO
PmL05raoHcoURKs+2tTS+dJndXMAXY3VxGYlVV+RerXkKP38KWtH0XcxZXJs35kj3rZtEK15mtzy
w/R6l/He1FD5j9xs6jrqhMf8GVqDhplYDf0dv2gZ3ob0sxTFnXHmtbocS9Jbt5sTkN7OBwP6QqMH
hTMsZKDQeRA2tQN6AVzPZcOoQwoF7gJ8sDnapsf5OAp6xY6iDX2Na7vu69GUaxQjQpLycnslafr/
/Ib6+ajVWLXysTZ8Su64T8JbNVxcpwfqeVZwAaaUi4kJEIn6DX4A326lPD/DSSlQ35GJKVvC9//H
2YYxYhH7y6KdOgPrj8oDLO7NU8PQ1F5tEIH2RL+5aoFY5K9/CiYX3255nIJp8Pj+97fki/H8cPfF
K3cWjy52fjcxJjXQMEuujQ2i+y628LvDKRey00ElFTZe5Z6hiGx4ERH3aHA46yHAdzSJTw1qUeoI
/2HVWm8yReJdtr/TRHJ+VNxVMyGlF239dXBnxr4reb6w38XFx8JFJ7nGwAmYGCBQtKQq3z9F3Sb2
Z0/9bwpULQpa9NURjhkQsmWstuQUQiMWuxt5ADxvfK6kMJ2aCstaQkgyoVP9ctGPwj7sgRWTbX/Q
iloy+eQnO7c4F2m6A0D6dZzlO2hhG3rHOpJfwwpmXfZ7G3vvRB7e9xkaOE2EkpDh/dCkaFLKpsWQ
KTOoYb6sJTzlGEP+7EuukLBf9XSbJdLkuhUPJ8zWSZ4hAFV+ZikxB5FMAhKqpvPB8+/poMokYMxd
AUe0a54NR/nMlsebnzhh5lJXcbvQTPIxnaXkB/y2wEBWgTmBEso0uwNoudzD4mb8Xb4rr0XDAjEq
maADN4T4DIn9fIZ1w4AEvGn97Gi+JWaarRCqi9KPV+tfFYVt8LK2WqgC7QoMMIE6MOD6fFlrlfc9
Ff2nqz/U3Y/IlqVkx0M0iaRxNKP6Wo6dsIvJkpEbcGGYJrRhPO0dnbr5W+SgVXNBwg0jJ8c/4aua
3T9sEbBjcJGtBHJob+hGNihy8szvMji9RypJeSU73hlnKtM9HmKWJBvKMgTiNUgQa4qnZAvWRO+U
PJMfqhHT48L333rqqFAhf1Cc67KV+3Vli+V6+LZ4/k5uFwU8kScX7gr/1l3Pp1vFB+HFJlZBf6vc
uYCkO5SHolIA/VY/KjDEPhx6QzMcoyOgjJlA7r/dFSQSWaPFx9T4LhBoU8PYDR9H9FF/ZrR53uIC
n97/6ChBR66E+tdScm3q+AMbUlo5w9YfaWlNkz2+hZuS4OgLW1SPw1OGGYrgvcuDGIoK3kR29ekQ
ICwY4QBsPul+9beKLGZS9/XLCwc6VDbleAFPMqRCfQadF3kUlcg6hGbu4bUuBakaI9wsoGUWiPPq
f9FEW3XOP2WBFB8p/+0q9ValdeKnJSeE6LktfEgdoKyw9ppF6BO4csFKtd9MkC+NUMAhc9PVxIwZ
EDjW0vjrJszmRU6CY8TeZW6D9YAV1kXZSQ0/sP2PU7apap8ON3gW4RXE9dCcQu+gDcqAFjOCoybb
ac4srishJPjyvP2dglRawjQlcqYf36YDCjoV9NsWGuh8VIWisyXnawE1f2zHesKMtZpJwuPnEN8i
wQ8WwnXPOS8iUoelyDmcxBsnhexaSdUfIDmuzZDpzKefHNPxyET7uz3aWZrQA8gYvgkqdb7Be4AT
tghFctZICNuXQosfCKC73jxL7XvyBo2Y6LoOEkAS30DvS5QmzK+reiVXbaNSp9AZQTAj9F/5f3ss
vpfBBNfO9G+/1Z4I8MqUuyLI7jcJ2M1T+jnV822zPcY9LMDXbKCevidMeF/OLXW9dg/RTjujim44
906/lwEPIMmKrz8ICI6N13aA59IrSkOfM2oph64i4BMhq98crB7/CfYzTU+d+rgzMVMSRlT/EA1P
sdhkyvMJ6cZsyeSCBfuxkLQbEz0k5peiW335Orky6eozT4g5mRLXmD07jBdKnwImRzb66W/fjjV9
6DCFiEysSPJLHkrucLL5lYnydz7fYTchLQya4boLKjf3S8ae6KP25UVqYv0Ff/vuSMqWWqnmrST+
61PsnKYQ78K5VjJH7eiJqn9KocJ18hvGJrqxpO6H/v1R8Zz4Q1sAKkERxqPww8A8jZ3AGjTlZ4tw
ex4l2Kfslmp8DQ+vUE/cHe5raFQXB+bLMMR3T32dM4Su4HKtPV6O2kWbZ+O/wTAe8N239r9oto1g
FeILBQHoWH3lZDmA3Kry8CtDdUhfRROh5ypDSxUjjch0GdcZvhcS6qImG3sCELGJFhz6kQFrW0b2
7cyBYEmqgdSlE3YjqZYQBww2MeM3UXBliAJ9MpSmtz1LALSo8lz/3W74kqrawrcbWJL+xpRqS/4N
NHH37nvv9Bknw+fREGbhKevQYK4tvKxzM4L/5kXx2Mm5IKcgYAn6o7+2QNR/XFkhmDAhYixMPNdm
h3ERJaKfDOQ+itb36JEzscuGfroU9zwBV78xPwwfiYHteKAe8HL1/KfuirCxvWgP2MRMnNLnRF2V
/sMsAefz+b7+cAZ2BKy2PgOQnYIoW8AxUkqEQEMXYlRyLqSGUWa0xzPE1tGw+o+TlWQb/klIwsdg
UA5942yNAzciT3iq+7jBYDSGMo/7/O6UnzXVl09JtYodxjAdUMv071np1M0Kc28pyATPlZwSKbCk
JA/P1/6siEQMtl4wg+m8Bvq/y828PItK8eSbpStZDRppWE3OpWilRzdvxwo8NwK/F7EncbzIgaYm
YHAKtIkhf9qZn2+rMWHZbmFAhoRvVBWnq4EQHKNubEwwc1d0QdwoN8DF8yrZRmyyfJeTLsG5007g
5TPOP2Hy3a4nksKjnejqGTRru2Dz70oRaBvnlwhxAEn1EPtMu2tAAKPY8et2+ZNYb8iVc+E2XhdT
mn/VjnqGLn6xm+322FJ+38P87dXLq1wZmImN6xNbxlLUX4zGwLE0EO4G5uICTQ9Dz4lOtGU44hEY
zUEQgo7JXSUPmQdZVhllD6jihzSaPuZDNR2dtOCrQC79asxYCym6fvHzrTUDtzUvUM16yhdhgzSQ
Dl0nGEuGVl0KPuR1nuNuxsj5Vo9EHxoo6eaw1SefA0dGt6fcEZiL249o2OS88a+ogTc0jv8evudy
rJcDzIvBQLk01BaKNXXNwtIqZgXefzE0vWU4on45QfIGwLUivDi2s4oDRphkIvuboOSVk/1teSyY
Tju14A/OyG1Vw4YpVT0p5DyJFa1LESUIS+9wISlSfEFvLzZIw7PRFCkiE9ZFY0ElUCYbPYccJAGS
JrTEQGpFRRqJB1bSpJsJ7Kg2wcmyO1cfdITgQwyd63GARd4sZRObRq5kzb3h1bpaKAl0cDohG2n/
JvR5bCuVV4iBlNCweniCvv7bXDvEAIBsNAa9Q8ky1oPZQHnhp4DCELGDoO08m/qOJrtNaVBZ1vLd
E4uybxIFHreTzkxK54rzkZo5HO3oBwQ7qYuCe9MubvMlc7+7d52xp4gY+66uar5qjUS4u2wamV+A
bjWvZTHfaOxngBC9PpvjOs9SMPOTqG7rl8gBnWRH/aLYkaAya1uwmr9M8ShiX81X780i7DmIUH8N
FWlekDhMyNE2DQio6jrZ9Q3XuATmqCimqGdIhGXPK753Ciysx1CRt98nMIcekKoUh94MvGIdRdba
ipqealqRlGDZJtxUJ1LOlu0lP0iLrQlyRdLLTnxAbIT5E0+H280dlWlKXUXX0mb9uCty+uu9eBAF
gIj3783qnsAm64Zc9G4RQQC/ndsg7pEE+X7sjBo/UrG5pSqMb5gwsf9jSOM8JIWno1KpG8fsXeoT
KIRiIxFkrpFGI1EdjK3AZggzZUFA0cY3rTrGxYcMsZCCPL5HL6Slv1NENCfELT7gNiDhm2lNiuRp
Uq03egkSVgq06LYnMr/pL0FkhTuREIoeyu923sBAc87AObp7PDcy8HUPBRq7h9usoBm3fZrp6Xg+
yzM4/nn1aNCyQ6DKwHX6Ont9GhHwHWc9OWTYwyjbJqB2XGG6xSo92N3VgLCEUkVfTXK2pYBaQqFj
ZU/vdbv6wRBmvX+IiWOoJUxH+R0eBFCXHUBTSVZxM7Up5Awz7Op+fYIZJDJK2KW+XYh9myDjCoG1
d4aQ4F+0WhUGFHqTLCYL9zRgSxe3UBap9JyR6868AdJg8cPeryfpcP04IsQdJ2EP+Hg42ouNQmkG
NVt1cWwR2iHpOYGArLBR6LfVDaIfbht+2T/VulcOB/jHUgkXLW/yeOWdqYaUB511y8st5A3eKPEP
Jh3pMV0hi55weAqaHUuumW0iuGuGC7yNOtb669OMtRD7pnuVh40hqCOZ68eFlXrlyF4VgPZSOZmK
R50Ngp5Edzhl6EQrJSpppEtlwQ1K4WxnqqJXZt4G2tAr2/oFoemGWkfWPN0kKFbPBwgSnT4eVJR7
plAV/iMa5y6omvvkAeTVttvUhRtYdbgtYvBqz8IY0Fm1Q0pIRYh/DiqmUBk4cX6W1nDifaxKkOME
UjqFgWLgO2LwitkvJC0biwyLcWOlhNP1QWef5mJCBJBQym/f3dIHVYbB344AVBoWFnAfbHq9kf9y
d3upL816am8clBn9zVtFgIF+lqbD5EPptyCaw/CU9+ttj7DRVZRShv0qgy5k2YUi7rHgXWwEQ/IU
zOWUIdMhmkMlxCA/D5/Uh2uazrkFax5PBUgwhtII6fihCL3ymlqZQM/xsdZqJYrncQ7ANYij0Pao
n+rkDnKGSwZq2bTaxfgpbRpdgV114a1/751xir14aHeX0IMo0nplnM4pMPhN870IY+sT1QqoSQYz
CAgQb8X5pAFkkaBd3/eyLXcFVswc/1PXrSF33M3ge4mx4XDWn+pEAVknbfLtWQ/kmNxtv3Zekxdf
reAyeN3cH2DJQtoyrmbHAhTYKOGL+XlCLtQpNNN/GFBuwUVw2hMVs7WRMoRn1Kjs7Rej/1sWZ2WG
kuB3tkhj01BXIG0+1C0nbnXhXnIEUPWk3JdqR224lo8fc5h5lVL6gyvZWgVlqHMR2c+78aIgMiQd
tJyo+x3UvFr4rKrPhXmR7kNCbDJjQDVaKeps0++/4DDg4PF3hEgTYkQ8i7gFajOgRkykAJ8jIJJt
XkzOyEbQUzXwTyP1xe9irL8j9H9XcVOQ/ei0gV/a0BjyOs4TwD2IvdONMBRl3SxQEitZGq+qAIvt
slF+NnGytF5oEq7se/48RnBnJFXbzqa4uOpYU4x3OHL+xObUE00oMUogH3rY0k9xavI9mdMzek+Z
THwvLu/20TOINiQcyfHuR7G0IgJIxdOQFrqjnR7LrYbnilHKWHGmXcianI7UNlT0Z3p4ZqBKzDXg
MpKvrpxjRKTQ5+kuhixvYWGkeqt2gPyQQNAOIah8CzFimYRDpOEaEavhX/Ef4mzm+zb3ytx8PrXp
MBQYMFcv4aL8UCEg7SoN1dPfroe2zCvbFFmZcvCVw+kzYKPDUIob9BV70+XG6YDeWZDxMCReD9EZ
yqu6p1m8U8qASgoOc6SCzxVN64szK3FeiSLLajHCGi7G9G06GaIozgwKXu8GTYQUToeoY6Mqpet4
NOVnv251rW+UaSZkAdoFJvReMHN7MYHKw5lL6xpPKH4jwU5NzbZo6W6FyvB+rnSPl0i8Xl6ebiYC
S/I94PfiGz4W47Ev6rZLaZCDrpiCtg4c7TKSL7apW1Ia+vH4W5ezpIriTxi944Z8TQpZFEE9rHqq
MahatBcbuqrYXgSsfjuN5MAjVEmzTPervQlsvE2JWmyN/kg8m4MsELtYj44F/n86f0j/TTJI7oSw
gcMJaWCqu4wLtjbwkPvhmXCIAMoM6u6WZW+Ffh2OGeJBMO2A9LnqZYw8gGbQU/3cL43VPUsyaYTE
fZ6rsIEedL5WUyzZM5BH2rTvO7en+JwDb+/BLmQ/xKjoxFkG2TdSDwBxgYx8pLyohwKjKnNfnZn0
RIUCKLQGvq/F+ulEsOgWV3sDbTEvMrGaPHGaOAzjLP09IvuI8OYQlj7zM2Q/uobzYyd+dpys+jGd
zqozIQVx9miwurhP3/mwc54ZqpistNEg0wTvGoR4acnPuRBe3ps134Ype/GzImhdoHEQJcOybUPb
UJamH2pCJ+Thz0s4U26ta6KbZLkvRyVTR26uLpy6ppKoQoYvxQCrzDu+vJWpQjl+hfo7jiKo2oVY
PCDxrr5M6qnRvRwH6QydLrsF20gAKQVBoN8m+VKRPZ/Q4qb9pRvT+HYuq/n5U9HUric9ccbGUYEd
WwikVlYeesMY+1a65qkhVuypc1NBf3FQmij1q0yytqjGYJ2BMheDYgZJcG5aqQ3kFla35Y1T2QzJ
dHxhxjwHTp8Kgrh5GORIAjupSxFzpRJ5+7bojw8x+03rIIhGGlnmNQ4CuAoEDQRb+bLDdrHstG/z
al4i5viDgIamez3SPSFyJDSBdiHzfiNXwEJDoMC1WUEZilY6gGf74K//ZRWs9DM9fv2Yua2e/NQU
6oIwktp0onD4mDrBbu9GYxnoyhUwvgJj7Hx0WWNe5hxCZ49AS2xX1+nDchOuAikmzAgp3A7Qdmgz
xbJudWpCDXOV8z6W+0TIhncls9xbyseA/iMffWcHf1WeqTiUWTqgWHCEVhG/2F8RAD8r9Jir+RYc
onGlrCIyTCF7ududiY4r7jnUm9iF1oah2GF5XJBQF3vs6yAn5LLpK0qXM+zpKdT0bH7UMmTkMfDN
RzOuxRbRd7tdJv3Rj6VOou1ocJbugw/zloOn2s+9gC+YQ9iOaG4FwsbjXPCuBAphpYbkLpuCHKVL
+ddEmDEfHscRWV2Y6K3FJzmuusqW7B9+dIev1MkPBwawkAhQYWhUEbXZrIePGEvzjDa8o56oOq8K
wOfYvEF3fzy8aznZPGUuVdY0tUzrfWdSoeWl/qegV26aqG7xmj2qt9nx+dMokNSqkbHPYwHQbI7o
fUuS/mTNdta/Tw7DmE3VFN7yzBFB9Gc4aG/gUju4IeiJo4JLu2Qf1a4hFtR4vE4BAl957SXlguYV
kgIWfw+WnBDhbMz8ygM34HTS8/je0RQMAhuw2FNt7Wlq0LcrbRUOJhjLvTF+GqVwyvJTQksNN/S7
5hcMtRjUImcW9dHJnTFWOgNcPKArFaNKFBureCuIRxOHeI3V9uL1WBhWo1xyr/SCoaOZdVcNBqHr
WCIHONh1H59uxP8BAWzpSITyVARmVr5ikMESrB+M4oXH40b74lhpb6yVBa+dAZJ7vLtI/q+xocs5
5zC7Tr6wqVaSonoKZBOTq/HEDKC8VmjwLUVfH5r3Mn2penuAU44ZlWl0h4Wgz7NFE8Ibmms9laof
8Hw4P2h7aolrpMBim954t7tZVDoTH46aYyQ0KD/rD8e56a42rDF3retf4QbkWjtbwwI1bR61Hqux
+bDKBcaBMJPWi8/H3qPJCHI3WPsT3fePoYQKI/vwXa6FAOZyhV8UCaFcJoAzfwu637WfDCu61q1U
8LvtRgqQmaP4Jx2U12SC8o/m63gOI+8zErZC9QGXFoDC1NB7sPfwEF2zd+MRK2zb2OYvIr+GrTjd
Sx9jV6OILFvYdAnExpsRBMQIGLCiM+0mQMfzQNPCIRC7uAEYy/SDY6W+RfSi5Bpie2BSUF0O5lmv
XGAigYIjWWOg1pOv2gMT9oNhjJblmClC7XuycWyocg1acd7GU/6xTAAOPestYBEY7s4E82XyLGkG
14Stm2RH7lU2f6IwZjtmqbCR5BcAOrFQBSJGo0f4dv+L/KbhgkE38z9Nz7POip5NEYjFZhnuNVpb
DxtbBPuyxdwxOI+NScwi7beTjkMZNw/r1so5H0VKtED3cRUFp4JzSyNWNp/CfkuYh12v9Qkru+9U
qCXPnsWU9StmSRnzKyz2aVm1Kvf2kw/nY7GoXA5fKbg8DqxGhW0sBDnD5t9qvtxaJ+XIuKtpb/C6
Op6BFjkjKOKghZYwgEl1n9/Dv7hMU5NaVwK6qadlgDqkmYiOAn8XDXEqWH1wyFTcWZywdHcF0w9Y
kcUWjX8CrWBEXd7GsNaf5CgOyoIEX1UEDUf2JNhrNIJmdJjGWbSpQv1ZEKYl0J89zKmaHzVJCE9j
89jUkBtsnOpEwMJw8XZthyCl7MXpXcVKIWGrmSNXuhWdUuuh6qeTu7AlO3wryoaZfoEJMaJX8ySR
N9UEmJmiYP85XwzeGU3TSOnvb2MLiV/Fy5nL1gvJj5stCXcnM+7Stzho/G0ngmdfZLQewTd94xyv
7SaEeM7JFbTXzjEuwcNe9jsfRwQYMy0hR+KEXprzvA/422H2H1Pe78Mglr6yn71JE2P9qsyXlJ7T
IKhDsHXJqDfjc6iN0hRq+WY0yx8i9DFw1YubARahC8hIu3JokQuXtt2UG5gkY/ig+VsHAiqPKNlB
+SzzdE5tMYB5/XaxHdrrF5PYhVYNfxOVPBYsKIEckeosVbVSN1Lhxb5gvKbi9PtjR0tR6cZR+z0M
+ycKhIzxqqoq99mIRJKYPrqlI1uvRN2pQ5+n4P9TmmQyjJpS1jCLFYuzp4nOAesd4J3c2dVAw8LG
2F8mEGwCYLnjaD62Zh/wos4N7gWkDVfHK1AEWiNeFkpkPNi3OhOFkSCn+FfgqnOHLOSmhb/BbTS/
s/hbI2NIj3TrQESkL2v/tf7pS8fuHyz5Gc1UzIIzKYihnyz2h23fJtVQYlCt6nnGAkMVZL1TsvPB
nuRg4QcygJIVPYG5C7GmbkR0v0pavwGyIybpLDpQu9cCCyMeq7d8Sjcp8inTmIMYDgZeOu0tPJqq
XoFlybXXZQ7fZr2IzCnA/wdn74LlRAr+YnRv+kHb9O63NMqwArx6XQpP0KCsHCn5LfNdLW0VQNKc
jS7hC3KygLR8JTrEj/EHT3sTm07AMfoeBTcvZkOJRI5j1xUBaEUOrz8aZ7bBUUL/le6I4733A0fe
hmi92Y4fqjR2V2h+Tl+U7wYM0MjhY+p/LP7yeObSXBfKeyNQIrTfKYr952wo23SykfQMtE9LDQCN
adM72yfbiCbrDYO+LM4RJBmwmw2PzSXA/zjaGH7p+eLVzeDDsktPe0h1HSh2JSqMqSogO2V5ye1Q
bGS9Zg47iZrr7Ma0i284lPhTG2L+DzxtIZQ5IPFQ+b52m60lFvdf9UKnxgpL+A0DjKCZJhxHhwQ8
Vx8wruxmjvaw4KEaVb3qMYHdLPNB6co1YrdQS1rKzC/jGDXMyLu31Xh9jFAzJKJF8PWnrQ7lhNyk
TvfTU6i7NNNb64HhGYlAtOBIPvgzF0cS0G4qvvi5mNP2szoIw1Nyr899D/mn0JaKQ94E5ZkPq1Ip
+pj2aM1ksgJue7Ieggj7eWCnUCkGXKuf/URrffPMVTcOM6sm2WPogM0J4ewB5aiXO6vxA3IWTyat
4HBvnY0sjabKXiFeIyLLvuC4b91ovwhnpcXSpSnr8m9ZKvuXb0EYsDwREAjk/6NzG1SYG4NcaH6v
G3+JqUK8aTlPf/KgsdppU0jr6f56W+PkRNDUU8TidrtNWiib71AwO621BQCkhuW/uOynBTkvPHMR
0qRIkEiV2j/GafA/iLSnIyo/GVA55uKJu6mkyV/n6MPGMGcqtt2vOHonwyELfcjUaCygfseP4eiu
syHUf8BO6NkmnqcG2zhETEAcgSNV7UX5knWv20489ucBIxs2HcrElAajW6doaT1+CXrGhTyV6nt3
qgzxqeuL6oPpR3d9bNRg7/d3NWs3DOu6jvpvhWf+vq1z9+9kyF7xom30ptBT0mjJKwYqjEoF2Edv
7gbuYdz6GAXXJV0XoiPKr0xk69sVICgU4i/F0g48zIvub3pPgn5uacX82je068RGahUX5ae5YR0T
Zpsi0sxaDGm9ZCymStm9rosfEGWb14qK6PF0lf5ssgxZeEQlzVQs8D9qIc3jIUcQ8HYRqBmJAJ5R
ZpWl+ojHmbaoiHRJIU+X32+C+gO2TVwZE7LuKmyd3FLn3wt29DMBzl9IVCGFGdvHE9nSV12UmYfN
+R+v0Zyn1EXNw0ubmUXj05coi7eH9iHzayipGqXEXPlSKzkBDwaFDrYRHyyDfOy1swGTH7YsOM6P
/YeCJ747XDcXcthTkjaZQuVFg5p4bl6+e9QOQRrYBLmxpDswXdXMY74VYYjjQTmfg9/OsjZ/0Jaj
xbtZTqCbl9biRbLYG0W1//kpQIvYGSLTBEfLnGRgBiiWHNKEwoWSfQfIS21FO0fBuIEK8eaOMjlB
YFTg2YcFF13vwtJCSJyRdYD2E208qvzqWhSI6lUWee0SxFmW2M/VPCb8jXVVeWUVHVFE/LTZysmT
V+uH2/MYZoiEKH0rFMkv7tZxa4ETlzVBmc0RNZe0/2oJ1NNkETLBbFm77Shzib0NHWq9F9c8Izd5
CEvbLl7uppiT9VObhHqQDSv9VIjWa0ouT9pRjZ0DlojpISj18CBfTcmJYxZ3FtCwJiU2yH3CaZJQ
JxLKlM4Ri37amOkRIYRut6WiuAqJgl6TxuD8KuErt55IPu7S3h+yXIoeaFfMJMeIDuE4bzLwRl3Z
Lpse2cIGmDbtGuG2QUPg/iqfdftrKhhgEys318REqcYsKwMOcxYjs0LE9pcPWGu8d1eWUV9Wquwg
sB1k7qyK6LgHXgmlZ8Gt77NavKsiPAuhyyEUwDuz6qbZQKZpvxrP4PA04+aqzRP/B13wCr7OkUA1
WrwuSRbUpYQknXfE8x5rWhxpZtbaSkbYVML2ArFyKMetaIEpIW34aPRLDtLaI8RUhePHL2Curfcm
RFioSI2Y+9toCxhC0/Tefuh0iArjZYlXHWWRuAJ0+/Jqe+Ukqm9ghaMZpvXe0aBkcADKbBXk0L9U
CRhGfdVUqwDVp8cxp4iEFMIt7w3Hmxpxz8cRCfe3bBi0U44lNpemu/RKZd8SlzUpXsGAO1qnS4Ko
sFxvf/DvhuHX5pN61w2KR5Kg2EJ6JmGE9BqchcmWw2SK0K9LSu/vzKRG8UYJE5CSJwEqsvoAA0GM
6SmIVnn941jfTqa9SvOsIMwVJDdFNS4hm+FK5DXQhqBwHTt0QupB5a0j2zcIB3+zoCkNNTKjWJrL
Yhn6Gvuz1TobDlKuetB1xQbkBQe4ZXNHTnltx+cSs18Vly5K4NNunnRBNB51qZbxOOF9gsUixtBJ
padPwsWJ9Q00fMBdzr3jFVMFTZKZwrD8rrMQjRNc9gjK/l7V0fiP8xIIKWiZ9tE9SLxOmXL8qZjk
CWhz2gyTgdYQvqfmx0kWdPCtm3kdCDA+ZcTeXKANWZryj+Ti/P4dNkztUk1a+A5FNiMk0nYdT/jQ
9R7vDFTRDRmfa7Idcs2+r8LzSnOX0d+aEYHLgE179NJDMVQlvKvuvvrm0RjNe9WexW14OX4OPm6W
vXbinHd2zbe8HUF21LtAG6gahgC0+EeQiwGyWfv1R0bV3wl2TAguLZWJWmyudll1kDdzUNKK049z
ECmqW+omm/0cNWOrH4OP0zv3EBEn7fBuZXpqoEVrsQspv962hftUEr/NlCoYnFVnX4U0aedbGy3g
Q1dUa2BN7G1f2AqJh/TH9Fst6frf+Hz5gnst5cf44taFmmIUa/wfHWPgoP/7qzx1oVPJZHNTYWgD
ribjQn7f14FZUlx495TImLlS+m7e6S2xD1BOfd91wxOil02JCtx7wgLWGJg8ucqfDXrn9RpPVau7
ETmn24TFZLyCwjQubmti/d6xWwPhFEr7WydL4O/pYCYL4RTQ7zYEomePMlEk+kSEH2RrOmW9/da+
9DS5Ak2PyT0Sn+e5cYI0VXwhpZs+E9F5oP5E99TLF2tq0WBIjWN/mQ46UN3iPBxaQ9mpW+msp8HT
O5tRmeQgHDpZp5eZhsy9lBsyzLrYxUu3TIIxxGnKMp9Jrcl2ObyAaEIXh+Ot4CGwYTI9vtjFscOi
spWp9s6x64LAab9jKtrisQJsnQeC3XM8/bjhbaig7pxiYgNvWtSf6prKKUtC6QRz2MtOxwo7sRLK
Wo6eAYdKHpLHozAqrdTSK2qy5D0w0DwrD4Z22EuX+kM6KQdhq7yv5PQrVVQPAUw7ef+F0Lo2QkZd
K869939+VghdJLZwyltZhTE1VLQKk/KeY9GhT9IdA5m5IjFHXkUDgjV1XKzCZ45LuwU+JzxPH9AA
Lm6az6WkjYX4RG9gLWaN6gUld3/odzGfkkj3hbZ7a7w94idQC+QlCbMwoG/JshiilTGbN2RZyv7W
6XWXWbC583dWeukBIWA+umRYQGPjwoa0JbIYuo0BBSccgAFJ8VZmjfankruQVsvQoGA76JyDA9+b
h2I+/G/Ix8PdplebRztMaq4Jc+YNzUbmN00ylW8lQEBKhn4uHrM+2feOmchP7cQwjNIm6m7e0mHi
ysVuxp0DmBWEVbg3BgTdeKcTBX/iQe0KmPtHh1K0FdOD84qDw4nJqT7gCmbRqdx+S6zH+BNZWMk1
ZGzyfv8Ch9VO02p4GUOaoBSPMY/HO0tmbrE9LTsqWS1zUOutrlWTdUJlkyH+atDpEH7TcQgpDfz9
Ssye8Qg3Y1MSE1SIGddrxTwatBK4SlwNmhCH2FIFEs/f7O5ZTYr8RA/nbW/zq2F0Z3oaVY3neaDn
ZJiwmtUpaHblmQzt/1qgxLMoA5yuZw8dZ4kIjMFMGXi8r6mRysopCAIvEcqh+p9E5JbJmKX1NyFg
T3r7dMcd03eHJ7NSu5R+o8fMmuC+9DsbYwSIwvXvdm2PlImleXM4BvMPyO3iuJOoZ9uLU1qI7qqd
uSrVcGbJX8CqNw0vbu03MIYUIj1zrFJ5hnrw9zOgxklO8AdXow9ExaGkOSmkxDXaYrkxj2Q+g17b
Wj1d4Dmj93raVdTJdDx7wGSL/OlYFLhPWFH8oXeh1NAI7qjLnjTMeWqKMvofInV6LF3jz9z6OSCl
478JKVy/YnE6xGBoMaTFytPNPxXIbc95hef5U5KfHxmGELBZ+8DFsS6v+WgJmgDKtFaSanVApwXF
PJbyZ4I9oL0YJlTgJ2dLw9Fnoiuh8ZHIDhKmW5Md/HKtCuRd1R78pXIWPNz9U7rsSr8jHU1GVJon
E196+sQmYz8Nnrv8UAAkSb6NHB+1SJmacyBVQXNIKli/EY32V/JEN+/dubvH+7ivCsypvCceggKI
thfInWRazgvz9CmyIo1YaDuoNylTck8gPegKB1G4bN2VC4KPpatxKpZiVgNXMMtE4UT4O5qe9E8R
+b28Zq4emh4cHVdu1EFZF4MTuln9c/Evl8l4pGUPS/ecmm0byvDkiKthvSovexw4xQMmj2vI6jay
TFQ+HqA95lWQn+VqfcAfd1aKFTbhp7Tg1z0zM9R5fWVZpyUAM768lUL0xfH1tOdz5kpUqiQLbErZ
XY1fruEWaD4X4S9lRIYPOZjxFdMI37gcjPPP3j2lqIPStiQ3ZzouDJYbqX1+6oDOKu7MA6y/U9L1
MDv4Jibdq3i/myjx14NeEU/apK5HFMvB00TS4vOZ/kpGh3eWUNo+8GhpYHeiftVZts1W4w+u1md5
hhU478pWVPYjPtXJkqUoMqzLqCKB63sQjLVSQ+HwI2GBk2twGKkk9jm4kKpbe2Z3j/xPVGBPmz3c
OoEhiq7HgD6hfJJc+Q1tvoQbMgkAmnjzSwz7jnmaMsNQDZrY5/NakP5p3HRUkmhfGplSrcieH/Lu
e86mZWZydLaFxmFx2zRYGPneq5LtAtAmnrWDgArDOYrtETRvZvkH5fil1/Q1yjnMLoMNBOWPGwJG
R62FodarNnidPmrNDoFxL5yD4J04XCo9RE4FrKreZ9xGKxZP5k6Htqi14hMJqAOKD+U1kIeC4803
s2qatNL1w+Zwlb7IGO2S1HjVO45udioMzFQ6fQVB8pwKQsKEt9HHhV5VJeV7XvkDqHHgTuIjVR5i
XEOnOmoZc6SYuKzpVdjhLGZOzecK4CBce/sL5TnmiqVz/l/Lq4lfd3rI++UjoImPEkCtyeSfMvFg
28T1s+FqNsSGVEOUemlE+8Ix3j27489dzLWpx2humRSrd6h39brzC2MAR2T0BSoo3PcU9XOrrTbc
TUvX3YDHst4z+D9OnWip2GDM5XNvPLEqxmIXdwfYG4EYFpDit0QUBuzJ4EmKCPFdNK4o+m12ErJf
zEVWImFWAe390V3ErAAtsVagk7TynMuNBlgzcLha4o4875/BxF+cbmsre4/CbNaKGmmzVEkFKYfx
uEPUEaR8+HOnn/wmNiCgPDYYlmu+aUbFqDzv7AMo500OQlyahOC/7R0FXB7bdKMBppiZSu1jtoSQ
wR1WilDcU8i7zccvamt6kCvMc0lAXmzutT9Gaf9BIQhxV1hb/eLmRcle4VmTGbhckLeB17a/rYdm
sTSAJVbSqQAh5LPwLEbmtXd2OrrBc5AAcU8/5hlT9NzmLFFJjDvN+1etxCaPP3PBh5R5hDviOlfx
4owphvz0qzEsvKKZMEj0epYlBzdeP4ZckYP8EknjPUQ4OFwiYaOPIgZaF07R57kW/wWeaKOOmrxA
9bqWOcZcJ9zpxi8dtFu7+xW+a/z7WehSfAnQi/AFkJwKvPwTCNltoQE95nZcoaKgT55m8mJRTNq+
Xb7uqMlt8n4kZOMfQ7jrZOxSR+OkqW+YCG7C0/Fc2IyYPZU6QYEY4h7rxEY+q4CF4+5hPafOcsDB
rLaDm8mkO3hWKSaC/cvY41qL1CzjIENWEhz0PlNgg7U74E9P5fOAhCzMG1V0pc3dji49671ku9FF
2/r4W+iE4acxMmAgaxbiiRbOKst1xFkOxxr+msqETDkKgMZm/+yWfF4nTo+XrYJ2GUIGebl/RTJM
zesEpbR+xRpo7dhqMTOB6zF9usjWuF44A+bvmUCTd2MlpFIwep7dAsWSTRLQrS82aiF+O2IlYCZc
zqR5gxsXNFGwj57kJmogJn3LyQRjdQ78GJg8BQWo0vHuWvOl7uagc/7wh/0GLnLvORNTyu9moRit
c/K55nQlr0HamZ8zJotkVp+tyHY+xIOaMdfxk6hpXLm050px13eX7NkaO8hfCgzXv2s3wumM5tmg
Q4ZJ5HWZUTK6BWIWIQ5zCU5GetDK75DFk7mgfnCJNC5kJQDd6uYxrPPN1fpOTvZpxgsLfWn93Sb8
+fUezEnVBDVoQfaL3/17mK9F76gEcAcIr3mS6SgKssxluecgVX1uxWxmQ4SVvIt2zIQCirx3TkIQ
scBosIPm0lLWiLUx1v7aJtdIi24yaJbeESlqLPz5UinccTVWnQyCvj+bVVW5ONgGermnRdnKCeE+
qAZoG0a73F+Y+pBUACVTQBcvtQiNhjzwp5SApEkbozITaOOMcmZn082qyMPIyi9mwL8J6nC5o1EI
2UQwafAzTfToNr5ngYSNry57IxxqS+QmRzcDAKJoDxEK3IL7VYOoDCE7QrEpqmOMN+B79Un382VF
rmDrJ1itZH6rz3LD52FuDKjFU9Hnq7r8pV7/GYwzO2ehfe8HiW2cYee2TGG1UymG7uQTHAoiGXMl
8r0qkPGK0r85rWswobItw0gscTBNZh4YF3IDGyICW253+sDrJzdkKOk1jyeJhBGRRg/KTWkzGTAo
m7aPM9EOFOhkERjxh6+/pN1xVhjg3hg80Rhk19K4/eKSJ8LlnpP8yhqvE2FsnQM4LfIPl7ENCQEM
mLzaHVOYF3MXCUoGj8seZXgb/Gt/48bNsDWCvVpnfqt55NgWoyd0Mcj9x0egxU4bIV8APjL3DmgC
jEpohnl6D3kvVzkmY3sn+lL5NPQgyPAfI/Jzt7xjjZ7beu3TpAq7WW1WONJoplL4gDMnsTVsujFH
L4gCUVdNhOvND6cjg+0tSVMYZIe59k0VDZod8FwtIS3L/+Qq//fWUh5uAOc9vknxv2aoStAIBwhm
xUaxkq3aJxbui7ntpr+m8O730zN10YeH/Ajkf2qsAEKNJjUYmrFwVxmUyixTTJ70d193+i+f3zTS
GeOjy+MdSoOI64yXwcdFq5s+BehcZDnx3s68ljJ2NMSdRpvG0ePzTPVJo8m8v96r1KFzXW73+EZ2
GquSwcbnmVni1HkpGx9PIHkQSBiIyw3vBYV44N35hTv/wLslbzc97vUkFuceIvEIHUXvkRZWoRd4
xm30Z29onxcfXX0tjAQP9+P4Gw1V0juvIf+d+ftCRg+dtf/Li4UpIVaryURRaTmjFNwRcfV28V3/
iKatYA/vMvNCZthbCVwrinhO3fW2eihaSv5XU8hCEBb+ReBBykW1E1iass/e3Nh383AxWJo5cQNQ
GMVfbxTUwtLsgbCGDK+OE2h3GYlzcr53/HVACEyh4YId09aoBzOcOc2L57PhrP1tZu6Kyi1g04Wi
v5ydSj/0cfJE8L2YSOuvNK3ipFiIX0YIDy6fObPcsN7TqkOWPT7tGVFBHBVjnDKQxt1aplraj66O
3cqzcqxVU1oUrw3dN2n4Gjuj+E/TUIk0oMuC81Kbqe4kA8T7f9pX2BwIsnUUyRi9phgMoYEQjmfS
AZstLNDg4IKbtxe6UASuY/qE1mV4dKdCdT+QPD5ZuRvln1CP91xuUPSfffOFZEOiW4lvdM8QPYjY
gC2NwOEWieL0vcrBRbx3IoRxVP7xj/nvonEuza2yCu5ZokvPUZdliFuyNFYa98bW+V2z6l0pn95D
2LJdMNBPIy61KqMAT5dIt7cFARxxMwz5iUGWXRuK0SPV7fQd09qLnxbJMpcTwbnDdJOQ3TlQy8M0
8iDkm/e46Oj5zBTpq090YpPoO2afyNs2i11bOScq/xUjJfAi3YYOe9CQZ22GOjcAW/neYTQAD/11
gQ9DWk9g99q4UKv7M3NseaTJfQVVbwkJ7mlqg79FYoLyt+f0lFphWa36DcKufB8e9u6EBC1A1iwD
RLUh+qGETMd8egXdVCXefniA7TclRiOQ+IKh0TwdllpkHQTxYf/MkaXnmxHPVARbGUqcHlAxWzLb
bMrmxoZ3hOqNwrvcJXlkvtVcFUY6cCu9imRa51lhfefbv1Bsy9bcsiIw635AkpgzQ+SPMNx7q3cM
i+pqPxKUm6wQ2qffm73ha34k4MFwG2sEoMOw3ZZtDMR2tjnC+6JE2awB9ZpNhpan9ZQBgMm4dAfr
LLfdFj/r4cE86djPxCnAzJ+r8qoY20+H6WMOozRSkUSpuguep/hp2Mbtw+bf5VIxXCXlPnMrEGDo
/+ngSCrFf1t+KP2oxHKn9yGW96+T8wED6MDfhgtatgYv+95oSkuF4kRvuageuioRZnbrn7gVfMFQ
zcGJbioVj3jMYsn0v7mQF1wteyIkaXKmtWTbLy9oIrUAAUqxqpNSh0wiC6O8gBZzWpOH28ZHSKm3
LJ8TPfDUbdAfJgiuLW+cn5YVvsdLMc2wUJwJcdKYg9+3cGa+Eiih75BXfhJGvUCsjzh8fpFfe1aL
b95BmUHDW43DBwO7eGhsh+yTWuZd5IDMkV2CAwdO//a/bSusCBsraz3RAU4Z2W/NTDGhpjLVpL8x
yAWGmiRL/L0Bwn9nUtEGqBlCXhlCBYhKQoec9Wr+QnJ1WCJXtnc73rJwEVufHDZ2PjwZ1cpRkrzV
q6aXM6S9Nr+HbOkWObGH+OcDDzqhM5qr5WUJqEk6zltKQJkMRduuTHfhm84ca9j+s93Imcmm06L1
z8P7r4X07G89Hp/rPkg3orpzHJ2lqs1yJ+e++QKqcNGx+1gIBtOjv/itlWuRKdWNts7Jhu9o9a1H
RQmTNM2AkaIE+6rtFFLdUiMai0dlCNqLK1oMFVbruateoMpVbcIRiSC/1hDUt6/kJKEpK3ze/FOT
0w6Wz+x8ukCMZ58m6SxpmvM8YjDgNpR3fRi0IQO/HaRd6KNAUWX//UoEbIBhmmzXa6Yzl6wylqq8
2nBZzI38VTEaJjs6a7basW1R15RglcMAgA7D4Uq9H4uJl3O2nb0z6pIGii4GJHZF99JQMOBrN3J1
LiMpMAw0GdeAV70QT1tQUQcQMv4qjr0DiZDXMuX85Ga6tFmlpy6qh7FbwHqqPVoE3xc7Lx3XkoDb
hwhJiyKMXe6+OlIgU/6tbzQ2abETHYDxM6A8syK9odPh22CJuNjV/NRo/k36LnWULSlSfLFHXAYQ
ni61i15YJatahTM4XN51mpDIS8AQhoH2oIfeGK0Dw3zqR9GDOgkeNAElpInvSajjnRSrt8i7ZG4/
sinWSkrSykBbUaekkVTsy2ShGeGz17Xn0FQXtgDwUk1URTtNZauSxjm70bVVmXS9MADC4QvPXL4J
GBH1WMa63tBMW6XnENS57YQRvzI43zY9/Kw2G1SnhMnAylh6rvlIZMH6Y/CHN5OW+hT1FexSsbVy
NQXd/r48IgjtpvivRchyfbkeWN+vcBXnq4xTomAfYIeYoPHcqJ6dShfo1wkyi7xKOcMz5alzTB0o
vxXEz4Z8iQ+3+B65puRXCE3auL/DBaSPHF1LxRrdIGLIocex4B+G5tuMEFfQ69vOap7CtcYtlvVC
2XGhcDIYVtYoZUn8nOfjYGLjlXFUhaPiTEZikTXvE9k3a0uypYIhtufReTjI95m02lFhMbKk5S3f
KE5n34WRaRjhoonnPh3P82poTnKASuqLrX/W8Z9OVGDjoLe8M3HrzszWuOt5y6VztEJkdQsHpro2
UEaEHozD8ggcL7sAL1FRWo4SukXH2eM5th/DAydg1734ZInGSYJjm/yZJe3FvGRueAiPrlyA9QNn
W4/RIlvonCCzMgiyStidwWQxJ/BlmsB6Ps8ScaTKBy4J0KoMym46sXuJFWuuVMvP+FdsIgVpM+sV
CPoX/cLj+u9uRzEj0GpPPL4B1bRvzdxalDPjQRz53cNTgr0oxSfjb3P9hZxrcEC4LpcrMro9bAah
fzsKYEaO/skUY5SwvQOe0HIZKCwLWVdmgv6jaGTEUrceQFUypzT4NlpeYRKO16yzxwnW4q2EaCIX
pM4hvfevJXiik2ZGVdC2QW8pztGEMFjcSfl8ooRhcScS0e8FZXWt1nRoDci98sc5gIvcichblC6a
OxXct9jXrggZZogm7rhSdyU3aWZ6g9+8W3VCL475z6rCq7IR1WNR7OCiOnm6neIS2ZsunmTPryym
G2pfU7bsET5DoVzbVLYQ23lghV7YIi5TsPdQb97ojnziS1H6qMvCYQLWaOoShjlFXnC+3D6EW+ET
ELP8LfQBhQB3xLsEmL621iKVmG5aP/0VXcjHWwayzoX89zNgnOZDYaeTJ/U+K7tPlOFD9bzenu0Q
H9Htm+kNDZLV5CS6iqZO8mgd3zgJW4mXxSL0o89iNytd4jF0CWnuKTKBbpMbv5XxjCMlt8H4k23b
uQwAGWqnxS7Q3J8p/VdOXOMZkbEIzlwLNY6IklIZFbRE/9jJAEDbPkDRkc8BU/xdkFY+lEptURgN
uJ0O7eukVLX4gm5MHPWxG7NJK8fAFoTqlw/dk1w2DNE4RPXsQWpzFgXB1hKKdU58tcu/paHGftWb
USn53ilr6KvTZHC/3/FDWOtit5ec+X2Mss8+vVKZvEyiQGRkIlwC4bD3l9v+5bJJpHxhLlOnMMZV
BwEn/8QYnrbz0qa2nCQ9Z2e80+fKGNVVs8Cr5/Y9nR3TIKqsICBF19QE0nnddUN5Llu1ebYx0Jck
ZDYYBRbnlnshT1yoepdoBnYkEYVxlopdUMh0/pzcmeUUyaO98zwsvn3hBhSIyqqT0xVWNqIj1T7O
V486+it3HsQS3tRMvzC1Fx6Achp9hbGpsMMuYvrisKmC3d742CA+FaQpNUGnAu2Se7RXzR5rhP1+
rr3Y7H50/0eZ8/A29PWF242T6MHeph6mgnUxyMqm8XCM/jFJnPMfuawfyVyt20D+u4ufLxn5dsN/
doHEA7ZKC7ge37GFBBXNQJ8tCjo/fKrtfAeSWPf4+aOBiZFqqOI0rOjB11HhMcqtatnX5k08sKFb
Vk10w6xpa0njpPleoJlQnV2XXQEeSuOQ7i7Io8rQ132T2Zu/x3XZh2rKh6HpoDpCTwCw+GIYVYnN
eKNGRBmmK3MAOz19veTyMwcebNnPVLdwMFYopIGh4Qk8+wzMLegGCRlNKnpuJ6Y9lSuzKoenMZNW
ZrMUvCwyV1jdGChnurLmFpQDhImOHA3OvSDUkF4oBuAQh0ectq2gBpFdQYrHWooFxv0EiOLmj5fZ
dH77D1vLI+Sh0lqb3LZF5NTjz+aHgPmb3Afryif+UOwaHarjKfQHR8SCQhBuK6eh3hIhxVTZmdGk
/qxEbRJJoInGEckk0PgZULD91kjkMZ1lqL5NeGpG1QzQurJ1FrdJMKZi2a0oQrJBdyzaheSYX0Rb
ZMRt+2MxeW1EgCAlbtupSFaFWN5QDc7xPYh5k58YsCx+v4WMaVGFaQ+fGcsuBI3CsHbQMJVvOanO
BaXJOFpaNzc9+n4st4fcgn+Cnxs1kqy1Mj8b7vfYjsDHhWo1z1CDBirSQsx9B2Tn4Ja+t4rEjBJo
sii61Lf9JeoWRxvP5ph373aGFCjkPIPfNbbapXhUUHcdQvBrUPrJhjXpQK7V0qZBwfCOVeBkhd5V
pc561vclGmmev/FrvOgwQoOJSvvMVf3OJfgc4x6xpX6n7469Ad/bgJu2fBU7Rsi8IMjUOQTNJZUB
juY/DLUFW6M4afkceDKpfNPHcjROadGqKUtEKKAb9Haq32KhGRqXnZS3qJgeiL5/HC0LoeCOOWt2
E9I368JLfqhuOrmZ9Q9Pe5GIMAEMV6fty4nG9aEcNqLfE721vc689yMyyRaJ+Q7HIEldnzBXMrt5
+suQYkvC/0XBOK6r4ufEA7sCFJYRb4C61SbiLzUPu22acVZvqnEIt3h5PJ5wMEWHR7gTzNMIqc2t
/v/8C8zJ+/enIN2Pgk/T6yq+8qJuULVt6CcICTX/LUcM4ZEHSfrm6gTapFo4xVR+5dTQ0bCVsOKY
jbhBZ41IaukW3NQJwM1xjSKbORmiwNoDMX5ePbE0pGPJGZevQh9/27Lz0A8J1ISEQYPR4yjKUKSv
ozaDTTyWG3JS7yJyq1IVYPXF55T7igMnFo7b60CGl7VKbAz/AvAGWu3SRJg7fp9P+q5MHyWAFy71
EV+eqoUtiMRdoO+uTutQfRAPNS0pF2g6s5RJRyeraguaOuqBSOjvwbaSCdRIonBZKEzzPr+axg9C
Y7sbf0zUTCq0yAsfX9w+54goipib+FtKzf+AbCW7+kkF+dkcxALVnxq1VJOHbJbfFXjTsttHHDBF
q8F5YEI8qzjVtWoN8/vwGAlNaptt2lvfMjp4ei+dyrrMuESFFBt2tuwSpV8nABDQLowXGeuvt+Sp
LEnIiWgy61sbcPaIP45831gvGzo+ZcKCddf0OGEAIIVlq5PViKOlus1KKu9lJMGcicBrh+rlgjf1
6lu4u4vQoXiftHZYp9HbUZ7jMRIoKGlnNq8KzFffRy6WCPRfdIguNciSRkBeqEwRSdWMt1MdhBmA
D8A7uhamivzmGLm39SIASrqs1gQ9iKTHHkodDyqqF8/O7kMtqustd57IUPYEWvJpWRX6zrdGRF4o
gLvNM+smI26sbAXPhXsFPJE7McLUGyjX5xmdTzjHIrJ73upaIb6RBRGase2F8lNfBF4mhzJLG4Vu
MeDtG5UxvCNptXR+ps29lo3tqL05OSShHkR85/9j2iGdRo0tQHcL7SzwVZ3aTNEUEx/0XfyJIBiF
fJ8meSsZenyq5oZIXhBuZdBoJ+qK9NhCJ2ThZRgRk2k9EQNwKpwq8LyWJv8GqXH/pT9WpWnxszkW
PBFJXbKD38BdH9IPaMYGIvbZyUGTuNUeBK3Ymav9PlvQL87V3V/lMqJRIs5hGeYQHk/Me8p/uiq0
z+rQZWGR1AS3XYzCkl4yO6GCeC7GbnFkSc9CmsMWoPu0AvH1Oiop0Qv4vaGuMi0w+KQT/ov3yN8y
WlEwa7GG6sjotnfw5/xkKWhz1NpLW7n1t+1EXgHXNhNZXNVMuO9e2K4UtKvXfJmXctpVqTnkTm5S
qQyTYUw4xLsKv1trjfjiy8nvQ426AUgvVKsmijx034oJYOr1VT2/q9ynj7bSG4TtO5gPZe6zwUnD
JstLUD6Pu+zuwInp3lDbvqRA1uAsnz5njBbb3BY1KC6HJ+seIVSBIdUgHDc5iOGPLJOzenjyuZY7
UOFhDlG+NpVFWYR3K7k0W/gvMPneiSal7jkofpl8UqPdE4Gsv/hvh5vwx77NW/Mqft4TQRTuSGzM
Tk4Hh1yvUhkxZMlpNaUO01aAynOjxlxlW14XGZxlIhs+6Vwe/XucFY91ROvL1CieJgP+b9pQWi+E
mV0/TrRHwh0wOYGFqwC0UNq37aFRxfzbCSYEIOUlK6JCrYxTvoZztT1NnC8ur930JhofGRO/vmE+
k569BuyZV6WdVegjnOHN1qt2iZXti5iQ5vIlrG9Lb/V9mNBb1PRThwMZK0Cp26+gwSEa0WlQOA0g
aX/o8F1mwt4En8V2p7LllxOLaKL8nG+TeNIN8UmUeEefi0pHvkT+vwKSyKPFPBGbPIOfv18MHLsH
Tk6g+Lox9Z4Z6iNX/NZ4X9ztFVDPhxnvGpApyqoCQCQFb6jeMMsB3+TtUVXHsqN4ojlxQm3v+B+h
5uzVQIe2cX4BWLhInwDIuH+ve8ngbSQbR/F4U3vEy0Zy1Kn1zF3QaSgi3X4MR3WGkj/8O93XBFlj
S036S8ZzvSvoFiwl3eYyAYbMoO4yyAXZejRALcQboKTwE7nnNUC39niWQCdn/J+sbMes7+2duCX7
Tiv/aqZt1dQ7Hw13rTFSawe1aLrcAV7R8k0Tekh4ujenKzntqyHQI3sBUJWIUpWUEn08sgmokRMl
rv6ynBfNe8ILK6xVOKw89cy3M9UtQscyBPScysi6V7n5W+87rDMr7+SybfDPmOq/ATo1Rxkfu9sd
UVQocHz6kQhYmJtrUACXZUprOIo4vvuWO+TT1bsb0tuq9n6CycqWwSYESWOqRdocrUTQlMMdEO/N
Xi6KB0j21wW6qpHkTWE3n0KPggCwaGO882WDOoC6RsjCewvntCPnaW0jV7ccq+Jb+EpKF5HIHrZW
775T8DgDoSrSZV1CQNeFCqeTuXUJjA4iPj3kahPfMIcNZfadQiDNEBwoZa+E8KbZ161YNgS9ath8
ltCWaI2CXIkOvZWSptS8U/8THpkaqyHuBEsYYwXF3JSZ6WbAg66WMDt7caxTD/Q+IBzZdFheTqJ3
qmO6s43dI3QKHTx422ie10wIfrtr9ii+LIZlRNKcTqBLhibxvi48GUki1TcQzRqVWeoJPfZmmimu
LI3YSmbv8ENyBmKzwdth/XJnzCLwIP1MIKrhUoArW2bnFoCmzJRxssf/Awj+76iW0hwzHnW2GxUY
RkS/k9ysqVCAh2Fl22qonnAGvI+KOlql7zi6rJmriJuWHv1uXW1P3saX/S9oDiNjxn7O2dFoHefP
wr1Iy/VllA+xYNDEJxsfjbockTdwo0ibYPuJXUf1SPnDwuNUoq3nXvfeg+0Xh5Fh5QgHxtKL9v+C
oomQGkgc+OIjM793OVDUst4COilNaCgeS0a5B8PU9exyIQBYhLf1M/3wcEFbkLS/96dWXUVhaeAC
9tePaYGr4IzC2lRb3oeO7SAFk1lp0iBw7cxATc59tm4U9GhLR+D97lgc+I2/8D/jEBfO8eRl+5V4
90EpRmKvv9PYAB1IWqQvyldM9wlOnOz8ApwczQjfUQSBBRlNWusUbqKJg8J9KPtOC1QSB237bN74
6kBkE6cWXG6fgUQ5hIYHfCGH1mAQeTmpJBEBfjMxvyxoMTgDTFabN3ICBnAhi2P7vbR31mttaVgg
TDDYeYLtf9pkssAPS83PQ2Swj4eSpmagxzsWVvtcUkccSQGVvlP1v0B/kviCHFE1bF/u4ywhVsDz
/pM7WbYmMixRAiSaHrd0GvbdMUIfaAouTfSakVEySjlyF9JF0Qe4YeEAPLS1ovAVl8glCzgE2997
uPXpWN/fhiNTk+G6rOApaVwj9dI1q483AK6cpqOUyd2gI+365Bjo3Id+FjgjqBg1W+63Bj/DU0x4
bz42VG4LfneKj1j1jE/0nz456ilamxmS2RHw9LBTElzQDEI7jS1MfuxaQOs5iN2XeeZxJWtMoxwi
kW9qhpOLY+gfYhzjFru0fclutPzTrvMAaQeCv+KO/uqBEt2MOW5CMS9G9gLvSmY8gQa+6EUj7t9N
BY3UgDX5EPc6QJXPSakFYOADGWQTs/vfxLzR/ynxVg8FftgtTv1hgafRMreW4VKiao7i2ZC2Kbah
HJtvAITcjZ5FgOaIlFKLivCYGuoeZh8m25Kz7Q4cacSu9Sp6wIxNit/tEd5fbO1t3f5MuxLdnXig
PYaIS8PM+wL9KAfkwS9a9WERHyPHHxRo+/C8C4HL0i8LhRpUz6Od62n/j4SL6DEwgg8byiuPaTpY
hk6Eawmj72TPcJx10aiH3b/h4BL7YKLFva093gILMOQQ3uyfIWTPQOte2FapFC8yw0ODk51VgKyt
mk/bxDe+QNfurePHJBCNGMkEflxocpAhbyYQ6bazdj2ldh6eyAc6zkafh2Qr1FgwmEKOMzLzs5mP
xcTmqqnyLYBl/lDL6qd4TvEvuEeig4qJgIHe0y1M4jm41BhKQYQHmofIHOVYflR12Gu5Od51DlOc
Tjy1IxwWTDnzVifFm6OZ0sEZ6q4oaw5AZWNc+X9xA46GzL9sJCEXKovQlvhmlJIbAyUq7V/Y8qsR
SiOhdkGqdeacPxPPB/2tdXrtSsoNg1n5eB1vKUmMyKG4T2oSDstd4yL+ax4k9iomiqjw6C3MIEgk
gNcRTM/C2MFBlhQMds56mXJSQ2zO3LmvdmSJglZehOs0DRvvtx6RwVe2+pHpiTHAh+1fdNRtkoUO
/N0wXr7W3p7jQ8VyqzOxus1ySp9qCgEb8k5nuU2RWFTfmFbk1Zqinpp/s56vlD75mNhWl4Ms0Eg6
96uGNt8PaMV5cJcJ98rj0UhsFKzlNivMmGciLHEBG1Phoa9APqnsS+IuyjwINQRUz1aKrhqjx5vY
irFBEcz/Esco+O4FlSNJ4Nvv33/uCeYZSdJu/TA6jLfQAtPX4OQ495QeVPICM2+m3BEHppSsORDS
y/X4HfcOUdevl/JuEsody2xOVgzwveBIVJOV3qFiNd88RSd+5gELzr2AGl3CBKACJvTiVgxFypl7
pxRzVGzWSoe5Vh4wp1biOydLx4B2fEBkWqbBygAwuZTJXwKh80Ln/iCGMQNtOCVpr52QM0QOw6G0
TQE+bK9ALsuqboEOK7cNVd+8wb9+Qs3r9kr5GiIF0veSentmwrqgAk3iQqU4pSexGiCjCrbvDnDX
3UMtQ1gJ2kVQZoACapNIfzRIxqsZrxjFFi0aB9Rspf0EafUTePUk+Fm4ccfu6rt3aZ7/zkRJkRc8
bQbCVVWr+ullCsYU4iJpl0ky5AVQy6+QugTmDKWIXRW0qX+ZIi3RdB9lMbaGELTzqOfLs9h5ruPS
l8dOeGItVVm+v0Lbtb3Rf/Pb7GqGVrFhOUCxbEOZZFUmnSTNHGmgodoC8OVoFcYzHh394hJDvD9c
HPKRKvIn8i8+US9YFhMGgBQwVz3BRvWcjz/sFpo7k33YhgDy9o7cI0e8D+6w/xyIYvs9hG5HrkM/
qg21ozxP8OxVOCrJO1yF/of026cPkJQV/waQc9KNE9IR3/En1zlQNfdM3Q2LETY52eBQZxJ0T+7M
KNWtexKw0rVY/lfyBj1fgC5CdlB1VKFJm+agcxyjyRsLREHqaYawXZY/ZE/L1JkZsU8ZHWmHk37M
E6U+b9YxKBNXCRr945k97eUWHU9pLyawxGqNKFgE9+P3WpBX5tCcmp0qQ7+8f+IuSx8t27cgzChz
rnoAa5IDjKoVMb6ZEOnANvaSoE6EZhLhcJ90LBPbD6s1vrahWW2mafFMufPpXoZhZZTwoAjaHvqI
milwaWRdqK1/jl4poY0KkyFYm1v0eH+75/DV5RGXN/SaNTPmYACx6CRsUMQARwpZT3Q9o3rp+woI
+YVFarWqGGSH69s7S0z5xouGGiF/7C3BrXEKaw8iR+qWzExkvMUTX1W5z7b/Zq3zrIr4I3+UC0W/
fYH4jPGwfuuVYrDrthSttMQhZpqOpyXx19odcAh6+iA3ZpGcWL5761p5N8Gtg3skAYsFyTvEOG5O
BXXpOv/O8OU/dcrzTFGmYftDKskFyg3/hngGGb+sLmMFLTRG8XtzEJdhBEMTVj4ijvxeg2O/qTmD
QpZqPK/0PIPirmC2cE61oBogEWJ4BzpQWECtoqjgO2GzlZEW+hMOFqv24zXheSNW0IK+XOK80Rsp
mhaeUt1QgngqbUaVBviPg/xH2rwPdefIdu35Ef1FLBASPYNPF6g2lP2eVVL4SggKs1gsy1mxloyG
t928xVJ0wXL7QLJlnpXFM8JuiLi5XOMzzJfKK2IYGPTzxHEXLPyFi0DqirrDAH42W+LlnrVFKWtW
FDEpizxoSNZb8FxInBM/wncxOypUrcarUIk89pwRahPyacPjde+pAyFGfpKhEFVGj8riRDF+hN8Y
O9CJe7231ydQbSR67CIck6I/STvveK0zFlvCS9fqNrHhLB4Ofk6nVZxN+gF28LS0hWOEY5KeT7tW
JKOOOdedzEyAzhNL6ZdytyTHCU6fv0pj1VeQsSQjOGZbUzxaaafiwszb5XjlCtsW9tuFBSG/FAk7
0r/BLKgyOLGnqNz08hx3ejGz3xp5j/hRn+Dm1fkncO2CJvLD5V3chAmE6yjKuufS9UT7i49yyfBf
CL3jB+2hMLpt1vMy1XT+/XOdby1Tm3z4RJueYM2LwB5jQkZ5m6MbAqm1PIEWTbfWCmUM9jJFMNev
itwLkNZS1fthbGlHTb0QP+9gmwuUNY7T1gKJLif0FKWxTmPBCdSZ2++myl+wY+RUQ00WgA8NI5AC
PrVffhePI0GFtPm2XcLbNPvtsx93EFRIyKT05pQ35uxrgyS5DIdxJ+k8lGe3i/LAaaCpeUvvFV9n
HeUSQIikjB47DuUSe88NTzjtb5FezivSEubTO9MI/Veo16CnxD4YtpirVIYKBNxji5DH5cIR5d62
e4TmWYrthehnUblMvRcrYA+urEw/L54cu0lRH580r5T2pVp84g4TR/14CniqRjfVksDOyWlP2RJw
LTmRQ6EIaiAdp8SU8uL6Mi4q2hQHRfqe2K2rnFVU7zCpwwMoG2pw9zfwBtdAhn/FZPG7SgUDrnQb
Gp6Vtv19GRgcqsCNV8HesKZCD7wAGtbkG6QrApnUkZLTNzCGrvSURosgFd9yrscPfFNpRrZVsF9a
tDL19Y8g1aur0dr5ffelqL0TsRnt6oFw3ZqFYRtEPIneMwBKi9PLTcJwRyeba03gwIwhnMx/WIg8
qJeXKc/rDxf8/H6NAJ4wFwjZcmT7WAgnhZT/XJ/frYAZga98r1Alq2fc1jKKgpO3Abag4rdALvbe
8r+/18NYlH6mEC2aA2uhWnwENZD4b+CRZHiDx0Ij15FPVzvYF/yeZ0vgpc1eox9Nf59JAp8T/egi
EIltq9ZwmUETZCmKZTOBesGs1wmpjoQPDCtLhuxHZeVpbKcOZr/XuYh4jAia2NGmZsEknrcxPHtH
E+rrSEOJcGv9KchTlx8KDUkTYs7mSscOUrnGxIdstqgqup8cUlQJ4/ko+9k/KvuURBfGH2LrQR8S
l31TGTxe+jPs1v0bejrdOO4U2PQ5QfKaA2Bn/9BA6Y0owsdfS/zh4CiVrGXX//o52GbfCluAuwcq
61hvPhHJMWxZ3HXc5idBbMosBDWSGOUgnRyRisuBV8P8ZymtlxfeL6RJBpdJzYMwoxcmQqOb1kqE
LxzGyW9CV9J2I7jjGSWm+JCLtTGLR2p36ouoXSbsGOc3Y37gLixk0oj5ohE9h8N4BBXpLEu6nPUD
Lm4a715yDQHew4ApaQTEXwwSRSVKMnagw5HgtIfg2jYk7xZ8XomSS2g3F6s2AcQB5jZatDxmyJu7
F+9XkBLdPaLyyC9kZG770py5kbHKZpD5GB6vjKbiM1rUUqvKiG+N/DRy23G5+1DD6Nczkfq0FAkx
u3X8janjqNlDXXeAS9PBiC5GAshrIJnD/apGS1HejKOBIpcNgCa9omm9TnXR9NV3+eMRpmx2p90C
sfFBJxxV+wWyEc/zY5M00vMSXiH/90c7+8LmyMr9LIp8Q0FjaJpGqiIncnrK5Py+9G4rrRm+R0q+
IldcoWIjhMLM7Xf7Qn7qNnY69WRYGaXDEe1wemaxUfKSyUqHbl+/1LRxrpt7gmuk5oAB8hIQNzmd
H81YNqpmWQc5WfZTqCNclwkPJsNlI68J5AWPndciG+QmHtzB8IcdZ61IKY2pgbZH8oRNHRKNKjCE
1Kle1O3IgmvZqqecUFg3Tz27+Zgz/yUYthQkZk64XVhxd5lK/sZ2gpoXoLYVfYUO7kqr1+EaTmQb
J0pqoLWQXY7P+vrQIDHiO1Nnfmrh2FaGnO4txnX19mDgV8KwSyNZ2Dfw2l1aMZ5OGxsPVQzSi+PE
g/0AlImz5Tzjq2YLojsWl21wAwQcgaOM1bRD19uAgnn1mtPmqN8TCu4H85vGy3j1Fg7cMxN+PnNa
zElF9nEeYGVBsNH1zNZ7L9jv5JFzj6Qu75+XznLXK74pu3nu0uSVXEDSbqcj6MayveQBCannie9L
g2XDNfmnfBR8IFYkG0XmQhfjtgqAVWWmrjyqTrF/d8xL8DEgWricSYFoxBKmOjfg0jMm+QfnF3GB
d2YargrY7gbiMGRLDDnayqArbWANKyHMh3Pro1JKkRaU7ckAGi2Nvu6N1sYUMCvJ/Z2USpfORo2d
pXapn7Y4Js0q4gfEvlzPZ3t7HVXqgK+qQU2S6hkhcpXLvszccZLrYn8m1rgizBg022v2/TD5s1HJ
LJSJPDlQ0H6AN1IJagfT4MfapopHJcPMhFFbeu+pfiiCmpAZ7GQP7W7BY91nixOpEUSi0E6+VqDW
YtfON7COjkBvHAXrFVfDbokD5i4QdW6UTvZO9NuWaQsiaZ27MMMBoDEvEV2IQaK08dBlYaPUJziB
En10IDTS2Jj+6LKY4xv73hsMTW51iXTaJ6yJXCUUyBG0nyzWDijazFQcfLYQZDLPJRlJwNznmNpl
OunzabE5u3p6njqMNlKcNv2fjM1eYi0+bkgFS5dUFilBO2TEsxDY2vil8vM3w1vvtzQbYO3qQm5u
YTFfzDeCcPObbY8L+CnBGKi9Hz7kMIUxZJ79u98Y8OEOHqCR5TIvKAb6YFGhdIfyGPQ4d2V9sK7V
CYIWDVccH61UmgYJsF2LJHDQByfucXgH4eeNGjnxY2vx8Y5GGpJjmJ2rs/W19pKrRmeKXVu0oelO
4RWuzJA3E6RbENcalr8LfVkrKtY8hbsAt+jX3W/qust+B77Q21vKRlZeL1NAj9GERmT8eQYxkaBC
gbsqPoJ+w3cEPYdCzueyGlt5ji0azJQY4h7sobJCoq7ybY4IYAIrNKKCvXrihsc38KggIDA6mxCI
zGy8/zNJROiaB95iQ/8CZAIFJhnBtgO051SEWrILV5jP3soJwRltYn+BGOk+ZVlFQxCsa7klByed
cxZRdsgSAGZn6Zqvl5gjGiegnV4xp5w5CPjRgw4UIa7zUgZq0sqsme/0RTWRtW5V6evssSzu0yKv
DpJ+i+PoQoSiav4wAPFKjxrQczMByK/cwNTjEPlsqVBIvUIF8Zj7gsT3rxr/HmDJSj6A40I4yoVp
KJUmIEt/vA8yAKHjDfiZAkCol++u3wrP6D0AW0mmeivuu60IWpi+y0vcn2Vow/EtEETwtRB2xCwJ
P1CIt/xyBb9e2+AmzRHqoEoSXTFtPJo7/2sss9QbukBiUI4/gMnPVy/ob7CFg/sTv0miL4TMEmGD
bgdbuTVGzw73+BFTDBU0SNWoZ8j7FXUyDM/qimObfK9TLdtA40dA0eFKIVK/ABEWiZ6kyeKk7f8s
hDwI8kjwgxtxL6u3sMSDjiw4SeLOyObCr/qqINMTy3trFflhqRf4IT1iiqZhMvFTeZISxm+jNSfY
xAElT6a8KEmX+whxB9E1D3ldmzTY+L+H8Rd1RTOPesLfQb3Feg8PnpVXtLmMjCH4JN8PMqthp+Ta
DbTxBI7ihbf+ZaS69RHJfazQ6aQ4cJhehfHZS7i1g2pNIwmUY8l/CkqQ7O2dnb5xtkxeYpcJWZK7
P6V+7R8ttWVH9SI9az90MSAUz0xJUwp0FCYq3gszB4qo6Zmo5Qz8m+/KM2SmroaL6t7QiaMggr27
nIC4PooEUVOmNLpRQigRagPQClpyjuyVvY6gljMphRARl7DiKP4mv1pzqJvSi9kAzCJLn9c1536X
Rnn8HuFwo0cmNxRcB7NzTgQJaUWDagziC7eCoZkGloCLlsoX96/qdhZAIPYfA9ckTqhZsxQc3Be8
/67JlKQo3bdZnrR4au2hx4WccFzvN8qg8Id0Nkr02Njv2m9tzN8wF8WKmj06lU6UIX0kEmN9U7Qi
XPXXGyFPC4vVJzEfLHX5CmDmAOm3ZBGVzTCFgu49uYOMA2JtBqmYrDCmvgED/vXPWgnyaH23aH5r
lab9cn+98jRmCcOmlfs6MbvALDq6vThwDSETcNWd2Ovc45uL/upCv13CbRRqrFnMiLBe2gbZ0710
ebpxOQbb/9Cd5HcUsImeU5L9DAlbHY+UcCrnIJPEKSN7fYE4bGz7bOkiGBoBNKmx1sldXc3v4gvc
rLia0Pj5WIRGQzfChROvig/vH3/WRNdFmjjcsA1KSDjw1m7DwvJcnl3PkLbezSUYaIggbgKCfpWY
QoFDV8HJpaX9AujXid/CO94igsF7pSElZO2PmkCerCsAa4ww0yisRC6VvmWlrgBIMfQmQDH6Lrn5
JlzzMCqbNND5TZ1aA6vsyQO7v2Ernp1VmGQ8PS2l3vpuqqjRaNAD6p7pqULJMHvsgMeqJakplPqw
XXXEaDNY5/DO4CZKiBk85ThbmRETPGHk8XV8pl1lY9JHGdxzC3NEEXmzo4yckuVCrFNb0VNTBSt9
rhUXgnu8+saSa5mgnwWZiebd52jXMkOG6f+v/HQNUCalaLK/dqbJCQkH2vRJtzwxrLPxcbMQ+E8b
XOGeQ3mL9HIhLxlXAwwvMRQXPIv7n+xVV6zPy1cPcR9JRsvrz8pyE5cjrfQ6OZV9uRsBiKWjCsUd
FGFAMADiWOAE1X95Aeo8xw0cQkUGMVAE4wDge2/4kV7jMhBMx+zfiF6ykjfKXaGRNuQDLGcPyYOp
+iOIJGP2Elr1gCE91TI0WVvvhIS68niek7MPk+kp5Gif3jmAGgBwCS/S7tDuvdS9pgvYAEMEh09z
ue1rGMtB49uSdutEv2k+0dP3pLPRJmQH0JVPTG0qza2L/sT+/Y59l9SmIM/8ysRbOfHZAKjPU8C+
e9EIl31wIc+aSurYiI8XNMF9NN6wcjuJg3wG1Fpn8vAcsye17S9fuhRGIMBOQU50higpz94S2Le/
ZeVkgt5Z54DbF2T/l0QFCT+iHCN2+iEMh1N7pIGRFEYOCA4ikhlWFPPNXvRNB7NtKKFvv4HunvqN
4LVUeSCKSRT/VtilaVlSCnzQRAcRD5fTBZMuzBzgSD0yhBwfqhwjxpoOD1/IP9H93VsuRdGZWtj6
8gPzsF4xmJkArag2VUMU+5HVuOQLZF87+3bXVfX36z8RLxk4oFYAKVqTs/+vT8CX+jNtMNRl26SV
8+pNvy7uwkL/P4XgGF8dFLuCG6kZKSxsfM3cgm9ZGGZEfkYy6AiwumwjDOPNBp9FM7bdGZAEN0YH
jp6F4raAOgk1Z3hFTuMSgep+tEQMfeu/WnXiE9ZNjFsXm+H7fknspN29gsrv2ZjNnQUq0871vVTH
z6fU3vshHBIY7xGH2613I88Vp6PusF/x7PLb/ceJvocEX2aW2H1laRpzJAOdr9JBI7cVrMx9Nxaz
eVXVZYC31l+gqgUrVyoWB/YNd8qIXeZvg+FZUA6mHLXRYx1tpKgi0tnjS0LqKIMd6qwVZEyUxIgq
TJT/+qsEecQjuhgCR2Gv2wBKxpDZMsqsu7PvGD1BohA97IkbwcLldCGx2iPen9lDxsm5M0DOkSrF
xiEMPj0xPhMffsHRmXsDR3xaUN47cLJ1ZVMD1dk2UT0j6hVSguJ3gZ6QkpWYASEYPMRB5JeJBUHI
kFhkrR+p0D8cAM/47b7jd/t/XwVUm0vq+iof7/6Wv2maousZJcc9hl8u0KFdUxNpm3GNsTq/aj7t
mH3n8eX9qbsb01gexZLy5MVBWGlzjU9PRXxFGAMwCx4P6oxb6XlkZxFyUAhZXjFWLgCL98iIPLRJ
m0PcngOHRHOzs/UZcM3Xf82Q+J2NxvfQCPaM4OMOLGCMvxt3wAIF6CrMa+XQvqJhyWE1FBz0DMVW
JjA0BmeZdY297apgL5XnRFS7lPYbXub8LDHMkcEIulAN+lPX4br2Smq8MuxrtkoFWrb7Hh987igR
AZSEpywP1aQIITIRVWda8H+2vw/fUaaRJlZ7ES4RiTOMdZWjb41k9z9cmP+hlJLD9VpNRo2srMq+
hViTBacaHO1LKEQMASBzewdK/ojDCb6EeCD9UWXwH2vHvG1kmpeVqCbN0cRRvXKBVmS16Wn69Q7A
uxOINKqMRXj7QxTsMKJawbNSWToCFyKEfzm7O9o7Iewvy43Pp9E4YXJ77Lxc7DkJOQSUnCLI5sXF
7Zm2KCHYXXoxROdPFNG8lG47rX9xzTho8sPr/rsaIczIbJ8k0M0Lrp9UeQciPkure7karzZMVkkq
2vlJfBiPsJoFRcjtCufiYPwfShVa22M+N5p/pzTepX6eMhS1ydt7chai/QLqhX0wSPHlUP4T1c7g
ujBUP24ZPAH1Gz4zK3O0UHSwW5rJJYWBS9CGzYF0RyTngAAdBzI/XuPg06DNTywS8CJVZiMwH8LT
BN+OJFACRe0P/6F03uktcHnGddzBBnzvC4Erw2JOSSjA31tbE+8wBEk1S8TKdFc7tk/sXntyde+q
owVBfGbKKPVvCpsatE1XnhRmjEEh25x7FjMGcioI4Fzru1mYBUm2j/Ycnzr3sjscxRKfmtNL9Xqt
NZN86zmecOC3irq15DBwB9jcn+G1fVT3X00xf0sRJkj+w7GJpyRR4PfB3anp/RZSJ5kSRP/+GI8E
p9FccT9G5aqNJmUGFup2lGxmCRW/ueM3sVYHfoUIWxyEnXSBlaB43oGyZPPmQPXy5TYCVL55/pcu
/4xvIiy6smpfhOc+1HpoPoS8lImV+yq8KFulrWBdCEVDdSxGZk1mvVJEqAzHtJmyPic1L8AL4QEl
nqqWFrkhT6VWaW4XNMp02Q+bs8TLu+CTGrKaiEFQbPW4XZcp0eyi1gKam/Hiz3K6J3c2hGhnqGUr
HiXc2f5bIRCPfFFbG7AWADGunQCNlXMG+KYA2TzFNTopuO2c3DyMyK+iQQMMcXF7Cc37SOvIxen4
ASiBwsTvxetIsovES0uzvYWwZtfPxFyoBFgf+gLQgi6sX1E1OilwXmILtFJLHDv8iiXxvHtTl6Ve
lS6UNqcVuTJ932sMg0RtC0n5k/2Kl8Dxyohx9ujjs9TDl9Lm5Om4opxfhIyzVRgngIy5qIYFJFdS
cnySndBNT+Gc7M768JegVBhmfTOvDgmkaWk79BZXdrVmJqZGzH8IWzcZsXsgOeBvZzMd+RAyKxSc
4F8sAGgKLCVAfnBldtWhLA4hvExxSIxJ71uWtDoFey+gDUEHg4q2gbTgugZOMUm1mjuH0jndRpZS
265Iv0/gOY66Br8Tx0bA8uU7VHtcpMXQJWzk1Qr13b2us94bvEqJAnnDZwfdFc7ii+02CIVgfYYq
W+dcDJcqi52TV1wsFB1+isWqdoABVFOfKwCTe5YiRdl0VSfUzDI2dGVGRL1JWluLYXprsCqOvavW
xZdUQuQRH3zQsAo+aLFYe3+xg6y3jFl1yOsbI44AHFeFo+gZKWt7KWMnvffkLpOwSbtcOgLjSFRX
7ugL6Meu9XTUB5izR2XguRB2u4cnfWbNaEGT8yNP8vMd+JOzJ9ltSWHL8JcNeT6LGkli5skHnvSA
KSbK9xW4KeXCoUEYD4p1f4hoQi7aLz3ihbhVvgSxTPymXHSRGyp3+r+6nTAJ+KLyYdi+YMB6Pbg9
oPBaVwC/yQfUtJsOD/qiv11DAddRGN6w8HD0+y+L1Xs0PH/Ctz5UKgdzLyVTamO9NeW5LiJnFjSu
Mvk1fkP62ojICcoHQsJXIgZSXy2w8UaEtgtG/bdwhGlnjXfW2PhFfhtF9iysbtja3m2mutRq2oUa
uJ5sKFf+9V60YobiJeOD+iN7SltfB0bJhwz+pO7ubouTL1itet8JXoOICWTEc+S0UNLfa8wtakqr
lVKl8xAaNNXLCnov9YDKdYhMK9fCiDom5m+DUXm/elV8EB6XoAdepkDRwT1XKC+B2N8ZycLHiHWp
xphfmCJkaN8rc/C4nLr2F40Mg2Drx5mAdJy32jo/NSKFSLAXNvCWST/7/gf9LHabfCbYx0trhlKm
2Ej7UcCjzK8l9jnvDtcbKy2sTcxNcCQa4aWsDZZQ/vJDrl7FIPoD135KmljUqmZOC1yI0W2yrP7s
Ddlv6Ihb1Oplqz+shm2B0wGLS716tQ9sC5SmdJwvULv4Fi1uRCQuF7qqx8uBjCrnTtzUOZ3alX1J
YSaF5q1tZum0LSZu1k0b1c5/Gzz2AiSM0s68OOa++wRxC8RHp5nsEPOLTwTiJ08qUal4HJlZO2sw
Ygh2JnprSRcqbKKJPeGjORLP7xD1KhgWDcB+Eu0NPb8LZIMwCkv49Gl9TY8RbrIs4RJhJxyPUro6
/hYHVOSLckjhwVy8ALBsVlGVBdDL4ryCuu0eyavKQClToDH96REDWHL10Sw6Y+vfcNGy99B8CJwQ
V9AZmu1s7gasA2Y4PVEtNfc2o7hkoZwTCE1i9A9tVyTPL1VT5stoysISzfOkHNkV8jLyYdSCJndk
5Jhmei+OHq/rNFE/23Nh/4zYej1OooHiVmaEvlep7UY6W3pyPt3dAV1j9QhMMYPppSGOn957O7es
Eli6AbrkIEH5BtJtjmYiQl8c/pJ6qQVVYg9KIcDaq3Dr9CkscNC4ELNG7OuPG0uJTn2CgQKNQ0fW
rvmhqi+OphVz9/q6gdrf1JpNpWm/blW9E3UM92DaPg6fTuiRCjT8gaeRYuSFe2dIyhnkPrt6ONFL
I7CHKb3Bp9GplQ1MlpE02h9jXgW1l6YLHQjemLBNMHxKG3sU4lq9h3Dpht0DaVx4bM523lP0CO3I
VIN3g0jpxHcV6aZnOtad4Mt8hkmxv7b/wHEPgVGfXWEFmTTybh0JDltD+CgQL5qSYBk+DukKCHpF
JEgNQxZjcRJfdWJs+7Wx+k9qw3XgH8LhFZQkJwhyXY9q6DNx3Qrrg65bKsjmiGWayK/QD7sfpVC6
bWoADUbvgEatBysBVx8yQRCzzHMxw7JDxzgais8jaEEWfKsOmIAd1iEkgZAPtK21hOoSqSf8sMIk
zaSHAkaAs65qmXsbGyCkMZpMo7Skws2FyFaiSFPba2CLImp4TC+VRjPkxBwVak9f81QSDkL3kp3Z
FuIQk2B0HjsSVDrORc96Ol1Ll+W4DPwKTY3mfULkF3K3ytv04NZN7uAm+7lJbxWLBlq4tGLD0H6j
z+H0rT4++wEXnsEOMEnfLbckKDaceLznjngfngXo/luDwbqIYv5hfsmM4fHFwcAFsYMNqGcdbNr7
Wt82mHrGVyX0MR9aVnXdDTWuOJkPIg7AzEbLIrzEyCqyR/bZ2p5hLakHapzSRm6lv4vyNTsMFxvm
+XVzn7ZVmg78R+N72beJodSRR3IqpkCsux5vUqh/JfmKdOkjGcD3ABteLNKBzqrZKbHlUaOoW06m
tOHvXGJRJjauxmga3TFXc2jqhXFMQwJ+0IpJkNIXrktcgqzMUbtPdPsLT2DdURqMUxa0uRheuujS
5xDI09r03GLM8ZEvQFDi0C9gyh3F0a2dVhSOAAE0kxo/GQeFT0DpiM3u5ppCExRhYoBDtI13dye2
A1lCynzjYMSMbhHvCeh1ZJ5U8Ur1tTds/fGZ972EA0EBkdRRUfflazwU0hNXvoZGH4XwPravmULb
Rbs8D8eSSFJMMcSJWuvxY+fHpLoyHEl9c92lcJrCdolJDS/t0OlHaHcK5NNSTREl1QXiOOk3nwxX
6qIYHYqkOc7eVtbfifoRdpxHqQnrJLNXIHK3+Ci6Ehs3viXbP6vEYjZYsgwpFZFT3APk+3f2nsHn
N7RWJaVkanVEpUT5T3BgtbFGhemjJqgjdLndiNRcFZxjwMxHxhejDtkuLw0pQVt5GWFWR4Ssr0Er
rnyuelkcATydrRKilp4DslzFBZrnX0Ja96QqOeMY9bKvMZquHngolpVVpdN9+B1Sdf9cSioWD5u/
jwYWsBrdu19ei4rfg983xOyy/bCZGG3HNLxi1LS7GHdnBuzDAC4Qlj4fCKRO6uqzNtj8YGPt66D/
nk3wzgJKClSp25P2VC/VEMBJo2lPlupqn8p0K8vdQ6ewNppZfFkP9svAtkTl3zyy8ooacNvKjNSM
AHehWhqM47avetxgNKkIAM+w3+7NdqlIbRElo7DCUqxcm9esEtZKhGcafFiWxpu5rRQZpdf/3qvl
Xofe2hT2gX8DmOVWcbpgW1Y4hIte1K8ctYf73RaFb4MUqHqamrVx0ysq1S9GWBvwvJtW/QCvlvRL
p1eRR7DV6v6dM7/IT7zjg6VarnY8WBROR1oY4YYJq3aGkWKz/un2lTT0RoO0dFf/AfI4Pf+3/Pf5
9unZQFSff6ZIRaKvQgBg2+kHg65DKP5g9WloT2XSSqiLdHymJBpthRUbp5eGeK80DeTOGkVSpRC+
adWZJf6lkS4Ww20KDtWU6cstocAsMwxPt2kYQQYVVefV+Px+l250W57Bbq+dYrlNk/2CwKw8rKO0
7GKlJp0JxBE1CzP7/doSFSM5xekTCZloVHpklyXOCv3j11PM5qSTXB4JF75UrrwXOYZOOtKl+610
ZlgLrBYTgSnnfSaSIzYGKth5tvj3cM6hqcKQrb/FitrHpngcV+11+pL4hjlcGFgBS+UrTh8dENef
agbMjPs0RRJoNpI2LuBbEgEFX/ejVk2e2bdCQq7QJOqdtB/tkXnFlBOCfAsn6Mgg2IgzQ8m6YEx5
yf+cYIm2O8dILfr5357Ny+PauKM9QhKQc80fd37Amt5Vgk03LJ/PbH1Wt69Ctx5HnZPnjwLsG1Eh
13z7TJD5stDvBTvG7R4nggDhK0WRiqK0XYZqjd6erfZr2Pb1HMuksYs0sp0VsXrghAubNPs79yBs
nlQ1mVjadPTZExhDsthWpppqoliQ569VmAJxP6UFh+/bxMrb8CvWsZnOsNskbD5Lvzm/RZxcAS5c
ZW1B5Xoi3Qe9GwR23dTrl/0XBcBPIEEiirmgAvWsER0Hzlt4hSqv2mzAMwVGkZsdlsKbqNG+qS+v
krO6W0UPkutaDONPb0vriGpgcVP3tb6C3MfeqFD9QKfrHcKpfussHubsofmAxRuaAHNYgDZKMrT0
fIb1vdgP0lxxoUGrs760LUReO1PYk3GrzNTYRaTu39sE8t05tTPPtrodDsN59+qlRDnW/qdJRxOf
jRZ6fvzvqJkIJVkLJtM0OBDIg9H/uEDH5Wso6j8xUhcG+9XaYaojZaK8oWPijKj73ueSlNAmUd2W
ysiarShxRpxr1i2pTKVu3fopODkmGjMEZ/0f0ezN83BEaeNe7LNQMX/56YmtpMAdLeC2EYvYovxe
rrGVJstfcmLWyPHaqYkGcVl9qwQKJABQlA21qHe0NvFitNdIpjGnMIpab4pqN3/OgRhT0QyE3Q10
5qeQJIjkK+6B1M+3PPJWdxfPM0TXmmY5raspvLhIGPudvCXMz2ab3tOasGlHm6SLDmiD2WwDomWb
xeylQud44IJE0frhgVlknFoJjasR8Iu9O80ndahlzPCqGVbZ3TOJ6ih1eSkaJhJns8BITzEEiHTX
dMGKK9HWoM2X1jUFifu6kcN9Ag1qfjcPd1Xv6lvUWv5d9zsUxDDcpS9xTa/z+h1sAn6TsRvU3BZU
VJV5ysmZaY6ll1nrTdbqazEFJ8nmS7u3AkcmdX3DKAy5nv3UVkvjOax7ddlqMWL4u/BNAXVKfZnC
KKN8g8etI9RUvHyqsQyFoqWWDGn7ib90ezaRM19Flee6Tkm6mTLSD98bYtCuYQAZ7E3OEV6hHOQX
I6IQh1GBsNAaPMaM+JZBhEOBjMTRkMUJatlUsbyTqY7YwkfCrL9bDivGTELkYz8bt5HJ3uB7nzh+
ePWgm6VHi8caiL5LYgpVf4EkcxlvKdo18h2mqyQAzx2PONaHMdep5bHuO2atZmag4qlHxO6IFJoT
h52JzbhROnsv+CONSwSzcvRAAgWH8OI8KhWhGmOrhFT+Na0LKnIjBR0HuHwnVSxMMfP+CxbuyDZU
V08P+FTapU0RhGElxjdA5tLDYrLyAgs5RzAsz+vC+347eK7N9waaIccJ2xRt0xmcg+bU1KmlLqne
izsyKC47srSYql65xrlOn4pXI6H7hfhf/oxwZpD7JPJ3nk1bi3z8dqBYirjRGdnbwSFQUM2HlP1c
TIXgFn6int00/WbV3gFi259nc5z2LPTrBLv+gbegHTuXwjYKkOh5gcO6g2uC9ltJIP69ClJkakvt
eH+HHOcqoUBHUNBPlhD33R2SyyWEBSd0q7tQFNFC3monDQrUMv2e+if5QFzCn2ejddh8yGdQtlaK
dkKJRsLU99I0HWI8Tupi+LG4RNULdtAn4Zcm53OorB0uPYpMGZRyh7we6kAMc9gGZc+dU20cGn0K
2eXl7B35HmvG1tV2jTKPvGLew/LlF30yt5Pb1Fm87eYGszuVNlNbtQ3VhWJsfsW+KBesr9jpwQUf
N30UNCTCn7isLWXo6LT7E/kxzALKfUADkGJ4lmZ0sg1GeHA4e+5N22jxBw0D0E2cf64878yI8lOu
3Zlx2hj+Us9lriT75y2Jy/s7oWciNkfz3C3DFk+//Rda8Hnc/outUDRMQCHDwU9OWgpOOzYgZoHg
LqSo9p4gqDdT/azBlifUrrQO8LaCu2qwwT1lEbfw3aupNtFVfpGlMGe0ZfZhIaWz2pTENniYa+4m
Jdkz7DCkvu/Gv//8s5kRj1ya6LI44la/+ocjX2ZQHlewVNFBQ9Jo5jrXVRqqeUMnYMK4QRv9F3kH
LXDC4lvNbytxPrih2bDat9ROvCGUiqap+oISMJ7mH/uo8W5WY98fVE4JE6aEm7VntS7htjDw1Mk5
JGVgEKhtSWlnhDTrd4dbrI5NFZ2GBM7EZSdFq6N4NZ9ZKIanYvfJ2CVMlnmDIQMT7iZIuQtuzqnc
1whLlwUFO+G+3bYDN6Iu5gFlPfHcB39ScwAUFabrB9xPjhnA50p39QrV5KLLFwZGIiUMquHQgKfu
g9RVimWHNgILlvYqfE633f55jbef6wvuNalhnbIw00D7/awihpM4MvWOzM5AN8PKJxJygNhxajWu
K9XfB5dalJRfyDw9/KPtNqKzv3YB9YjbqXJSoj5lfEtG8OctmhzllcmRyRTtJ8xdHa3nxYF2walm
Mf3PrIagvshE9Yqqdn31UPkkQx7WAHV96BAdvlguqkYw2/FJnTh6DO4SI+tNkfQIy/b19528NiaT
d2T0JCNFkgd3PwWkeoUDAzUmtPL8coNc1fjlqafOa/3qpbNlPKhzEC69Kp2CDUZ1gLMn7LjyBXPU
fyjbyeskV70yPmoLtmF2ekJZWm+LmDxE/PSlAFZ3EGB793aXH1cyAaZTX48o66IXMUwxXQTLcWU1
DV1jWoMa5/5dO6Yu3PtR4yuGyGj98YuDLQpNNgt3PPvY1GKhwB7ZwYY60rMcbPdHbtaoQA0rI66l
hg8YUwdyVsjBywFEG/1oE3bes/BPoejwFREBudI41mJZJsIbjMEOZM7Q/ncvUox0nDfhyRlGIlUW
otXHdVItk9b08SSR7v0+FCo01K9BAk6WlSUmkfXCKN6C/TpvX99jddfcnpVXNaJqfik8dn5GoHGG
qNNHzNbRdIztf1c2StVESHohum/o9t+tfQhdwZQ8SRywE/CCoCigQeCQRcErC8TYJtieeUlPcBWV
GAj9982Cw5oM47ndrx7+o+zrtsF6U4yUtu7N/GEOqs1aZFkMxmAXbmoA2uxUpqNV+vA669qd0sjl
FE7UH8kVcGT9+KLnz6WESThQ0HiocCatvB0xKIBsz+ND5smoAi00E+dBTPbdp4UlYsHsL0yb2qFD
rgFE3uXwN66SBARZkVq8q+6FY4JYG2mG5sdDMl+YrWzgdv7GTNaM9zybv4deLnb9drBO5ngHEoUB
4kimvnHuX0nwNwBpaexSdQLJmFSdEZuV3Qpgaf/FVvQYvJsKLRgMFgiVhAa6nRL1AFoIHe6gu1vj
HR+n4EATnNBNnUHny1pWpfD//R9a/wacERPkjT+0JdkIssx4ieCVG7eYaGBDpa6kr5ntVNe6EyDt
q2YcIEeprgjj95bD2WU91Dnoa12WGy1z3q3HFapo/XD4EaFt1LpbAt6Q3u6yC0nu/fXbDDaGIoUS
jKUUoXZE6dfFZ0GI7hdSIzeYTD6gj8hbAoCVPiYa4eGDrPN4TxQrJlM9epA7baDDIY/MqVwqmope
BxcaxqT2zXed/xtYpm8kN7ZekcL/Fxqy40oHZoNUfBrU7+FW8v8VgJuNDgY3ApRxJCzO6ZhEV37W
gt9GF1WjFbHBHddertJ2v0nTTxIJzS6RbhRLe4Tpe8ImFN7QLXMNJsMFEebIjlNJ+2gFqb9a3ghl
GK/IlREgZd6KqLzNqyGzVSEKPTP8nG48ybx6IBTbx27q7ZoEAqMtwWbDAq2GFeJp/lUJlYpJOcdR
HU7SD6SQgtZ8UfFpEkkKaKElFpenFcSKg9g+0nGfYfVdfYFiXeFlXNg2i/sp9gIGC84gHclY4aIo
uycFfm2KYODa0NdEl1Z/6LdU+Pd+ZmZlDsEQPnHGYSw5J50QJrsXHF3YSccEjPm+9Yji6ChN3ZmE
A7MGxnGfFLR7Qy+s7HwWlKRnlzaR+G+mdN39PXa93CK38Fi93BMME9OP5kUGnKso1TfRsnct0QPu
78rTAkvNuJu4agiv/MKcDbSuzIVi0wJC8dE0u6wBwIMxFbrOTIV6ptvMGHmiA5iQ8A/dcB9uBVF7
YVI98S0+C91SyDVttTWv6RrJPTbpdgoUmw0EKo4CRKkFQaV7qZjefAWQ/gOuKzke3bU3FvUp8T80
myJDGHWcIzylqVk/+HLMenAL03yEy9EVZuVCvuYio4G8ILsYxwQaQLEJ3b/vKnug536vVIRkxzha
x3nvbvfGDGIaOWCMER2QBdJeLZpUkQaNl1AzEI3qJYJ+vkt3nLQnr9fuh7KptjIClt2DrRUd5TZX
wMoTJhSjuCXPp8Q9rlG/Nr1X3SiJK1ZiEn2DXcQJ04dz/gAJaKzR5jUNIZJr7I70c6JElTjD4j+d
cLG3SWGm+NKRASQfeiv29tqW0U4KlJpwyK4cSkwpvnizzsJ4H8WJFVs7WnGlyeoNB04bLASTvtsA
smKJRk7WdwuCeqryXe+V7r7IJmuRzytivx4hqifqzUJD0BH+NktyGNSQV5p1NWfhk3hMZvc1LfyP
YeKz5OClB/Lms2hYh0ocy650NRiFztJzfJG5krO7EvGNb7B6Kz77cDz794R0cM/L5JDlHaF21CkJ
KuWB1PWLmp/6vGW38fELiAnxW4VlwdeAo2Z5XbcfaEuT6E7JudpVFu8QpC4MmTXRD1fuLXtM0Kho
gideWuPvRi2zD4uAEWU2eBaRTMmZ2RYKOdMNZRkbK9Agp7E8p+ISBvQKbL1qPCKG1kxwqdk0Aqy/
kmG5GHU2BkBhkARowQotrA1phzEHAO5PEYn9+4kPk3m9DlBe/BcdbQaCwInZN+TMyldmArpq8uzz
SrjEu756iocuLxMRMWaY488j87iSb6XWqjYWGX97Ic3p3/vqzRzoxbvOfOZvMeqrUC2t9jMRnROv
3wJfbjUzjQ8GZ5uyHomFboupO0KhG3TNvnRHM1hQfraC8IyAC65C3YCFBkT2FcGniGGawiwQXrEP
wWHThVInBQPtv+ZhAaYpb26qygK64z5VphTdqEF77YmjQsWDCtyQGC2hk+vd8VqxEQh1wXbqm2KJ
ND1MhbjW7qOWUeDycSZfJz9vLsSkbPaU2i8t7iEPJUHmxuTW/HYZe8RiWC0V/GApqB1L/crM5s8M
hOaUHAcPnZWA0KYRrBBdbFxEH6z7unJHZlRPlPTKlj3yiBV4BwXsyHYi7QjKmUU6eskBziIvjmuc
q3NhEglN5BKlkoKlI2Yhr2uNUSdY6+3wNHJMeZ65pFkQNCQxcTiAFPik8Gb6URzlkeh2SAbyx3fl
oaOqliHM+cSOLTD+QN9HYxUzaIJEudg6b5veb81oc8hcjqOjlAzyJg+d4/wuTstkUxashudKD730
dTCBPBdcB+rIfWhE3kx9fTb+RPLDvaAK14OobSWxWyGYRdqjQ3ij5RzrfNrkDIYDRRdMklqwtUbG
rDLem8dUd9lux5quxuOJJEExBvUJkxVv/QiRvGY1dv2C346WxXWnDB5pmyVDEvfU9IYMrd3+3qvV
ECVgrp5+ZJjxloLXt7d9HpXpHS+rj4h3nu7G74nmv1qMUI+qbx9F4txm3qNrhdwQV07S08GDGtP7
bfiLBXfhoOKbyMbQ1MWef5w34PnhakFKwERXLmDx1tfSalDWfh1T5vub3alAZPItqo6odkYg9fAb
Ti7h9u/rU8gTNAqAJU/dBrn3jV5vGFomYgM5R5Q1ZYGAQBBWGvxh9a+/pf7C7HQbTcAgSYlqrUDv
IG6vriXmtDop9N+VlYCwagG8tBJyHdPDykmzTyxagSzLvLLGtECqK9yUB2S451X6msNR5oFRYKkq
cr97wz5+2nwMwi5W6OF/xGFNGOBjj06pbv2OxReXh6RwUVWInyFUK2W/94vaqnL+O7shpEzMZirJ
s2/zJV/j1dMywxMXF3wqIWZ9ELGSFMbWBgIxVHKL6GAWTijPzcktoSCkrVAan3EzPfrFwc5Oj3DG
82KUjNQNg0iMzrSOkNb6OpccozWLsJZ9wlN/rrwsCiKuFRKkd8accO2H16Dle0XBc+CcIcvnQ4C9
uIKkDtmylR96f9phiiYldgNY0SB+0uRkLgtXQjb0U/hLF49HfYLUTdaoO4zRcSAhIbYB9kmaAi2f
pq1qbjFbQRxhsk+v9R3inh/PlYfPBRFyeRCob2xlo98P9RWCRex19cbaLaaM/YVM5TDcTgh0sWEw
9GGIPxsMoOOu5aJ8JroO9mtltAZ6ltOqFckjx9d+ThONlt6nxP/8qE6O+6+nZVx0t6pQGmEe7cII
pAmz9CWIAzjuDKZ1gL/TbuDIqQ8TiJTjd3AIq4tqtgpdp6+BXkxj12105h/4IHwZ9y56tQ7k4wpt
uE1SLg6finMsvcA0YbXNnb2KRcYvoEylzw7pVaNEKh43vYnuKE/4N6SPB77lQzhPgKla7ERWs4mh
qGuWvCzAoAGnaiHqMTsIEugf7zw5YB0py33MyXdPvXmYvQIdkrI/wy4pj3Mt9oS3IUMjDKSst18B
GI+ViTrgUadVXIscfI0RHBHLY76NLwNVIK5X7CTZSHOUlaLDj6Hn778rq/35k2vZi6LNB0aqw1vj
7Pe4sThF/KWXBfvZqWZlTSBw0esZNSZgKxlvgWufvbHj7OoAVWkTKN1Nq5kzz16WIk4RyMMyW710
zYCfAFQ0adrxCQr2j1ba9Ku4Kw5t+5xI05oghaKSHFUHJ4ZgDXgJv+Jkug7FgK+zKzyhsY0W+CKe
JJ6cF5OGX57mTYQOikCYvUyp4kjJZi4f7HwlrAwsy0+v0a5fsYQJd/eU7JjXlLxwOP6tgdvoJmDD
L9c/RiPXgMod7n7rg5CwU4ZZbbgSq4Uu62o1dlja/LF6NfFOjfl17MPCjRQm6tvPNQMVEZBZ2PYk
A+l7t0MFopjfLL/u1l8cyawBq7TGvc70VYBhUHZteLC8qgz6wCfAZyzeToqBXSHoyd+/Zvm1j3bx
ZoeuIB1Hy6jBbmkgk5lXA+JUJ1hxm/cWCpOiDqQoFcY4J3++k0N3BZS13R4ahAPO9WajfsNNfuxW
igHqgwU5io4op4mO8+TgKZ7pAgjDNjSSA+aFyCsS2EJY8z69mmvCJBuG1sUi50OASdBZ7HxO+vvG
XyIf4chNlte16oGzW7DYRR8mQcNyFV7PqWPm5Dh+SxHFBW/Y5IlMtbe52RXdrn1Aj+3nGvgF148/
iN7vwIrLpGx/DZP8u1VJBKTqUoOZwEjaStN25B2MUBF9ktHGR3tOljf1AZ8abVcx/pu+s4dw9+Kp
DbePRIQzvfcw1oW8Zi/kFVC1Zqkky82pOQ/g4DEq1FB0YJibFUlu43faaKN1YhwrNkZSnbcC/BHL
Pa1DQkk67VGEOaP4kHEnjH7smQe79iDtRxkaHm8sn4RfsuRX+9LN7fUez0YS0o3CK1euXutOPbpB
qbJaJ6vfAORIjjuwRYZgpJZf9V1/wJB0eG+5t7PPw/hu/1ROrJB9rEzPHXqVy8mNJHD+WRjS/pJA
2Qu69YOR2tEO4XRZl3ieKiKZAirBVyVYx76bjVEDga9wOI+wvV/pemAl9L5UUJKTvisZ2xlAfEvq
oLIstGtAJpQmBI0GHAUoMMnz4vToGGX5UaHH+0Or20ojYtVmT8HjUVQyuxmiPS/Hsc04cJwLHbYO
2rZoMl/XMzmA4PXUJVoOGR0g+cwQMHGtpjqDEiWu36hSkvy1oGugXjYFZL0K+nSEmYmBt4iZLZhu
QXX4DPdIghmnFt5PO3FyYrnSQYNeT63ap7lrQw+S7tXGZT2u/OeNb+I/+MmmmEEaO2u0mRR4cpdE
aB01YgYJvN1TuEYYrU4FknJba+M10iEIYJBmemkm4neYFIoIiqzye+6qNpQrFNIbIXbtu07TVOPi
oRx5VffaQvawlac4VSmjrh5jSSaKm8VsR5BWnIRLorj1ixqo7hWY0/ip2TEWPh0WQq1W4IdLuzLm
gxAY0qonw+YR+XYLfsiXkr3Nh7jt3RSuIV59R6mXFFfBoD+/PkJh+4DThq9E3s9q+cozChGouVfx
xLEWyhTtkt5NVJYyfCnDe9ElzTD91cYtowoa13QUt4GwrfiSKSsCscpu+7MhgV4j5P74v9Vm/frg
IpduaJR5GWYi2igT+yRQfsfW91c38Di80fF/xJaFnFswHTOPSnWUFPTjS862FCE/mQksa8Wcgnrc
XnXGjdRxoU+7lcrVi4ikMPZ9eHZT3eXt30y3oL1aJvj7pkn/CIyodLEt7lyjZAXi7VYeqlXVFbg5
u0vyw+PaxZOcxAFXDBpran6TdWYvusNd3zS1902icCH3qWypcS+9L0HPLjMojiCBYRVaex51FOUj
10+muqmipC5u/6r3AQLoE4ViPadtd/suTwLWQEipKMLZU8ggb9f4trnHq87Fozn7whFYdfjleN8/
rD2TV0HYWRKxh4d4+ywSzTHnhk4Am2hm6El/pxd2NXjN4XO+Qcv/3N5njcyv9wApEmvuOnLnAUuO
fnVQ7CLUAWW4uWEHW6qj28xRH/6gMtNh0GDMfyAOpBSyKMgZUu6D7rc6nAMM5dpMdY2y27wQqyR5
ZxQ1DbXVszDxzN6I5XgA1ynyyhS5aWbYGlLIpVRr2O2mlD+axVUmsGbNuK9VSXIG7isAfNOaYkiL
nCD7fVjJi0N4X63JeJlihbaaCOtYDuVwLCP5X4XQnziK3UlfPPRLGjTLweRo8ACfcdZOfnRAcjsn
ri4AU9lDIIXxyQ4W1Mw+oyPYf34YeP9oDVUd/cdEZ8S/wwmLa/bodAy432VKl/4YnB1AdDxpEmTG
tI74jnGr026gAHwD8zZKCD/hAMs3wUC8chwOFK0X9x05UwyPXVRB1RoS3tGOq/5PJpCSBAxQ+5iW
EvaAsQetsV3XCF2qY2aTY5FI1u5CFgFwopolKGMPwVdUp/QIUCscH8UMQLzx3YCl8k8CxkCBXHts
QDbPMPdAqbLUSqfqmPhgRdgCzp8XnKICRcqnmb590tmArmyrHNHPPsQ6GKQGO1SNSk3MPU0Ustex
rOOBGfq2VnBci9ztV4iFah7IS6ch+aUanxtOcdJeoMJviFFEkfwPz3zuybnkZm0B+ToIAz82lMNA
wiQro2ZV5aKF6kCnO4MpGn0g9azyw9PMmAswddKYoDHAHj30S/mSwBgAUkq/wSV2pChNv0TMrico
7vc8I6g3UVO8PxfYpqOq4qafCBghK93x+nP7ETDZGvJk7V6NB/Uwzp743s+2pysLopUEgW/4BkAY
S/zLbhwDhf2EFdQEWBt7RYmESbULRoewUBiAM+DuxGHz5AIWBFxsq3Bv6t87pPVehyHmm/PRN5ge
RC8W6VCZsu87k+/9jNtLhf2OeGtulj5H1kEWOyMBwqAobBWrtAoDmM0vlSYZZayubL2z4Gkg1g7G
Kl+oGr0UgcGEhfPFxyakg1b++RJh0KwHBc2aAxPsgjjCBxcFkCOwmV2i4EEtZHvASmkUvyJtX1jI
iLO3irHMk9au8WHNJPjO7SCTE/Uh0UjWt9yY33F2ZIgjQd6PXG9ew5fMWvRAlHJyWjAE3lWkcL16
Zl21XpCYm4Q3ZHPuBDXbnAWY8k7q+4fpMmE10L7T2679YIp5TScWuxY4SimbcR/HbyVPYCxSmKO8
jMieNGP+YjK1VBoPfZu0yTAyAOLJ5Qd4hJ0HTLuvHHJ8Fu3M4bBBsO3p2RFP9VxKAFCwbwHoaGy7
dwWbs0lol9nZDavaTeeCZnQsaz8u2I6RPOUsAHn0eAIT2KmDXcOUXDEDcfTbKS1eqXLNU/fr4NaU
2KNuomdssbif9q5Mc0Vvn/BhVeBdn5wsIRbLx7p0pS06V447oGxWlYCeSaXBwcHQfmYN2hW1hE0w
CA2NQvZAvquw4w71/W5lq7lEHf2wRQVriHtQEVnKRF9KhY0aigPooKSIztDOyL0qOYjC9pAhSXxb
81wrS+3QnhS4XHb6n4cwNJpbUobUGGaEAlyYKJXMPIbrwjpIGV85rAryRvZU2JwGG/cH7hoxeQbh
2lOviGtbIrZ0vwnTpuNd+BPlQgPqt+qnBYFlg4miokizXlEmFJkrbrf4pkGHa9Qy9bUbv0De6mAm
8b7K7ezQEiz5Z+YZJSrRPqjvEG9sk/DzJF9ySZQ/N1IknVbmJRzhS6Q1ZIQ8PmJ4BwUyHYiALUks
kRQcGXyALLyUXjewWY1d9M5mR/1A8ZrjAeMDM5kPmf2ixUhhGzaskLqtYafXNtlFcl2jfeNzZ++u
yAi/d56UTTMc+tCyevw3SkhSlMxv0rnDmVVAOd1tIkw8gX8xfyGn3QoeEcTXuuR3ZW0gC0wYicZM
2zz92qUMF5jpzZcqVT6RzzhYQ9VxUxR7x+Kn5jfBaEjcfFdiEutXzWeAE7AZpjuQXcIZDnwH1iQx
VugOEPamQd5EQbUkfJo7ddXL4pbzRTOiqzc6WYy28+yMIQBS0jYTuWemBky3sQsKM3gcRtJnLCQB
iTEl4ER8i4nkH/xHUUENX1wtRTMBc7xx/rIK7jSOvx0EjUPPJXA7ZHh366yR43ipk+WvXe3lnPZN
gW329pB/8CrWNdDpjQBh4H1UZ7JB9r8QC572Fz9McEuRJ6yVAf3fUtlrqx3Jc2QZF5yZyY0tHf1m
0d9ek16bde7HMwGp03nSeQl3DqPcltwpd2xrirKU1X3mjlwRyzLJWTXIKF2wMlOuISUq4EP+4zXv
ICM4wL/SLP9M6zEHsn8eK2LgIKozQ3eeHgpHlHK7QABdSC5tSBuiXI1RhVJsjstoM4MxSA+Kokll
WQe7q3beG7En/K9kvgLsJZIOiIuFgydNp6xvNU5OTNamvJ6pQqLOsrQKEFwEoqKQDBEnX0Tg3DQT
G9oLtad2VPI9N4rdlr9k4UIiwPUVo97cMzoVCnooGs4k7cvPIaBF3qJS0iMsrE6SOU6iLdbyb+/Q
NLdIugufPdyjbBrn2DYesZ9GDavIejpKAZuidwLsmDJbN/TxSGqCoB6vRUuLK+jxEiLu0YQHpuwt
QD8mpj7Klzu4tjeKEDalOSsWeJEeTza6/sL8vcALOKX7fXPeCpNoyoBMNyyncvZoU5KBfAP+RdvC
m4ZT3xOCalwdie7Dy03GjrD54CKKaGhFaIOljVbQV6Ww5Mn4Pl9Clo+IUmQysDI6B+stlOx1Jtat
gf4sMlFsmeJj+dqEzC4eQeTArCiYeDEecKm3NgMXSyIiZikodSBnErtYibRl8mN8A+BEgntkdCH+
WNYr5ktHwMXq/acDrDFslnzivy2UVTtouL0VewdWLgRhTW3dWAaNt5N6K058aRFLWttn5jBWngCK
RnTgmSxUvCDFX6qYBTpQPKHG+da/8DKrzfiYAYTuAv7rFAe2iVsf4nCU/ORtpZcPcBph2/HTN3j8
KCIVLAUSmFlHmUiqakJUiKu+J1WcX5EILf0C+dJ85pmOClu8onpm2ztMctJ1X4SGhbwk+e+cD1f6
LNGcBGPNscXJZnHxEFTso5YAGt8f+OpxCk5+d8K2SXs3nNYidbUCGj/PNBxAlDZ5yvTvDszfcW2t
v4bKk+bV+0uh+2JKrlqWJHpkr4o2sU2lbBUbj2Fxfi/BWAE3XUIHI05WoZZ6Vw6BVqnN2U9YJNKx
SmsZPDsS6MKAoGkQ4tJLZhZy0QUInAKCQpMVdW7cCAgFKPigZ26OoDT+rzygTyP+TiFbbWCZoMzi
BzuGacfGL2MYoe/TUCfDg/iSKbLF2CxrQedTHB8o5+h6FmrSQsEbyWjAYRJuATZnzZkxVOFhpe5H
uYBvIzu0ezRhxtrDwE3rQGAKNFkrWoD/keV0NBKXjLNfw+Cg4e9OH7Q7NFAFNzT21r1ACfAI+hdh
djVaXrW/ZipOFcqW6b9PbTLKX3JBLg8qrx2HUMV9SDww38yi4pHR79FGC+4mztpoip/QeeAeymFY
1Fk5wnka2xkxX+RhRVlf7cNPHsBah9ANvyG7YovGDjlTVbKL7X9z+px+cpJXASaR0j/mrhOsDWox
46x27omIJNAzDycRqkW4q6mIc1+HI3C6RD98ZvC4OWZlwgTWuiBmCDSsnaW6J2x4VC8AHJO1XSgW
V4aDInCpkvm0r8fhVc14xuu1TZmAv8EjiYVaWSdxHKPavrbTPc18OHF7bpooS9CkglYeOWVe8pBv
jsjQOLHc6kV7DdUC/+KgVm5qsi/eGD9a2eTMG8OLriYpqKb6xvyL4e5aADaLBvRgHxOTBf0++YK4
kvtXt7bRYp4KDbFcFiYq6lWXQbCR9n+RqrJ1dvoju8DGaG17kqM5RT5DIB+DQ76TGh7ZZw3haCvG
/wLjyfmkKTkLyyZONb7fuSsCD0Apu+5z+YhIdbhxPxVTwrooJKW3Hl2S3vgbtDkh4K5mIWr8msRG
3US87c3iGiJNd5wk6z04hTTQVvNLOPUX0ufkJJGLEZnidU11wGhSuEPb/ONPy3Mba5OVs5qC9sUy
1Z5zBZA0t+cqVRZ9fyO8erpsAwJ1qUyRD4tZ1V0y5TQrVdNeFRAqHPWuMCkLG0+Oi8kpcslLOyQ2
lMFbSZModBLQKlUUzQms79dyMDqMZu3R+uxrnxyRhL31ZGmvsaolnWsudsOrxfBelbEahsvQApGO
h9YfCL4BgNXjQP40VZlNcJub8dAchM/GDePfGMdIZ4rdnid0/rdKxY9lk5U4INYpG85VVQwOeqYK
HdCXTw5Rny3r/G14kV3rXBXMiEhqu6TC3GQW8qTGEnn/SWQDOTJa/NGsHwtxdADkrk+zM0J5DE2t
rqFLb/zdWxAa6G8tKheo+498grlVfAdXPe4Wu1T65zaGvw4zn7lZX0moZVviEuhF9BbhT1314FBS
UrLqLEpFOXn4pcrXVRZyPmb9tdKlssG0CHYZPWmFS1zoZapMog19ujcxMFOxWZFdg5WVcJ3qJRyW
n5ENLUEr4LqochcssyYGs57x8AdnJFkG2k1BcvQIzNWh07AjaMRLun0gB6al/LmlztEZDhhyNbI7
GpFE0UykS4zvXvuH9ANDqvxNjQVHQOEpwiIOkucrjc3mb+ZE/xB5fKM8PTAOdDbZqpY4tlfnm+WY
KVuUwIPkBU9InhFTbQvzOp9tHeHhgTtD+uPHbFhwVo9Yl4RRKiw9nwkuECus8Mbo26aqYfIv8kur
RcRl+zIbim88YNMXWbZUpRxick+/HzTfOYcU4VF3zTVe5XyBiMtFlIJO4qf9p9TPMFiwYhU2Zhg2
rg+grGtAxDm2utWkqAj8DNhtKQC83z3U4lTxumQonpfciveYTwubJdP6JNHyr6oIU9236FMcZf2f
yQ7Xhyq9aactK215PfIAlVJAY60sLhKb4k2XxEPcsvNuUJrIE56bntEFbaJwV0SBsDoIudMERFBF
B6TogAuM8pqOV3Onk3P8Bu/c0X2zED3e4S+oSGcxqv3TgrI6zEFRkvMJk+Emc1qld634QHw01b7r
ARaB1Hv4rxm9+CDexhbSRyudMm6Rui0UySF1FSyOMiSpU1aTGUPJIkMcuN2/m3quE9nGn+1g2e5H
5sgOzae2QzRdAYcusy/ZENpUDp2Qc5/QaCBvdZi2+n3yxUN3iUE9M3aAZNJputYwcJ1/mzvrES4a
1y3v6h7NjoG2IdSFmAHDHlZfHQ3BNkhNKa7qHHI52U1mC8Z5X0K0dF8yCdKgYKZc5ee3m07W5dql
oOKRdBQcTcEKrpMvJeA7W08QkX0D6g4XtFk7bjAluCuQZxRgLURWBqczG6AADfYAbVCzfAFTyI+8
QiP2XmOq1J1yh07v44jFhBpmU3xbXOM43AZ57Zh9Sc4d71amEtlrg1gWtkMbi8gu1uf0J129+2f8
yAk2Bvd9kkAB4IOKLdYCuhUUB5Uu+XmcqHvuG/XEmIPXNTdDUZb+YQ6xT1pQLiyi6WDugqSSZLWv
T6tbEPTACxi2ZE4G+Scvlf+5dJkx9hHoWQq1yz/b40iiGhQrGnn6KYom8g+STyuYB9HFave3yLLm
MZfmjwKbS9OY6XEykXgwCvbuqgEzMWIT3CJNVl5rvf/VX9mkIt38N6cTuuoS4bx5PVbnfarZvU1O
5BNc2VMzLw8wFl83lPvqlxJUrvUWMazyOEsWW3/1iCu+vg/0Ol+64pBGpeU9mehIaNp/Jo44lPFT
e0AcXP4lMQ1MtJMMzb6fmXr+DONDz1kurym2/JO2jqisFxIa480DIcbBcqV+Fs+nWx4zaxxKuNWK
I0CBmU40uSNc6C65TrP+oGMmqLInnIheRUno0Pny8ZqIvmgdXEar4/pmR7jYl6RzZu6rSvRzKAJW
WISgoCXU67Lh9YyC77Tran5JAtYHizOEZVTreMNjHbt8dF5zzySLHqzwGd6agjqjKoCPYYmorD2T
UGP0skb576nP+j7uccD8lVzInycwbKZh8Bh1RZHAD7GkvCboZRm3NvwNPQ4Wql1vDUaLOIN0FbIH
pDaGGpxNASeaVboo3Rp03PzZSvcnb0d0kzfIguTWKCDOc/OF2uY6DM4aFPJ29fExtyynzYdFC+67
SazTK938sqWao7jdkJPaTruf1NOg1GbWbSBAOhDOYxQtAmROZqI+5f5Rat80bi6dNO35iWXo3aax
n1bDhnm5KN/MP3h7PITi2+0rIkRvtKXKjTzxdEFjJ3a6VkE6ouwuptvvF562VNyr8tmA6UfFKBt9
in6jZjfDBgxRmHnTUUg5oEyE21drjXdFFFiiTjqUOtdBTIyPuvSd0cTuWr6axA0NW8MgrrZbQ/R3
XLR3PjBco91PUi9k8CDdJMPYtnJXWhTfVu0+g7A2eOX99yrErKRwbtlvDYxZlU0gcxEFDE4Rvm0H
AZUNP8zslz1dBHwln7/JrVoDQXeHI2rQ+LbFvcs9kZu0NWpqeQquj1uoQk0srzphiUDrzz9XtG5Y
W+3rcsBS4ZCJRsnHbie4gHftkIuUT1AHB+LoAzMW2GkEDm13dbLAxTftGK7Y4PXyzTANdwpJncBc
CDahy4NXZCPWxn8GOVsDPcy680urxdjM7NRzN87BsNR/BVYgjaqYJO+NsRKPgzUaVx+n8YwyzbmW
G/8K91sSFEkPr0hPOvocfRU0Uu0p6HwGscnUGHg9dgrFtaA6LM7BuDBOrOV3L+DI9AHCVYNcJ9vo
oCQ60QMHdQdAU/tT7vC+jq5FpbA5hYgR+M2fJET3ZjmcMSDSWpBT879fzPpFRYASA9+PDY0a43Zb
O7Aw3pliRn0ZHpTY0qc7HxTbUtsLmf/Qiv+JODLwda1UXZzBr39TfCX+ahcgyePs8fM69QHs4ekH
J8F75vWRPmyL5bqenEJo6a4NPLD8+yA9GqFYrm5Qvog7hOwB4l0hvHCq9kFA7gEOKld12egog2cV
xA6hfHUBr5AbUuJoyy4zYnhNNzBBYW7fz4T6oQmHfS2T1nWxGIap5BEZSt1OFgSFcR4zVCC1m8OC
/eXOB7L+4eeQidSGLxMBa3TBdI6eUytcx5ERARbJeMeqiCNU9hG2xytOqdSwGsofEbukpyGpbEdJ
pdjBKVaD3JtzYZeFWr6ie6BhUgA9xxkc91EfBz0YCBKrS+kvU1Pba2+clfVPz1+vuLVLoB8OxyyW
xdzknDwwm0edwbycy89pWp78Koxa/0bt6Ia2+42qtxMr/rGYDVmk/c8L+/GwAukxHYlYWyAveObO
fK1oToPZ41MdsadiiYKnemFMegCwQBit/t3lITbzuz8yweejViGCnUW/ePu483ce01Mz0dviXqjf
mMOOfstvsIOREHCYJbp5i9ifZtRcAd4hcdy8ssWQyz5+Lr2kMQmsxq9GkI6vFzOwEme1sqY5Bv+V
DGPn2tbsim5PRp4FQSNDA4XGjPEwP5Zijj6n3vNm3q/qSY6sw9AJQHbqbNkb4eE5h9SIkV/9LOG9
19lpDfOLaGzTUK+BORVU4x0s9/s5s4gi+OrrP1vhqsaRZ4yuJPh77p/ljNzIUeD6rcBVw0SfkDlT
MrAiskQiExIFKQ1ldbY1CePbghuyfpjK91qPWq8UB7crJpzxkSQ+w5YGNTj6hh+4qAdGKrlziVul
C/JaMvjdMvTqOpdSavd0LpjBK/y0b8wjJHpPx/xprFQFTSzECqdIBkOnNc8dR+GefCjhrwcQNsp1
/qyiG56HQWilM2E3poilofmibom9tgIv4tDbQ3EV7GGIRchCGK0f8+/8bAlyrEQNoLLUr9cCBWLY
A63R1LS+kExKOx0JUSM3uqMrsj4pkNWdtcRV3lvtR8MTyoHYzPSkgZS1ooAZ6x0UXzJ7abNiyCAR
wUflDckHBly/KsVDsdMz1I9qpw6esWea/M8ToKipp4TEC/sYsigEXxbTmJT1Pe6d61A0yHirGg13
7kfjgEMUVjP839900A+qCV2BMBlvvG+K8tuS2CUtCj6TbVhNVcEX0QBUt6zcJBIeTOOAWvvWD8yC
0UksoTgq64QSGfr715GO80q6h59kT9ACVmx2LnIQUKg1Om3BYYBPoqE2QFYbsRE0JAbfP9yUz1zW
5UCmI4vTRxzM5LkfDjTh2CM8Cjcy8FmNh1CAxOdsOPPWHkla+Khpk24Xw8Bh0csyEkKs9DxCBK6C
JVr0DElpI4yeZ2FWp9D1mePPuo1NLAEMnQs+iRRjiVjuOH2xwoYtRWI1/mZHDqwR1sAxRYA6C0DU
FjNj0csrQXWun4iOU7XKcQCSfIYyUaGYoETgbnFYxp43PzDGodNK/RyDEkXroX6pIS1e9jXHmB0q
ry2f3jgQCalYEDneGfH7j7RH8XXDWeEdWQIimELP6qBTAr9rcC+je0hJG+Xal6PrPb8i3e/ux9le
BR5BreiSzgs2F/8ViO4yCMgPptrRWzkq2TOrI6UdtHsQkZMP3MK/W+jOjx/C7XRbnJgQ5sahoRhF
vE5gyTbMWcMQEaOJCRIXpI2YhfGPDBam6boAdgvQ8mt3gGzdT0Vu2cJ8TtAl1xl6w+dtNvsnGpGq
MYqzdWip9Hez/S4DwyYx+05DTWU9s2bLk0DQHVe4j6sDJMcQlUalbOQrZ12yAInE+XWpCmi88CwD
CCTl3A9PYUnLWowZL1DSBoEeskurctgrSKrD9GelMWe2kmxgk/BAbk+U5QqlVHebTvo9JqEyvaxl
v8Q91jHM9I+59QMOXz4KP5AfCc8/qz8vUEaACTaq5ypDWiKqXyTqLLxkgZq4E17PjWfmtnTBl+J8
/Qdzy+5nHb/RK+iwUdOu3gbvxJRJp9Sjzf8O0HuxhCjcSFdkCNdjR4hVVSlrFVLueqjJKesRxKCY
BLYbUWdFtWxtzIV7s8kAOyJIGBQOGOVsD5jFVaRxyMDOGxYG7nkJIL20+YQwrb20PGsfCsWzfxsJ
Az8cAGKgXqulfqktScOblDimwzfGMdDPBZUKxf23nF+6zujtHQDhocd3NnYaFfTAg0jjInBPRqNH
0gf82tRYaDAl4fZgUDhNGsjvL20pVc/80fiVbxvR/YZDjAV89zOQNh4+8/vD6CoAHkjUlH7bf4Qk
Pp0HqjD/kRAIdrA/qm8JTf8SVdLlnvNhlBRjzNEEIAIA/4/78sr9XHzI/JK9fIbb64raMtpD59kS
tY7G1LKS8LTUui8+8+lNqswqIkzwbCDtvUNBPYg/KWxodiXGqH+8icbhSx+HtBXp8/yN5LEdwxy7
jF2C0Fzdoyc7CoEQ0ubbojrgFBWPesA38KE3tnzZicj4wzgEFWbhYsR/Ky/FMkjHzvSBx5MvcAq2
QzaZAY8Fb9lJxnx9GE3PawSwiAAbpoOhwSYo19DmNyiyZpOXsuOz5TJjRr57LvLsomluyTxaVCne
abUMt+grKgq+L03yasVGr9+rj3ERDhi71BhHGADF8qlWMCLjaUoJq6tB8G+fG9ss+NGbizdHOnVg
miwk6y7inY+fRddqvrmjz+NIoLHyaNNF9HAbveov+RrnZxI6bpAT+SFW5qJiBtu34xYfhQQqc+ut
B8OFrXUkZiume181qSDwlriiYvG2gHiTT9YdCfzmYxCPOk6MNDcCjm/mGH/UIAFN/D4eAmDLjOTV
b4+e2UUIiJPCOqsD7kXwwm9HlAAgY/tRi4sV6vKsYrCkweIiitlQNY3oI2ipjGKlDbwvct7cAYvk
gYbuR1wgMAs9lsT4pVdl4e009K872I6pa3sdmJp/C7fROqVmNLZhj6Oqsr5DHbvMtYTteJqolg2f
0ibLsgFNDleYhHgKSPxpjOic7nR9oV5bAlAstXqC51GuRydzm+UurC6z+VCZKpPWcvAvJY9X/yre
eqiRcPXMaMOqmhbO9Pp1Dr7CuO1yqj2Z0UBg6E64rxnEMlfPewnYMkqhkB0U9vfuFtZX8428gM2r
OTZ86X13rhz9zTRQG97NE08mnLq9jjOJLag8TZXNRMTESynVoEa2wa3hpJCSC61u3tq9H+2hqN1T
lZGJtjoGxyfbimzBXZ1y32V2sZQcfObsMWyeGlx0EXl+0Q0K/ddHsOg0MaNe6qUgaGlvsARTIZxM
nngTRmNxpSSoaFFnullJ8alU2zVRwyg9LTeBTcrDvHwMS7k5NandAdRUf9VA7tsYu3mRLaMnI2yY
i31isTm7wbqtFT/doURQaDNjjsOhu1flN6ZNyMCFr71JiDDNQvq6R6CxIHWtpPh0tutQoRarUdRv
q3u3bYVj0uUU8p8fFvjksH3nn685oOQP6Q1z3T78B8nO1s945kuJh4yjkkiaNz92A8KW3Z5ktho0
Hm0g/5nNCpgiMjrOna/PzOYUDE2BNuaE4lUNhUS5W/dG3A8z4l9IvTUYv7F6BYF6n5BIDVaANaKE
BM619ztOURu1VHdNOdR7XgqPAfs9Ts1+HHsdzF8ndoG1BzBfXttqaYka2kwOYZZAT7L/eNfiRcOh
De7QZ4ioQn8zqPI2iAQicElzPE0T1lRl+Q6diVEjPeTaiPT1pctT4SYA2Phc7YcrsGXf5IW3/nTe
KXc03cb8DFyBt4xRfTtR9TCvBkoXIpgNxWuYZQPnZtdtRB//JZaHv79hrA3AiKQreLx5ed2b6afg
XoeiDcRs44UDk6h/q0GvIyLQKP6D90IQ0BIBKgq1C+JOFEjB+yPgZbcuWrigixrJj9yuo2zZvlU+
sROkXNNv2L4UMmSxFPe6edj1GH6gVlBoIrp4vcadOcMG1aBSZ2ocAPW6P3dgNmdVOcGUIX9HTq2u
ZzMmdsSi/XppccGd/wtRJTvOGIlIkYdXMNz+4agerWvPEocF1spbF/zaRU070XpfItFaLG228O5M
j+GGRPEWFzjDOPGDdsnsKl9kKUxVMpqvHCn28ZJTmTxvWPNiu8znvKCL9kXBJ8PXegjz4MrSNYxR
zn1xbiD7+b2KLxHP0P48gH/RQhxEIMIRr7EXMudO3btCNH6xMzkMVbpODbexN5NuE/99AzRnJaqo
3ovx0rHy/WW16Kbi5Y/GFLk5XcATqdpExKmcW7oxphLr9YvTVJ/FLAWmMowOZqoA9P9ENYkGUwoR
aYPp7t+AaTN2wnb22RWGpe+PlUSGl5aBEUm/dl0UIZ+UwcQSjr3fM2LfdxcyzwN2vYwCHjYd14Q9
+dC41ZEEuy6wZGlcafe9z2a4xkdV158aHrGLJonqkJGCaoUzCbt9xLKjJLr29JFpY75sdNINZrtd
X4dBuDhw5C/ecXc4uA8oeiKTCbKHjgEmikgyUxSdfL8P4YMkTF19+Qqn3NMHMRNoG8tdmnJOkqBp
yeSMYKUnZzQ5OfALOwv55uVbC7tjL4/xmcbZRoWYqCzAVLWNkpcivK2bnX/y6Jnr7yVuuaHR02Na
xgXNBd1koUnMCKGIaNYZQPTBo2b8qO8iTS+OOYV9KPZGbvVD4kAVNHXX9klSU9J9MW4NITFHjmQ2
4ppDisPcrxQHB6ZOtgThz53iwH7t9jDVVWJYOEornMdvsdv6O663kph0m/xtEFmhCsZgPO+9a6jt
A31Vr7Aaa90zIFhiikXK/u6WwmZG0uRGegpvZTrrLWwLVxO1N4LgFpyS4P+3uBM2vL43h0H5KiWL
tQsa0Nfj/IWY5dbwOmzleOmrKrXvMYZqQCCku/HTv6Zi3FZcyf0PFgnHNFmfZ8QTA/By3Y0xtGoq
etuG4nHf4UkFFKQwlwz1c/2zb5qGKYZe0qUnFz0rLUzxKRIW4f7nu4YTL554+1osXne8e3wKc7ve
hEg2DfycvwkapYAxfrvdISj0XLiHJsjYHmG+2bL8OLPAFFZy4/6i1r+Rua9TuprRy0PEEce+apVO
aivdUUlNZ3OcLKZOzHASJHyXvX3cLxWnObWYreVcq76EmkG4Gkh1dbN4vuSJRyxviRfWSLOEx+ZB
OB15YeARc4/FH06gQIO+0z3mtCoi72J/IFEQrVbbG5niAOC/Ly1etLhTNwymtfGv08CSk/EGK0PK
2tBDiImr8RrWFAWryttXPzcnsNh0P63S4FEC1MKRKtqdZ9QgpUSzeLm6/j0G+MVSen+4eZdKpIMO
WAKkZaCWRI1tb8tQBq2plgg2otXB1d17WStnyOjymBUhDPt9D++8X8+fZOUdEKVw+c8gSw4mfYnp
tFYDuaVPT2pGuHxdc2hSOlQU+1zWo1aJGJ3JRxkNRWoPqB/Br1/0UoQ8XBnfdcnGnWVU7etblnfh
WFnPqa2zBYsdOGMZsXGYNfhbUTHmC5Ymld3OSh/KWksDJk8iTnZ0rZTU8ohM9K/gDsiN35hWDhqO
vCVaO6VlVVs/qarJSl3siIXyF21d6cyy+v+ppG2AyRRseKAr90jl4ciBoxvre0MG0rBbZHPtj/tz
G+Ff3gSwb5JV/XZhysz/KdsL4J/gi6pOWioR7yaC6/fn+h4jGfmKghh+a2DqVAmeHHlWWpvZwlPU
XkjhcK4VE2hOuU4giXl2mQXrcuLhi25nBtzjnQmFcWYukzYKDFqMDFqEDsc8X320VbVaijmfxWq6
aVgsqmNEGPDUpc658jUxMxtt9+sS0fSWyj35M/OEeeiw49LpRCKV633veTOtBrUHBrjQ/8zbvxsj
5u+Nwe69nabX3h9IoeBvUgx7Jm+vPRRc8Tt0jbVioycFWXwlbDVws12cpOAVBCbwu3EVfZi9Vg+i
KUz944W5cfZz/qN40qi3eSEjurR8/S0weXMtqKzLjcT/j6v1U1c/hM+lkaCStniWs1ZLkzkvO0R5
8umD2gM1vMmwOFSbomaUpv/zKHmRzTPBVJM3agw4vDg70lC6YJc1HSHL4NQVMEBi+GqPFxOSKEr3
/DqhY2j47FrpYbd6Olt7oMO14jvgUxM+ihKxBWhHI8SZmVSUUpSmXJuioWvCz6JkT5xFeUjcT1uj
zNPAygwvuM9hnwEIMzHqruqYEIkPUJB4FARu+vE22Z7bI4UF+sUbNZ1AWRXYTaTn4V1r5WNNmY6w
g8Vc7Y0nBRj4yAI/SE2i2Cls9l7chmvFJ3XGpPBWU9RA3uGcuSya+H7thap5C8ACJWMgruVzDpz3
PDeuG7OJL0M+hgwdNqmJ2qz3qoCm4q8Fry4An2ZjHp/plPGqv3nY56hVBDYxzcZOrFmfGVPujLt2
xShExWXjTNXghV5zh1eX2UPKTUo+8OzArTgXW+WDzLTY/8EKlqBOFQdJjLrt3B9FozIsoCZX2wE0
Y0Icoo8rxvEZB7qNLNFSEbziVKkFC5ZUAgwL1Yy363wtNyJO/hd5n4e/8PX1iUAmgI45zD8AflUJ
gIryy01i4ZeVmdG1797DrGRJ8L3bg2sZKzghgzZKc6E/+PHGtqrG+oWKrviWCen0dVRyakqOeivs
E8diw3TCk4CvHPZ1EC0OMy4DfhrtRuzp1TnDhKps0TbgTHI3Y8qZng2FdUTm7DKR1xsi1Datjxeb
dRdwufKyw2RTzgYJMlz8qkM1ET3eVROXgyXMX5d+uyQ14frBauXUxSCyMDnzX7MxT50gVP6y1ciE
mAzlHMXSUF81AYfQjZdA0t8T3zNBHF7Tmb8IVS/H1G20I34MBeL/IGCYonpbhQ7/3G3VKNErM6v9
b5INHoZbiHcg6kh2Bosf2bXQBLV75C0W9CmDuGwvnMLt3fJfKuxR6UyeNU15yRXpl6tCTx5+GXZN
AqNQ3EjcEEA2qx/zVVxJv5/Dm0eKLj1K6Q4dcCLy6hkE5Wp+Y9Hch1hZg0Dp3E7SFo6SYWxiOYOX
LOeIoovo3IlQ3mkfUDppDnXmttNsAtWRLyo1JlTQSIoK8bu5cLxmAHdltNcTBUqCNuv9X8s8tk27
7nJlaFV4sSl7lbG+VP6l8A9OJcOMy0etwdSMaVRVAhYZTe04qjT27QGvi56Cs4nwWxlHlifere78
AWchFz4x3f5Sco13aQLbI4XBZRKh2PGstNw7eVnvHLfGBd3kk9vK8RQd6K3n1nkM0axQfAGhlaYS
2gHMxtYZeD5WjPmj6efIF+/K5nMktm3CgdeasVChxRZmO7ExHOlVRXdF0Kw9h7/1wJd4m+I4aJ+F
QxoIED/POpNUzeIehJqd85c2CLIeuL1Kiae944nu1WwcIOy4/q8P9ckHmUpyKWrNBH4RJrwMwpA8
f2oxHhKmefnYEfXAx8U+y/U/MM6OudHs81NoTeEQuMHCC9gj3YyDjTdJV5tqbI6Udwock20QvwO3
Ga9Kv1p0a6bCdYr8pX8xygm36bn3HxSUr688OyZAMMTyM4O7Of33AH/GnIYjn+ftweJtr879CfmI
xgpnOYFyQLz4xYyzLv5QC9xCwx5c5C06rSOo+iN/7Gv2jerXpzCsT3qQOlPrTNDEr63ko21ALxkm
raW+d0vGrp1GN8bESKlEwXwHOt1jJCIaM3IPWM9luh/xCR4wvoCFpgmWtHKNJUHbaHG82hl7bkEq
r3f8qfLkbDAa92vIAnBmVAl0fRk8E/LxlCVTphiu3nC7z1AxfLXL7WDs0jKcwLz2Ib40jwus5H9q
kedH3s1/vdUHuS1sJyf1SP+B60nkdroDpKU3Ux4CkBfjG5erhiJ+YRjN7eVhsaYB16rQk9ho591C
FV+vuFfqrfllmjxamFY9VgUc3rIbwStbyzS4F3bAZ1yTZ+4kzGrE56O1SJdKxvfGRydoymHtX1F7
5nEMFABlcscqzT+zfcUDKTc9w9hVXCCIrEcQZ3msC3QDX6myc0MWv5lBPka7MKhR5N4Aif1vtsyM
aCsWa6CE7tGekHy71eMK4TtVB/ZjNTos+MVVyqDlaG5UHcjPrTCZAts/cUafzTZKzNSWueS2q8jv
FQts4mCbKh3UR83y4NVd4HXyXd7z/+IFAXtxpg7QvuOpTkFVp/5GkeHVIeBZeWMRbGj92DwTtztH
ENlePR2vu/bIr6HEUSg0TLidHN6UXu4+VbZwps9Bkd88QyoqiodvjitLaSznqxM1aiT5eZ/Lp9Ig
Pwwd5qiVfP5W/YmuAoUIPB9DeMhmQ4E2OBLGjPtziKhF9ZZSx30rOF92OPC0MI6reFs7XINGWso+
SwuP8OjjpUQckJY4WzlCYms75Yhdx9xO6XJiXQKXCNXk7uRElvAyWxfVXzRFmegO1PJVFG4DIe1r
wPbMRHlN8/i0BMa6O1+TXWlSdW693OUVDlYdgOTWhb1J5kIdhzCn3sX4tjg2ZBupGXEdAlhLnF4v
ROMIOIY0OSmfRMI0k/oS1kWRYFZ7Hj1QugH+OugLmxDfWLp5KdewtMzrQmMJvpN3j5CApdZP1+nJ
Ico3wD30hjWD4Ur2xFm46S6FP3F4akQMh8GJgb0OozJj5SAnycZpoJhHhpjbSf34i6ZMBmP5qPJn
RnOqzYDCDgHeYenCqIRFHIY9TymGVoPEAHgchmUWegnmUUzSruWPLdcuamuUqRZ4GWMYUSgQ0+8f
d+r8UubhnDV4pW2o0DqGHFkf3XKoAiUXrXhqyKRBXmPtXSgdrLwPT8MU8H2Po5jXg/sbgcNx03PL
cN+b5YE8kg27bIWHYeN7VoYbC7vI31ynuXo4L0U0DclmCOhHWJvHSN2eV2IRXv9yQtTFUeiMrVE4
rsMvKTVg2ZFp0CecDsGNePJR1Bx+7nLE2boacO1Md110Fq0E5WiPORWNeKVOLSeTimsTsx5UC72L
xC2UZ13XYyFC0OtHgDvnu3ktIz/dV9bTjETHVm68fdYVA1o2Kt77BSvQnrvgS0zQx38VfVYoH7nV
x8zvXRpGv6kqFkm7/PF5Fev87hs9czaYL9dXBWZ2P8+Znu3Yn4lj9IlwQpjXEIDLV9eJqGkSdXgm
eNsT8fT50qBGU1kIIkDUNmT5ZR0RRGryeSdEmx5OWdn57YSt+kNjWasIJFTz1UutuwrytYQD8GNI
hceAFLoiFCOsJgVT/7lv5kwAERWs2QiVUlNUdv5lIlZfJgrtGN3LRULK07Goo1oM1ixIXvoFLZF8
z5PWkl8X0BjjRXUDzCtn+VfXimln192DqgU46QB1dM9WWEdFnxXmW8OROD93rV1ID/NF2Kq5ll2w
wX+VpusKTa0a7f44Ljl7kGTpaV4Gx+8yvfTHThnQ7P1g5eTJVD+qt/dat4FJ0FoEuPTeWYHy9SUJ
P/nWlp/oRL9E1Riom57WMk5wcfzUIM8RhuUgCVeIUeUTuDei0p/1by0iuFw36+Ed8/lH4vRgI0aX
kzO25gWsfyaBQ2jKS3LGVfvqMgQHvPDAazFazuivfbw0WQNg11ugA/OGQ83bZruB+8cq/MVU2qJY
DHXP7QfBjppFFfkQ7H3gxUEkHj5pLW2QgMsQw10O5xcfOfIJjU8ecKb8I8LvW3N6vq6k9WUqfhea
amkq0VnecMafWowwwuvs+rvfioyTSr84Tyz/oYpY7Vf6eXoQFZA/UZmYKHsFXPAHupByuBkQPsLk
TLSbQwcuYHz1Ar3XLnNdwgjeffX/IUULinXw1hnFW/m+Mj468bzx0vBdP+jhwWZpxf8Q/nbgF0h4
y7T4LDjIZ4m54lTqf0W0NXApbAcLsh5+2/UOafKyVKsFxwjqmbTkPEj2TQcKkm09yi5FgXiMAZ81
l88FbOGkf0VzGjSbpOo4Yfi6WSHLNgXNvGQcVy/BsYVjQFX7zaxuVLHGBmk+h6zhySZPYeVQBbqj
dOvlvhvr0JjjZayz+QNR5pd4NBZQWRIOtdFEHRjtNLGJD9Cg8whWZZ8y8s1Q+Xu/muHOkl90jlLB
VRsSF+M9C1mJuOmeSt+xMUxNJvUMFmUOZcPu6wui+OTafhgvQbF4Un0ETSrFFLtMMKNiUI+KW1sC
OhLOeN/8xZnZ+2wag04R/Ldy2+lEgfEoJyFsXhlymlnIoFNqOSzGjSLUDR9YEqC3jGgqHMiXDc8D
CAVvtrMAWCOpzNT5bZuId8v3P5Bgp8zkmNuJki9RnrS2Xuk9B/NeIIfas8M0LRMQl5ycZShCCn1c
W3xJTNrPdug36u8BKaNIiFESHrX58FsAk1/Ls+RoFCjTHcaa4pg5B7/NBd1caS46iMd5std1zuJf
oK+FhIUWUL7XZq4ojxN5hdtt1FQ5/WWVdAo5ZMkhdeajlD+G9NgujClMT7XeTR2acBFCgji2Hxdw
/BrWPZR9wPJqSbQtW0vMnfVjpir82+E9tt4/yxybVlr0zHWMA00cWbP2dW+9f6Gp+UO/XQTpGp9I
piAJTOEea7Vf2QOey0quHLWlee1dWJgJoxds9HV3dqLF0BWbQ1nPg5Z5Wr54jXRj0uhR7aMpJAZO
LNYRATZwfmq3+FLmWr0dezAzLBB4Kfj5a7F2o19EL3AeFknxNCSoMumYEXzzB0i7DiOymkiPGPpY
xvIyqERA7PzpBUCuWP1mFHL91qI9vlgjL1jM8v5tkFrV7nIoiNqmC+fzBl2WCYqdUCnIUvn7B4t2
rqC11W+smD+HTEas9hWVQSiTkd8yoXSjtTdPXr8gzFrKXjEYMH6YQqda20JzL9zlG0ygUOIp22/s
0s6zphHBfCXTyJa0noRQ3Boab0ss95SAuxt8jaqug/MsFBRwB35qK/DXSxlzGMAJUeaHn+GT1M/Y
gq03A1M5FJjBP8sZ1XlJvPglBsW4IIfLr1HhUVsvYBMRx8WCvX0KAKM30uKmWMQfXjM57ZdhBnyr
Sz7BmRAElIY/1sb+yqwccGCC/Udtzj6qtDimHHxB9Zb960UjerH4dpChWB6l8nGx5dt5N9ojAj65
GH17OLfdH6oH4ZvZaa9ZL8aUPpCR0aJVjVSHzDKGn1Z6faJs3OkMnhO54MS3uCDcfgb5MUtcLcIp
maiF1KjafRSunwAWV4WWTABsnBaazPlWsM9Sl82qOQ9fk/JxzQKLqZRdjLsjJq165fpChzNNC2rg
mGgPsyd7wvsumQkbKV8se1IVPy6tvk/Axf77XsGctv3Rhj4qUznxoAyPg0/y8DBgL0Q8/YpubN1w
K3nGGxNZByxP6a1QSLp1PSTe7DIbTaJMcN4gfLsvHfBBW5LpY9bkH1TpZbkALxDbN/j916N9kbgh
bnUeyPhcrPO98VO+KnPAIbVay4nCQZLBa7TcXgzRZf5wLp/wIXkY7B5xCx4iFwXxDV9crphgsMW3
EvW5hKstKWcwWWDi1qk02OsDyDGoORQyQsf5jPumzqiPXX2znUPdjoI6eGZK6S+h8BBawUnZPmp+
XxPmn+xH/+nbxIqCSVW7AR+JoMNJff2S02eVWdpK7B5YYRD8P52kFA2IqnTDnUZYO7Pskd+5cY/W
Ig67U5PUrfFA8OsNfRlp1EVXzQlmWWQgA7gUdqEY5PtXl5M5bQluQ82JRh1+bSWDhrBoiM7h56BP
/CR/HHoGE5AtbC1gd0wBbhp1TkVb7sfkSNeRSf5+MAG4TCLRWse1aXGxrKE0zDdfayBwdFjOWaAq
zYFifSrl850qA3mxLR5n33XLKbZubeuKzUtJXu7/01oeSEcGiQA4lUwcKCye96md1Wrd8Iif4WC3
ZTMCszbOpIO+T55sTdlxyhi03m5AOFELbw/RFv6nMpMl2PhWmN/5+xjtaoP5lx+zkhqHyRglRQkx
2Y4ayL05EGBNDYAUs2WaZxWb79NrCReWpngd2+e/eGi6jMnOK4o4Noph69K4bq/FftF1A3sC3MDV
UhJNviAVCtdf5HHTRKEVYdgmxDLf46Q7SK2f6jMrkBJTPqFMPrHX9n45WEarzSqeNFpZ4KHmBHBj
sWUwHU2ME7RWNigrk1iOCjBPWuOCuHqSQCMilPw67Mh3zbWdOR7gCl781R2dOKflb26i4QTSEaVl
577C7ajo0KZkUzGKG0dx0Ykw//9UekXQuYYT5mnsm0WkItEZUff1iPIcDHYPiX2D+hR8btt9+OB/
K7I5XijCDMWjRuCrptMlUb7z2S/n0boy0ck5JxXVB7nq6xx7sY5ltu5mV+KuP3Zbpkus2Bm/LxIR
HxrcPu/SvG6E8xKf5Aqw0cKO7BnaF1rDQ0M9wHIuc8MBI9O/e2E4l+jvsoOUJS+3k6GgNwjd6JkY
Fx08OsmdiWsRQYT2UgEfeRd2zzOkdG7nfQqGU++Ih40DAB9jjEyCduT24TUB6OBbErX6b+kgcAyc
0rQ5s8rb6g1XHUhMhSx7VfwixA9DvNArEvgnytxPVwFrNEXsG5Se08P3Iboo+1uwIBFotWuRI7T6
9pgIs6uXTqKUNoRSeRSXgYB0Ghj0JC4esP1fMkFGMB7mko1gmRd67w79/gQXGzvQszGGcL8oYmQT
bKXFqx8TylZMvGFDO0uBFn4WAcwjM6Dj5+nFl8J2BqrM9xj3bst0bkWaVeavGg0g1CPOjwY2bQbi
pNnasD9xSGZw9IQzzJMiIPNx+GyGnYC73ExRk3BnXjGBxaRghjTXe8CJrNY0g+yJd0Lzb7JE+CTK
R+fP89vW2eDsHE6i29+PGL2I65cxzv7dga56aB1hc7aoLPumfPX2jbHitb05NGeWFwQaxw64UYtk
AfJ5tr96mSAGBGsVULJK/NBGp+EUJmZvmqKxEAvVdHdL1p/icwRTM4kFjD9te98lO7TJ9VQtI1Zp
CTltJGqC4XCgLYPvp8S7919Xbktl1f1ZyNa1aBWEZpeNmth8fOUz+ws1j8e841gTVqTqdFPNaCDV
KWpaw62VCNCprIpII1TUro0DYlnSydc8EYZJLUPvyhdf/2q6JJdZWACKuRO2KC6GVpBGqyyFOWe8
fH7GmlJ67owHyZGkO1rBRvYfWuCayIBFujBeD5V4WLXE6lpDKmi0xDmBRg5b0EsAh3H8e3GuiFZe
NeNnCur02aRTkEv45ySu+0bsW+9j+XcyST/COZ2K9QzJSLE333RVhLPydSP4fBga51F2M4Hhx0gY
k65m53x+SmSPGeGDZjJcjHwKlZ9x2ba24cFJ6eTjm3Ajt8oKmEK5RQ/P4pp+yWCcR0gVkU97kqu3
xBrCm1yrjNDkzbqfir1vEc/eBUnY41MMKEQVxyGiu2xAAZcNqriIdJa17E+ef0Ls82SSE6IxZ/MR
XbuM1HCRjL5SXnPqVwhc9jz8WrQg1xOwWsN2dYP1OQqrvLYNoJG7yd8y0YRLa29TfZH2LNVFQM/f
CnuM3+HvuKKvNT1kIuwCsRH79wOPQJw9KFQ+qPDbKxolWL0YMAPgjnrYoxGiSjy5Aa2Z/qGrXJSv
U7mWIYF7fthyx0LVnKQOhSvZyvjYVfXBethWoaYuJYVHeWgOzfb0ugi5FIAgexmvxj5Vi0Nhh/xR
CujZknF2QbB0rdwaCrNtd25Kh7HISLlVLhDvPzT6AlR8V5q1Tf0SFOeTt4LQctYF/FPlkFACzXah
ttDFJfbVRnsw87qGOopyJ8ozyX0NU2BMbQ9y0Sb9EEsxeT5vEpIvWrD1yBGmjDLKn4sDQq7pG9vq
M6wihJVRwe8Em//QHgCq5zuzQ6kxB6aaFpqh3pYmf5FVAmsUfpJS8mL0AzjvIKO9BwdN7tjcUiUZ
CZHn+y/lw0X0vNQDpld+cKN1K7eL6eMKkjvuPFc/WD1eribK6djSgXEk/13Eo45GmGqAjQFK0c9g
eMMUK5UgKTgA2LwVldx+2tL261oc4SljCAWLP/xsrutlyrQVYllHIuPTi6KRVPdwfh7J9HR8uZrz
eZ2CxW7pSTaSicDEDFOPRIYYxihQ73tyd+iKmkbmpmV+WUuvHGnF1L7LJG4x+PiJdJPLx3dKlQL5
ADBco7yPhMC0euNsBWVrw71hK6ay2UGwJ0Th/twhHnyVd06b7BisnsGulk65AEIbsKmZTVNUr0XH
asJoU1VaezfePMvvBQL6ttyD/dhEJYkEFifM62I+Ob5IB7YPAVRU4tttMs95YrUCj+Bknn+H6PYG
772w/bzzTSKFDyLl/ojfpb32Hn6RzdvN1HId9FtiKJ9RpOM7mIaIenu2RxOqN4YrtUnjf0lOpwFN
qq5v1WJ+CdpH3hISRL/8qY0NmQA5OROM9IWDUX2iXvw+dSMLw4MJaHI31GyyjcnulaKU8xCSysTU
tvmhQGkcVLOqqeDEgpNbQEqtDedBIQSZIumiIsQ4u3wPEBvLlSHHkgxRwYAfaWEcYxmvTi5pnClU
bjwNe0vXzs9rI2zXpuEEh/qoELEylKlQWC/imgshVHWiA4n3dg8xyow8bbA+k9qSyhqZKIvqf1JD
KaA6eGWjvgBADc6I6YXU+cJFWq2Wf9i2oE2J/3VSWBsYn2G6migPqgmNR2q36CjJZ4gHF5EWS1ep
1go+J5ve0JZPRnsZ6W/+Q1Qbo10RcRHo6iRbGpsm5yjgI4hQU+3hwKAOUuvw8Wxf+E9mVlEoI9yp
OzaJqwyD/1ATGVDSaOEwcSer/gkqO9TBrN0JzP5I+A1lcvzzUdtf51S8oNq8ApQ/lBGAcp0diOQ/
a61ab0t1aBmu11ctKuk6gsPiqUPu6WchztQgSobiMM8VvxhrJX/Zyfdkv7SjBtvXJS69fqyrSubr
tgn4kzgkTr8GEP+4EwIvHOX6iYLk+VqGS2uUa5iSMbZvjVusIdjGWbD8/ncrjOeYpyeBlOHYGZud
xzK1c6TME9Ay3Sg1K7upUhM0oKiS2RfeS4dGRQ1O4+iM72xbvvt1+shzPTXAxJYjNMkqpzsCrmuz
I9QTS0eZvPlyslvLF10nBhRilxg6liQ1CYhYUtiD5jWfpKnhLXauDDH3d+xXyG2r3tCvBoHmqDaz
k434Ud944OltrHIDw+P9Ix1LMPYBkTAZ/773tPm9f+i7Uj3c1bgNoNSwY+muP4MECTWSXHLbBDuq
bXU5g+MlGcFpe44Vu7iFpJtyoPr/l5eTkkd2+mUL+SJc8WoRM/SDXgg3jFHLawO1jRhx5yKJQ7qK
ftjihZSHG6bFFHWcwxZLEpdNmgFqfnvofyCmzCBTUgzUXoaZilocJsavqz27SDcapnTsDbKEpOP6
dvL7tyTYO13tkwGkdR4H/kzo/0zQKSXTmYqcUwQDR40XRaNGYA7qAOu4z7qquAhVEEbhT0NoWJXH
4py/EnlLt2YKNb8HxhZzvGoWtCuKBw47+OQH2P/z/XsCLnEsaThUeoAeWTi1B6vJUkkCREFA6q1D
Y6zLHs/ldrlulg4rhMhy0b5lcwYXLh7pKgfbGWPqpMI/L5zfJhN5cIWmgbNZ6wN+PJR82+GJ8Zpo
FA8aQpMaHfW9VDeasM0BpaaCupiVVaoqIbiubvoIE2pWUmmNCGXxbeADPwq7uI+z2CQDKQbNvmd5
nTop7FnkIWmmhutgAdIGyhso072H905L5/3AbhS6zDUyQK2uD5v0IBLXgl6LgtxLcd5NSsDSbn8A
hnJpELdJQymZim9+k/ta4k0G4GHXNJ4nVyhBjFS8ulCLEP8mnj2kBvmknyYXvfiL8aBFnDX54dpF
17htaqr9WMeuPLgEEk5lrltPU7HcIJwHTcYZSvWB9JXS5SzzjLjRfQKDxLryVV8NJCwX773IYUyn
a4INd28RorKEHdBOvQLkC9gFvljvGa4Xlea2lDHGqOmfENeljVOrvprAh2LcQmBqbtNM5N5NLV0f
05l+mTSCOgTvvUKjq2HPXhaqSnx8YbrolHAg0YY204jFy/sdDF9twZeMIzspwW+BpSAbrROHjsgM
Ba9tJ4A18QBSTNRX2AicOJVsFecy2kDLzpuwHT1VFd8Yak45ymuviNuyF6JyU0GJrxwSH8Iuam6g
cqhi8F+zp97mj9l4aWUhOoAMN66ETsTIHziL0htwWQdJsGG+sJdYgEuoEozwiMfyBZyBbI1i4336
moCaBmmRZhGS96N24dePYpqewobDK+r3wL3pGiRReEF2cz3M0R10Owaxlf8ZZROwxjx9VsKRlYdF
DLqF5A/BrI8rFrTIiuAjUx23JxA7aJkI8dlzJAGKVMgY7D/VK6rnv6w/q2XmUZqO8SVHxvpFL1Av
+0En/phR9R2DYXaZ+WIOG6v+BJCU5sV0zxJbTvCz+N4IxDueaBtiQbTTHQ1ZqBgIYyNcG1d4FRoQ
VYSyr3Azhj0vSNSUu4s0ji3U/OOb4rpoI4dp7qDvnprTAwIY0PEt3Wv/JQmeVppNZRlf6Evptc2j
OPaacYJnoj6X5q4Y9xqWyDuzUeJSqgFpqPRkZBuiW+IX9jtjbVKvwhg0/nsAN9aKSpaz46R81idv
chpg3PhBUgGARXRyMQOHjZN22iiWQcL6oRGI1nWMmu3xvEcVMpf3iz1aWdpPwsOTHPC7DQwZyBNo
mB866265j2h4nrcNm1n9fdy8lkYiq65MThMMBEzWkm018KfgwxTV6kn6UTgn44Bdh/NF1bi4ySqa
E75xcrpvuRUPGB8qqytPSS/KU31Yv4zVuSc2MWcsVbIOcps6O0+87TBohUciF7b3uNfSNdpCTi7c
FGDbahhsdtDUdV86tmrcWMUZKfTauv6LuBu5duzI1NUfHAdNFVS89032bIA0gioeSD22Y2HG7idN
UsJO7Bmbxa4gFo77PHsyGBglX6RYbLpvysOfsaSk28oQ3gmrs2/uw2iORER6WAxzuUt1kyjYaEbm
Kked1beNCVxtIbqwQWO2LMTavrHIlnidkG85p92vyJsc93t3g0nwy01fniYgFbFdgNC0whKa4xFH
nzBXv81iquOFb4RA9WA+vL0oOCz+RW5uikP/PXvI6AukpbRRD+qoH++lyfkaEPwvgdKeP6G/ycbY
r+lnl15pgox5O/g/zEQnmeCcmI0eXj/pREQX0OCUZzRNp/sz382GX29HRRxIOAZ4WXP2k3jbS6jw
ecTtXdgMJpaZWwaeGNcdzcIRwEQF+bZLW+pd8Qh98HEpcvrdtzsOmc8dogEgmYDfLhWKpINmq799
bx+uTmZOkXoye8jOWMTGh0DRuGNpcjMk2bBLaWLPvhe4OHEZRmbUHtrodo11UWdrwqJtYcXUwtpk
TsNallCFv20bychOy3xzuLG2DUvkMFos1uxgEvFQMAZKW1FiKFm4tRPtJIdZjpfTGXvvXQf2mQci
wwrOwS/7g0py0CjBdG6BbkjfdIw4bpHYt2bQ82LoO2rEpIz/SEEAfM0rv76bj4HGLVJhBVE9bH4S
uskwl9bjEswJMrSjkeZnRDUEArpp5fzul6lHkYToZaEK/p9VMPc7qsLVQ5k3+kXu6zP4g1HswtKr
F0+Us3SP0nwHPFGTiDf3NrNAj0Bu+VUQ8sKxr9+E/2l9sctUYoCpdVHVBrT4mwwN4bfRrO3Tp7Yk
+NomtoJqjaQXV0M+5GoY4IcHsaGEadNajW5CI5sbLQcCQ+dAxynV990232JrACDshPCxtOdrK3mm
JE0ztQ383kppk2U8itUQ88GX8GqIA3dak1JAzN7F9/mhYTZM7wnNf/upKqwB4Yny6p9pSWdoQvck
SAXCykFlPc9ev3jt7QRhW8SDOcraakYw4V+44dU5/KzcBrNDr5kaT5TRdmMhj7sNZbBnKnsUGte/
Oy6bOtkzcsUQAaiWATh8yqYNOV9I02fFFLTVPVXRn7/gLSWu/NFKZBVm4vPlHnoV+gBdp2lIHS1e
GY1JfBIod4TdNsZizoeUjE5Bo56/4A2ngB8B97owK5yUd3EIPoKXLO95L7NeJinAx1t+czQdvDKF
iLjObIVPwBgRxczALDDZDIAAPUkeIYzLYxuKHHsPXnxbpAFGRYvPNhrFLzSNGqcVg9jMk2AiS24L
7U3AR1tp0uG86Hkui2DhiIDnLJdft1uBJixh9I+ChUehuXqpCO+hHY6UE+a1S23ib49NfLp50wnq
B6yc6FafKHepydkAFaPdfGC37LuPRsIeFULEZy9tMUp2sT4R5iwheaJRXPdp1xe9MZnT1UE2LMvT
pHyix3pYvodCMo32YuLMt9PeibYlzlsqUsJYjPd4ErW52VwtxasWGRsFpfQn3SL0eJIWvPjNXGir
5fweo6MywCg/ggz279cpK2Eh6rLsQ0omRUIESxPF9mg/orXPHT17zZjLeDEfrl8YTT0dSGadTCpU
wPVGo65Xx4Gqr4lj1JO+Khkn/mJSK6c/2qyJRyRsao4B2c8H5VUARK/9xLzmYhYctWU0F/IeWQxU
D0QNliNQSU9whQ7Z5NXErC2ImyFznTADRj1IV+BRoSu3qQehDMqxp1yfm2Z5iZmMb2AdumM09RLh
AYS4g190ApiZBgEeJjoYy643XF8e1hiWPIu3mNzRhdUWmUIUlogC6bMwBsIbVeLJ8rk5RJiEerX5
PWkIN9bcf3zBbwpzE0dxHhjbFjVhI4UrX8GcKbyfxVqfABilf47uNG6qa6XgbInNJ63pGl13v0s+
Xf3LHr6pMizR+bdppbN1MSoXzrhtIUvoMN0ZTiqukSAhI/axgiaphO5a2Tqs7SCY0LSODySsixuq
WMS/QcuvlbAF6+Fx7wiIpF5GCGT3RmtDQ2gzOfYwwOHdD/ANP4Iyyuv00iS1VriClyFBa37sxjZz
yu6F3bFS32XhlbUQx1/iyNVOVao1hD3wPGOriV3PHgA88OirU+KkLAMNRKd6f/wgzVeyguKSZx0i
vU23zk4iVbVz2Koi7IKv/IHXuOfrcnllMF0ei0qMXi/s165dD3UgEhk0feOuLjtENk9msEJOzdWF
rk7eqg5v5BSYcpmh0hu3ywL8PJTuz6eGkCfqEEzKWXbL4CrxuE2urvCk+EoMjjZQkDbO+5iYfeze
ptDQPcRC8waWboFQhq85Y2cdIu2M9YiHdYCSk+ulpsTYlO3TH7Z5IbjmhvNIJQT2eMvIbynl6bHV
xXOuOc5CUA4m8C+FVWnV4KvK7gR2vanuOycrFv59y2QtzbxUvfbDtbJCltiklhDeZMTJeE2jxP4O
ibLb11uXmqookfD0wH6m/Bztz8OfR8DeyNlfTYquu8/o1unX/UUBR5j+UKPmOS4+z/LlfGLPKVDF
JLGvswJANv4a0cTjra9bQL0lsPftG5s5VbOh0a1LEJnjQzuXil5g605SrG37SprtLFiUxMk5ypsY
Sd4X3A6yuP4uwc8R6GP7bQZ6RV0IDDbVqeCuJChJMWVCYXiEpxIDoD5e8F1jHmDYpYRgiKiShWK5
llXcQ+NKAuRO7ALlhtlq2ckf4YXZeWPzmGr+qIKyFQ5EGgtXZ1k8YfUBSrXgzKo34RRFxwHFMj5Z
o67bs59gc6PERCE66fLWEmLn0yZ2KNQWUWdYCvo6fFgS07AujJc57UxM6bcxrGPoEsOyO85hcE4n
fV6JpnXWceP52xtpIotmz6hpRaKwoWZgaWuzaEVe4UGGvCERw4S1fWJavomp9bi+Dj5ku636OoV3
hsNkHLMNDhqQ5vBwHBCIX5g+fNGGmYjYg7eu+KZfMYz7uihnNRAouzIxr3r/Ab2TsfmNihOG3vWP
JCBO+KQYdLme8l+hmFqVajwNRaJvyJNF5jmZNvd5jBVHvS4iLGo6tSQpkgp87H2Qa54oVoHn5o8J
LclID51clDG9rundg97wacFfEsgn7i9vJPpLX3qHYZm1XZs3JBZTgTENBOyp312kWOLt/PZYQOCb
/xUla9CyaE3E8ytoPNnllMAA/GiiHBKIrDE51/GSdGfAAux2Zii04zQBXWFqXX9x9V3/u0A0ZYhN
CDnkGxtC4U+DaJRbfb+hE5uzITOh6CabyG1fdhaqcintdRQO7VdVRxwtgSbFWeBstEPtHf0wSnDS
XRGYK4cosNLscT1QR4arOnh9lEh4Wj7dpMKYrcdfBS9mJqN9IUWFdW1X7ZZHpmPnPP+EZFIj20yb
jDbckW0Q2J4mCfc1Ko1jpMYdJ9u0GnxDXkm3aPogHPmfnndLdbeOUkBpcEkiIgqQUmy+wEG3Apzd
yXCeSFgZkXBu3H53bomU4cn69S1xTItY6YanNUSxuTr1+GJKDAJbyDPsuVmiA//Bumk5OVizwXtk
0uOc6XKYY35lHdrNn8nIEdIO6ssNyQrDV3+hEzm9Opl1VfaJxgCM1aNuIxOQZ5fGBdbdeEoXPPGY
w2C3BY9YQY7vyFpQ4FS0yiRRmOH9vREKjwIebOTaDdlmjw9PFdlCsOpRo0tAPv6Q8VfyD3lW2WI8
al0UG1rHYivp3yZ6XvIUvPQ1ojo7tdpgIwKpYG5FOeHCvVxFtJmRROJUQ+lMTm4xsVEmr+mjy9jN
8CTJRQZDyQk6qOfErkWKAHFy8rvtBk2O2Mlo1dYuEMhQBiq34G3cB5+hDwj8OiVuzTQPwTR8chpI
j7diApu5+IJy62NLPQRFfS+ueyEa8eacgbJpusDMwi5TOE5g++P55uDCINdTCosHmqPMtjxBl6Ep
/I16gpeM1tC3ekQH17Ip+0uOq4dnEsQUcvEz9Q8n4Uaq7PKFEM/Y7tfTRwpym2iCQzNoKedjydeE
d5s6bQwWgVN7Hk9uDQ2YWMxKf/tQCASHTz84P5JnacFJ6s3dmV3iCXViUBzzYLupdfTkRAzGp4dF
GPXW5eQT2qJyATnto24y3yfvrZmR0o4vMEHQ8UnLiCMy2tMsuroRRX+HPil+P1VrpdWSIY2xUhUU
9qUZtAn0ParXFb5AD7l0NsS3PG/BnE9XoF076WRCd3bEuSX48WzLzRnQH62f2XYDfG5Qb05l9EqG
CcawrUFPe/l/8sNkxY+yrg7Q4WgDSJnUu2Y8fKXGhUiTgVWBxjGeOSe9sNZLYN7FkcJ/Pa97Kcob
TNQLXqaONCoK3Ij0H+Z7TuMaoI0u8E8siu0K53coD3Dd2tFembSyFC20M0iD10rkDVUWXbLAAL8V
wRQBQTFUZChEmcCKJBpU3LfUFJ/5d4Bs6XnI/xs2XM7IFa/5IWmjWGAL/bFMHnc/KrQyAbIsUPlp
r6tB02kAUVVjHKwE+AbGY5q+c4yiHjQ/SqN5IuqApaWZNzTb7idYeykwQLZ5XYuZ+Q6KtqVYJiK8
j34luwSrB5HiaHI8Ji57iC9ubQgJ+JdgafTbuCk/U2OfqZM7liiE6F5mwR9xAF6UL42NK+UEO/gC
t0bXNATFO4p1HBDb6HKMsUjejnyk+RPs2B4fngeQVsiRFBnXOK1boe35sEph+lF5+oP3rG0Wpic2
mdzjIevMjyxGHlewkNwkQYPffQsNWALWLzjja5pFmDxdJ75kMRBfE7hFW/Ur5beJfW35FonE9zAC
ilhI9OyfNlSGaAcCsyMbnEoeAf5BqJmOQGjS+KakOzTbM37x7PKkEvLy7BiEA/XslcBd6IRRa/ib
LN/p2PY6LbjhgjC6/JJUFKo7yY3lNIGglr1ZqRbDWwJYNk5F4/z0uZpBTQXL9SOsHpV51wQ100yF
nn0hGrnpJjFOeetDdoeEzAT/gnpy2pwCzYftqYMuwsYuo+IXYxT61mIsPUF60Xm5ToS9UBQ4ywyB
2OfDZXXfaCVu1KU1pxV8NNYi5gRhlU9R3pOLTLEBmeJDfylOa5UWdzYiaejQmS19c+F1+3CBoupj
3hnG956exiKKkPo+AtenbJ/+G9cVHj6kbO3jgBs/M8yBAZj2CnFIRj4Y0LsudK2o2n4eah522flr
P1Xgxn0Y98pxd8S4x2Dd74dK7Z5ZPYvTllX7xt/aU9f5bypwzabF9OpRztcaNDqUbMfpfnxQfJVN
I4N6oZG5FxmKXNpe09RqudBYBjTInh0UcPPLRzZZUcJJeoKg+lhUSkFmoAmZSfi1MNb7MiFVipQX
sTTO5ZM+FML4WifGFkZzgEoUE4YW4ubgr7bWCDWaQsQnPQ3l+MmeHL2oq9m1myaXtS2eUJ/+LNNk
Qxaxgt/R7h6srxySRIe1oh8Y+4CF6ZTDoIzAarBNdmI5NP2TGjTwntqW1MVU6sQQBnpdSRelmT9P
mkhhhdhf5FF9DSBzQ8Rzr3aqhysTXfaobhLafFv01Yn7qnbixL0GongJW916Lax0WeKbHQE/Pilx
YBoJWlb082uCnNuZnkcw501atSPAU9pKYGJ/SGVB7XsE0zangcches2FO3UQ0ypeOIGlLKVPYx4v
lE+7ZDaQogFOjWNEEjbK1KhTIiiYWvQr5vHvELJwfiE+PlYDIPOpYCr6uj/NWSWAg4BCW8VwmCPe
5lVAZ/CSpcsgIaN1903+d4F+JvXrN+hZHjiYpoIUe39HjQOhL+qRXbS9FgKv3NDocc3HerLhgZZo
vCVk81Zh1WI263uX18LOvYzYPjlwdoh3Qz31sP3/qaBXb8nE1N9kDxB11EMW0aOXZYTztzuOWGek
WxsxfBKLdVwkXPibK5f6ZcPXSz9wgpTbTY9bKFx157/NjH7Zxokjgr2qJXcLo2sKSU+lOBo1e/J8
89UxACzkKKw7XbdbeJab42bm8pZJX6eNBkBE3vkLqZwEOqWQIymET0kbYx0oay7CWCT/kEbaP+Lj
QDKQ1DEhALHEPLiJd6Nu83e+FWGUzQ/KfAYE0yj68r5v4kZObV/feCNWHsZhorQxELosA3TKJ6wi
7SMeEiUTmQtf7KDvRzKYE4TWo4gIQaoOLp5dexZRSXFbkjXr/M8wiI8SDy/9Unth+r5d5eXYelzD
X/dmz9XpHtxJvfEL0nuEqJwhzBimBL4So3FY7A7dyqAnjhyNePF91+AR5dLHhvSCM8JFKSqLnEMG
0btsRnIor9R+DUeh5g0L/I7VsuZ+oaW+nxtT47OPQ4Cr4cmj9QGLWsZbL+3akmOyqhDDa/IfP/HC
uM8HlvKEdx53K5yUTqc3z9YifFV/zrU46G5dmuc2oX4L25dA7l0vu2vLoDFkFS5QLhR0C7b6RSaE
lFmwnBqOX9XNI9Lkc5CJM/oFZ5/KNsamwI/atpcbao32D5/Z8jYRL8LhqIcRXU9ndVLNhqM8EAB8
BXxzGftAbMXI6mdhBMim5qS+fEp3gFfJxXWhiNTUMRUSFFRR9rrKs5cGwNcVvTrSwu3O/0WjbiFj
2nbN/TaNTyTjy4Abk7UilwrkFy5hK1LyRd+LE6iwimTCTeBHSv8CbvldONVN6Imbu9xKJaCU12pU
H91MHz0O7J1Wjbwh9njzdfLkQrNmrb9+6nHtrnS0QYwpnQiKec3iJa6l+Mkql/Ut3xBRudBCcAwo
skOW6Uswl6atS/QgqOk0/bZJKgAyUv9vTJUGb9O0OMXHPzn6wFHLNCDOZDslvPPepDlWQT2BQrqf
g5a5468G+vtGY3A7DNOGbNrd9fEC/ojYDFgmF/N7yh6R5XgBPCP7AAViPpBz6CtJ8I9GnVe7SxsI
z2oPqwHxcwxygwPmicKiXBZZyEhWkWiyvkf5Cg3OSr18Mx2EVxFJAzzbtOzHGhXMX+kdCt1LXzk0
xmLTqSQJILkcZecGSPaAd+jNCjxAm9/IAytVPkO657CHI8IQAaAGneYuog6VW67irPoLDfEmOxq5
FiFfyZxlpzWrlDzVnCL5OaKB7rg8bwZ3zN6WDNBKpvhCmMKK0x3tKpajz9PAIhL6ziHGGt/82oLM
+EfqNz1dBScHgMij955fxXBwTm/4+ALoUWnR+VI7ZuLfCe/ftlezLAGJk49N3UuSivU6oz9OkzWr
fWZwD/ppcUKCUgr1/UIYkcnN1AqQbugf311GFmOLyPJ+jzmloD6Ns+orn3flNv8OQ1lTjMrmKLCb
PRhMKyjvAXjZyYoziXdgioIrJiYILxq/A/lm3LcYM5BLyszQIJITGFQ1s1z/7g/dt9ofh+KxUNWY
iC8Jm2u9ccbHBq1TXJM2ukI4y1LcGXShqRt6OffPfoMj3Jk6W/HpZL7PFPPZtsK6T9miVxryHSX7
6FuIqs+MHacAk/2CFQ+PXA0WP5nzF0HcfkrH+HUAkLH5ghE45B8lj8yZ/uOtiBHeLzJUbuhjsHoQ
EiF67zCDiihyGQ86MCeRNfQaN3gGx/BNGMRsMqt14ksSPowz7XQsvfSfvpUpN3LIkBRFnjLQNxI2
le84U0i79l2kBU6x1jI7UZ9bdG3uOMxXRVtC0hyavmlMCB6GSE8On2br09rgtpJN9CFj4fPKIKOg
T/TiLaCWtT3jthwtPxT4HNzXHG2Ht17fE+ys3WcxZpOhB4iv4jbW+7MR86nYsZujH/Bfz92NaMxg
kFfTkRdoqyVL0porHM9aiaV9ntyPgzYh+ejk9w4Fy8DtGO5ulnBk1cxbFvEWPSo39OIwNfpftfym
LbAu/vgDKz70xMVPdfX2M4h+Fx2Z0TnjpzREE8ICwcSF9Ot0LxfjoZ5YkytwqpCtTGn2GzM0+qT1
AI1+qSyL9EEdk8LYtQ+J14JJ+j7zG3hBjj9cs+aCNOzN6NQcz5zakEWsD5GRTkt7F+AS2zzw8QIi
rVUj1BS7esA+VO5E2weYJePXeDRq+sAGWCrhIeJYFV47tXScxMEM1Q+QJaIZQG5Em6vzbPQsIfY1
0IdIGXaWEFjVps5vwZsbPhshVnK18GpEO3lmXtmYz4BibwM80yDertq4RFBrP6d9gU9ltG9j8c83
yoWin+sFyjbwv/nlMDq/ErDZ1rYpIJ1M50tWwjYpmg1HYUA4q3XVsnHbFxQYyycy+CB3fbGyCcMu
XEI7zby5TI/dPE/2vtE21yT5cdDsUu/+WEAjm+Qc5BdpDb0oWAR04Rx2SW38asiO1E4akIFWZ9Ix
3bzknkSgKyd01EV93MjhSUOt8vOWwQBKicXY3f9Dqwy9gVswaaouqrBGS8JmRkmVeeHAg8U7jIbU
j74KC30g1UJyQgFzVSkCiXMXBGmSScQQaQSrDVw8R/Rg2yfT0KmD/kS+TrJqBH68bY5yUz58fwLr
oU9bVKsQLnxmfLqGrdmcV5/7vomxhTsYyHnfk1kyaQ7tJqfiLmE6UC7W1uIv1ugnWo5klSlMIVnH
unolG96kUmw8rl7SLOn+UrtRzns0jdbbbjSq+qgte8KTWFhLTRhDAGy8GKr4gksPC0l7tfe1fG3w
kgx/6796NHFeh0/ASC/lhlA2jpV6X3TnU/ae9S7gT7cjshvsKc/69JxxLn8Pt1rYgJHtgEQwl646
GtIo5+I+XD29YvquaQfl0SimzjtR+sMygrNF+QdN8JneMtNUABK78Ycp9/FR/8X2MziDOB9LIWZM
YQzTrKvKlha+GleahiB9kp2GVHstgNqrJ7MLKGuA+zZz0R5RskM0h9dOhJHexrf3A6mCwJ08SEco
tXpsviwtUMUqEKVW4mv88ZRwqkzK29J6T0x+n8Wn/v+RXeMjl/lXJZKYlZNvV1RforuSSXKxajtB
ZaYZGg1+TwnBbgbNJ5ZeQqUG24U7VvQ+CNmIH4p0wPoWDLCbZCHpdXN1FUVhwewOYQi87JkmcNcA
REd5Cq4NaVgq1503v2F9cCXra+eGnV61L7adNKgsVWZFk68KNm4beX3iYw8ubvwMdgBTaZNsw6XU
Oro8TRPf0X1sE3JbqIaPtbOdMlGZrUiJo6zU01M7UKdxYZSF44ik11QfSAe+/ppWwscLQBILRsdb
UUuVpckRGs7tkzD0PFc8t3c9pDU7T/12DSWlaAW86NIxKOQV7790bmdzCq5QEEIGZpDD+itzj0Wz
9rG+DgnoqWxuE8Y7ERb8RdjA38vOCzkVNvCyCHWwUfgDpY4HI5zl7VIUe/hcI6SMJ0jA7p7gG6nT
opt/hdavR+sAH0iAnrSFfN9V0UN8E+b1QIMUxa3EfyEiCoPHlbRWvohd7dC7AuyXXO4f68CWQ0em
cgl8MWXzeEov3KWOMJmn+zGyRUTTgiqizyDS70KCP6HYjz0NHsx3LdnGNzE/cLMrv29kNS/CykmE
o2YDBKo0yUFK0Zw1CnJ0/KntBOGBbkICnJj9zPwmahChmLn0L2kQUIhbOJHJAqiPFweJ6JJSg+yR
gGcDjxxxVc5G5wQvESZFr5H/OPwbJayLyX07eA/2of+dxWMPb1SKx2YA8461zZnB9hsHsExd8cFj
+7KPn5kczsd0Kp7n19xr57bm3vL8ywylCzB2sDkPFuS2QbT2+fXhsaunmZjSgKPtVv8Ex0qRYckB
AKpYlvrLGEOEFcz/IQc3QTbFWUbbWr5pQBEzmd5qWii5M62336Pnve7S3i+g4zKy7cXxyUJ3bFLd
59Vj4vLUn7o5sK5gwAzs9QK2Vim2RZ/PtvJVnlBr85pkTHLS66F6YZ7ILSQV/Juxyh8rUasBzWPJ
G7RjPfQXUGD0tFK54W5E9qXIz4mO9brHMqJ40ZLj/zfZfmPsh9PVU2oxbRQjajOIfU1pjpTqNotT
W/yyOwP2hclEYfyilt3jvPAJmsrSvSEh+5BNar9V0wPNjc26LV7kHolJqowLoSaRJVOXKxudehlL
mYPJflhrrLSlvApPS/4/STXDCaB4Wajc93DP9oVe4fcVcn65Lz1ullSdj1OO4tZyh52zMOi8zjdN
YeskuzpLkaDVAOaxzEaBHh9mg0HV5M0SwXpQWxsWEheL/ShcwwYQTvrBrasI3ySzZ0awUfGR38ln
ml3uA7OJkU885HMKSjJMPVur9h7UxjZqVqOH6P+X49VTtn+32vpEh27XhrjeE2Ngr85Bbsm+YVG0
xr4SBZVLqjoMyqP44+qdwlR0BEJ/lVuM7nRsPPxylrt7Du+3XmRVaAetmtkzHjzyqUNCkVwkTkDv
v+GmOsrp6bo/jgNRexx1NHtZY5rTAKIDzQTFVjDeuXFH/LlX0YNE4YdGEN5JuZeYEi37ZZgx94Zc
LI1VFM0zKfGFwOGcnuSvkbaL605gGQHMa0RoCiDs6nK/MBuEsYEg6C6/cPUkXgqRXmoLbmguQh8E
92EDk5kDmHlVHa2pNthnjWkVTLVnNqAx1yKADQ2xrbDkkcTNbi1aNW3j/JCqZ2/TUGVDZIMSkBYr
hcUTMFU9Fn4xirayff/hn/D8VBA4BnTnF3If9FbwcUQlT4mIiPPYWmTVX36o6QkmO+NDKMYBtwfu
6Ra9Rr/SCGAp7CU2HFwW26NLo/T/gEekmmGpq9T/CL4EKsfeaY7RQWqWDOTdjaCxPPfQtQpdukon
9MasrQIyfU+hL4JZE32Q2DOtMTr6lTIXkkeeRHkbALs0aV05zxwhtiURYOP/lrf57BKPOoutAnPw
dwyQwSDAg6IHqgzrYCMYRW17Z55ncLILFGh2FNQXV2FaQG9ni7wnbEZErPZrAN97+1oIGmyRDY5R
YUhbGoDvEvN89k7jFTO7e3GQaq0fUKNc5s9qx4+XdEMDAz3DvYQtVCTUANBCdc0FdO7bireVd3KQ
Rr0FSXr7XDgybxMcr9PyCfTzDe6XFdVGlHapqRo1D+i4RGnDhrXpdMSUjJnClGtFm+koifdKSaZF
ENgvJJI+62gD+fIkeGCeZ34piFhjSL0b6wg6pGhsU1+7qDP/bxR/dj5LHuhJMUw6pDcWAgEFFqRL
8xCfRx1lF+ioCibaZ+2riENDfNjAFyJ88ynW+tFKBA8Xu/5owyhUBOv6lyrBI2qcFtSETZ4U48cp
uoWgi0Ep+iQBTfWczDPu7rS4CFiiWdYk4VurS++w7nTd1hPvp96frU8xyQMapoRX5DNPmx93UQMI
HqIP/eNGKzW2aWgjvxskZU8rQWu8CjHVPi7Ovmlt1R4Acz+aKAs/LAbPa46+jI2zW6tnjMmb6lMk
lpPoYm0XFZ997WPJqlJi9Sml862UsZN8SN7CSgZlMkYGrpcpcc8TxZKwLXLOGLDTUAjcHUMCn10T
MtVMoOpoGJCFVTksAbOu9qu5S8rEmOpQidHeTNKnp4/lXMmOPxZYcoD+UBNJRuRxWLTjlX8Y31Ib
d1bH6lST2dLSyUEId4jThjrUzfEQP5/t072NFhU+uoNeZDcR1YdLghfE+v5avnfjvoHlF1wPo6C6
mxEeK42yNeCGGPkSyayemwgQ2BKKfcTxqWYEcw7iUktWR6fUPXdPLSGTPB5S99s8AatHdkCrqVn+
VU+yZ9+9+O4Kh27v81uWi7Aw9ZI9YjI29vALLNiBlL2yOYOuz3mT/UMlPU7GnsYFjXK5Vdd6qPCX
h6rTjz0IP+UNl+KzhDumjUucT/Y5WZx8XiyR4ATznvDIWmzE4MK9iU9+fvJF8zrLSmooo83ujCX4
OceBSwV90m86m7yr1+g3TfOwvbYBpj+O7TRmCkgxBRcVr/o59y1+2TJ2aRPnKLu1k1x77WrblG37
x8UKsJm/o4WjZlKGrS95Wm5jM0EhuOavmYtFs9L3jf94ibizeM1EXaR2/LRORaizFxJfcN+tEFbN
VUIDjclX9/6JYPnNOcL+dWqokZ/Wl6BkjOmi9iAgj4ITYxOSdjqyuUW/KL1fvTK5U3QZZey2zBEL
n4VR31B73amyo77samFHeQcFAjfmzkc5aPnixSHpVdj1iiI6cUixnchgBTQ+K/nLZ8WlMIzPWDjc
Oh7FAixCSkiA33zyFhcRnD/vaaZR5ilcixcxYSwsRXfh9UFlcVIbAPuF1p+0E7DquVW/QG+fUxGd
zdPFNGBarOhWT0us0mqEyC7+8kj00SQrbudUoyspbxajkrv7MbZiiM3UxspH9PgAzxkidtsLTb0F
KrBTJbAgxpe2qYN/txftriNcMX/+bZ4NVleo+FzOBGdRFTZVz+wGBfmPZVshzYBb45iO5+0hcx5g
IA2gij9gp+58/OL2wmG0HHRV6ukqXDozqd7z4AHnaT7l3+1nJZ6bRofxS57CqwAHfVYDCIaOVdhr
6ftyhEg/uzvhC1NR8IH2Qc3hawG9EBN09cGAF7tpeeWWPH27o1qcz7eLqmeHIzh7ZhK7Prf/E0JM
lu/6B9NURF8o5AxNMv63VsTT2hWgqMCi0+F/EGyn6nX5ByxnCUj76xsy/ByY28iQciHUYIasmUG5
M3UNrRagR1jNFSWwiEqndkBudJeguxHznbXZa6tydx/mTymRgniUKocdaMgiZNFEeJakTfgYYMpv
ME/JI2JqukfUoqQT3tAlDS3Gb7kZtXp4HvHAqxkkndshww8W/+pNMjV4DZtvNxjkA2wAz1GoL3Wc
y5PhhQU6LKZWKtC75su7XlF81xUBFzY10qBKnSURFOUHmlY2goqW24yKahChRc5uKC2IxSzdxBPy
gucyoS63rA/yDx4TIabHZ5YIM/Jr+/MzrT266N1/dKGW752Vvo0dUYGWNkE07kVLcbbso6BeC/oy
FkaY+WzVlMJNhWCuIl9+RHGRCHk0nUOfo6sgM+Zkuip8OfaPP7mdGA+7Gde/aOY8vmSHhB5yUJ2m
nHfJJqUNmYdFTeLfxH/BVKueeor+M6h03RIgidFmxCjqRK72masltQcUmbZD9tkULY1ZvsUyvGlQ
2eYcfrxb2CIfcLLp+dPtXFYkkLkNgDivyOnpKZ1FHcw5Z/pTsTpWU6KiaFIEQ8xwd8Lm8emiCKpX
gDr5aQw+3xdai24Cf3SANsUfPvsjmnXzNy9jFzDVhZItFitG7RWvenTvVB7IMYl3JttKOBY94Oja
hzRiGRNVc7iIj1MZ8xOn9htfTh8gEyGfoYTA6cTsJBdFZaMC7kxnrXJgA/tz1VaTZxeaiipIEaie
077ZTYlUwUM4ACJF7lhqWhtw60H1x1DT//UuZWm6i0F951N7k1YmvdS8F4BLOgb5zF1ZPSWnnTrO
OlMuL+mdZOsm49qt+MTqWmWdLMTkpDOJG5cU2biTRiX/7htV1nOWyYbJsiegvXY5Pb0iaklLN9y+
7GcVURFh0lqMOuswh1qUZPr/tYEXFyOi/u6kZhtHS95sB4e1HWL7copX+StYR5lxFQdKWw7dA+Ai
v4xPZHcdrHhgT+jVzZnMczr+IHYYr6t4dtTha7dak/AruE4Jzv7v99upoJ1N73UNDjiWksR5pMXX
zaFmiE5Aj/ba8RplHTKBT1Zd7Pe9OOt9/LnFg1gb56skze7DxupvEaDPYPWBympN2iKfKxXH72z1
zlS/D+6d+p1nO05ZJNRKTcFlnktVwOGWRJ6EVTN0Cdry4LfE4MhSPAwqANtdyZVY0ulTHHCj/ybv
pzC6K7MK+gy1uAF0FkET/j7yuLlAogayCi0caJAUEp+nOVY0nSOLYFNs3wp29v21QPfD8nZlkvvO
MhX5DC5t35O1sF/+dI6z4P/7uODaEjQZMcODBXxbfSkVfhIvUi3+6Gc0ZB3t+ApfU1PWUwc84XER
I9AISiRHgYM8Oz9GF8JFAksf35X76Ix4S4WLLYRrKnx5S2sCR7PKGDaUssigrvQaFQ3oXP0XBfaY
2MnXCRevzd8PvGZhv3OpQ1n1lHfHpHa3pHvl/3Bp0hk0yBmldPFxWnHInxnj7V0g8cvTL+SW8sY2
ootFIJC/HPV8diOSxZ+U48jsJCQsInGrt5c6/KHRgb6xsOzhalc4ObMPDFqIDE1KCJ+IsRL8h0Ir
P7C/vwSlPCOnT99KzFKTu7gdCL1MvRo+jG6y0OjYYJp8dSi1qOjdq+lKj4rWpnLNLOkeRzt/zA/W
G7+Dy9BvMIFA0al5H8hMn8m1ks17fYVtqd7xRTWifbZSRfcgiTF15Rb3Xh2rs2XpHE7uQl0LBGuG
QESS3tqWfuqxMpdm6GFjmbJKeG+7/1KGGInRk6MpAV50Uc06AHw/zR1iSsRET0QWwb5rEjdQpWHO
eflOqiZ8roUt0brO5koqY4CEn4ccxx7KoHRBiWMOzm7vr0lormjfETeDt6S4ApnIIVRO0eb8P0EF
Pi7o9N9MQmgVgdXKtlTXeaD1BCI/BmYwxlf3haMkejSkoo/N0XIxg83Y1npaZPR5IqCpLjjQ7riS
UMJXM/tK+IcL9DAMEX/Ragu+i+JQ+GPMqzsFcC4pKK2jJkg2kXSwACAyCD1Zy+aHSIbPxlvEBko3
EXpstHcTP/GRzxb0UlQBsIf6KRzYxs0g5PnyYc+Wo1om/CgvHJKBDcCvniq2M6eaGcUx3fMpNEK0
MOSqlFGXovyGiTZRnsdM2NnoGF5JxzKpqDbk1HJ0WgCP0uXl0LbuAyA+DXC5ZJASu/WEYucuqLjB
ssgPDUcB4k4hFH3QH00z5Pg6ykUWAML/wAKSBsv9JVDPLQxY2NayE+aSI3VRv4teDnTESumr63lw
BXwPze4xB3vkEmxndCi0UgEpgOlFt9F0/eoYSfTC7APvo3OAHubQWT3PgblcqpmF56IxptQptJhj
01iopimQdxhzpC4timbYrsiiFSdYPwKjzCfaqfuy4lMPBR2lF6eJqbwQgKbiE14NOiTKDXviNdCd
cv7pfDvT/pgUeziyjV/H2bTNSpJGpfr0SEVhlJTeBWzBVMRQn0BQu707W8hGuS4Y+N6izS1Zeb9n
DD03H41PWWzosMbz8g3F4KXvj/yMPKhM4/gfVGUVyL4qF5m/lPYoBCX2xmU8uayfoSvVmbffNFCA
9EMBmmFurCKwfMnobKxyu8unWzeSEq/0fPHWX5oUoXyYnHjUpesKZkxyD3MqEy0cwjeMCevqnHGA
GT4LLR0Ja+MPm5YGI/hNGFGBz+KBP1ckZKxZ+H+koCgdqvIGZxfa+KATm3AVGMxN5hcVeDzrwmos
z5+SJE1da+u0iLP1OAMERNLDYGgGi/XuCiwotfW5hKCYoPOI1Rj5scAfte61WRRLFzm9NDOeM5b+
SHbQjI7LvdzH7fG4yoW43d2elwOPFbRJL3miqfTI0AJqS9DvTWLh2zKxrW7HKBbPQ5HGoZ/i44xN
3xLMidpmiK/B1iu+IecmiQ6Vlv9cYqsCR7jdCmFwxzFVNoRDKS5qenyi0EMSwhl1rTTycMoNdT8W
211KhjAUym97f4VbC3ZF+rHlUnpwiWqEIc/pb9PadC7XeHPWbaIHjN41jTn9mTdbcv0mHglt2rlU
3R1A2ZtSDXI2mW7XwbGbQRfFnoFs7miT5LodTzGxRkC6MwaqM/Ts7h7hdXI/U6qJiew7yL/xEuoL
jxSYU6mAecDcf9ZY9w380W0bWkjJN+s51BUjqffoNqFnC5e0C4nRJ7rj2VxcLE8njT3UzM4NXuir
z2z1cWCxyA9lsL/hWjDuI8bUr7nDd/fZ3+1bvQupqutXd9S2jWOwItrtW1c+QtIrWT2y9wWyGdQE
eR+uhbPA8tGNJAcLRWKCdVkamNayT4yBlzklfVcmYWIHeyv75/S6rizAQLse5Hn4G7n9zXQn+fMk
qfEyvkyaTTa4DALyl5r4fEng/ddMnAyqOsqViiibgeWzHyDX4rHn2lqtkJ11bBu2h4iAtwRiKa3f
/YYOMfvjpxXHYo4ic0tMRxqHn6yXCtvkeW/s7oftsyEmRVmMHMJXL3ExYTOy3Zzfau0IGPrewLWx
3jSskaWZl/aurkCPxBU7i9WLi6WzWw6T3S3TDeuRSAPl6bVnjl1u43i8F+0WZDQZqAK6dQ089wMy
m8AifpWFXhzVGk+N0dRSmNV9xyizBzEvBspqy0RKlSxATZ29C27kXSaAwOu1Ae1l7/x/WmRf3R46
x/OEsVjEq/jJ74nUOMwJyEvwJD+Tp773werbPTkrHTI9kMu1n4px79vVpdCBQndLDxSW81qkWRyY
XXts8/Jd+cvqmHmnCYLcD8SWJN083Iq0cfNfWTdYB6P+HzDpEowzUAbli/ZVsBwHu67XD65syPf6
Vt3UYMCn2O2YO7EZaqLVxwCArNqKyBmGos4VVU7WfkbpP685wITFIY6iiUoqipnf71S6vRLBMbi1
XG+DoG0ZcRv14P/n38/a+7vZ5A8/5K6EfjF7+/F0YK8+1fUOZDxC5Orz+s6wm/nfe3tQQ4+5LNw6
9YgVrSllW2JjGjgkfvi8ORB9pe8A7wP1IRci9ytnLnooqkZjwSm+fv72tucCqdJk3Agjm3jaImT7
DUWrq7G48xwBtRi5KBaGsAfXgA/neXD7kPWyDCreVowanOXkGirdncGe0/sQB+Ks8aRapp1KUhsO
rQEvbgpficlI2vwAm43R6Bts/Esew0MchWc/tBT6VxZwvR8g/XMGVEOewNZA36VUIf7wlKzmdHUJ
6cNMbA99Pxjr9uRJFIumQTM+3SES20sGAQL3o6Eo/9/RZQSDu4Ch21lK+ujNgSMsyO7PR3lJHWZ5
WmdTU8eRhY4tjHf/pxzxua6iOKmJl05g/s8CckAQPX/1tTP+UwqlsTeG2r4HLRKg+PjKneC38Et2
SsVMbslE78ShW6k0Anz2kyDdbpaGrwou0bWMAzzXZIb8fflr0g/JBYBiiW6JZ7KNKGWqf5YbH1qq
LETln+xi6ZWBkIcxwYj1hnZkYf0nOUJQNwfTdhYgagOxPGGeWQRDRCOIx8NGDw1YuKLutmrOEnCO
Kmb6MoObiI7JK8vIyYuzJzVE4VlBaxj/ymhyAWKPu5ir7LFordxyZeXZcYQP3ROHiGPoXS+JcG5t
6qdvgrn55TcrS2emuGzHHI9bCNG7nAZ3oE6+lIFKndcTWes/SSnb2DyxzGLrDOSPBoMAoeXgtg/E
cnqJOiTWUTJlJZnjUmLpSapSk0NooxRCC+jySr6o7KzI1YMGqXGsYfAI6Wjy5al8MVZ1FHB8DR+/
bydWONePa8ECTjuX80vt9gSYwIKb8qVkCeYHXIGE5QFlGwEFOJ9q825HIxqKetgo+N+sesPnVG/i
CKtSbQJYEGElrRGzJe7YHJG2zYQKLyt/i8dV5LeXJfs4KABfNB7VVMulg2bPeB3Q62XeoBXvGOu4
dCZNCEWSBq29c4Z72K2ITDODjUPqMFI/4oaibJ0WJAIaTjiE6rsMK+gYWbj0hwzlHd23KGSrsiqS
fnZAHAe9RrDzbHlna28PXDqjupWEW9n+FgF6KxcnSkwl3lojqdqg59CTfbPoAPc6ArWjumq1mDJU
w8kir6E1v5N4cozUQV/csxaA5PhUddMX5327u+1D2EM5r1RaTE0M41tAvsR/cexF6Lz23ZId/X7v
dYWvxZjBwZOefM4cDq3qPyQcIp3iiiJNaRkrBcv/EGRzQtZmB8/yoIkYJhIiwrzeC4XozfFyjqPD
7v4AdzSJFbHQP1pHxTVWYZGTBGolQIMdwmQD/3B646wgjJAEm+0KBGaCTOBjWpXFUiRlmf65Syoq
67dqtMrnspfArcmAYO1oy38dYhghT66TXUxm157rzM5iKUY/HEEPU9MvgLTA4gVbB30qj0r3jCmp
Y3ZRaUHala7EPAXuc7NWmb0M4o1nEJKNzdCmKf8qvTQD4x1RDZYNEoEnmePzmQgCPdLq2G0gEW0n
wCRJMWF2pfMIGJYORwhObl8mYD5L7RsW4R5Nq0BwPzBkRTEYPRDt9VUHOpB1fXHPZHAk1np2YY2s
M/LwwWjy+bbzPEgISqlp2JfoedUSxmXeNZEU8dWduakw/59cU+MKw1PIhWJUftpSxqz2QGJBIVKV
8w+XtlFDpNr9OYhfGFQk5LPD5ipj8stsCKqLjpCX2/uKfKK332XjR8mH+A18kU3iE7WYLDy8p9mw
/8GMVHd+3dAdYTvpPIqsShZ2l7bkyOgctylwvS4l+4u5Drx+qv1SZ89UL1zT8ce4dSH2eyt7TGXF
eZpKzQs5LUWiXfMfWLVXaMuUisv+/cVWTHHc22PEKCA5mCb+rOt1SnYhS2+WiyJl/d4qQmgKDLmU
t7eGDEBPYLuTD4uujlwpiknGroveyAV1T6TjXQwKzoc8cvLrEhh+vIAaUtXvnK8dSlMGc0PZcNjT
SnufYi3CZTW3qSA+abN9GCu1bfpjxPHc/Df7RdRykOlc/iCHQQILxapv8gjz4qmqV1nXWG1W/1iO
Vvi8My2+KH6Pb10cN5OhfPOACHltC5uySM8XgVAAZGAMU4qMMNqujPdT27Zja+EucmFxTJ8RylgZ
e8s3WafDwp0vhSOrb09Pp5/ViaDCqwYWnmpPQO7eBiwraxWhMBl08fYuKNmYZLf5tzf+185UCn89
4kP8k9R70QarOTC5jyJltObdfp5jxpYQDPglCrG7SvZ8O6tb+0ELAPPYxaUel1ZKGUXh5SehV9rb
pUUI9ZU+gEmQxJ4Kdd8zLKlU8rwsYdoOOhgN3Z8/tAIoq1lJdCAklA2Z9na0P9kYx+vX/CIPyE1o
D0q6buj8j5c043I36LLRVQtmDvyAXalsoEco7or6P1C+5d5h5FjWMZN5HgOi8jP1w/ZJOEPdA4QL
hCulSxG8cBYzgMW5gUlOci2o8/Bl5ofw0y3tqRRF8PKN88MB5jd7JijDptQvvhSK5L9uwYV4qedi
Dxgtb83fFe38FFoBpLBa7IYjpZLvAV2mzFsyfxg4Vs5ZBxKgddK+mT3F8tjYJrs5hZgGQWt7UTup
dg2Mq/YTmeOT/7mNNXRalIgjTKkdfPOFlAzrhBpIzOcGKl5K024HFmzsLCrmkjOhVo0AcObDLPMN
JgbiVFBhiUefXfY88lBtrpYZfRhUZAIgoGDMRmvxeqWtkCoYwH0lOUKvf0zKNaS4p6YJhhhvdRWi
7ThugI/LnqLD8fDrSTWTUy8+9Li4H//JV0Qk3Me7PCAYpSecEeeb6cwqFrL22afKcybjSRcHnA7T
gP8MRva5A23ldfQGLp1hkp1upwDt16OmeWdaaS3eeMo0jpM08aqY5+bBDqOSLDuE24YvglyBlCDH
iT0TBsl8H0OYDqF4eoR68Yoxxl6tILsGPtrG+MntWDLEeZkgKXe5cnQoEDdSU5+6BZjqn5pCjQOV
nKcUnsZ6qSKwwo7D9y+Q67wqmfSOOsF5v5d7Wvd1/0BXmVCQ12anx0a+Txm+4UIXgfBCQmEF+rQc
saGA0L/0P7kZGh2OFPbWebyuj/K7+7rMaVKtpgcCeIE0uHaVWj6iB1cZ0TxEIsm45RsSn2eMuvsy
moGgZiHpB8rlBCZ+yhtrgZVd05hglrS0yQEdQ14HR863zi/xkyDusmWS4UlVM/LTVb8I1VaPMmXs
44yCH45ZG99umnDHp1BeUnO09Bj0mqAdeQiBB2W6Pw9obaKPci01okhK3mkDEqQBocCDL1jMMZGU
SEaFV26n2C9P7ROy3NT4X0XSUuHY3JHo7x0GIaEYTN38eSCHLlf2FMMpSZI+PVXelc55DmDgfVbv
rMRD7BNPJnwoFTQVpMJ/VyUkT/cjaS6Hdyyp7vNnbuFjUeAvc+1yr69gKhjH18lJkrbzAoXNz6ak
CEEZ969BG4wkL1X/gLqKDNb321ZSdWGkS32FnYGyO7HNuwu0X/mdN+KdK2lz0jIgOq+Yf48E+tbf
Lf3JUMeOz4sjcPInO4LuFASElNMRX9RnSIgidMQ9BBdip5OwuqN+TmAM/BCLF1BT5i/0fLg6+GkF
38aJvpikeIiM0uR9ZauGDqxZBMwsNDtu/JbxcgLUZ5W/t1XOoY7wgsQ6J44Gv+D235gHPd+qq1eq
giyln4O96WM25BcPjCrfu8nGJ1xZlEnzPQlNdRu5ZhEJ02hsts96WG7w4nGE2WfDJcUsEVbQNPJ4
CAhqH8eJXpwmRdOa+LhP2RWG38/1KdBTPBkV5zmOjjg6Ut0PiegRcPPom7SFXB/UEHJQS3m8j+un
8LctS5Irm9oOCMv+LXXGLZpCMMaHVtb4i9SXIaqrRrL83sZap9BzbEpkmQIJL4YLrcc+1RfZhTLp
sl5BmBfPGnWyRS7rDNalmAdR3kWCSuXwm4gXI84yatJXooo4z9vPcUgUST1evuia3z4UzGyrJSA4
r6p5hiiLYf1VU/ZfOj6VhrWttmxN22sc6U0I4b75nlqn3cXlCEoaqNuHbjPLjk8zwwBe1ge4S0Un
tyVZ+DiuOX32KxflQb5MlrhUyeLEPyggv5zCGcKGexI6FSf0Dv/x3ob8cFJEce51SLsfKI+I4tPr
lc5/S7u/50CHmYlIQ7Xsy1finAbWC+3EQ/LvUVt7rESZuF+NbdpRVSuLiQQH/1+0w2jTyQF2cAlx
QcTUqZ/fQ5ztEJy1zCRupvITaHGLYmnvZy7w+SryL0+XIQF6oZn/olRSRgcU8iiD+eNa3pkHpaM7
7JDIhlVvsLCH+p+jn/c+i15FdM0Bkc6q2eh8w53eWzY1Gd8cVieLQHtZQiW290PGd/DSO+Ycr2oS
KK++P999KYENNGfhbQHineSVFTsprfgaFnaT6XQEcNBgv8MCJFUDC8ZcqJ/IFGBSm8lb+BHF6gho
a9aKXHhbjxoeowGQsZFc05f+2XKy9bMnfvKSLXAL+HpIQTcEPvzxPOTiYVF3tOSxx3SsdEov1W5M
11pRdKHrUdYHkoJkXA0klU1ZlvuGDXr5p7CoLaHLF+2M58piaeWJSHbXf/ZMuvKkcCm2ISfDJDIs
tFu1B4VTiLgEMXeoAe7QiyVFggUkdngDbo2TukrgKw93vQxfLiF19g86FVHjZH8E2xmIgCB6R9NJ
70ErxeVT7aaTfpx6AmOVKKofEC4iO8atmY/3naE08ZLONHCSu9KSgbaNCpy1JS9CdocP45CUM+68
OPJ3DHh6XABt4mE3DSMU2g85abwtXiuXa2H+klIWX8L7a3I7bn75QD2YoYX2R3T/RusuQzGkey2o
Hef2ziWERUw8rQWs1lAn9EbxgG4rUYEiOiuNbuiGpkW5GwL7AbAMLVvfW8tojlYNPlk3vUmWqAbZ
FEu4grZMVxXKA/fP6asRvyG7Y8l7Z22KCpqBcX52YDBbLgXbsQTGC65t2NkV86r4FUgqhRoYWb+5
v2exCD40ZNa9jcS1elR0uqOAxKLt9GH12fZLXBRn12IzvB0hNrJMYH1MlxYOdwAPtEm9Qh/tSfr1
2AEQI7wdU8YC/Lt35IDRoidHNXN3WpLUNNt5V8VFKCYOLD9wBnV6B79/K5szRDjq/SIVlFMtlxz9
/Zpp+SxaWjXr+szoaJJzGOomgA+J8/N6pkWhu2gAqbe67KaYTPpaTkqdA6Gl91YD3PBAGRQRO/jN
yzv4fFRZ79AN9tzPeVlEzqY/wIoIEIfPOrSKsW1wYlRZ0c3EYl/6TwuFokYRDDxMHScFJKMCHdc7
ojaseUcj+eUrADQ6h+IooqThZcN5GxSduHfKR72Bc7I2OjIifPqFHYmCNb5DOon8QgYvzPYWwKpv
K7+XNcG+8DnklmD3fRJ6j0pdfezVm3T5CRTkz23E3UCWQaTnrH4fy3fkOK/OGeb9ajMy0Q2wZWW9
b4uSpMH/hKa/pyOq7ZhprN5Qsqm2nf4dqrw0Vc6KvdgTDMBPwbAuIFyfyoKs+VlVLrr3/VYbNQLs
bnIItNugWbKNq+Su09mZ2zpL+3U5KHmevSN1ZpdA63SiSmOjChM+/mX02bRlODi7+adyoYBOUU6a
KZjBOCGj6qr7f2cUuioFjYXGM/CcvIgUCCSIKkBjfrvm/ZYSrhDiFenM9dgkyYcYIVsh6ypFU9mF
9eI5aY9amFPN41H/LAgO9nPa0FR4X9vEuI8rJrXI77WNKxZ1beRci9A734AgRG/34jwBt7qP3xX2
WHnCPwoiy5ZnYlLIg/65YgNchmTqHIsma6LGreJnwH8jF0DXNBLL7ofFbUNrzuiWeJgM36M0sQhu
TpUKV8FQM3NySGkreyHS2Etcxuue0tXKH/27oTWoVIRa8kQHgw32JQJsaVv4A0bnBu40QLI/E41K
+5+jdL87tBVNoInhSnFIc8qITAF+eXrr/yj7c3eu+ILOIrubQygmUQ5e66RBhuXc6aZBVLlpGFNb
2WP/iuaTDzX41W1XAfrOzf1oClebiQ+D/6QWGf/GMI0hgk4tFt/8u7Fyx6DhDP0QbFG/WF2B3Lll
vJfcc0mSw19uNNHDDxZO4mcq5NTR2XuSxU5c5E78lO3c3BsT2Z4W2tkN/ODTvB1V+FU+NuWnC5ID
4/jlOo63vRwnoYtWnxgHWrFm2OIV8bbS4mfo/qNnTbHUxwztd578rHU2xZZzQbmj76Gr9U/NxUfK
7B8XKrTSfTyxwQ8CuAe+4U6Dkg+Tg/ie2jiDx/Aj8ToES+0LPa/4DimXTHDKpQr0k3DqlQFGmsus
f/gN3IjqAnh8Xx71IclGTAnsM6Ygke6JeKlEoGzLC6vsxpsSD8W+g72YrxovG47YYzZ96EYpoAKU
u8fvZ8yX0CWXvcOccRX/+xi5x4j+aGEkOPuG7PkmZBwFq2AZnq+iSu7QwckFco/GhILJIltKYu+V
SyLXHLzHwdCSE/FoEZphBT19kQuOw0UPkdczYig81Gjr0y6lL+QA14dlA+Llsw8K8Ulkzp7HD5eh
A3U4hCLYCxbokEq8YfiXPZ0YlVoVr9aXiUw3mVIef0KfLgOfG4iV6U2l95t9DXPEzb5lC56n5RP+
zVI+F1WcdAAtpbNXZaRPHo6k1SrWN4nagnSCp4pobgtOzuQNsLwQUWJt5YtxX20RLMDtdSCS7d/H
V5mM7bzDtkOti/7pwIUNVgdq9dOJouNArpw9XyxVuC562Vqvkxn8n9hKm744X/eppj0LDrQUD4wO
8jYFTvINRMZp/9YopkqvreKabgKxzu2ZCgkCA90iOnJgXcRRrzow7Ejw9mN/oCy1+UTuQBCOfTuD
0FgY1pS8Y9Yqg82784gQqH9HdjfiIyREN48Sq3ox6ca/vWzo6gFgeGUSDrizNQP658PN0OAnE5LW
7/xRxy21kMbH/X935GK2cJRV6/U2Y0/g2znTJCo6N6Lh0Af33y2UDhiHypJZ+pnXgQCgl1dtI+hY
wul2Kvoz9Nrq8c0UPb4UfhMD4M888ECyVnEsCT40tKmwk82StEHz/9Udz1B5/iKS4Dcz2CHPI/Lv
YdsWxlG8+9cVekt3eDG/wNEEbtywgSJgnHngAvXOZ9+CtmProgb9oFRT5Aqny/E/63F0oGJwcE64
MWAlhbPROtfq/L1qmUu/H1AN1BX/1/ZCDJzT2KrDd5fzrP7ecVLrgCEXTp5WTQls7v3ogLAJoDn2
fFmO+/Ni3H2tZEJ89v7LhWJt8+WgAfmjX8gajOj3m5Rv6O6TUKdY35Bmjx/WR81NN7aDirJ5lgFT
791GliBHrgwJKLwc13ZtWzN5tUDvHJBCs00h/YFj5F6QVTnJ8wdQWiIcRduUCddlQJARgy1wmDXG
yfPjFWKwYzrEGTPRX5UgRfOYz6JUHSUPZoG+XW24SU336tXL7HANzHvXEZ5RQUB7cLMbaB3SIr58
72fNynG+9OFXlnIlALG95IFBwPkErKqOYgvF8qGklLqPODyVLP02C5+n4zTm9q2KYNUiz6RT5EvT
D+53OTgNJAiaRRGeO3DKdMNRJEOHtGECy2907EaxC6BflEKPLnfvsX1Tn+hhQvL1tSEmsdB9XcIZ
AY8j8YryI4AQDjZoq7VHk0aKSdo44Kt8kJ7vV36m8MBJC5XWs1JOFFP2mV57zRNUhS5hLEUTtl91
rBDSYzWDi7OROVZCVJkfhOCxxP3Y+8uTt9kzJd3w5LUamW4JOW3CMrb3Qis1QtHQeRPCaQEUO2VN
WzNtUe/tG4KAP5AV3ARwdfoQ3d21EmnrFlIqGHZQ12UkEES5PiyzpsgFpa0t2QXLC03RTWB7Uo2G
XNJiDNlbHHby9mZnTU4IUzC51wX38JXZkHbanmTAlUbN6G2JfG2jbwzs4Jkv2Li6IaK27egqg8XV
9NViGJNTyGOYY1D0b86CtF0eao64QFKbzyxBwKGKOdQLdhXdTDrvOx+2YNDjusXaPfHOKl9hpAY+
ew4Th3p8HJCZEF3gCxYPmr7MafQ4IYqJqXFspsn3MFWoT7dnZIoFpmyTUNH8dfEL5FjNdNGds0Wj
AspSUvzMrTlXIPCvHKT3TpJgesWoVCn9VSkCjWDjZf2NhL8utLiGyTg7J21K0TMltDhGUp40/2qE
3a+YK6K42I4PlXo2mJC8FZ1BMZLLb0YPYEDNzo1j56Q49dxCV6dQE+MiZNgnyWUpmXEYKtmxGVIs
Qt/aP8sFy3Qrr811CHx8CuPJiC92/HncMr3ZeUhAhfu3jn+c0OLX1i5bxlr10lNYu/DZ6UugHG1i
nX1dzqRxHt3wKnKeaPl2zqFMgZzgkXTF3+Vdyr385DsMwz2tgqAbMDNwZb9Vjz7kHpN7HR4nd9pP
N/OdCKVq4lGCXO2N3HdXcO4OZ/CjcibW5spXnW9+4dPOW5FFMndocj6tJpm1Bnzbtqy7T2N0Cwsp
P0KR+u9NSasq4Rby62o9ww6WbCI9QfeBTvkCKBzJKA0jO8LoRSQZ4zJ8mMT4GMgH3tLJ3+FZUgq7
Ji0DztvegftAfDrRizO54qI86p2JH5SvNGmAcKHXi70h+ZnY+XOpj8KZtBYCg5FHABAGFfGrzy0U
rBoeiSx4bGW6VtHo2jPjlW7O75eFlNmedYOTEJO369XwIQoi5lWz80itAchQjCP1EB8tWDNzFRzO
lVEe8ezP8Px/P9DfOnyj3GxDon7q3GWrYl82u2gHggLyNhS4s1u8xtYMBdyS7VGuJBnvHZA9ecNB
G8OdLAGZm6FnfSNCvuhKM6SDHdlzZ6N+hAAB4zqwSwHdy85FVNQ5I9puZW1FGXC+W5fLudkS++1D
29ObinfznNNNrfTCDFxrJxg+CTy+N6YhpQ5yHPq6BSdWky6JBbsJCHUOwcdR9dV0uX0SKHd5sFgk
1WY3w9/PT+Eo2rznhp+hNl5ENqUzIdtZ+fkLToWzsSz/nUVB+F7QE0akU0EPpcs60tlaf6IhCCZv
p9bfBZ1uComMD+S2lPQhPK+1iU/xcgKzjsQ5Alx+UI0qV9akaWowhNqDGPb7Pu1/K/+GKdi6a48t
DY9fnzwS9tlrntYNkFulfSYho0oidKqAEXI/h9+sjYWSDUouV05UZa6xSVjZqc6QhR20OGvzx97A
Ze6J21pxRvASeNJNn5h4KyWMLuyRpgSzajCmxrclf6uA63BvjaW7+qqTrc7g3xE0P+FanQV8UM0h
J/f6MP/JL8aIPpY0n+G3Ut5IVI1USKgx63Jn2lsn5I5JEOp9ForfrKkHxmTvlT3v3PNUKnSxpAZv
w3CcDUqNf7VbXWrOi76TTUKlpui3oBQMJBeHEI74lPNuOrtbE56+UaUZAbh5Iz/OB+kGw6xq32aX
ZClhEfvMIzJlEOlkT+F7s1KcqdDHNohxnNksGtrseqLfKsnywk82UAc72wbQuoqS1O8827y7Bq4i
9RmeF0y7HL0pQ8oqcqSiRndx4sTvnVwzriN9SnpusAHL9soGEJ4jIFNjI6/kInzQvHGcmN2c1mHV
HuZ+54gHTqDsBoixqwSnPI79kIfoc80ScgoVWtDHXT1LazvX0OjLPKZJ1ERl9Xb/+wRDaHwDrOln
C0C/rQu75fJTKGfdd7dUf869ys6m/y0vutTLV19TEqBkwotbuUNfA3u9ETIRrm56t4YYZB2pYIJh
KCk6NmVj/XOPcYIQgOFXE/aT8Vpi+KcRRh0ijAp8Y2aeWXkXENC/epRzj4kv22+arUcVqy9RVbQt
e0RbyqXLkCqIqHC3dLBh9H3aVrdBaijk0cCGfXG0eRosPs/s35Omp/HvrMFdY83luBVJxgbbz6m2
UA8Z84EhwQ6iCrEef6Fm2CIv3gUee0qM9QcbJA0q9wy9nEaQ4rpm0PKXfoa06VU0Lm7w9D/Ei2Kp
dGz1mktIZ/qYKgmhC7oyhmZPtt76q1c9rsTxVJOV6sv13in5AaBrXZpuo9xwrkpnKa4sxwq1faQk
ajNYAbSRsZf4TCS4kOv6wztEBsavIW8GlBouXo/ISZuHzpW6ju+UAlxEZMrtvBQ25p51+B/aaNyb
YMRUpwVisCMn8BOGJgnUBxADnDGVxXEOQ8iVbTbq5YODw+cGiXd1SmwuyhCJELK5IS3hUw/4HnYk
Pg3AiMxgKKQQv5/WxDL5EvaELNWv35CCOWLzVH/M4uVc6zbrGW7xKhGQhH8d2Z0AWHygA0v+m5Mx
rYysOYNYYtqzafSmEGnTfNyebLsFbvbxOc5/kP1kr69hgGxUlXL+X7WXl51fPwn3Cfiiq4H2Z//4
0XYxSdLMEORfdcqx7W3CX71EfDTB1Os8dFaMH9WH0rKCNRMTyDa9OLC+wXUdx8V3fL9Bm/TpsGIV
/gx6T7/vm+43jqI8xpJiXdbQwxDPmxUu7k0S1oXe13dmtpLVxRwxjTQt2L26zOsnkhBEOvaBL5q6
V6YXFfV6DvFbDOIISg5pKpymHliwBmdzv4niT+KeK4mGhx47eO6jXnFyRKCu3qGrA0x28TpvybJd
pYBZh6EUKvhn1Fwzvch1i6dOAAQF8rZfLLXsxJcNl62/Q3LZCbkAYW2BnoNYbO6v7lPO7Rx5E8RS
Ckzmm6HzwP915lsd12dJwtExcdI8351uRSh/F1BbekC18tTSxZJDUPvj9d7wU049iisH/fMNHPd0
llIpOUonLFWiZgaiJM3dfuTRWUqH7aSuRiJbtpQqwL4v2AgyNGtQJdjVx8vGc8XpUq75gyu3oZdH
WYWT6l3keFMxxO7INRIt3IadNlRM1zMX+ThEHTmq5tgUWwOEW6bIo+xf+/ssLF74GY2QJkRByO7C
afawT/mRwVxjujYGXOv9tLp1blDQfi4pvCO5YO/h5NUUtvsx5uMBqLcGPUrHm8tbcJsB3NsTln7k
r4OJT1HRIt0RINa+Jc1F2JTNpYSjnuqBSSal3UWh6Ioy3WJWa0WDajYboscMTnPjReUaM8B6+f9h
sVwki8rl2v9MUSVy+FowqZUTBUUrLvT7ygnp00qMxnGhKYux5TUM04js2mDJHWj2Bv4KLskPMY8y
0/b+8qqx3g/x+Gu+VVQammgADLYM+xe7zk7v668paoklltSNPSgCh4CjprXPlJ8czSN5ptAW0ZAD
XlPi5XPX8YWc3Wc60c07e5eNr07IWzejsbBZ6AVsDkQYl1LbOPqva9gyVxecQLPUYG2bkPdl9mA+
WT1btBjvbqs6SAAytb9PF/o9GJCijcIJI8exs44qn/G4Bk4qMJ+KbIXUPh8e4sF6NhGVnnoSuRMA
EwYDB2jnJOFdMwYYId9hkgkvxaq4aAHOWInGawFTEZcFSyOrfCOmzU/BnCm5lr7WUfDeOFzqqoWz
6dw/cvmIm2k39FOF9S5M4vpm30CbpnZMg+2uKyFk53iwjoZ/u4XFvKTitOwb4+wGWXQH3coPs7Yv
uLKiZTGOlrWfgfXeArzlERrsx0GpUky04mQWt0fNR+KtGMyLQ3MaxSAh4ZinWOehMpVOOzwJXzP0
C85T5qosZNz5SHhn9AsUfzd9ak+oeeBndEgyj7GveESX4O2E/+08OJipMh+reUrLh1qk7XdfmT9L
GrFwAR+OSNqPEhUab60r6GB7PKVJZHwE8agW6GMg/MuXyu251fr9zm9mF7OtqUBrPIimAZCk0sc5
X6vhwpmTkYRRaCXmF7xi/rUR+PBp22MJN02gcplMX2ZSob670SMPNy0NmBbmLvajfctfLJUZVdt3
+IeZYaVucNSJ4Cf1c+gpcrLEIKcoNRnQVndU/ck+vFhCSy+7UBrV1U7EBPT4UFtRiFn7inLNQye/
2mjXJWoM5xmVcPpgx9XEsE0PoIxQFVUTsyijULRzvAFvTEzwJZySQ3qVEas3KZKYEHu4XvNZiq88
QKQTeFYqT5bFsKvh7DIP/gEaUMxVXDunklf3sewagiJ4VLne3K6J6Vkv48SR08Ezi/UbGnrZ20mv
PNvM+zeLix/eONDSa5vwxum9f+w/NsTi9ydPHdMU6tkAvrXxY/pCDzdmY+fO/Pyou7H97MvCzhG/
5n62No1062KSzbtIRWH/L+44oHpUQk02hTVEBiFYTtx4q9NyWbG27N8j7ty6WuVgeGCnt6iBuXKS
JSP19l0lVYMyerZlYJGlPMED0bGeUKe1+lc1LGcaL4et50/3AaRmlYa0NtoUPH9Yq1BGqYbpMl3e
s+3mTTCy9UAB/va6oAz5qz4R0la9eS7hJF6SsqC2NXDnFFpFDvKg2iXr8ma5rRJYoPiFARM/fz68
j9UD8L2uZjYWYR+92GTfhCb5mN9AchPVtkx7TgGeuuPqUFJbAf/UiE1D7l+aBmfjA77k1oUbwrGL
7MgYzmQ54KTdklDDNmU69DsAZm28ha3wXqF/3fildy4Voie2WzfvVI7BqLcwpmz27BtOTmNEw7bj
eVR7iGUjg6Fs1fnkN6ls+e9B5NBbQhX0yVhqV12oyB7nBTq45aAyCCpi/yZznTJ1DhJiyzWk3BQw
O3u7Cmcj9R1UTFTY2/6/B2q+v0JK0vg/x21w0fT3+m1QoshYOlALmfqhgDsyM2wUiO58uZnespZA
IgmtcqlKkJGf8bAx1poUZY4q2p5nKHg2o4wOC4/kgoO1ZXdjhocjTsY3m2agRvflvtWh/Nparw9n
88GzH8jFyiD1JkWVIY2vurxDTg8ehG4elF3RqpjhU0gmW9+x+HlKdHPOWSy2co4Vhg0ycn1C7JGe
e4bY0dyuKBWnHQTxMeruTzfjNA1Cx4KmiSfzdDaNK7kMOzcAgzhME8nM7PQw4FCgztStMrXWSv/6
cW+nKvTUjJER7N77IE3hfYGEqJs1dIneYM46JlzJgOQfjVh/40rnq4g06bWXHXC1zMn37f5c3p7z
yy3Z4/jmI9CGscgTlGBW99N9oVxCsWgVXQGWDeZNmPoJovemynkLye2ro912a9vrPEoe3dC1MQaG
VFkiCtFFQ9SL9tH9ZJQI5dG6KNApxmjbqeUL8Cz6FszF9beZLkgaoYKqwcKtOVaeX9lV4OpzK1uc
tOO3j74Egxx1IEGvZJ+nc0WO557AQmC61IJiaz8K0R8JsuXEUZvyO8ksY6PceefnpoPU70d+Oq8c
BPc72eJPGe4I2RQbztioJv4bz9w+hiHU0aksurzmlUKc8MQcpyCpvtY33q8+aD9PB0AWbWuSnLzj
9py28CzjJnJ2C2WAhjY8orgSb3Bg5esXtbul4H9pvn7u41/8Q3jqP+vNTeov8xZ9VM/rWs/7qZVY
Geccev9A/6cr2phOcvh33SHQ/qchDSmaXsyFjWJ2GomdZXZwHWejrmex/O7FQoR/7qCS+DihPavZ
Wn9p6KN+GuDLdVNbt7dE7GoNMYgf1LS5hvl+q8Tw8+vGQX9aUtwV3ley2CbSqYBZi5xQYFwZq0MG
Luk+0T3BNy4gELUpkTw1HzPYVETWSZhUmrg7edpFl2AWbL1A+4aRulDy+MCzy5EtiZOdeNsfshWL
qCBmp7dbs2Uu7Xmq2+p/Z1kRBQq3TKY8nKrdrDjtQKPBoSYFS6vhBiGUWVpSt0EV4CwiIu54NwuQ
o6ma6DM/BOKNTbjDd6uDMxZfeDDKf41xIop5X0doCtDdAwuY3Wk4Jr7KvjtrA7xzngafvFOBLm/J
KbHmxbAmQFfpRHtqnlFkwAuvOJ4KlWFGvgcoPtpiVh9xDrzLzWGtIOmr24qgUKnkfm0BBmF9R5OP
QWt3Oqi4Tl8jRihGyOhUmHqOgfKsb3NbYn+3uy8Cp54Oc2HUYIObnkJhAse13I8x+hFX/UJHzLus
vcNtVKR5f284HyTduzRF2NtaEgTFjsTNn6Jv2v5EwZFDrcZSAVaIS1SP5/A0vrrSytH0MnipADLh
yziMLw3Cksm4gUhsOxz4ivhr6RWHXKR2/WvxNaSm9pbucJGYj84bRinZ+onTiunX6QMbJZRW8IYC
wvjPjb+KWjNyrulmZIJeo9jFrShSO4bewibUcvirXy760MqtTebUgJ+mWoes9XtHveOu5fsIp8t9
CcWbyb82DrSJglxFpQvNgXF5axrraHVO0YuPaTNc0FBtaC7ZArFLg7Je0z+/Uq3UHCsrjdEyyt4+
s906zYA3w+VWEiT7OVoHjT2Zl4+foXOd6nn0O4wDTp6TtHzgMZZcmsYEUF1E21cdJvEen8TmzVYR
Va6qIRrbYpqDidhrVcWFaUV2NfOl1Wtno0Ua59TE4mCCwdHRz65NqM9q9MqJ0Lg1jzoigJmnxBZY
u+egeDfvtA/Ng6xO0rt3gXgqjWLUBHrB0paDspAqmk7C8fmgBgjzwe0lRGXK09JOhNQEMVbSewEX
OSqTv1Imt2W/E/LvIOsOx4Xn+kw9KQcpLcrNJj56EFVggbZ8ZZtjopFpnzb41hI7ttxw7MuUsUQW
mJPo8D2rQ8jiaLpYbN808gPz0sayw/eNNjJ/lOtrgz4IEsk+8bV+wlFQzeIizeYhqEdLyPpZsx6I
ROG71g0RDDZH9+m1qa799X3w3vq5eZ0O4PUWNq/q9ZsTtIRPdJhiNH0fzNWoPafsELQVLhHLuBu6
qBf1pkhQnSVBznjMoLM90E55TH/3SvCjQmVFwEOOGxxecmhmm0KNOnpcaon2Y2upPtDSYsqi22qG
U2I7dKwg65rs8uSU62nnG8yytNZTUSMDbNGDoXqx5/iNehL9DMXC1L1t6tdUuq1MmFuJd/u892BO
OgWrJ/PaTm1P/1YlCYf9MBIU1H+PSqOa7Sy9u9qD4ZCi/T6pGN9CQenyHCc505ynAIvMJYXdFlcd
ugkqICAtF83q5z1oOvEMjpZSOvkJd9Uwdy+Z0GVjxLxQYfCMQvvaxT6iL2dw0Bz2mnZncXw+PEwl
tSSMdbFlA/UV7xAXehVscnYiLC2Nz8EXPNokTmS0D/q1YwsQD5zFrorIsh3Z2ObkGvWCTs4Ipwhe
3qDl/kqbWEE0tq0A2r9+h7ub74T9wxlpyr0oGJUixLtglaQ9tGPNJPiWyEm9WVR02eJWKR7p9M6b
JjoLWzbTqFSYQOHrvx5TkWGYY+1pc74aXmSdowqV1MKvE6qfJxsl01wUjjNpRlElbra7fc/s/R2k
C1bmv1fea/OU4cJlpPmVNUf+3npSXBj9vSnUcuOva/F5n6QpMI6n+z7E6C/wV4N6evGoYT/4f6aj
qKIvcoV6PnK2DA8Ww+gpRyWWs7yq5DOxxwesPLLPoskTE3kQ+sVUrRvneXi5dXUJRWU9/Lt+yz5A
CC+bNEBuVHIUMczFwJt/5POYiXkduX9l7EuzmJFSwTg4uIrh/EbFEk8ulpZSJYQPM0GxZzgACOHa
HXTe6/ZsDpptN6U5qUa89duKD8Jxm/ntpW+iyAQdiWJ394WjfcYSsp3sBIqRrtRhKSan2xDsUGFC
LnNARVrQoDh+iy5eE2V1dgMnbkPJY0DFVadphTLgNtAzbIHeXuWLf0X2m9YHPUPJL6lmSffodPtg
SF97kdQkY+T0k+OORYW60mrkxW0GKjyXLFKfdbeeZ+Fl1nnJcUSIrvbRWNF5GMOvjdHcxxv5Y2x9
6ilesWFEhKbNYV/1pokQ38IIkOeuGJxMEZOZtkz2b5QEFP5f9L5dQ3YWS7/ATaPQTHsYBaoxHez/
CZdtNu9oY5NAufxLALVbh0q6DBK2iZ64VgTw44G5DYLpmtP5P9O+13fq99vw/i8q2ZRy5pa2aGfa
GtZV0DA8lfDOwbfoY0GgRwQvPmCiCxInF6VZJCnp7zGb8ff0sj4DqMIJNRtjsSPfd9jDw0Rbor61
GaDYGZ8nYAoSUqL0B++DHruZm1grLVlLg4OacyuawStd7QTt9s6VM4+Fi9RuEzcJ6nvSB5KjuucQ
Kl2WKHcOAzxCq7u3hFDJEbMARac4CyViIn44PNvF6Hji8RXL3S2thSif5DlJFlxzfv3H81JbiEr+
SGRWyvcdoOiwdNNGIY2oxilFI4oINj6aONAAOWz03K6AMVz44zMl61AK4JlkWYAieDf5TUZ3UQuf
tk9CPTjY+noeUKB7j1zTZaiOKL1EvQR5rPYktnBvpo0dqrkbISbuObQDZwUHuX6bHDyRyW92fRYZ
42V+b/whBOfe2IaTD8fhH4fFk0RySJyQDlKi8fjSifilqYevulCUfLjVZSV+dij/7s4FPOzHRUXl
kbWWm0gdu/D7F6Lop4DB+4xf3/RwBtkTTBpH7HTVKNHg3cK0yLogtPwZuOtWtg+hC2TEpK+rFGFa
NutXN1q9QD4XJzKJLeVaHWAeX1viujG122ae9GQtk7VsVt7thjjTKkf0dHNxU60jT4otuTBAkcxt
/LVd8ezVJecCtZVanRrkULPC6S+2OxGg5vqCE4keNWKGDOeb195kx4nq0jwQ4uLHZDClV7bLMKyP
qg43IIYBQo2L4lzKcKc4UR9hR9XFe3NjHVRRXZoaOq4KyHjABaGbIMKAH9t8C9j59QgSgIE0Jcvd
kUA+QCMCdiv6RaTJJLRm9i6/DIp0gvcMBtp/HR8crQUf6X71gYRLki1ExMIXJpWLbsduba6HwFgW
yyhiMldM835vOTyLIDLUaiGL9pqaUjxurhjc2cSuwCVtT05gSwLvmbuSFpt/e/v6ifAXFo4cK9TR
Re+rkpNXhslCzoa8A3V8G8vPTrHcQIQcrTtYbIfNnZgXx8qnP8EmqBhXbwaq0qqrQpF+63Y1whDu
yAmjZP1n+jd/+fmVpl8o9JbPwbfDdUCU6Tic3lYCMnbBxGu6oRRmmqfxH/R1uxbhkQufIxYCRBsd
Py6NLvLYWO11IXErs9od/jxEe3RvUzxP1oewQnnOfiQlEdH8PE45QhTOLfsqDhEo9R2kOmnbwzva
9R+klOAz+3Iwlm6iG7w0ENSUVhhlKCK0IS+dYxtyvpmbQqVSuyyYK5beIbSXQbeRPaM80+girAgy
YOnZbNhZKOZIKEzXoDCGhkc/TjG+cUxP6GC/DdAjA/jSjkamabdYyeMwavb0xwAqRhjTsn8jQzVS
rm7KxzdTdHyGz7Jf0qxKfQ2nu3ddsmYEpfmXOqdy+fXMG5J8yTIOjmIGBgQvIuutYc/8XGjyL2qP
giKoFml2opch19HKoHpBQH+5aRwDiiyKniLBIuy51FRXzuFAsHzjpSMzWNjiT5Qtgm+6JAEti7Es
aTAUglafUgg0lbqgZxu+rG05Bjf+f6Jnt8vfwQuIDco7LhIKYMaFhPiTI4pJ8MySCza9IRZOTV+T
CSHa7+nwdT4lB68M1mWh7jJ/FzFGeBFW1wkaWt6LP7fMV/ygzmTIRvjXBd3fPC3lvuzSQw3DpuG4
K6vZa2GnA3in/SUIH2owDs1Qkb4PgLx2rWodT1EQys8Ew2EiAenDwY+1cXbO4wmlxQV7Ac5jyqfG
nTJ5gGrtlIORSq4q3/i7mSsSuTW9AtT2NJGHMVDVdBHj5GrzIVLLlUtVNoraYXjbRpPpB3FKtpgD
uglMSQJF912A+l/lnb0+AwofjNh8JXaVfBPXull5CQnEhNtP0gUEmvMa+xcgW6a5fu/Qe1e5daWO
ycuLf6YHfR8P379JoeGV6GwK+Y66FxgiizY7qgvVFAtRtQca9R3rbxG7F2tLzhhWJFK4Rytyv2IR
g3xY2Wk7bv8swVfsZI69fk5qwyxjH8qiumF0sBoNGcHugZVFh6LeoX7ICLmMwzfmzDKbh3LW7wwJ
YC6b6fVKqBM/SC/H8CR04QBoQba6CHazYAJ3Ljvqp1w/tN5AMSyDOrUfkZPb0YBH8ZoTFAAV5iBW
ALgRV7UAP6Ha7zYC5MC3C3DxTWE31phitR4PuGqlf4RjXqtwRSCeWWcTaJlVLCSuEUdP2bUGH6c2
6mcWSkxrP7+d3ILHnWsIcwawmE2joNQ8Hv12dt40Dp7mXOLcoU+aaDA4UYZN8Lg3KAigYqNEbfF4
pIItuOH+Cmm7+Q4DDdQaDoQmwm1ZyPC6m+YddyZAnWYbVXsnk8mShzjiMXvBACqLkGNJIMRVucFU
03eFCRu9lzhXgrRVDp+jQ2nP67WVlnCgErEYV+pyGrOG3QcCawOZealljXc3DsLJao/lXzTuYAdJ
pHhWh7vuM7YVpIPFa/ilKcPIKchvZZowpmO1WbAs3NrGdNIuzWWVU1qlUDjOuOJG8O3KlXdHjY5D
ocl6chNlVlsHgAN7t8pOOFjmb4m9XqDL5ybSjHmJ9reGRWgzspyZuFWlC+0D2EX1lGEsEzXjgRg4
IGDGtoAyO7J6pDLbopwx/TKJfLGIdAfq54OoKgJyoPfEydHFbPKMthU1qRxaEboOcqneEOtufIF1
712edpy79zu/VHTkyJ9ZC/f8pqIo8VW9rkX6NqbIdfBXa8yEqiUua6nhPsTV+lVhy0nTWia9TTH8
VeyzRNymXQSIlzAKAWYawvV/jVcXn6EuLZse39KvekLyZ33d16AlTR9ZPZhgTjc3NgmBqdgc5gsY
HDNqqxjTytO6r2haaPxyHOqQah1PY3Kkilg4So28oVEmFC9OVB8L//55hTazGIKIdUXhnoALwFwY
2Y6wKyFRsFyHbO7bdjMZzoH+Gok/uL7waVgpmhOkQlwgpAByJvbUpYTMLKcGlUdII/cDfI9dXOKv
mcGYdZXP2vhZKCRAQ8y3iSRL/miUAfeCbOVd1x3pArb4W16CB2cWSs4skgKq9Kvo36+ddHIWCCmY
MkYx3uUBLC4zyCNgmGyq2yEJW86641cG6UtMVoBit8ImYz0eRYeJS8rNdVVgFNiVjkVEUIlVP77I
PkAwK+stdJGZ3UkYyJyZyISf/fxf/gb7Mih+2JRNLUdPEfguzb5J/5NyMvO3z/CFQe+gSNNbBDbV
VKEEKnPyw5gAua+K6Ll5/FRQ+t1oQlJEk08T0wA7OyRR1H/pWJjEhg5Y7hr9iP6292SqPaklKHxz
ugO4+5H5bcrYu9HpFrZD2E+3Dmb4VF5NXQ4gv2mslhaIoLvD3t7hWRa5ozYsUPZeo0G2b/3eIfhS
l2jrccyoRG2KWMR+ZqClH0kWkJS3W2rcga/MoRCk4ub+2hcbTd8m5qGZAvHCDUGixGmsneRE7T19
BAfTiRY+J6Wqylp2opKXUYiL+dbNBDAw6jaLnJnaYUOmwEHI8ewY1qC3jWxePU8ID+wRBrZBtwam
ydYy14402MeCgqvsftScxMD5/+8WtZtOkw8Th8qReTKDOql7/uH9YVeKxNgaG30uL9trkK8JYMdC
OUD0+NmaIqiQKEVd8x6Snd5s/ZgcBAbAINBcos0vbJokqlaOFMUrRmYoIPbuBZqMe2eOejxov/5Z
4ZBsozMFZtPYNm0nKjnxwp8lv6vStU6Lq5uPjJ7eH4komfuWSFbMPui0oYtcwiCQzs7F2NAg8v3F
eLLHtl9SlDLRGzfKqq6Y2CpV7DYGIrEgTIdrUsyZEm70aF/q9jqMp9u/MWoUlWDQ/pJr0zH8LWBZ
Jtk50ZiiKXvU/AnWR0PriqZwWRWFZzOsidKPDC3NAWhmBhMRhrdzUwMMMZYbBak2yetAisigwvHq
HP2hWlNsVqzL2UqYrG82uBcSYte5R11QHKyMXVzKe8yTwkqcQ+DGqtEEhSH+t31+h+uKtNaLcD3a
Vj2VxmSppgWstN/pKkaFdnImdmIIMJtkl4J/ndRMB2UZO/3hr1rF8lnDB7HDQHcXF5vgmgTOd4oT
0MzGsgeFWYpgQdYmhH9d8CmzAczSLw0sCriMjCRYQM9FQ0NoGJ38hFIJcCIeUyLFxZP9cOU5P/mF
8ZHhcQYHzXH2sOakKKu8tnnFrVtNTwTL5JmCZCUs/w0dic+86RCTYVcQTPfFbal6NKMnmbvS79ec
uJ9eQdYNyS/1A7/CRfyllzyjyPv5TmbtSDtTjg0IttPdJcTlFh+hFSunf1Xib/OzbV6tHn1MOsAl
gm5VyoDIuxvGBqqcWP/H3JJl2WBTg+QIWGXvDHn5PKMKdVmIlpftjXllbiqBJcEzMWJ6x8A5VPV/
MyuEeSKpySgT03Hef5zf8BQnH35p4dW+A7ptlYH2GwqtRA2EyYhXfa8xztv/KjhTnjhWwNP1DuWa
zbWT4P9bYCjz7mnN/7RZpPPvV84wsGJmCiqHtxOqC2m5M27/m36FHXSMoyflLMys13jDNm8rSHFE
fQwM2z2x+DLXDPyO9nl/KI8tuMQmSEvrv7xMYQtfrJEK8I+P5UGOsVSLjLLYT4oAVfvuQRiNzFUY
PUantkDQibaAajYlT4DZ8A48vLlfmGXEnCo7pkZqcIInBWpATXEdLl3lvwoDcvJT1C5rEJw7qNwK
D/+8i8aMWkwgkq7vYCXVqdKKHjfQwrJ7jWlh1y4lGVJFfXFjTvRHByCwJOJcqvj5iIZsI1MHhYqh
sQKugUgEcfAL2UjrRj+XABRmt9F47qSxVicPtbx49yeqSfWZv1JAV2VWa+TlLvAZoBIldJkBLoYw
C0b/Uuri69QqBXjqxAK2TsqJsGRZ7W+pdgi0Ws3KgAy1429sa20XFkhkDehUEVxGciqDPXFYJ21N
tlNF1acjWAYbWTuckNxQoP5jicQFb9sgDAaChaO+IAPRK5Ld6M4CaU/01UQ9zRYnleSUKMUbbu60
AwtxRPbs1zQRyqf7Q9W4HEJHrxB/OECobLIqTxR2F4Pmzrk9HjQSbJSM2RIF07yA7bK9y/JWjOTr
g3b7Wb3n4IZ0aK9aqKvnMvNSEu3Vr/AwUtjq9o6m3yYUhigfImPjTwyaplXlxYUplUcyOa5SfX5r
fo2LzOVUpYRvVecmB5L103rN2/BuVjbRIo5GzO1MensD5UcoWAtbA4znUphUfVIdvU8pWRVHBhM6
hRtnNxD1zvGYuBSeTn5VxplXI5p/6Qk/cP8pt2SfcL9hdj5v9vKjOCBJ9KSLiEVzR2jZq+8fttuR
KFr1FsVIweBqbqLaGjklJAGC3GoPQXSqDkcMgQduRjnRq8vyjiNgimAjEke9L2FxtEGZGujAazze
KBnVusQ4YoWNyrxuETc65fFxRlkvu3tdebPtNvlPS/nAtqu/7PhmtV7Ci4gIwbM+X3J8DkLwEKau
YxAPdZ1throHJ+5+1vOokxXSmVnMrXb124GSBIGqtpxm0+BzwE2f45ga9tZxgaQih3Ppj1jiPntL
thHiapSObBxyrFrIJwE/Enwfp2tnjG6bTM8AeNL2f7GTCIgBXSOKLUdBG+eXl1CaUxQtYjOvu5fP
QgvsuI0yopl2IRyIh7xEKrimaOzn/wwCexKmpcaTSZVhtaLziuACI4xp7PbCU3pckICneBl/z7rx
X4b2PhDzKXdazVUc0o3wnDTgTdcBFuehaGic3nUbhfF4fZ9LHNMNRd3zKfzD/s3Ycpq7X09973V1
SDL8pBfDeakpTJn3wWrtPQiZ/g620n2DSvBg/IESfEHeFtXtuVz/uhYOvlDydDAsRPOj2j70Fbsq
azo3QGTp0oDmT85B0O5yoBsHYNoPDCadCuNtnV2BWFEzxgg+gND3AtenKaIJPh0m6RhIWpIRSH/e
cPAwmKbF8Xe1SdFVoY04zVBiVGIS9pfLzRWuHXuaVA4OFQZC2HgcSI2YoW7m0ND8sa/SOHIloVy2
6caFEQ6weiL7ormC9GGrx6l38FOmO3e0Q8DIlPGaEOVYA0Y+sAeHCj30x81qJd4vhwsWG4O+Ok7O
8kSP+nXNzw5Jm+521Ivu5e7pniga5fYKhAcRKSEYoXk09JK60LqeGTrd19LkqU2tgNBx26dyXGk9
Ih1pGRtWTcGrCcxV1Xyk4pOu9PXJYumbkZi85biucREPYwMWTQf58OlvwxIhURkWlnu3/1iH+PWC
DFBi5Rb6tC1xWVRcIcdJcp8rXonwIGGJNTP68jMR+YSBAsHjvStmZkGNx84nih4krLHj+oRMSxLK
joQ9S2XJYRiAuFFetHm5TQHJ4BVOQmCMtRDxEduNdlTfRP1+7A8A55gyX/NcblJpyNZUPN/QpjG7
rHKTq2EqaXumNrXr3sL2jDUa3nUlTfPDPEmw7abVoADTzdRp1pxSSo9weVFNgWC2sWxJJr53FBJi
sloSZ6ZjnCR/FM/a82c6uZNTz+hYtoUzv0xAfh/vLIZgL+5hAMyCAqRv4ZOkx/s/I4m5OvJ/mMjS
73HUhpCEgrwTKYeTI6n4ERIgAwSoMzDS2ih+Xbd/6GKrqwHj24FgNucQ3xYySOMfG5zCFN7Vy6ur
6eSNGU3h6m1NR0zDz0H21uaV7qGtERBj1L+qzsNuSGB0SQ5cL+XRGVYRUwxGtb6gzmOOj+i7MC3z
Tlfgp2rOUkSTVub+7PbNXR1Ecrldepl8DhZhs6cYUFR6QIk6lDpPLguJbsta4q7lfXUlpk3uLdGP
HUvm1rybcTb5T3coUfsnzg2XYMO9+iEQhPcT7t//qbxz0mP9UV9h5Y4D9YrPeUpLb5DYuU2WDZOw
BwlVZUx0xfu3ArUPVnkDKlbBqUll0IHU6l+YfMUInFjz5kYM68yd4RGdUV84wnaydqa9084gBUq6
jKav8LRMyQnfWzvwdZBrl6IaVGsksqHifHqlnX0AR6q6cmlW+fLlGpMVkFbAUPDwgOzhzKVDKf3N
xuVxM1RMAI0ePIQ31VOdqhMt0XEzx+aMtfdNV19XD66XK3YjhYPqdgEMfP/PTtqmiScV4S4wp3jx
W+P8f8+AuHuR7Ig0UPnKHpd2LOK82BnmJn5y/kGPYhAjio944nnTDIIgxbvHkHLjBaOhJ3axgG/M
AAX37CH2eE7Ksoi3QUt21T4N40VvF+bGn/8TeS20Cb1ankFdwQOMUhXyJpLmrIUDNhc3682yuJ0D
1+btq1ypK78LEHFSOHQh11y2t46UJBxcKtKTJjISQfVtCU3QOXPBPJBXfwuxC7M36YWcsDuQ3T+Q
zskJUnnkLLs89pIWu6aiXLp4QaIynvOTLvGy/b6gCirkrarw3BntqFPFKVU8AMcjlf8qdArO+2Dl
OzcJiRQXxVlO2iZsso0ccuX+IZUp8iG5Ijz8n94HFmdNCLDXI5qB61ULUJ1Ypi75z8SVII3O+pBR
BvKRCV7NAd3qtpcOQRXqkmHDWuwRw0NpfnqDPrUPqJccP72Xth3BPZySGWIoLM6pSBN2KQN2R4vb
BM8NLTCkaVPw15MoDRdSyCk2u3zIIQHW8D+K3anB7/vBEflR+hTaNzlW2KY/AlXG4nnkuO5HwAms
AmdbyLPDTBkDrXiwUf8pe/+BG3AANTvzuGZb85M/q+2759qcBBnpkwMzH+3Z7LIVGm5bVf7mtDUV
sH9+2/5jkpbZUV5Ux+OCjh90wxJ7fh5p03YrcKok5QIe4R5H2t1vWIYJxjAKJmPX/7FQ/B2PwNcm
XI3ue044gf0/0ihdDIrGXhpyn9Vorj1EqrdmKP4fawsoY96woIeUEBQEHOHA6NJ7FI+tInaHYDlH
sId1zNe8DnQ1uOG61OjcTyyX9TFUIyweiSe80lH/hFaQrDQHCQ4mBPvPQUMdX170dU2y2T/p2lyN
tnsn6dIxRDu19jfi/S7rwRdzsaDl19B/zA/g5TkAWEINBIaiX9BDBTI9TCz66MCwp6/usvYnsM+P
0ZryuCANw2yn1WHGXjQM3iaF8I3+zZ6qKe+WEU/ldXyoYAqucMpG6JlH78Aw3ho+seHT/YnKADVh
ONbVza+738NKEg+u54uz31HLEm00Z4jvKC4qd7DV9Q6+TEeQdtxHRKMy6iHjerqigx5zO4X3iliO
NfxfOLVLmPX5S7X+HrGMCl1+71cKOPJAyF9eFeIXspivHfmaqQdSk5KfmT2uFd961nxDIQacxBd9
P9/gotS3DM4OgVd0glQGNGhu88+lBy9fDShWY8v4M7SYwDx+7DwRgZmilEdd8gFcwmJbaTiZNwuv
uvuBmao8Gc+5CZTl2SDEdp3zerU5fytiDuiVQBYxG6Ep+T8ZI/yyBCtZbYhpbnV6hrNQwZGRqvpO
Vy+NQcA1FZhVvpbu1PXeOL93HKpnLRcQxCPCqBasXMD4c6sR8aIdTzHaV5tfyB1NWWdIG7qpup6m
Pl3h8EoM0jw72T6nMZLQlMfR/X5+vWKZXSYfzVf/pTTNGKJjHndVHLJ3bCUbWqDhxb4Gru+aCLYB
y99DESQur5TQUoSGj8LioX/tpbqOvCvd2r+ijhzdXR4db+RVRJtOCDOlxEw7+IWOFzPKEULPrUK0
d3nPbt3C1TpWqS1J3aI0WT/bTTZORKIGRXPGjYRy9axZNUSBBn8JKAMJslPai234KuTAxvKJkhI0
9Wg+1MnV0n62L4rsrSkr7MfiQhoB5lBv/+n6moy3dureMvvCdUjLPP2BNwR3/cxU8dk4ARuozL13
G5VSHCgO8JYqN5IlqqgJB1W8eMDb6hFI4BEwS10bG28yytMCM6dcSJv8d2Z4U6MoZwR69oCywyFN
85lGy0u2YGISsBE/oy44DYp/5pmSueg8GuDa+J/l5UJ4RjJoxaQfvG1ceOWFTTsiYIvJgXqqa8vc
XHYmpSQXskpzqS9obP1YRK4+WSp0PztRjswRtVt4PVHczdPZNbvGA22Gy2YymRNrwVksyPOWdDjz
MdDnXNVrVTc+N7r8pDO/X135ANQyNLvAGqdxj91vBlCrwm0ytKe2+/oR2VhLZxc6FRVGhtZ/tb4N
3kCwVhBh9pFHsZlKWakuda/U+ZPlBmHBDmltwpDzSOcFIywb5DDPPSQdmc7Caih9J9jYtZDEico7
AZI7QL7XO7iG02ZiyauiSV/s0wtiRHCMUoH71S6pPx1UAVPI/tA1MpVyTewsgUrKUzL3cexKvs0G
BMSoDafAiBxzjIpNYqwCf3l3KPci+3CxobESQkfZGlw0rTPgT2nI8C0vRXPZxoeb+4pf2CUzIp83
G+vh5tLTCHNloYq/fInRz9YnzwCcek3YXtLBleyI3vgxoXTnsfIr9YSw/FU4WImAsEDIik+xNYq2
Y5Jyf/4MM5Sv7TtBhO3vCqj7etFlkpKyRwzio1pXHR4xyS5dQMk1TRtRVZsi7qlSbT61He7n8VgK
Ma69b+R6s2lHeZfnH+tIFhkJKM95Vvd/jsJr6yoq2k5nBhwLDi+1uzEawgzuXAjkrLQ6E4d9a3DT
ya4gZTLm3OAYqDcB5MZgetFmg1WkqPap6cRyqOFdtd/tii4cAPdjvjIQ9WX/yhtdbQOVwMixGDiW
9L+XGCiO6287Oo+bizdYS0NALNXP7M549iljEusfXE0yh9tSgf64FO/Q2Of5ESGK8kWgsMFntlA7
iVXswmZiHwZpNdsJ9i+qfoWx68J5QSCCe0PXlfdLinPTx47xq2zhlL959HfRcZf9em2veDgVq4f+
CF2lII65Cs8Rr6gZTOLj82aKm0RaKb0R2JOhQW1lS6xsMD4N8UonSicQcNs3n5FCTdl1xIA0Its4
qdXP87NYhH+tSdEr7iCuMytKhSEdifbE1LHrL2CsUTV99bUJjAuyUsbAtAYuOSnWz2IE4RZCgu9d
KMxQil9SUtld8aK4JKQCZGF9ehHI17UpEAxd3XXgYetfX//9wMv9PVZd0L3WnRtVxwEZ2xaAC9co
KZf0ymAijDZAYgFkMVf5hIKh3zuiVtSP9H7lpSJsGThYXS86WRRwvk92v7rF+vsK9Yeg5NbR3td4
DTLXtjLQCplzqOmgZgpYx1jR2PndSGM8+BgkQ7uSRtotAjAbMGCtEPlPUwbh3+LwISlAhXcUftOO
7xDaWe3DHwHtOneMLPl0yLn22/uSp83Tu12RqncRCaVUWn3eJdiiB7m1l6y77fBfLvl6nJ09ikHx
IZ8rS8qwTBGp3zwPcsdSYPvZTN3gCkp8NcL4TuNeCnGsEiD0fw862fHrYOAtVTgPkOSsi1D72YMB
WAd2MIvuA0i1l/bb900co8LxToFw9URAgCRNsoSLncOP+7/t9Mtqd1D8ZPAkqN2SBU4iJa3cXnvR
kbtqZPZ+0V/YIqlpTYpgUXfeDzR5ezKlvafG6k+xyHBbLh9k4tvziBxbULe+/M+tUJ1kjTiiFhnd
TyDsvKhsIg9v1dw4sOcvBY4KBsGIMWAdG5DbZjYolk6Oe98boHrD7TUQ03uO8estbzRMkFfOhv/V
9G5h24LlCzIKK32rfL4LY1q00Kt42GpE4io8wU69Z1xikwigaD5Zyj/ylsdgQBDwzZlD9JvTJ9Vt
Yr8zQIml1/OJJ50aYowo0HSSWEvdDAuMHsbC2qDeLqjkSQ+FCfCdtDOTs5tXArHKCGtBwkjz/APL
rguwSXZOv+luAOmm7FylsSEyb5gCppYlRF/VAfwyqS7AsFNmK2fDxrjLDqCvcxZkVuqN2v4dEL3i
k9C3GvXsi3veY8Z5N5LFzJsIORKeeDQ8X9K1CXQGJXIpK0DEzGCgs0lGq6Ca+l/XOQj1Cii9y7cb
5h0tJmNz3URZIH/9w8qGINoblOK9uwPsnRjTUafMWZOcg40AYcUYJlTmrSVAsmbg8rtx0D2QQjbC
R4g/Aq/goGuICvsiWMrE3yDCWtCOdJGYP2PH7b3TjniHyCjgAvThLxrixIBBuAleknd18m3aKV0l
RYGYXbCiWP21Us58tvHJGx7WOhRCaw5ZXtfxP/oxwpTJMgKoCVi+5AtvJchUqIgq4IKxT2fOtu/h
ScC+RTz01aF3r2zE6O3jMpqGjBy3JOcV2sEoKHO/KKtbu//hE/iD0lFAuowQA3GMekB8ZgK0z9zt
kUFU4lsFNiiBnMWaQO0MjnOUfjZXM+O/tX6liG+RaVxttxaku3NB4FIl8Be1+hk0EedoxuWb7+R9
gBc0i6KPUm/tNB16AleZS4odPREU3UtSHRH9cFFtTj8NijvkN6bQckkuOQMBzPaJXHWA5wZNNpjm
XGyS5QNgImClhiYK7sBzVrlC/PbmNex/8Ix+Nqv//f539Z7yPwlhtrm8+ZLFHwc4nWqSQZXRYnHi
fPcFQlZuHSxYjw+UGoCJD6aV63dBxULztXwy7uZtu1wr7NLp3nTc59M8yA34WPaoiVcLy/9WXd+Z
WaK9SNLulp8F7VIW5xw2ABxVlMhI0zBgAVpVXeDO376YpK3pz1rjDREiEW/xB8gtK38VUCJNp+tO
QZWrNDauA3LIIecIAsUlDX6U/1ecbOz0BDHWpm+P4PzGwHCJ+kADh2NvVyxp45TmUIGqwh9I2V+4
tj5MuSGMOUzc2bNcCwWn3lS/xemIc1rGR/7tJL+VVQYULQSRiDOe0wGjpVUtogm/PCqSFqMKZMO8
FHVvyKoTarpZh7QNyM2dIEFvdkcbXaa0ngoni2XGqRRFjSAS6XGxu83Psy5gDNpEbjvXqeDOhbj4
GleyCi9+RG9zVD5qA4bxwN1azhkUow0UrNu/qWlLZ+K6K0Nlwwcpx/P/rz8flC7Nl35NhTnRNjPJ
s2t5FPzPwBCi4GBCkWpoiXASm5VWjSc1GyQ5S5/mLHZiFeiIV3rkddafpfnkiHxrrifbQCQWIZeI
+idoTs7Aza6AXzgk0hUYsmBC+xkB046AfA8HdDCZuP6CicRc6cWU8NJnTYxYxQBCLS5qLcgoOtk+
3OqUBqk1vv5Ed4pFuRu5gGzzLRPf2P9G4qVcBm7+Mq1LsgZ6uyd5X1M4H4MtIv23dY83/CT+WSwe
Fz0Mf+FxR7F0BVi5O7KvL6kkgwkLznS5YrXZZhoBc7VEPM49lbUyyXsDt0iP+kqUzICU2oFf7GBE
TlYiDTd5mHzqp3LChv4IZLFQdN6CPDZcT8JFi4df0NyDB6a7v7Wxht/f5BVEQtE2VSvSBLcLjebE
bDds+ArJFt+WNccw7/QG8EAAMvLwlsYb60HS4UYBKfg2oaiaLiByM7/3TDzbjCsxE8dghYIrXiH7
JOqRl1fNgMT1S+EbZqbcoUfwhV45Wb3hf58vnjEtq/B3Wu2HN1tHw7Lc3j1rR3zFMOpaDxGw1zI2
TB4wzAnvTtOPM9tsh1c+t0nrimlfj5W3A4PwX2h48sf7LzB8wHWKJQ66iEDxG69H1VQPHSqEdrz8
E0WN3IxC3NSxnJLlIKq1D9UebIBrhuS4fq2QyX0vMRT52c0ERIfS/uS1AdvHbVmwl/FgZDx4xDKI
UImzTsQn5odn80SM3HHF+7B3Y0goRRKRTmoH2UAJ4MLmtzRjjyuxl17pHAZd7yOzgnQLL26uzOAT
K6MWusyzkN2x1mff0J15tQVIYqzJX8ShDu1MIoK4hNZG5YZNDeoao/tRL13JVxMCaEKOuTDaT7TG
pgpGQEtNao8o2eGMe6mCS3ncfIm7rfTYopJRiuF6vmnP7uyWz6Iye9HkG5t+FuW4fGXl9FCalUFz
iFl/G5HzVmH0ctzROgV4y741QGFih3zQlfZHN2wng91awPGFO/55tUfqEKV3PV37hB/AGhk7EZBD
nhWguFUrX1tQETY5tauXnKPoBRKQpaoImR01EiVkb7SyPIO/qJAstaJ9rrsKj+ilFLg9+sRDfC1q
gMNULAf76rzkkaFg7USuPBQNKLexrm1Uc/EcdpRlarY9h3Wnh9FyLJgkjh4fbgYEmpzi/XsI2nZg
sWkcoK0QvqarjwCRyOFGVUjsxG7kJbtRg4qXpgURyW+qrhOUpjMziGkuQ8j+GEhUlH+m6obG3sVf
hMiFP4XhKT59BbLlRkm6Zz6foO5JkJfmY+qz2Hj+qT/hOTay+O5zQ5Y/3y7PtbJI0jGqGOC4Elca
xG1RN+HMvQS15KordCLnf69fsexo/y/Cu9u75KdijHRu3UORdU9kQyyB5o705S4u8rXVn91mEwC9
0L5bE3VVFofJtBcOLvZQivQSQGgY5nae9RaZU8WrsVvUbF7FmGfMB407ecDb7eWhFxpnXLgGkw+3
8yhs0uWKA7HWK1s3fEJVnyrOGY71Y0fqCAKDh3s2vjk7bMTpNID9TWEOOKTkkkoxnyL/k6Hi1ZzF
oDWDy3PEbIV0n8wZOu45djXcK+TIQyScU9sVPWWVFXY7GwivahI/lLbAgu7S4uZLQBlRmgv81EB/
DNhJnueeyFhgs58nqiyJf+RjfmdJcCoyrbxVfY8Vnw1xWjuO9mLdvZvEixVR1wQd9DvlhvaRrTO2
QpI35wX/l9nljd31CYPl5nyjqLHT4cqiOwg2rBLQf8/1LxWKd4F6PLsmimQ76CRndNsSBDNYH+jz
pifArMnrEcER2fnhbK9vAHq5Rkyr1qvGUXCHW1RZNvgytMS7x0ydi1qGCZ+7SzKkAyS1yKc4IYtS
33Z4+udmVtFy8YEOyrAXpfWYdNFI+kRUhLSO1an7DsaeRZEJper8QK96Sxt1ygs6jwEG2DX5Vhyo
zTL17nyPwP0eCr4PvCnNbKRHBYL9yodQ+QwFzRvTrq717er3F6Pq7uz5AGNVI9QItMvulVJCBY/8
aiYn8ddKZyFDQo9kTUfUBTaEXrM0qmztbg5D2J7Oi+AQUvnY7EDVWTj+1cW70UQcAF/4PSuWZPc3
ZeAm4zuyfTg6QRLr4e5tSbBX2M8SmVd97AWFvHlGiq5BnVnjsLaOBYjlvuv4eKuZ/1zpgWoeRPhF
bQAl0IXAdmx1+bmB9czBMQXDiHExL0g58Lyd2YdCIS31ybS7WR+6U3zeZLVcGrNetvZ/rAXPCthY
QB/8JLx1xkugJ4w/xj5LasTwLdyX7tJ7pMwYdrnlIVkiBDS1+us1dxprCpW4LJUhgVc/cskJ4jXM
qzcZIhFFno1qFMXtvBZ9/3dDtxYyVB1uBGHGdkvr3mPS9suhyAQpttp+ZeJ06/oAC1VzmD8V8kLZ
Zv40Eo1rLiKdHsBluVaDQOcGI2bx7tKNzWOhTGF0ormQFns+8JVlZ/KV3GAqFOL9C5NtQciPhaG5
DULielRL4msIFITaj4Vzn4N2D93ySufGBw4OQOECOFWNyetxvBB3IsfbG+I2NjbVUzkQNqO1x9Hi
xCJVhTwH5ZyCgJzmpeRmlfrOWHUtH2CDLbIm7MPZvwL7XDX+w08KcMCFVYO8VCP193o0ZsRGtT1v
umDDCcevF6WaKOtb0HgPOvN1XES2vq5KuatzwJyUwVdCwL3aHFlFAuekrl28jaWcC8Z+WgU7ucrD
JP0eKFjiPe6BjnNYDHWTmzkBr5bGPCcp5nfOKXQ+W+BPc0lcC/ZlBakfAURAcbAXfg0qukb/jNGq
zXiKas0sOd8YrhMN5mxoz5smJ9sK4z5GJZb5x+R0OjRvZH3ZFd+J/+xGtoX7GtECX3t1nts7maey
AUGPsSVNEpyRFxHQExo9poZp5PGpy7HXcCgVCSSwuSqjysu9kx+VD8oN8HX8XWStcxc2DV1SgnB1
Y83DX56w3G5AP6kddv2WDfFjgaBWtzvtHoRtj7MKuiibFckPLnE5vqPOxo8SL5eFjy2Ig3/8SbrO
9gjaiZwkGs+b8J3CBcglN8XUIw44x8GioBMgwmgg2/kRifYRvnCekX1RdWaAXRe7W9lhITW+0M0U
qPPO8fSxwc1iVidU9tBIzct/6/IB72zBslXQo1WJ2Lz4zaQL9NiQymexNB5d2fgUCXv9ZE9Wpbd5
+lljxom51cCb6u+gWtwgsl/1EEs1Yx+40GmUVKFYS16I3nhrXPb2y/4+FJzECiEqZidGwn4P+t+/
phVNcjgImJzxOr/PLK8IWt4kkWqK2XZs05qr9fkwzfNj7Se10qGNByB5ew09VFMpqVweT33kAXcY
9izprfOFtQ8srzmSrgRoj7Z7bk2Y1JLopvuZzex5J8OAHMEIXLhYj5Sn/GbJ1D49jO2TyzO0yh0o
rDFuLvsVrY3FqsUtDImPKzwuIlBbq0X9hA/Rdbfa6mVMcuy3FC3BsZ+mnMKDsTgADvOMC3dEKHDA
SQSpmCOSWRtz+WwaaI981t4roTiV8mjn+yXi/6nz0kW6gYwflhmOTXf2Znc7YWflgqNR9nTwKd21
ZYITZRGiEqiq8AXmpMLWI2r1T+WcX4Q9AiAn7HxfUMJLbtJgU+KZowCu1sASYuU23LSFoeSePxg9
7lOpGT2EUrpOVj558Uv0rSwLbJZ+mGWSGdaL9f7HjhYKN/RhHHCrveXItV6cqdcLUZHJqR5yXk6f
QOSLFImXWa7wH6zgMlkW9fgyZO3dw7C46IpLPRlKS3JWuK8SAVYBdf1I6pgYA9JM8uTjh+rc9Mje
Fio23so+DgVJYhUMMMU441YyIJtsYQcFYI0RbQ7z43DhY0Q6DuZi1UYYViaEkkiaTS3fCdBNeswJ
cUIvogxGtRNwFe4qo6GfQNPtpX3oYIcp2ibSzt/eJm9irnXvb0y07cZemN2pZUBgGXqD7GcYjOIk
yrxpmrCxjxLTlrjJrCLmjODsHNLkMxX/IBIpyIbiNgAVcnf8nfJcu3NUpOPUQHhHLDji+YtnVofl
5CHEWY9vwwNaBbowAWNwOjpnfyKyxqm7HHCIBkaqbJB5if+DJciq+d4QNsiSBDJN1AeAqCQkjqmz
fYTyzv+nxpQFfPSOdQJvgwIRxlqiVpPdpg4BnxMsf3E8XBAihCLbmihwAosNTtEOotLNMw9809Lr
FAcYpJzDbRwY0gv1TVsJa12MEYN9UNtfTqS4GDfwPyfAfAoyQT4HVSROkDL75RjUEqs3ecs66nUy
SPK4AdLR7cGjVkfUrgz7jQXMcAQlvDmLh6/V2ftJ6e0qN1oKNRFhi+2f00xbWXaAfmBxOa3mY7/G
WPeXut7hQoXYXrxp0Qe4QQUZbMWVmEHf3QK9VEpkxixKPNEW3whHpVftOS/YzaJE+uwinW+2Uek+
2fbkBEVUYyScw7BV42sc5t/dIn82opTBUtzR9fmYcrvjewr0mPowxiQcTwJCuHXJ+96X263MfxI6
usb2hYF0U8N5kOD5pqBhk4te2te+PIw6k3aq7CjcjV+kGBcwFAykoYPugfzIbX0JfbHhgNCG5KdZ
1yHGFqbRBCDMtJGw5x592tkpvQCy7ysbQzJAxla3+q9BIggYje/X9ahx7MWPRuNBC0r2toFIi87H
BMM8oLgzv8TAnBa6PwIhHKMSlh1ZlBK11txHXaC69slfyzlbHMk3meso37yC0c/xAqglD6IrNpIp
zLKjZxJ8xada2xVnjWip7TaBYdOFVwOw6Upgq1z62WyckaJL3o4HZ/IxcN1CuRLRbfT3rZEeG/u4
SVX3HCzAbVkAXN5M/1dGV+hLJ5sQQLnTSefH9ej3MryV49NEx/zQ3dX20VO/fyPdNbLI3KiMVwjM
7MIRfyqcKl+lM6xYWFfK6f90OAgoqfhFtpRkK9fgG0xBpQdJ5woNv3wOOcc6wvCpx8uuvHOAX8Oz
Rmh0RkpD2vbJos2qq0u6RumPwh69HRUoSthS60cHj1kWvtHoyons8H2IdBrm6MJ1pqwz0DaSyHVK
fRd4EuMpDfp7k6hswz2q+/cDq8I/YQDaG/h3Gob4lfbsk8pMZ10oUrsIv50fX6o4BX9gx2atXZjC
IG3ZTFE7a3QrmCJDt4aEkxRd3/ANk0jmEx5m81V90aywp3IsxdodA1RNbqWhANUIfzTVDtikJ1eV
tjnkVYKZrHvnNJuFtM9DFK4+IJPuoXEDB/Zd+XWHUlQ3BORerTME6/a5QIAq4DU2g/7H8srNtoxX
KQ0YNqLFweHmNQwywuaLT9QCEPJhNbIvdIlS+U+idx8vib3415hIiaYMv9QvrrTixMAv7ZRC8R8D
RfOvbr9aZvv/YZRUFtcDb4nzPM+9e2FFs9WyVXSGTIwgxHR9cih6wPhJ9IuWeu/Opik/5idPwbCd
yEYmBWz/PMy5MPNtYg9UD6Q/YaLn81HpCr506L4yVwQQm9nyohNWOnTTnVeUWr2Wr7DsXduZopUT
K8SsgDoyUvXZ6DzcJR464mlULFWo+8BTolJp6yjZjhMzopisYfm8HcV6LlVJL52bvwUueM5UZR+i
m7epZ3GHzYjim2YxfLQSLZrD2Pwkzx7+sUDcH7uVY5A5fmOMPDv+OGsXYHM3StsI/h/p4sTWWykM
enSvFtUxfcde8Euh5VFmQBwJwKTR2d1Q+2SZCKN+92pJVz7Ni+sSQcmYdI1iPnUSXpxKgHNpg6HR
xGmoK9q08YDW/8JXe1hwB3t9KQeQaOqEBjyL+5lkbIwGkis1sIr6v8bOod6OJ/1bB/4IWBXAMCkL
nj49+MaFO0XemW3bMdW02N54i6qNAY76KU+bD6QObhFjxOIdTHLjxgTT40VqWJsxvjvfUPYn1izE
7tLA9s8QHReCh4xzQcaUlITMg4l9xOms6gR3RBNHjycg2g+H0JvmEJqgjWhb65ANjrHmO5fDb8Vp
eR/Fuk7Yd+t1OA/D6f2YPkffuyE5SIwRH68FiiE6EKFFpqduDEMcmsw8AII3BuFeydzSYF/pASE7
l/TlsitfvmDoS/qGe1eAteXB5ONGgSIu/ZehTLsBKK5/s60JVUKpuOnw7RyOeJuMiCilYMOPiQH7
IWCZpfweElmmnsj5awdg/uG/csRL6joYiPhqhubBsRCTBbaQP6Sn6AxUr/PgUAErrwaFzMe0arg5
5Va1g3xiEOhtvp8CApSgBk/9DQuSljecrOCMq5OtSP24S6+sYniskZd3fzZm1p0ur+RnKicW/mOa
VSzvjl2U5sU+2OFFAFkyr1HtTtBvn5Y27hhg7eNYBgMJMj4+JS2YBinCTwLJ9+vO0Xw5GL+wLTWw
wpa09EgJvV7hu4q771iRSg18rjERSD0HJC8tD5XW0RSPC1a5FzRTHsudcs8ZgvrZNgNTaKf/REGo
9nmJizax0FTGKs3d6p2z7fyiTAfxoGSQhiCv+QmVhdbdt6qISuR6S8unTSNA8+TMsAUGIrEf7WWy
d4i498Tjw1+ElfGQwmj4UZ+new4Cl/I3aIN/mPwovgqi441137xRGHOiyNbskTDf0WhdcIBGDmyI
5QBQR73VANutXeOJfgnUg6zF1f4uOutbiteOXEaUf+h/BHJZHKvR43D2bNkmTdMw6wJgkTiIeb/R
00ssterJxhw1c7BHlSXH4P7gyoIrjzhjyAJ3YMRyLQT2mNhOiCehcrxh9eNWcsGJAY+dl2WGzNbl
OaYdO4xiZIZ4sXwztd5pz8e9sIoFIuoP98go2l3/DISwu0i+lsT0GMX/lmEn96LEsxKyUCSN/85u
+gjjitdoAAFoMx5dlEdrQJI277iV7m7/Fph5qwEd2SahJGCXSSBXw2sXcHaVARCGyFHDAIMUoLmn
llgLBDmJA0VGOv1X4GKHBONhRN1F5cqF7CzH+l3rLSACLfXUq3oUYoZMY2kViHqtWISkBINhD0s9
YKyzePRDHOeUxsY/aXulZe4Gebogvb1w+n2pBWONlTQlaglNXjycHYx9DWRTcCE5/+wOjVKtWnOO
1nufkCAXnzgaH2bLHXLOJcH1+mkN5GGzyUH7IQQmgVlpGSwDBjWBP0nEmqo9ViA8R69OJnnVquUk
/TE96C1Bxphx6em/PJ5zkPuIjGasnLIhjwagcdg+H+4KkJ5CsqIReYeIevg7wW3QfuXjV4NQjI/Q
XxoT7h/fYx2dXE0XwSZuPTaKUJDGAToH0PC4Os79IX2FTHBHNaLNVvL9aQ2gGRue86QaLkvLSLPR
LrNvwmdJlVNYyI1Z+dC/9xe0Y689oDcF5LJz75Lxj4iHJN8pLC7XPCAOZlXbd3IoyeagNdPkzm8Y
hUrqM+k5Kh+GCHRrZSnEhLY7gxb7OaFrlXKfHFFpwr/FctzV4jXRzrT5OR9iZjMSn5kAw7yjwqRo
Qb/vtgLUQkF1OdHtmOFoCTST/Ztfw/yFSdIcI5DvR7WAHWcJVs0w2wfhxwPmOvrrdkhnsPSNCmsP
e399TYsNShwZZ+pFh2PpHSaQkIa+mG9s74lWsW9tqZJ/APtjpxg8EZqCrHvpYwsZuv4NPotnVxfh
ND4mtVFSRJvy7fC/wScIvmLhdgnaJjkp9wX/qRCKeWA28zuUEkxzW3yQYHLaQ8ujfiK3+489vLUX
r4/epUKzM0SLLYzzgHOiAf3Z/RfLF9XoJG7fcRpKdDkTwv4/WphTm8WHC/DTsO/qfkgwKkNOQZ9U
S1EPkRoci7Y5XFEfsu97zcg77eIKHAsKLjCYSt8+dcs42kaHLJzAMPgF4WCB5rLjaefyFZw5Xty5
Jdd2xe7tnqBaP96fs+J/tdrTBBRnHJ06me9zH6qabrffaP39pYGcfmEZdjjG+0U4r5Taa/57Vfmh
aXKgQLB+e+slBHv8EzY7I0NpABEzonyKECJX+Yw2kLj5iPNUA1iVCuMuF41pdjO/hM5j7zqbDoEO
4avfXuPbz2l/75FDqQo7vnOh0XJgsVWShdYkI96vlQDmy4x5RXBSHN3XEU3XNriVVnLiwVzIJMEm
NuOT/jbq/+X/phunA9QFoHGo5prKlnd6sD98pJhTOyX2RpyxFEiII8HGktE9Nle4gjzSqF49ZEeh
LEwHRXmPKFliThyOBRS3T5q/LKuTaVyGxV3DI+MwY9UoydmPC8D0L6u5uYK3tNyTRG/4Jo6K6YTM
dfF/nITfrvrnwde6KHjS+8UtDvbHSeJHBE1f3w5TtqcBwDaAmy8Om+7RUFA0UTlXy364LToGcTb2
LWT918Gm7g9U2zeDHmw8bTIi758bgW+DyNwBap8XLMUo1wo1hL5Fj65WvYWYD88SOccLlh5SRuDc
HuVeOb/LeU6E4dvc4ZHZ3Ai25N7dxBDTYaBvIBHes7CLRFGpkrKQIq1MxrcvDOIEBqFU5KJgZ4If
2OV092JwyBBUwk7BVO0lR5lgJ8XkCuwrcMJ2egJliwOCKshippNbXb3Aom0gHB7DKafHFmEyK3Xv
L2bo36gxVQDRsb/vB26iDBJPdoCV0UXwiPsbNqEgoMt6tIYyGFWXjTPWEZ48y6mg+A2uOuSmT+1Y
9UVS7vKV5pYWqsFB7FZoW5kE72X5KEczfxeEp2hqZ0ua5WYfATKdxH8BR6EkrO4S+tEl5YkMKRt5
TM8n5EVaVdevUCLwpHMgcP52m7krfnf7+DWuxCQjxLYlLOHUTCiKEV779P7TiQ8/H6I2msxoFlye
gd6Rx4A8pYR6XesE0W7N9payNC3eI9U6psUFrxYIeGwiQRzZGIw+UMJRir3ZCFpv43tHDVKogXWc
hF7tqy5mVmp4icBC+4FWW+j5zLTLvcokK5uhdQnADTudBT/XiKyWq/IeyFw4FBKo0T7lPcemqxVl
XMBK3uMIME6Fxb+oXDu1Z2pcjd+vR30+k4ArVGhTuzQQgzg+ufNcNC64rJjEQN9WnvX8T4SRp8ee
ELF8f4Cq4ofLYLm/XkvmHl1gMHnDLIZ9gVZAYAaq/e7s1hDEgJXf5Zh35T/iVaOjxCIkTLS2jjJI
zlCaWaEE1lF11IVHk/cjHPN8FXk9suZi27G1Kcf51J1b8WUjcBB4zhGk7f8Roe0yAqXnAmcrKA2d
Wnn4P81Wlxd/JkhEp28UU/tnCcao8ELOraEwBIXgX0KgRsOcYH3mOZZNrWlRv1Txf/+K5qAhLhsC
WWMD6cJQEVhuocmCOOHV9BeOGcM0UvNCBwxmO8XJ5cEbfS8sh56yauCmtj/KH9FUTsFmq38JdPc2
qMiP2gxTH0/ZnTQzCod8CtJej8k+eGVHmCvuhqoT5CJpssiX06wISIeveM1CA9XsbGIjJSViIYlu
IribKlqCTjPmyXPvJALmd9YMnOXKLZ/r+lxYtDMEjzuRmNymSO5JsbIhuN0AOzLB6zdtdKOL/WvA
gp2CqjZ40esJuRDw42zTQWD5Ns3/ECysTzYl8j9hqrtHf0B6TPKA14jg7ogHcTS8WUbuX+jnOoU7
tY+IadRhe+5rjCB9/iejpoXqilDn6ROjHGVtiwOALCEoBcx+J27DBGvU7ldMTtGDrIo0nqzGTNNW
Vb+YTw3Pwks35210D3LkcTAdFaTtvxVZykw8WB7rHAdsJRmYKubmbxFm7svdP/rFKdKvIBjsdV6m
WLL2zQSKWuXSuDRPoR/B89XjZj3tgWRz/BTgV5WFACkvumNkpz/hCuJWYQV5QbISpSPznkOH/J/C
blavxW1XTlFImfnBGK6KpB6PujkRoY8Y8JtHwn8SzgvMo9UM6bPy10cRAVnu/SzW0v6GRfwMPqRv
aeYfv0k6V4aWJHf03cIyh9nmMvghn/R4KdN+7r3cKEqCR3ZGEC2gO2ZUy/ZPfi0aQTs8OPhHTFyI
ZWxMc233rJh/4tIWE1hNI/oO9akQbE4J71O3kDGGug1cu1jRcTgLokuEbPnCjbCZjZm04bH4vOK1
PcJWWn+0MQhKHPcY7YqZT3speg4sIJlif1jMniFJ5C1qrXQh1JECB2mOldCS6BwZFCG+S1QRtV/i
AqtZ1QT2eBsoIJrXSI8x/SHdLC0lKkNKpMqMjQs0FIGjWlSyJuUFlRFfVNpP4UL6ufSfhWdJ8sh7
hXn6pnKz4gRMFMRzR3pSgio6jGnJOydgabEhtW+pA6p+LaZ1euRM4fG7YFuudi+dDilwvbFByuBU
ASZ4H64xyJy5BnFAjr7G67RGUdEF0AaotTQEl1KqpofMewEqr7Ua5dZfBBOrE6Xt5j+vhrIbLI0M
AJRXe7QL5pljjQD+h5me1OeDZHw3NY9jnZo/RzLU5eaRWUOXTIvR8OB27zvyPfd2Ft4M0XBo9Bg1
BPm8BnCwSk8RNaXXZcZJv2g0InEmLXHAREi1o7lAraS+BulzY/PcouxRYq/M4x/FYTDU/zBFNosl
zZqIx2SmFeik7ALRJeDgZQ7ADrloIhCK5aGmkMMVZl+mIdYJSwNQlEjK5aVKFNECypGdVgKOYM3n
EH2Jq76+gTF2i1FebZOmO0Gii29MQzfpeuCZHft+rMibqxo46+Fj6yuQ5yfrUGQHaOrFeuoTADDh
o3fDLMfBptfUYV5m27cN+bGOA70LxprhGGtALyjWDEOe6y4EmcLsZzDqIYbVXvieq2DK6UsTB38g
cvQca0F7lFMDUrGHWju+jBdfwI3zdDyM/YTLAqP8zqYbjxGn9JyruvLlnOGLjk6ebIV4NAIt47EY
Qw1SKK/GHZeFY9otj/EfEJxb1BTjxXdCM5usK1/r9ejuXpnFQMtMtGGiV2KiuQ+q5WrtYLLxppQ+
9v1/zYHl8x/1veuLN1RxjwbG9+G7muyhscaNjSzPK8rMuihyhtQKrA3lyXQktsHWKIgL7nbNL0GB
Wj6NeKDuxiR5QfzHvmg4TJPLTmI0UvyZt+rgA1y1fSLZCs4JLcU2VSPHnZNEUY0w3IfVrq+ZZFjm
dxNg6k7ly5VZ/DhBRBW8YVetkDeJkx2+s1P8uqMGLeJPxm0/ma6SOwmklYerun+7xd6brUuzYR/t
2FMGklZ+yUpXtbR8/9B2so+JVI9VSsig+9MxoqFf1W2/pZC/7R+oxF3Whf505RAH9ot26VWVgORS
1BJRyOku/iQCqFaOzUwELlBt5JWbCcB6KK1b502wK8GOkibusLu8ibacSD9ZEfP3SGjt7QAuh8lX
0+NvNtvuMovHMmj7BsOTfHIcV4TFVF3zw3FIj077njgbnkaA5cG/DeSCjxG+7Ug1BrRN2B/9x+L5
xLdPWDmWlcsOsSa03/osJJv4VQFjOo2ckNtXqw17hU11bWMqXMzXPdJmKJncW/JqjEEUpJeZJjoF
wlD3Nv6v9fyMMhqhUec3SoWQbjMpFCky7sq8ZQNfQy0fBYO56j4FUGGPhdoDz28vSk45yS1Cq96J
i8pBHKNgmuzJrxN+dA1HXsQ/iYRjsI2dXnTK8gDkeusDRrG1WcrRuVp465ESxvcUM1ugVyhUHOaV
FgKvzGWWxL7BTuYMfzNRlsb6OXBEuZ3UOTMZchX028thphHo37F83+5UYLGEyUZgEf3Tdf39PQLF
11rd5lfOdNjpvrfkTZx/wyTNVcZfATAO/7cJusBlxAcI3dUcRATQAchZ2z4A4lMHVjm0Lenx8Iev
T29aHnQFh65bbIXYX05px9c5HLeVDRP2eUrWfUyg1svbuuJEfgKoAlPdJg1FFzEzPVXR0OVCJa3O
FljXe+wzzxz0m+3jR0pYyQRQ+ylhXj5TJqJDXcFLS4UrijzhHw33bXSxSPdcKb/5YfqLvh137hdZ
P5KVsf9TS86FnulRvt3rs9ldphXX9N0OlJFVunkYt+8BsiAVRPyG0p47EB2NLlYC/NzKVMc0O7Wc
LOuMrNFADQFkEz3Tu+7VC1BWfhDZKqHQZ591bAH574Y8KdPPXJUUHGdNXq0ETIdSEg/FSKXV15Je
KyV5l68Rzu0pQcZgBWafQPq9grA2v2noL8PWPjWbxYM4JtD/queh7mNpemLuV0N6XGrrfxKEwruj
bUbNgD/gNwawVbLLwrMjKFpU7HWTKGLmgRgv1ef0+i44mDoS3lLlTthtLZaIIeDNFulXW9BpmZdb
FB/uCDgwSOCyMRJUN8e40P4By2tVLpqXQqtHN16spC4slNSjgJJ2PIQR4dAZpS+t+4Klz3KhTv+2
cPDGq+UOvlntLpcEFfppHnVV2sdqPCRIlbV5mcI7pNeJeGy1gEZQNGuD0mCuZYXqgpd6ykfWNuCL
dBY8IqJoM+nXcT3+g2p/EsjevYAFkkAWlgIISh+7ph1BmTNJZ4PiQ2pk1FUQelmyQebJ6ZHfTJWe
I6TBapJXk1zrLYnubBbykRW5RFbHEjFBQ7VO3eZhXbPqNpcRmHzH4Qq2PO5kveFGSAztefcOPCW8
ZEL76AshCueo9bGZyJ6M3/i9TlfszcULDHhmuR62wKfVJF3aUEzGcC2WNPg3Kpo8pA40X0eRjIZ/
9yNCcDcq6HSVlO+PntxN5urN+D4PXDjRWJOVJQ2WHJIJMmeOHxGNys07gwy6rf0Ij2d5kODnXN9d
IfCWh37Jki7pBfB/07LL8wMy4liFNs8oEznG0EQnWJwvMDbB66ZA0r8aYi4cGmF9ZH9pe8vSHKQY
EtUX7nvULxYyX4ByXoWzLDo6UpuqVqCUT0hhQ/DKRiTJ2zMeMAeSNZw6NsREhYCfCbNNeYvlHSsk
P7+6GQibPOTG40TZmIGTbrByzYClCcN12wrw3pTjePTDDqj6SM7JOZQ5xFYpwwIkh7ftEySEAN7+
xUiHmEM5Irr/eHrRi6KqFXkfxC9St/K8En9oMXiNwJODdsZWT6qRHHXIFSroLF81k7eB77mFztV5
ZjufZY1zGJbyci/lIyaPLmf0zVhhdwErLZ+0GKXB38uZB4nexPE6p8XYD89Ta7BnHJwDFBCm9j9L
8s0gvIeE0H6lpep3KZLXT32xOxOmpomDiVuQF8V8Fw6Z+FvZL3F99JOs5S5TVszm3TMqCqdlM7HL
6zaLjcKZOOyne/z1/wlKZqhS07T6DcsTGIYEbuP/2gGxsdqIFB6A6WRfu7IFwg/10V/db9GMhUpp
RJkkw5q+zsCkSwUm9zFnu8R/teF5UQnijFITt8lbMTY/kdxgnl/8BxzAX6CKZ4+V8Eh9fj5teedK
mGAqo5SrU6TyVh975Rmpl7vA1iHNpUXIZ2sQZU8cXfCaAUIL8MAaVtI9zcFnSl75hCM820Zp9Zyd
g4+KNkexdUAALoZIPMypBlDpwlbgck3A3V5NLQ3vu1EcyMUoEqI5RBEiaQqUGVKGjZ85O3ilZGva
AAQdSM9HzdYrA9dKmQxCxWO+jMIsCMZPM3n+lfmHhObvlQOwGeWAOub5x97Fjpzm3+JRUHz4CuD/
IwhP/EB4ujXb69QIw4VgdAnQ3Eeu+fnGOfJeLFqqjx3AepLtLaou0kL3T8f92V1mRWGCY0n4Yp0x
INP4jl8HmmG3gMHY0jkO74xIRQvmYHb9B6WVuXHLa7yizPYzIjFJw9leB9xv4qyEtdPNCvK0PdJ8
hCxu8msijVUY8ImMVlgAjDsh3xCuHQBHY/l/gUc/yLuszkMjcggmym3iFP7QvIax3i5hMimypLVJ
6+TWcKzdgOhFkRYptQU0xYdQUNmeUJ5QZnEQ2T0AA9ee6tNEk7Wo3xO7jEWbMZSGwvMuTVZ6K1S1
i5r/GG5wLpSYkkvZFK0UTNBqhC3ce3NyBGzx505GUsXH+5WBar4jP0SdJ3n8WtfhODbSad4pwvEi
ZkNWCq1/8BdykEBrfFFQS7ePnt3uUIr4InO/AaFAr6OHq+/E1K7n7xP7hI+Wa5fxoOFHYEz/HGQQ
GJdI5w/m9m2czLmbwTzQbfy8l0uRB1eeiJiyCJ5DYsS7YcOxYA7X48s1LtV0yEHesRHx4/n4RmlV
lzSw3xDZY7QwsPBwgIQnzbhtLQlToxalBRGTgwzOA7+mMKAKsi/xmPNgEfBX8qSDyTZV22bHwRcK
Nh7toZ+DWnTG4R0SMbRYsdwGV7Hl9bUN6G+V0l5ZoY5Sw+sAIR5G1Dp+7pVWT8avscq+aXfowb/E
o5KWESnMYcrTFJHKa8qKRZmP+Y/zmkXpcMA6pZyzvBLpp1UipGMUwGA5I2vXO9kqWPgv2GhZFZb+
OY5VTLP7d+D5CTgahgU5x3wQdFzEM13oWWrm0OZfu/K0RZRh5qCT3SxQbr8eeck8FKhfu+ytDIrx
ObJHSXTtKIFgpVgylIzf5uS8q8COHi/36+OHGx4q0kwUfTA82F0yy7HVNox4+ilK0wG8z1AyHQDK
SBvuTCUVEsBabezUQs+cc4ePG/73Y7U5/EFMZ1TMi81Mr6beZC/GZ3RGA0iYveiAHLrxNBfp3hFg
RgbSYW9d+7F8p6ikV9YKWiHEqrIwDqjOQtD1MpVfGHZkuc1RO6iYBs7Odo7/ylmMIskWI1Q4BHAh
CDLqVUDb/X3Yx1nVNu3v83yfUAkqYgeRXA6gtucbAzAHkUSAOlY6mER9V86LOijAe3fb52lmgZDU
USysIt7x4e5DzHVy5JUuD/jiRwWbjtWWUsy22ooB2j+0gfPWLCZ6minOgvW0iw/Esj7NzYdLMJim
3lw26ZYdDkOfZzVPi7IzKrLPzEB3Su0YCsLDsEUl9PbxzYdjn6IqkrJwAey78cFUXw5sl5ZcB+km
L+IDScJJl9HT7Mdn29hfmQ25Rm9PAiHR/sHHNh/oCoFBuDzz3MjqSNvQIRmd1qauWcErZRN2Z92s
/Y9FDOJOngBddrm8KwxdfrGMGhpcULInix3EqAYK0WKz0aEuVEcICn/MNkfpS7ruL31Z8W7zwW+l
jyNvxJeZetOZwpUxF5siReKPeptMed3I0mQwxr5QwlfU0U+Y+ceMGqqJXmaZ39ipSg5wbIbHzsfU
vcLnQHGuCiDSh3sFtRidTwV1Njr77M7FwKUDJyz54z1DG74El/iTqEXkAMCSjXACJgoQIHygspcc
BId9IwPopHJtwEGCiE4UfH6wCAQ1WVwdX+eBsEkt8pBty7+ilD5Y8WUJvoc9AogSF09+jJa8HQz/
1E8wYQk+3PeraENdBN9yT0XJiN6TmRSJIbek7qFglKVoH7vdgfuQju1OSBq+qGkg+MLnAKtFa2e7
KrKFR6AHdts+WOv5oPcyLb5sA+V/WpCuWAY4RFEUeAf0kgLFQ1o51zWDdxFFtQicW2LjP1uyVk5m
mXdRMT8L1Gx+jM5eXsRGZYkBx6efBGyQOVmx2EdRYgHWgrqOZmerX3XVyPQIyKMiNLukwgwrZnZH
awPVi+dcO+OS5KT+PAYrAZT0az5PkoHqwhzYbNBr+gp0+ygcR7lyw6rhi5VQLfq9Btr3UsvaIVSN
82l4XBcfzNw9+22+Khg//rOJvEZ/9QIp96X8zKg1N0f2jTVab/FZKjH+Zb9Tsaoktd2SH2OzesEn
z1IBQl3XkMw3urPpITtgvpmEd+HE08/18T4ySWJczL7OCuxd5V5wxL0mu11yDpVXt2n44vIr5di/
II305Vjy2jk19Ggc8nJ4w+zQpD0+zuH1aAoe0zloHKlttWEBmJc0zBR8Wbtm39obGjWji1TSYJWu
tq9SlwUuidsJrtUgEBSZhdKZC4K6zTURXo9FYl8slKihK94vc+qq0wZBfSL69Tkedxw7EFdpY6UH
1SRGLZMmP+G92yHcR3/MiqTaw8Q581WpM4QmDvtyiS2/+Yn6Qgbvf2Uh4wn9RwWwpEkfC/8rFt8Z
kckJCcPWYzuDQwO/gzEVetErFgcRD8R5x2bR7lMih2rBMBEWD4qPOKzZ3lNkGx5AsP5mTmOtumAx
d0wAMphm0ir5WXuk6Rqv3dFDYirnHgM183bunbqDWIz+wOj89X0RzY5ggpQUqnt3wo2INCDxHV0W
wwDA/SJ1W2q27yn8twDKsLjZsSDC4GC76AL0bvLer/pc2ruX60OThXjcvXIXQwGdD5bTOdh6Vb9C
jIE3W0yg9qYNfEt8TPbRnsjM1t/DsxhabRVaCVLkydWmcxpS6JTQTTtpw5ACfyLvDAhU/ss29Z/n
GPH2jP36Ri9Hl4YE73nmzYJLFI5v4FKZ9DK1NUJViZtmAVFWyJoHDX0wpKi735MuIcbolP/3cH2s
QbXnUlJ3VFzWZe2aEzQ9ItM919WlVhHYZ+IDaErEuBW+bWTfe1+G3nglOthK/9FcGKkO5i3y6Auq
yW//dzWpSqy/SgQUV/RCNl5Nag5W6Bt6DorC2ga11J1ziLb7VHa2fMRI7Qt/FXB+OvF7XH/bX8OI
e5gyb9HZtpv/8440IQrgY9RJX0zQ+tid1EM6g51FiZ4vLTL9B/clRzfEKxpcH7p6A3WBUnP1ILPL
8bGr0Rs9Bq24mqH3YTLKDWDncGgX+jYrv0Z5OBUNU0FEr8tH0CKqVd7f9u7jYS5Hr9dsJRZ9ztCa
cqyaVJYavKG2NgWHyQAQW1JbO6UacNKKWMgtROTVzKJDQ2azRA4UxUXo34McQqAdna4Wdv3V3AIV
0Hc30N8+zkhBxCb6RC8kqTz9tPcpdljDY6JthqdPa/Ff5lhSJlbtRyjqwiV2xy9SE8VEr8kXuEFx
9VJwGFriqpQVRIkFIZV02VYzdnMMnA+FKZFCE/TcYiCJTRJIMs+lGlsUsxMtibfVau1+LsCSDQU1
kIpTBpc2nnSfAY8TqLPaqNvyqyz3BpxnGst0SnaQAJYg3+AhBJfmUIQu+YPkLyvA1Ihf64bnnf6P
EBS7JQKQRcHkAGoO7gAodowFDwcwJMaTo4LvdvMcQpPb598RDqul5P8BKh1dg/+BlMPWb4o62rOn
sIR25ex7wj8rm9Gtll5wSKLmW/rKU9/xT7aXZTGClMDaSxJsTkdr0VcEIshF84S4mKA73u9NV3e/
8HXP3syu1sP48G9yIG94XskcVF/rrt/zayCfDoFzMBWSXJsUutqBPMXTu0eIIVkC5IGuTdXDEub9
hxZynrj9PWstK3Z2u0mgw9zFP7bSrt42G1x50b4qk12FuJ1tZ9kvVycPimlU3c7nSx2D2eTfZ6h4
2SJTFv8Hc7cuTdyl5xyJfkjVkNWsYDD5s6LEgK+fB7kPqtGNSSY1XMcMBMkzv4zf0cJD8RGKR/2y
u0UtiWwTGNgoJHMpUDuVW/dvovCU3bIcdyHLqx8BfVW8mB5MPNC5EaGTLlRRpF6yy8NiqGM73PSy
ogwhs82j1pREY5EcslBZUtBoi0n5KMcsGHpJriYRKbA0rhePFDJFSYetiny8UqFPGdbp6VqbqWVB
jaDZMFUjJUYvdqZttYURkFeZBEDDxRsA8r7iQVbWhm2mB9rr0hoGuj0OZmY2Jdw6vKSBEKyf7OLU
Kyx/oxexDVLDHCb55e/Qkc0CMFI4DPZC8LL/2hsNBTKPq+j0sWz+mq1oJDgsmtXJHsjAUopyODOP
ioEhuucG6LtMZ53o7rExrGDgy6xQb5ygwem5gdBbIRRrpTQs1DCuHLqXt2y7W+aRF1x/UMkRKnDs
hw3VUx1jUvpzA1slLzLE14POKNrZ02fxynmKiIHB4F0iQygJ/jGzuGs1KdG2xwfoATROSyoNJ4nF
oto1mj352p9qqgOO8NCF8G1HTxfHlAg2XDuzaV9BzJY1Z8D8vUEfVp2E/PvgV6zIA1yUdOGt691V
DbPT7WZftDWjrEGt9eVRzmBrIrkGj6pKCv42o0pYwQLcKKPjEKTK8fpdsu0TvSCvQLHupgwvIC3Q
J9gEKyUSQJ+t/KrWt+VgHpAQ6kEYKoa8mamSwmw1/4cSWF5EKhCAM+dTY9eS3+fFifpTRxsLLV8i
IuLj4P4H9sojDf92+RrsQNFR4eTRRTtoPS6UWc/ehtPQjpB+/SFhPYs668XP+ZrMce0YfkBgkeVI
aQ58uiNnvH4U12dRSBPImiyv3ijoAcFI7gEqkgCEs9Og2fUNbowomz4HbHF2d7azdd68rRVOhGOp
5enUMBdkStUYOZEKxtfuvsYo6OsDsTaYwp3NxKj8dbglwjH41AXoniPobW6cNvbNWjjbYoxqDAWS
9rgehdALudSOYkjzett11+TXBSfuT9kZR7Ny4gqZU8Katr/XzQDUeuSfkqxtLRfN4HFFhnJBX5QC
WcIvoX5oStxEvguO70mAgPx0iAfSL7wJr5BL85ni9v49yj9DLSSnNb6OPISHAqrz72mRFNYUDcsy
cT0d1VyFhIAZvrxs8jPDTHHKXz5IAcjP1lTpOGpL9cyUhOonKX23V6qCHauo3hpzq05SqHU7e70y
J6XyrusSyRTzj4ofJIzgpqgcE6T6bCsdFsy7SqHWKQhtq3Iy6RE9tjB2Vb3PmdjeFEWgv9jxUtRU
TaMU9BidKXhCfzmT5YjBUe3YKEOJwqTpS3Ze3tXE/RMKimjTTNXCFpn5k1Fjrcq08+jH8Q5FxJ4M
V5Nv9W+cQPGD13TdLYa2hhFnVRdyKPHttCoiwlo9DsuiDMlZFt0tvlSYTZ8GU/GbDgrIP6MQVcfy
h3kFOjtQ2vTwW57HiUJ3NRqPlFr9YEVF5o3RkTlvWDWIqRBFw3+Dcj1OZy20cwBgml0l3yzpgtPJ
Rldbke+OxF5DHmbiWAPN7aRAeVd9bRUC/PyYu3GUo5VJTBFZB8AZ3yIT7zGOlyMsTQwdU0jt8c5p
ytHX6yJqEI640QVXXJIWvHNvRWv3QoAtvScKCrN9NIdjdjDJrVpGAJcBZmMFiTy9/ofPdLJpcahu
+F15SPgrwyc2GPsBnjVcINHw9MLChRofPBhgX0+v0rq+dgECNEX9h1lFstb5X10ti/90z5g8ZX0k
8EUg6VWYWJuz7kuN5bMtIONQhtepRwX63o8m2ypljIx2FSMg/Cx68hojVqiv+x3t4w/NAby6QDJ2
FcHlgi1ck+mjv2Uu4u0ZgBhuLecWPi78w4NygFx1a4stUIrbmWcMSt6RRlXWIwr/G0zKb9Y0Lpcj
kYnhXDNnIT8nVpcs6awoeQkKcamu2DPjUbWJJB/a/72HOz9xz+aklEMqL+K39dOmMOja3rbwaLsU
6XfVPkdDp3RLNh7c5L5KQ4S9nXmhXMwcTgcoCPwvRONDN6xT/ptEglYQslJoBrU4nbBnZuaVNatn
7N9onMothGetYbHtoKfQvLSYyDCityEa20Io8d99jJkq0UjTliwrwuoC1FqqgtboiTWZa3nkXt5n
QDniCRhLYB9Ha1a7zjhVDR4jx4NFOauW/1IYpXLxuffAl9VvwLsTyprBj+bo4BHm/mLbo+tXQoJh
LWL2KDPZ4W7BhHqb3ANABLcmoiHLjyxl8Pm4aE7v7jtuPpfvk4r5D3HaPdjYIw56VkrAWJTWE56S
5q2SN/DVFVGfpLexi5eRBQxazP47r4ic88gd4rDmX+7PQ/RO6i8mYXV4tG9wrbVmecPDZotHcAFW
GGIAjpxPdlLWGW0waaTrsF91Ba3WvlBMtrfaKo7zgDykdV/aThALao9LX6IxCodVvmC4viONaq2P
7/GUk5dvDXoUJ+JOSeeBSMLq2Cj4+4v5EEKR0S8jscDUqFTYcd0tPX99kZ+cPYlI69UFLQ0Dg6KV
faWApxhc4dYSwAJPX6sBEu3jMDZh+JsfbFUFUzfTUUJ5kQ2tK2sRmhL9OCQIYmUQVY3J3byAeW3i
ss/RzT7e/d5SszTxtvSaZoxUmOAxXc5oDMObdadoxjfxv3bejI6MvRY0DAkwlR7UwtEd251G3Da4
VQsvCGAtmpwDZ/X6dRjFjEeGxUTojRxDgqWatd03aiHZXqCQWx1gji1RkxCuVidMeJg4sPxahHsQ
E4vKXKI2ZCBgrStZnGK5veJhKFLh6Fs9YypRiwQWRf9kCVG/BWvRT3x5QzhNBlMeIIoK4MJwwL3t
uTd57nVPIbv3TUBBsLRVIYgCPwmORj385pDDOTVxd2Ncd3am4717aOYfax0e9PEkiaUVRGD9GG9B
lUqI4mGJ3Ll4Fb+cStW7DiNiQpEdPRq6881MuaOl5bH4IXryK3uKYhEPBVs0/3BZlUO//MGYv8Pm
82hfzCcJkFTD/LLZCXsCP51JHjCCjXUmQCiNTstcT17qVLtwNLo+4rTB+IAAAW2iXbLQBD5ohhrD
bVMxMnATI+Jhceoqmt3JN/+GpKhSnotvG37nZ08nsgtKwnNepiQI/9Zvqb+dTsHMOiH1qLdAPz4h
UpdYRuiGw1tnWmpc/yMaq0HF4VhsFl63ws4j0T6aOKJgezPCTxSbrKGWuuwpklCuLe1pLnlkUljm
RY8ZBIksFMrAcr/PUzTPUftAFTQmK4S/4GhREkCPJGqVSMz13oPk7AhVNRL8jKopCO/NVMzauNoa
M1QqcTG/Ndb1Kpu0C5KBMghiQ+QOKgG0iQZRp5T7OqxX2+DVfdxx6FcWmT0RCvPV1cxIXY4VrjrL
Wvn5QhvfAhbE27qikDvPiMKWUwd/vXPmamRh6QQcYC2+WnIRlSSWoF4FtfdeLLfUTrhFJoui99rS
a/4JWN/xV9Rraw8c1c1yQhPJn9juaZvxSIWOts4795iiLkXhMx7s+RF4Ea3uVJd8nPWxq46CczLj
ssfxfqvW2EAu9o8h7hFN/b5QS7efDP7juqAddCrRjG67Bb7bFSlUSoenGG3eWTxkwcPkKTbtZi72
WuIPe5NoFJpySTNr9PyValsP5tA5DfILjZF8+jmq5+6qD7rtuJBveteoVy0frq65PKPksXYrGK7z
KDQp5PqzwVRWEJkG7JdOZ45v/cK4S0KPH0e+O5Pi60GRMsM6IvUqZjPObUQsxQa1gdd7MOatBisG
fpQdMXzoL2/6dIPASHHN32mSEMP1UyeTF2FQZAM28vuwqw2XtdGA6bQhPZqbtDo3kVz9vGrH9c0n
wOTEefooHL+0DxlqKnljY7CmO7nchtzCCRIgPdW1DVS9YiHMNd7sDGQEysOUvC9qw5/n08ZRsgQb
wCfqTKzQKs/DqNmchFOfjwMr12fxubvhInNSP+R73oLQO9o3+knTdv5aw8xRYzbgTV81a485TaAz
Tzzp1egQNusKCob4QphZRKJC1/tV2S/aa+3M/4dOaqjkPMf57IPoUaGbiiVLo+oq9xw3ibysXD3E
zM6btlXOaemgj81jP7ZeAHlgbeSANBqizeVyUA3zzrkuQdTSoanyG3r2RDIkmKBUqk0mQbQrMZoC
kdaHeiHMNjPQSBhffnCl49MuD/2KvOdkKx5FHWsYdJ1paoH8lEVmUhCWdZt1ST/jM491Qe0n82ns
peDQ0Xr/HIZOafCekVVgAKlB+7Bn+lFaC6wVFNA3vvhtb86RV1goVUOkWLQfsmXnfsNv0y15wJv/
bR/sYEBghykGAq313mXCbs7jns0Wl9MJYio1OVE1ZpueLlSUrV3fzrnB7SKjaVqliOXLg2Yquufm
3Bw8wwuRZ+rybo/Yaax7Pl9NcC16n9EsgQZ5I2dH3imKJpWzkFqUDAEs3h8i+PAyD2tdMtMUwxPm
4+48KhtgZ37SG9i9whiFfr58WgeTZ56HoF7W4+nDs3Vb7T78F2btejftUJ6YfzvUv67GrrBJ15Ud
YxLmGQA1nCpg2e/PDJM87BnZvyHgLxEMGRb0jftX+MMOVCwlWxsGM+/x0+9yoEbkjkm8r9oSS75q
NWey60qLk1XDNCP3c979ksUd6TaC0lYGH4YLgw3Bufkyd1EL8sTKINeE56sxuleXZOhxVVovlAWo
Q5tqhyZgl5Fvtt0cVQ813pktBGB9tieB2bXa3Q5SXrVb8OzDjlo8k1IAuLXZbnSq3JaPDLkQ8byZ
9i62GyO0tzVYlbOtFmgzFVAY3aEMb0/fRDH3GW7Bksct3wb7TM0AtN8jD0jBY2COQUEoB6b/6klm
vglEUquZgrVftJX7HBX9OMratdVtGFG4+0g6bN/3cW800AlRRjKfEfaixATVbEQA+pB0U9KDgS+F
d5viVGD6AFBe9U20Ba/z+wrZQmjHM+fc+URoUz+9a2EZNu5se3Nw6Xj9hs/M1jUQhxw9Xupq+5lb
faGZK6mMajU3WAfNlsrTFBr7bp/JPqcKnXYkiZIQZOyFXUz8tS8JbHInFdNJiU2uY5r/FvWil/Xb
46jaSPjf8STSBIrC2h3CPNpuPlVLST7/X0hYRGpEklfpDfIhlJOpydFOyMnblG1keGxNpL23srMT
7fIls8QyNHqU9bMzSJ8EQSPyXahRWJuSxu1gTQ6BBNruZAxjkbsqCExPG25UHLDmrvB3v/9hhO09
KZbsuMq4/wcQK7VVmDwjl2QFd7mqa5vmEPf0kDf7JHuaSYo3mWBdkO66NG8IR+iFKR1DtQunubE0
5vvW/7bZR09JkmQDo4OpgZN3QOYvyfQuIFR0XernKejb9mQgPKvaqKl40+BmvMAlIEVVxlEFK+vu
4ugZXRIcPafVEgdLbcGXMYz4UYeupv5WThnspKEQyGTZvwk9ALy1XHxXJGzYK5xm66PQKwdYg2W5
1QOGcgeVX7CpLTjQXcyjiRrN6QtZyzkMu8A/diZajJhdMPXRex60C0+5mCoALrSk024tir65MKRQ
MAlCnuZCnmOSQuMfbz3Fu+ysmtFvZ9NsGx8KwfAIJFJZkaNTBWtgEt46pq4tN6PjPCwx05pnMnHq
DWILuSxGNqlPcgD4VZlPBhffG3o1NpVjtu5b6UL0u9JKYpG+D7V9eq7kuylvHA5ouz6kW+vICgdB
tg1spvGFBbgHeiPzGQfVn0iuU4TUHiItMMGOy3yoiL+iW55BztMWB2aD+8eJbjly5eU7tIcb4Cmu
gBATSaxtonKtdQrAYo66rbtzn25v66e6hwBGiT1RUjYYlEV7qa02ADBAYApGIMG/D2uyztpEfkTv
O9r335nxzPziKWN5zcQHeAhiWWkhIPLU6KGc9UDPiul0oVZ9pKFl3XXPer4xl7vMPcogbqNg2odq
2OgwRCHSa766Hn2gm2cxH1qElpoyywP7S6xPaeK2R4Os8e1Ufg1BsxeqYs42xdfgp5qs0BHhTwVg
nQCPDtsYy8o0+F4iDN7BgLn5LiSiRdn3leDuz0XRSNJwt645870aOAm/tIacVWbBuOBQNwStnrrC
3F6rb7JyQigKWm3abSkWSkeQ02dn7Rlw52+g5/adWEgyNNCMDlSEA/hk60TPUSFaCwfZL95Ia3Jl
v7tPwLD0SRMg2JpZdnzb0VbieiW+S880Jz1GqRQDuEt77XR7TrQs8GpI3n+o94J/C834CdzvWfr1
MOOXLGj5rNeIZc9poh7Wcofo2tVqsOf673IDH74BCYp0p+LyyK30DGOZu4KKCmxkXVsk9JRUjGVM
R//aKgJnpx/s8QNHtmDiLBbvEaT8aYn8Gn3te69tI6G1uIFiEZoUrn4HvEwOWnWl9b3+5rCxrz8F
1K4nYNTEfNkvZRo821dL2jLZUE04gPyCYGPPMgNgNUH5tBijwGszV/a2XZZhDno5oMxmW6pGebtb
4tiyEOnv8THz6j1gPGaaIDTkL/pH7GcdX1ryFZMg8W6gyFZ45liQCSd3bRUzhaNJ+Nh0sUTMxHMK
bmdRgffLsZwXcxY7B0RoZCn474MjUQLC2g6GmnuKGEw3FL8/4XIocRITdwHLQZvp5onfA9GKzLL1
bTk6F8GGfkQQNcClOpe+10otVSGdsceNaamQcxQep71MwEPEX7giMsfJqJUCUjZy7pslI7Zd6hUd
5BKKqw0qO7kuJiMdgJYY+ebVfRo71lfPtv8ZayFJ8fp+qQEJUwQthVeckkpIKyQ0MiVFJ9JI7Z2d
SGifYFMLJJ5mET70UB4Ce86weMYZDf6+HmeA29QhFtk1O/7Oo3enPVeWuSazHHhJSO3whmGwOQN4
yyePQ5+Iet1ARznAfSI5hMIgv7acg95RbfU+1GNWymB0cBexyE4Bbquu7Am9jJvJa7uAWIV3yhP9
LjcSqICyRrR6uPWNvgHrGvp6kvwESHOONcKchNIY7DnqNuHFjlqHbU4PoOZhCNV7PxTWlDuV4oeG
jmcwv+VAYFGnMCfBA+/BLG0L2aUqJtPeyDKKWxcLaZfSLM9Ds6adkm0lA5E+BGMJUncWu1oYJvwz
e3o3jwac18B7D+eNiOEzIbojglwvWNpdye905T9CCqJfnZhsRGadkMapz2c4u2yRipobTTsG0AmJ
pIr9WT0c2VvZwIa1WlriBddONIpneH8QGJXf4E//8NgJI1s4eEWQm6zFGhi54zMMk/q5beHHjqPt
LiS802/pt4yQCZPIMEbOfgw9a1PcfMdCqp6O02hhP7mjvyAf4iYq9tRAEzmiigyMqY4aSsK/yAJT
qupSGEKmE1TKReVcbg0ANvziWJ/OVnH6ueQOd/chiyqoYvgBVIWeSxnCEdWFIY8CVWYBOLsrBFMK
EjWf/UeY+0b6V1QA4IZy+k5yGwgG8vgQrUKNPjF6qX2l0ArDkpuC/o/1S07wxqxJcGLDqNnMLnlp
FQ01ua0Jx0CjXRkmsEmbrvi6z8+ZGa/MBNcM2SBGGkVxLGbmxMZszgvgp2L6avR/MdTaYYM5NdTN
vTGLmneZ/lw6Ik/N7AvBmHOO0Egv+Zka/gyB3B8ESFECFCAb1hioc9j1loYNs4ApueoL6I6jFpN5
x6Tvc+5OSXaJFsPcmyLgW2SfCobN9GbToasIR3fZwPcM+Tzv7M9ueXHgFsZYsxZCo77mFEJyr6Xe
wWyGV2EpzooFUoWUln3xClqAPeU+VIjJsJmIHibYA3M9IUILFbT0w0kdPvLkuVTX/5kvd+isIwkN
nt44LoaFMkL+ZZbZmOi5WTkPb9FR8DnupGH0bZSYRQ3bNLRV6qi5aXbJ0xXvcqNkd2K6K77XCIgv
b4GxKDAad+uYSbQ8jPL0lcIA2CjlaNAP1GnzfFmApK+8Qj4NJrfLxy7GDLuPNmDPqw3rWnkqAj0B
N1ZpG4ZO688QLUyHEWMlDMDnEMwQjt93LLxQWLg2ZunqjEJRFz3kIfAFTnu70uzGwQgVmUrOijEy
MDOyJ3LXr43ZxRxyTz/v0n8SatT2lnLDww4HPSbN7X2Btz3g6OI5ZbrFWrhVpUVNkMpx2DC6RFmS
iGuzpLKkJxmeMqCufrTKZI2V8JB6WJo6ZEiIrf3YPe/M2uJuw71YF80A+R5pL+R4N75IrK+f0Fnp
z/fjMZc9jwnqv+vm+cOyjASXVDdps9NeDWTA8vgOcH2+1rQHWc81tXT+z+/+tb8DZWbHd1FfP9pP
9lpbrjqbnNrCN7cVV2btpooBvacL8iV6ZSGf4Mp/qXxpPS9blD65F1jKD0ZR8NzLqeP2yJzSLftD
EL6HWW4Z6xjFwxgfuwrQInCvI77ABWqRjjnTOa4lW4GuIYsezThiOx4zfdsdigQT3Lv9g7SI/Cph
2iAielmk0g2ZqS5f6d5EDJstHyd7F+MH8tgNrCg+C2tuCTDnvjWJimfA83b59NOaHQgqXelkKO1/
+/zs1QlJzsBCaIrVFjtBOntSBvW4FiE4iZ5iiljz8LLdLqk15yQdVwlmOF1D8VpLv/gcpvU0T4+C
Ycuaj1Cc5kLIUkypINkPqrBtezmtqAMyylfn+gvDZsyMs4C+AKdujDv7CsKh40g998jQ5Gcrbckk
BC4EsGmNK09VS9XSJhtQxuhA4816Ip2D8q/APjekPVSHh9ob4rhnrWef9DFDgQG4ZhXZQst+2wxW
snauAId081+PjLBDfOy+PiDRJazUK+JgL+InEm8pGJaD9seCaUTIxxktx6adXbNiMbYDU1hSP1RQ
pgmcJtc0KtVp30tAiC9koXmvrwGteUMLR7sa/oGLKvf9OaW6kVHzSnFD6UljCOTbWkAT896Ktn3A
ktc6Y4Dv4AfoPDtPJ1wBPI3n0YOpIH9zLfzKVM1IcDpVDCtRF019ObE2wunXfD6ELaU1jQOin0Ld
UGLTYheNwVdMfRotZaRm6Ch00nRLhV1zOBvO/eOFoAnN7sQcycisPwx6FzSgo4Y8bEXFsTVIK2to
oiJVbpOoNALqnRG1z9tSs7h2FA9iO9umjiPjqbSgb9dU/f3rWa3XxQUoJUUYECrmrYdKUHZPJT5W
EUW1PMgHtjBWKpfu4lBtfmrdUpm722f0lVjp/IQqgjQPaUiWuPYsT4D5kTcVb4trv028LrNDWRo6
IkyMLRqCWGMRlsIrggilrCEvgcdYGhHR5DzLyQFG/n1990ZeAEY6/Sh2ku/XvRMBhQvxT4ylfRCN
O80aDbdQz3aeeh/3b7MtZbCoiULdOblI+gsaY4VOfR7CUTm9MWPUOj8MHEotLU27WlcWvtymIW3u
MTGHLpeFMMfWaWZGauLjvtYH3WEob4LDysId72fFZPdu3jcpZJPEkPJkWDwibpxyVxGr3YK/EH8n
Bmit2Y1zTImGSTe/mHcDF9RRzQnP6whIrPDUoMsCiEdi0yzmO+xosJOhxrIrZ75Bh6ROT9/hQWMb
dBdZ4ZkajJCdiqDS9ubKRQF/JvReeYT1WGci4/GjLNR4ASKJccV/xu6wlqzJgOobLvarpaIN8HMk
vcTDjx14+BQrMgVpzlQfAYmDTJG9gpY2GK4BYcyKXKwglr8MpUaDfiV209OGIqIuUxzZAkNGTAD+
IgOVjiG6T/Spljgx/07eUxStc8XI0Ef+xjWM8AJsAvpZDRV7eDpPLWstigYlhRaJ9JkjEwE13/FX
42BWJXlo8S0i3ll5rVk6MH9L61vAmBFghVZ4dlNDx9tJjbnep2UDsNx7NxrpbCEW4wyKcVCOqcAd
Ete9yFvihlDtIy0uqh4jKiu3zvdPEoHIUyUAPdp4RmdmB6zN00cQrBEjLqkRkYExFufwbOGmkZ6P
NOUKOQDf9Dl7OljxHqufpXkZdEMh919w9J7DvQjLeSRDqMuikuxK/XWlsn0NRM6cwgZP8lHyL+QO
5Qz+r9OS058ePO9zVX05/c9FwTWB6RIldhHjyvvYKDNaofFedcyNEVhjcof2exIaVgdjips5Jj7e
5KrMrYXjXna6G+sYy4LG6j4l9TFactmC1NDaJSUZh/28vIyh+MHcAaRxKcS7GZfy8rjwJGpwqqkE
HU+A7KI8tOolUaQ32GPW2H/IghKRHS2DM0iN7U5dn09Ei0uPgS+CL3qpIB7AcnneIjRtu4XcO2KH
AHrC6Zd/UCe7eOu8Y98eUygMNm0VTYENUxgob5bPrbPDLBbS6M0Zs1Nkxctamu4SqT9STz1QKQEY
3xl34V9RNwkmZxBtUD/35QJIHdLzoGfDRVeJ4EI9Njcl7PoLFqcIwy2m1nQTsFOvjdLctyQCUvCa
3C5skcdkW6W7vraji20Lf95oyNMTHNJoulKEpksL/2sKKcRdP5x1Xs2hKN5B++fNoqC/6icjgBmM
SeEmzHtWRf6kmUaihhnj3DlHIyMoAEzariM6e8PS67S3yNJn7p3NOl7qT62ac3R4VN6V/44dCRHr
HFz4oQGPAQihTipFfBCx+1nFJx5PueVoLm7vT6r0zvwLDhtiuPyrD53TM3CH9XtdLhFA+GqGXdJF
YBVSGAnXI5gnZmG4TqBqFtmEEgGDI8RtBVEyGfojbPRrxGQX1B4kK2S6ZcQQp7bG8O0B7E5mRzVs
8a7uTx5UyLQPYIGpb+quPjL1x2nT2Mxi9g31AaRN4EB5mqDHlxK1Gfb8wRyQ+gK66mrF29bU0o1f
16d4c3r0uJ+kZ+PToVRypXN2wZezGcfmw3n9OSmqfs5cm9+Ar+I9QojgT+XVRtCVQp4Fif/JJpYl
q+klJtzdoS23nJNF0yESZRH752pK081Q/rMLaA1BcSz3Qatu+rULkJKliWKJpiO8A7hFIc3tFRlr
KsNYNE7wXUDZvloFU5KI/9ykphWji6P61lummges2CCoOrGMN48tU3yvPV5Oi1tuIk500UqiovBL
HYd1Z+65iE+k+DobS0pI0i6zGc81bJy7IyeVDnl2G9W9rL4vBidm79WitQ2A4EnI5RbMGfJm8epv
5m48o30cOHISGN9yaaJIod/VrwPiUROSsBKx7vLHiMaa3Nsj/W+xxImxOs2KzU6s5Rv4/C7fbUQt
3XSVrUn1lMCUnWKlDpG9+GHFmRiIY5cC7+VIlSEtvXstBss0qyide00eKlocKAjsW91G42vJ56zG
LTegdpa8AvRQ/FDaX3tMWjBXwMh2czYoUc/0SbgcV0Nuc2Nauwzkbaoz/dzAXMQP4w0zAzUoatGx
Yrk9AeA8mVTza3P0bOKoUWCLnq67ZDRJJxgqWQqPtt0iDp6bX0UK9HWoIGipfpbXtNm0V3m30Pmo
1c5MoZJ3qoR2lXomshMKGzJ6h6dru6tSOcEDEX81nJM1bKvkqHkI0eylCPavK5Ph5eQz/KZXAEro
JWriAd7acAQ2MxByeSlyXtPQJCCmVIUeaaYIZ6RnDYvdYTdXGn47f1aQXpWkOBHMvivFhuVzLs1b
VfUsMV9bDtYgwHgHs/4BnKqixQ+WURw1yYqSOp5GYL4faKerCVc4dTjrmf916WxTT5wXr5q99Osi
D+Cgv67LbZgrgsrp8gK2DPDpvEZosArEAycAcS+BiZx8sbaynnEKBXj46rOll9rOJAyNz6LVIuBm
7xHqdINJpiMfd6FZYJ8P7u1cd+mWTUcXoMvdPbrcSzpEdpydQCTgLFmdKul3IOXHB/EbrAWVf8Z3
BmcHq5f4Pdlk4+YlONmp/XzoNQME7LTfTSZ7/Fea1LYiN6iI3lKbKcxTV4pEUbNi26MTlbkeNjDS
KUBd76dDAxc/2Aaj3rxe6/U/OGNF4yMYr+PIaneGb24BV1/qNXJehp2YTvJVi6zkdPpqcmMHKNRH
DcZmou6gjHJGwUVeWaFog7y5ftwBrGBI/BztwvKciV7KGeBRv+z5HgWMPzGOyE+E1A7KM+1e7Woe
jRIiAAznmR5iA9ZtX6YWp5O1BocKdBHfokX774gRx9HEJq3rJjSZ8o+Eou1FOaLhd7SKkKP/1s+B
3OZkX3as4c742DDt+43c2dJdU74W4rti6BKDtHZA16kcX4RPLgp9fn2aKuDM7Aehmv6GxHw95Oet
bueTJnnG6SdXE6t3JNb04orL1ZWsRXyEx/uzEP/BvofImimwJy+Tp06UvhCJ7jfmz11MvYTb3dWk
9ah1GqFC/Qep25Fepo59JQxga1IBONHwEM4DNiPIqe/DH8LtNMV881I/mBVIOpMvwtFn+abTwEO3
BOjaBEh7ZDnMTfOAktz1hgZOWUEnshWFsVE5GquEzQWnT1496mTxPJ+ATCALScASBSIheTSIiEas
C2moo4cD3PZ6zsbJUKT6meN/PjPWgR7FJgjuvT9TN4+x7GzaulObWTI7LCaFrvNfn6AaDuwYbpIA
ndZgS3Wp+klcM3ZhuZNOKxsqEUjtsBjsCjiGygU2MABOqaq0KHa3Txu+Iq8AlCnJmIN/3Kr2xFw+
r3R6TGhNb3qxd6egwPiLjxc8GFJwOGeJNXNaO/V9yTXBPf1HRPmDLD0tWzeBPK7wgwOpWL4CLpRE
L6/IafEJjtRoRBGQDfw7bLHUa/55dnHzqOpFK4iSx/prIYTdqjtPWTzODxm8SDhSzuiHk38KZQUQ
Ri8xplefVfu/8j5SSR1jcGOgC9pDaveZwSP9wvEOwIPsbZRUFhQK7UXRpvZrxfILbXH5qaE5XAJB
fqjxbEi8RypvuaSFvS7knvpmACSyYW64GBpkaPP96wyDutO0dnJPUxoM+tc83Cu3Um2pHRAiwpdv
K4xCIan/bBOTxYrOeCDTL/47boRmIt5wMwbx+HZyCCYXlGCNaDADxWzEA8Ss7WuJkF47ibmRfuVQ
3TO7IeqnsPueKnE1VradYh70dSQOKPVTbPJiEiRx9ltJcY/5Y4Qxl/s68fdviATynGxOT1j1qklB
1TB0qXXGQw3PO36W+1kpATf12rEIz7l1FREyfRStuRb/85LADiWdSkNyPOYODXA9mHuh15KkYZWL
3lgVTNnC1GQtdHBHLpiBTKr9DfzARADNd8y3e1nY59Ci6bEBlaqwP4vbizu9gf/WSZNYAwhx44Kg
b1hjNQkrvCY6ZLZusJMyyulqhHTUqUZKBIWnYCEYex1yV6VPvUaIPzy4o38uyk6Nl20Adw2NHAmA
b1AeXg/lpHFkGV3SMsSriY6SQA/GpOFUwE4+bcSHoTtDcwd2DxBRTgzRf1zGZEJoBnY7e84naZmy
y5hjF0JpvxuoGnz9ub/mk2CauLvEgKtpPbB3pcihY8PORDMH5SONtyQ9+oPAeRbAu1jx1lbQ4zcY
kpOBa5kaBY0Wukk1ThVGLQVD39CUM9/ni/5GaZK5WiTl9hHj59msWqZaWT3QU0Q6JV4U/k6sKFYy
+8L6NX+hnJi32N1QSEPSUzz71Nh/v+ksfljQywCWODrjiZdTvmFjk5nZ8kUuIimjsxVve/hc0Gc3
sNHn8tHAqaKOkgNhuVLlcRlxPB7+nd7OUTdUVISx74o5yA8+f0xASf5S2/kFWYiM8TtTXI0fGGvE
9RHGGFY2fR6EJ8pG6Iwq5s96CUKXYf04YFoBLMVlTCUnpXTw1+NLxRLfS6lSW4JEq/B0VqJCnUvj
yyH/erYrx3406tn5DmWZ4z7jkSxBt0tD+8BnA+7uiQ9yar2U8AkgyZst2uj3ltkBE8odOveBu5EG
s+EuYF5BQcHzTAa2Oe53/NS49Xkl0hijJt7bRINMGsbSXD1AO/c9POVSY62Ybr1iuQ2yLBcKKdI6
nwojhTjSBU4E+bTZ6TENSp3zdKo9VJe9qf3qtSTFTtDLbI01W8mp+0bwUHo43ltlLHrfbwShQS6w
JLmn7k8wtB5neKI2tzHDhBi4+GX0fd5BMq8hxXNXnymv6O0U38Fxeg0hlH0gaePmM/AhVqR0T+bO
eWWYp9StlZE5fJN73JxvgJ0/iryk2Yub/lACVxnAS62Hb0WrTQp/B11DKK69fNWRhxyDGEo6qt86
I+fxXT3DMd+pbM9zHiyQA9WseKj5isH2zv3mZkKEDPRlFEj9B4pm25UU38Z02v7b4zhNDLW3ujyI
jWmOAXTiGmkgtEIM1ZcMzbKDA4zoDbkqf7iufWcueMc+KJrtKujDgxXvNdpPbo1g5iTQGJByWHFv
Tju12fM9r/BbaJPe+DqzUssx1c2qnP1hq587OiGLX+mx06F9GRWtPttb51jWQxSfp49lrrbM7m6M
ARqCY8wXj5mRD/veybsYpJtZ2TMxQyqH1LWrZJf8nNAznwkFaStDKQA7xVgw35E/2Y8IG222lMDB
dPnPaCrbMHK+RhB8KAAQvUJLDLLr8kpALMbqzU0Xcv1G5yrzfd2QL1f2lR5Hh9uiIOQ+NL+PaByO
WXE8bQxPPBZlTPI8bZI9C9gdw3FKwKw6TJnYME2Oxvyvon9WpHPx6NZbtegD1DxhFlz12wwGRYZR
SFdMeRptdv4WLp3V5+nMn1VeYtadnNru4jz1ZOGOvqL8nBaqIJXhQ3C2Vn0rgAOc6NWAufPKKvZv
bR1GJ1DqXrUChi9Dhj1XKZ707VjSztfHJySFuOAGIya1626sR4JuNqCpmmV1bXjlSwIqOmGXodpn
1/NqHVXAb0OkVVtXk7KfUEjqTRYDHNrgSfukGKJK3y0rQEROFsanmbiyW5wRqhKdj/ZddWwGoEug
YGSYGtJ6m1HsllfzS0TX/vUieUTd/4aSF7rMRov0hgZGEGEBUleVkRxubsjGQCGABYzbD6+joH3D
KjfAinbl3193c3vp8sqWgsNWNQZMOc4vxk90LGjnUzqombSJVdL0/5aeBaC4R+M8U6mErZ5B7+mA
/xJQ7yymJDwCLGkWTz/JCgivsrA8ejtVjCen7qY3ZbtaBr6R7NWPHyNQCTxYH1JlfP371Eg/bKVX
L7a4ncH0PS9BvRl3XrtYRSpLK1c1OFNxd2orb/A5Cm5CA7pYyXrN92m7tbCdPx2Nr0sQifVxyi81
dlFSnofKXkp+mpNkmN41m6cPBRN3x7A+LwCGo8u3Gqx0t0oI4tAm+PRgVSYfOF2q6I8GJEsV/sCX
h5ApZsqtljv3T/BsRBBDAFtvkBR39wuf7wcfbwNC+kSrsTWIq+ZWLYS6oNmZoTS4/9u2/CbbKWBJ
HJMnDEYf2oz2AWwHZq7GtAfAgChSg/RhGUTb87gaBQJ4pjgXg4CdHmzKweGe3nAGcuvR1Xt95umW
QIQZYL4QtA/URUGwGiT0jOLm6M4j6PTaW2C3MendLgJkyHj2b3XSElbzWZ9OT1IzcPLlop7cquvW
jjj3wQjKXrE+0nnQ+HEA/XFa35H9QW2heGc8cmUuqs2ytpQ5n9HY8D/2+x59amRoutPIL09hhDIS
soWgIPs/2DQVWgpCruqqx6lfcLtJvHvInf33tD6ILnyxUs0QpW/b+GxofEF+S6guo1C4RQw5z+LN
XMQ+4XyBwI6oNZYTEtf+C7aISbFZIUUdqhNdW4h9Oq96W2oy7GjMkSCkR0A4UZZ+64Xtl7oTL/Ht
jj0x7BtC/b8huP9xw3q0VSWrHC6F/3qMk5CGg/jcoyNgJB7o1MVNamcppusZxeNy2dI30WE5HsRk
eR7wOaAOlUNVyxyySAZzrpn9+HZwrT25zj/2bHi7HrK88MUFL7bZITIHEN+SfJtjPhYVRiSRCxvb
gU55Z9/S3Cxrsloa05D35DUpM3WZSU5SHrpZMFPEbOUlRTGrBJhvKfC9NrlrneK8k30YVSAdwnXx
8SoVUEmF+rLwVHt9UbTa5ZnVsk/Ras1KsF0QEyk4c5blDrTE9djiuOCjg09I6Oz7MBacisL79DCo
CQKp7R7O9lCkoKmdxBCaRYgoyuDzXQqwTpw5X2Cb2GW0gFWWlu9TyIWVGIs3KLxQMGL9+jMknbuc
646GPqx92cuh3Z8FawG32Lcrr5gRGcLQsMIx9kAtB73Snt+cWuWoJ1whtMWt7ui2eXfiTZvT7XzX
8VTy/3LklporZNp/Q3+zgDXaL9meErqImi8ragmSYQPSjjEl/yt5Pp1DYl7lfdC5x7ePqHEbbQ+l
H17nwz+Fe9hDkqUA+T45K95Li0DD6TV0XQufR5eQM53c9W4XMvA7t0rtiV7xMoalh5PIj+J4elFK
FegkFPVitCFzvT8sh8GuR5IECs51vf7E6jCRlZkY9Zk0A4UcHvql5x41SrE7mLjTbnM2Jx3hIENT
4ILt1SlmB5K3ZYy0OOJIDwTeQyFwJq2OSpYL1QC3mDCDghYn1BVre0Q3xRteayyLqf6jupLKHiaW
Jz/6PUu6CNrbQhbl2XtaDLfM46+OGmf0e63CYDUEBOAD3mYJVcD7euo1LrIURdzLfJGVrGG+CDsf
g48h93MGRCKSFJKrsucIFS0jjMDZvVCk/h+Ax9PecTNGcknR1lDH3v+54xzTpNlVFYBl6nnr7pjg
fosgI9ijJ3/vO3kkkdacDces8/qmfD/7S8FYn1clwTcQdZbqwYLAjqKmh/A462Ea4AAq/53JFD2k
zqQkQl5vhY2Vi+q5nqtURFPimkStrZlpjHe/jZRvD4iIQe6v2ZK0XzX8jREeqhTvfXRR6Bkpsvbs
vCojEZ1k0NM0U9jrl1wCt25Y3z/EcdMa1W3Z4Mr+Q6ILpsRV6y9UGgOkjnz/lUvJsPT6DAl7fCUV
fuIeRxl75PQnGTgwI6zmJGxZVg79dZ4KDnqsDpIMyOANKTJU6pIZU+xoe2cD0VHA8/RMLAf13LvE
+U5yCprtK/VdRZ1/UbpxAwCj0diBdI9XXS6FTO7kyqp9qpP32uqDaTi9B3ynx6Qax8cu8qFDZBow
RYIolkidDGYE/+a0eam0SRmSA0EQZNwcjqjeGyOPbicB9Ut9dZMzFxQaExUStcNQ2OF8dlh2qXGk
dd2eIUChsM1206Xo9wTj3iuv8aCTzsv4gyHSYLHLNcHcCv15or9xc/tZQ61lnPU0cVIg3FFdUhzy
Jendq2CAnEs716RkeqFFzjCRdI+h9yj5lBYqRddDEHt0FOHEiUfQdzE8g961vcV/OzpfN1LAVsHn
L5bFPQIhw3RzPLzGbUVSVV+3taH78kuT26x2IJgIuaRDZri0AkD1NY5xvHrRdS0mn5L2OX4UQe6q
iG0XIDLtc/ybgCGNqxTPc4nIfoULwUK09Kt7HF4+lzX4i+8ZnVXICZXScwhsuHpakZ7uGOc4pZni
AqIu1xx4VsJUWYPcHy1oadtki6JeJVbIBsicnXF88Q/KD3WBg39M2La6N9AYDgwN/8+iYTHCHzWh
H6+16Z5gcfc3TlpZB4ZiWkXl0D1KFi0z3tOEoS7bbSEQAR7VJIHQ2Xmh9378wKAZPyEOJKMmT3Sz
E0bOa9jbTBgwFxngAhXrH8hF+q0mq1uNATfHxihhXlKFoOuCxkPd9f6NwrZhXlT6eYoILh3yrn8J
LmtT1WaH7vB/VeXD6w73xxpc0e0vJpUD0k5Mq8QzCZW+1DXk+oYl+oYNUJ3ckojxe4G5W7NKXAnq
Nsaolwbxl9wca2Py9TuWJLuiDBiCYsHtigFxJK8FTTMJkq9bV6IgdVT3BBCZDudgZM3IR4Pzmydf
cy8MTrZmb9b0IX6c0FSWxj3tBGGMUNPWlAim3J3soXt+myGpEbImRjo9QAfRTrhrdCyp54xDjBPK
6W8BBtkOg28uIk7IvrWqHzp5p1oePPXvimQBhVVMJNABMFgfIB6kAJheQiZrdPJ6xsKriPXiMdAT
E5HuiEX5qEudmagHCWrfdykb/DesliY93YRS0UwmGLvkpCpMusjYYEO8YjeNIG3A67rjQ9SIxTBp
WIWfsT83j1/pnu+CkHkFkhjA+I+ijFrIYiAbdiSPXa59iDM32YR4i5BRSK+vxFI+bnD/03+j8zZ1
cs2FzAcGlUzz1YvKtqzaXoby5cUBprwg2kZ4WkLVJXvrNkHSB/o1Ix2Z9pgRgzt/gl74aUC/Phsl
7XUQJEzpLlFjWxLJ3VVgThCLWndxtVlmTQKHKVpkeA1LFeqNNX/5RP0BCF90bmlPp7JBUMJJpgyd
PdWPPHbaZ5lh4Ewcm6+9AMSVFhaNqJfTVRlYF7BITZuaapaQoEeT9SzOTlJt56tQ4+U2ElxYyf0Y
ppainwbHt6hTfeQtpjhCKRzyvFORWweRpPIBuZ1TCYa9+QmOhUK+iHClABhs1F31bGm3SKjPpFRS
6LXKaTfI7hu1UECBpwjKOdOueB0aALErz/R2at9ZpWtUsvjuJY52kpe65z/ppAYL1YQP1WO+Ldiw
WLRim2p7T/E+qbf0g0urfnEqn689Zzxu4YcGuMzB7YJFG9tE3wHs7ZzSqSaNXK2+jJFk00qqRHoZ
sY3ATllYmgojE43YlxphGLl4B7B6FGKNt7LxifUhUuMU0B5PDigaDT1v5VZHeO6eId8qkK+HJa0n
ZJFuun4rjrUCG5iTV6dHcui2xORPHHyeoUkdAWAoGDZVRHhMccTk81WLC42GQg0AlCk8HM7AIn9B
dAHV26Hvwz4660UZiXuEUPbj0swwOziwEi5g2Ua+SrntQ60x2MrtcGXJ0x5ha5nPSiPzdihth7NT
KnD74HEZ6xXZGt8rypXvKMDhjJCnLQe3sQDaPp6kS2oDleEZluz9l8Ec+yBlJ29+40LVn2ETl/fC
rzBuWYS0CA7tgXw3k74TlUugmJHizRTVAm6vW03p5X+aqM3KM2DjyFN0smOE418gUFQTTT/S4X6C
PeVWKyCljda7S6hWXUI7GdaRgQJPuwk9HBq4fpdOFlHz8z+zApjl0UBhICrSsXCaWwVLjo5XUaOL
/8wlFwoNe4SbJg4euJj5VBYUuQwsYc86BC6TbGsE5GHEeFiZr2xLiX+KiXAglC5yoRW1MumLZROW
+phf5OblczoQCWZF5s8VlIubcOMF/7kh3/8G8D+BtwG2GOzaapEAq8mITWhRKfNl2yoM10koV97b
K188pP0EbpGJXDLuelsJTSafvt+lRQMJgqUgyDH39+ktIhgiEa+0jj2tN8B1OFiVCmPhq93aeAA/
qP0cG+OR3dR+0ZJj5NYpevD8XtU7rEYMbN5gITnxko3I/oBrnqlV3l04uzqkfbinYTBqlLFHp4hX
Zw8Cfyvk0VqWtCD8D9j7q8i4oFHRi/JZO3Zdxtypf271bgn2rI71ltdAAh6IwmMdsbQyii55puHs
RwuTpbB7vJe3XMRNIoLu3X/6lfrDb+eYDDcWk3C5L0izdD7IINvnMPD8rkz/+isSllGQPe7yOhM6
gQys+4T0kQLkLZ9c4CNurlzX5QnZOZg9Nr+7dtL/GEGjC04sYzF0R0IIBG1f2ns0v9TEKKMVVEtQ
uQizDSz25ERk58g99uxANUkW6mVYnR1Cht+acppSGfDBaGXrRujj4uPiWJ1//3knbuEaf8t4xoFo
kUo/lryv0Hoyp5aJDmtVZ3dnhNwL8M4y9YBphXWhwtlQfJYjFBqJM1lrCfezMHKgViUxtssaxy3k
tvyOa6wm8OlpJZCKPmvnqIZUkPg5HEqnoCw3+xK9qgtSAQh1nXZQl1dANDjQlNhgvzgZVilW+E1A
/BaJhOvnNuHtiCBJcacNaCWUhF1IplzcEMUKJhsnaSr+dsEn4FooLPZA3Sa2DI1q8wa71dS73L+s
GZrbtyxiFaa1f4Yl06d5/SDsSoehe26zfPz1Wl4YEJjJoAOclWxntp21nFX3k/7bfUwumioC6ePZ
wrLwGdgQdBnBCThxnqBcY2RPUnziz1perNag4WNUiSTrC9iF0ByXkHhb0M+DmjsOeju9ljHi89/Y
WqysNw3VhXw5CaTpAboANjtniB05AaU8L4euwXJKhKmgjZ57Llw2vbeSdYSlgkIw5coNbFcJv2Gh
iiwo+r+J2550b7havMmukIUkAX7ZPzDxTb9YIU/B9ngeJh0OOkxT5D6jX2+gXvMR4FDhX/pKefZx
r1soxcor2WZwUwbreoevQmS98CNuEOVODInKNj3R9mMD27n5AXs7M98hxQ7SGVzeTOgQO7OrS5Cf
g6ufQqFnqwj2r2MPUbx4QMrU9EcF23kbOt5G5BW3nQ4xD4JyrUdwhlOxjYnTgGNzb+OYJeQMt6OQ
Cshf5291vwRNGfPi/GU9aShfe7DFRxJF5pIFSsbKEghOkCVa1mZDOYu7TiJBTsndVH/j6cyInDmp
AHE+FriWFFzEpAh6rbbJ7vAeizDv7Ag3g2nBaWAqZJvCwJMsEAP1E8/xnU3glRlyR9l6cyyYQArc
loo1gsGqKNabkaSN2H5kb42ZDFNEvj2S26i6dTvUrEevkbmTxKd8gdpSqpc/S65o7RRllouMX8cM
yTHx32DGqK0e5xrWnR1Fqn1bV/NksA109o7eagsqDlauOHtvAw41nalZqyieqlWpaWRhOsVrsN1/
KgpIsftWTnB+tNSdH2h2cSLGe0ysle7dqeYYQOVgxGFP45HhYnoWc156MnNwfs/4PfQy+mWqFXtk
9wxHM4lhpQ0kG1Il40whkhtXhDEtlYqZMFqOFQWKncz9GN0nZu90aOFbXnBheem/HwaR7cf46jY3
BgCfLr3lA8t82QHK3BpXIBy7+STmhkMtP6fp6JpZ7BMj9eG3U9P9JOyVOFeKrshsal4xv5Tuxgzz
74rVRJwDl1KkaEsXptXcb2JxNJaE92/msEeCvKATFDT8r8zRUp+JPYYsPu5n67ZWc2O+Qxuvn9TM
EyfgEEORaDAzRbrD+VRGfUptNv0dzdaZ93u1yxAofj19qyWAr6NNNuZoz636Lp7nDQLxd9gTiq09
j2nnhQSkdrNa8OQQOpfh7wIfuPiBHA/fodqIlM4j9ryZ0E1uqNAO44+i2Le4k8dKdbfh9lCXZUqO
JwPTbrsE4M70PWsJsepyd+W2qyuoi1b6kUySNp1FmftKv0L5Vv48A63Qw809LbRSUbbU6pqoAd+3
riREDJZeKjpOFfq/q8LdrybZMQw1Wpd/HDMGrZTaNAPu/nQxOXOWsxYbz+o/MmtGbA+PWICVjNLP
+sU1UJ9h0+qOOUCm0FYhsdpGx9kcqdrN/c/d72zCwx1X6fjWICOJbixhLBmIbOamxrYcDX/S7tp1
hTARF+8txEvxBtWT5ZYEQkJkpdgWkVs5oIzomUEyeGsiSIgfiOyA+Obkud1Jx6R9yJYcjWs4d78P
Lzh2Nc/4l/dQNETcb8oCb+1xHx/YJXaH0rL08nqHYAAT0qVZyynlmpGkkYrF1Jq+dgqeZcIWO3W7
F2hJxtd/zw9xKIfqCb/CLqXATCE5Ay5ezk9hENKLWoYN6bYVuB8Mm8jL1ZQYVBaIcPJ/+QJ45HaX
0axVhd+08Qgg+mcc5/kspWnozmI8lb8qva+4ITYgoiiQcMU3s7GmFYXKtSpo0gepGWVboiglCXBL
nSWG9OQcQqUEqRiafKECUe72nnWRaXD4afDiz+KRelHL4g1ePs5Xb7tlW68c6RDoul+JExCnT0aN
51R5qgOy3Un/QaCw+DH9G+LBt41HLPraghmy81uA8FjYQPWSG2GBwOhLgyeLjoWauCG8sNzOqIpf
isz+lj+2VmCBlC/z5Mnm6W6j3Iy6fg7rQSZp+j/azB5ozKsCGhsgbxS2Xy7dWkOWWETWb2/uHqEg
eDkaGOiT33syr8HLf3AoDncJrz3bAxBPZo51GqsRWBzhiC/qDjOOBKP1ib2MU4fAb4StfqfOlxYp
Wi2UxDFgUpHeTIDGGTxjIoeu8AdXVhy9DSz1+fLWhQg85vAmoWjW4/9WevIVX/DpdQl97CXCa1Bs
cKm5ZMDr+Hj5KWGo9s1947H40SVx+HePzz6u1W60gLcEuyS4TfpSzM359Wv85pGPSZeBbfU2r5qF
b3xywVpMW5vs/Gf+z5xUBMKS2bdiVRKzCjGnc4FVAr0KXRCqqhxkPs/Cn3T+qhVO3nicAlC3voBs
qzORf60Y4qHkFPpGkCX4vPkVA05q+YgUB85NrnwoVUuwwS3mcEqZE23vEpXURoD7iPcaMzrcGl9M
clszuyHqPUdOf9xVauRcD/p1qulGxNerB2BgNNCI3HDMkq7aUyf8TfJQ0wPJTBS0xQQtxNMxHfMu
Qnvoho0U4Lr+plsfscujlmdXszNlfJ818V82lroczFEoyo2zgpyfgN67fmvuouHs0a1oaGeR2y7+
j4v8HR5otSmd8fipLkdO4zAPTn5Q9c/6MRA8ArRgFPAEb/bYIk3JXeMTnhLac3sOI9B99ILVrkCN
ykHf6UYcCoDBAPMdEXWMHXuxF0zEXVjr0Qy/IircKOLmX6dyu2hRKPUI3ijrVEM5SwCLzuq9Vz90
rF5YCN56LRRda++Bl8heTq2wy7lANpbpYD4zh3QYV6JspVEM8l8XHtAhvD9hMGnjVHcjjdMTuYd3
7LzQsKcWYA4zYl6BlQecpRtCSdoXElMV7QoKfmQiBgqE8JYdoynluqBIoLI7aGddWRV6AmN2eJfv
VNcBR3w0/DRUoz2fLP0lck/s5NQBuSjesGJ4EoL0IIGlIZE7HbnUXx6tPcgjGURIgazEpvGpT5kv
8NkMM2M1whLdrPk9KjzuziXpWSGGnHsykjtcSo08XbSv8L8kr2d+AA9yjiau0Fpr73vs93+WuJJk
CparNNPWDm8DQUhgfVYJo+VENH/Kh9lDYRBFumqGNbUpNB2bj+ei6Yi6YTxO+Nd+q1aE/Rlibptm
9wHjYNLY8hcSkBa3NPzVo2E0h8UkDDUAMOFYaU535P3mTEXHcCrOnVwum2W/ZaJgYcFQE0zABElI
zjD/j7yuRziAZIBJ9r9m6m8pR9fLqGUmrxOI2C7zg95LTN2zmdsIsz55zqOpdUMNiYwCWckqpeKk
xtZWSrXcv0c4RfglJeD5bl7fmqj08OCIzCcwyxPM5V5Vi7La6rG05CzaqWT/jVQvUYyRNm+vbJAF
X4IR3rwOhxecqSDxn7Oed5A4/zE9iv5rg9b9saL1oz6VisMEY19hSYU70ZnPel9dpkdFjs6J14Wr
hoVrvjVvL/WL42yQe/QlYRvzGJhmLve4xfjn2j5XkpNesgHSvLCD9+JusbGg43vGPOKHoQUA4G4U
iV1542EB2xLZWCWmOufvL5ymMRZ7alMaWU8q1QjUhlKHYCwNBmTLJY4K4v1xGmI2fCAy9mpa/daj
WB7vJqGyy0kOJY+xXHjkzsTAU1h+HDqR1DHGajHzpSaXFIoN7SpW1eKISWP9QDkc6t+EEmtA1Om5
b9MiihH9yq1GKjH91O3jVnvhsxC/QNDEh+sXgpzGgq7ThdgpXH61DvyrLhjx8gytG31VcZIWA5QY
MpSy7EfvNdZD616KFr/4JQi7zBzx0/d9fkQmLn09r330cSVlGgmrtHobMkUZW3SaImxtnVA+ifG7
ShmYtjhu6zhjMrKPCT2G1xmyzwVK5T61bZOU4Rbg4nws348QqPevho4Wdues6Wf0JGQTHp8vtMaj
/eM83IggNSrRxJpEiRYIA/c19+mH3fXW4vPVJiLYGqm0bZ9qAvAoeFdKW3nxhmELptiZFgzaxAnM
lyQZPhKzGZ973PSKHfuHycmpvbx/WeEQA6a8H8ybDZTK6Ig2jOT2aQHx51dLrQq7oBw6wUI2bCF6
wP5d771Tss2QfQJ1W/135sNJE7PbN+ml+00QjmQNZFDYpG3ZrnzC2SD55UeAdu0OFFt/jbta8bIT
LbMTU12B3/iBGwrykJH6t0iLOFHaQdHgOKNQkBcV7Uh7/zex4BMPZ/tQZ8A5PH/MMy4MSUMMefIP
8i948EV4Vd3hkOEzvP1srNHGhM2lW/NVmrg2bBhEer+f5R/hyah6VRaTqcQTaJbOC19ZGSBW7eZV
Vs77UQKcT4rIAvucGAHpJn+P62G88SI2tGqF2xcXFFn5pijg2HkZnfjmAXZxV71+P/J2xjzoICXn
IdAARZU5/mkyG+4XkZXy44cWC6OClbhYRxpTSSngtHW5uGYCcGs4rDnFHR6EMMeYl0pLTJEYYRKu
SgnIyWlk4/XNPigf16tXh8ImCA+UdNB225zhEt2Xc/sG1puPsHlx921OB6DFO9DFfg7lbbiJ2H/k
v53Sj6ex/drusixj6Jq7zCOIdZiQ3GJPQV/dV9bLOU2k05aUP+cdFPAtiXiQ8k0v4rD++VYSZccG
A1quPSjrzJMJFZaMj4f5OMhbNDzMX0k9Cf/x5wKIZOYuoWYrhVJEdZjw34YqWUKE4aqBnFxi++sG
huIWYDTIPKMTq4T0oXbSQYHa38LyUAGyP62zWgDkGLMX+a3IhGcRGfzBm2+XhdUM3jJmGujkKbKj
TMr8qbh7iJdJFXCejWMUVNO+lJsNG8RgMK6x3Cr3NbQT2X8wIW5HRVN4sOWIRq9rCGR6e0ccIpiE
l1Kr+DqmWDeT0d57eteZDfQZphT9LjT1n13RJIWOmX3PyLn7lCLttYxqqkZrnCVoiEmMt0DsFS6V
R+fn1Hz519E/7tWxyv36xTlPtoyW555KVCFP31YX5VWHWxezBXif98P695CDgRGM8xqA37k+sMZb
1ddzyh9RkxUHvNhh4khd7SQxEzx47Jta5p/Ai3RlZQJthBWvPIE2t5bMQBUL+8qqSM1iXomiuR2m
TIahcoSMrZOLEB2l3nZavg/++5u7JWO2/fy8IiADYx+dOC+PEaAk6bkEo/osznvuaXYWoB19WjmG
VqDW2nRA4E1Ksxd71UIUo4NDgBB+bBVr0j9E+pt/bcA1fPOPlcSLZfFqLZHwe5vfDfC5fggDGs8O
DPjxwRvXdi8+hBgenAIHfrqypyZXPUuZ+XGZNx4MbU5jujFMlB6Jkzle26GBuKkzMLoasH813lr3
5kTsINvko4JyyZ3k5tBWQXZ2++pPf3d/NkPm0I9MU/XP459yD5nofcxcT8IxFjsRU+G6aXAMp+mQ
Lsq5noJgrSz38fLb6GYP2f44ItmenXhXywoBz1xkxYc4SC81m5KLi7/x/LJm0JX+9PzjYQtbcMpI
w9tHdWxeOMvxbkZeAuFn+OfiEruVZX6o1LQqhUF83tIptbw4Kzuyo3OkAnB95bZclLSzWiRIw4cO
QtUaz/IwL9nboWqGgPCIMwgEDj4AmxlPb7ut3DhuBETI9khdU0KpHUCI8ZZJ6xJ2GRzyD1A10T0K
d25jm+j2gUmfRmB7gEqz6r9jdNLhPu93gF8AXPa1sd03fv/mtwVrW3kWX6Zth2fk0TNLBrHfhj1y
Ve/xyebStQpWl8BetnS1NbXQ5i1bwpsoALMpDJ9QkmI60kx4tYSkD/y/0K4ntAVcKd6OxOKCF4aF
idBIkZHg/J3IOmz1NF5NSyIRYy4Ib8CjtcNN5sBfig3vXwC+QQLebCMltPW23eOCbtsxfw8ohH0b
cSJKjnorzvZRjdbndBsvS/1qXXNWK5vpz9oP7ff1aHRbPYj5DpZpGsqkIsbHU3m6lneYoYkAGpT5
Mq7i1yqsFzBDiYsljKTdejUIha12o+toVPrX1yWshb1/8/TokMgLrHCRT9de0xvCfyxRowQKhqdm
rqnLntc1oVWFgBpWhIprtXZPRiKj99BAyusRO3HBdLGwke+fvnpoIEoXNnj3kui5maryVBKhHkLw
DrmixUMaT2xipetcI6Ao5zEIINTL6tVYFMct+yPknUF3RjAhghYqigYwYA81GVrBNSV1HggkQBwW
HSWhSP7l9O00iV+eZTNCNSTAk9X1NecLw0bhulAM8yNGyElezzRuMeZBjdU6+rzUwUGH/15mzYI5
y1hvyEumph6QwXgMJqPjLr2Qoe2pgYg9X6YvtxrWkTEgB56LmrokboJE32hKWHwMh7piQDhk/L82
fSLivbSCOoYkBgQ5zBV9QjUhJBudz2XAohrCRRWZjLxtwVO2nTN/R1HDlKHqf62tkT2oQ5g/NvHx
QsxAH739hQcG0kmepjfy0dN2yW+WZ2CQdtyu5DdiwGNER76b/4Mgi5w2AUQq/KqYkVn2BM3i2j7p
38rI+weN9BwvcNDE9DcdHN7kssnw1tj8DV4SBES7qjOmEUQx8D/5ZwYNQyU+9ljSxi5PJS2tG1WR
psGfJhfFzmt3nGdMK6rAnihvWF6eax/YpoID6qYWho0mDPo20nzrLVCSdRALdo/xyDnX3E1Q4HiE
AGxxiRNlPZy/qCAAto1VK4iGrEVIL+Z2etCgtN6/HULmKApjEcP8XQnQPoMNeNl3LgnxQVlcZW3F
r57WR3b4ot1mKeBwqAEwaO2ANBP/WYlj6L7Qgf20suu+TyzDeZEPGax/Gsk3VMhvOOzfOIpliAZW
wTKClMe0icUXIFghQI9TmUAKX8AydpY2mh1g9JHNUWne/cGsFsuDERjjqycdTxTkkvZ+cmlkGQTo
E2ugnU+5U3UoXtiseFOGsEdnOoZwX7CfpA9UzwDsEjlTN0/r/QQrvNKytN36Za8Fx+0tN9Utmby3
wyzuIX9BovRippVns202QyiHgELLzYAXX7JkwQsaapA3Fpb8UBJZXo9Df7ueZcO1zAISndWoazbs
dDZy4xSeWDONs9xXRm/0n1CUjGqQq0R8TUMaHztXKykQ+dvwxlHU7SubI4nlV2v52ogUp+RPlj1C
khkcv9r9IPBR+Voxpq74Z+4hPVvE28oO/71ZgdOIAIp/navJVALaC2QRlHizQHzP3pPm9UsNe63K
sDRJ/VbesssrCkz6jwbDTfFWHwfPkAotdBcnV9no6diKyOO+e7xENQCTRf3gIujeCkTjFB2faeI+
UZAbUqoo3UlkEryROMbRL87ebygPLj/olWmBD4C8kAEJUzO653ZyQ5jM9Nq9fVTyD4eUnurY9be7
Wf0chXxtBaxX9OnwuPdIM3+ZriptUzbTxwSF7o4FyjoXWRaCTI/AffvMbsDikletktS8dpMvOoJ0
iR4/7vHomQZYpMYEDySTLtraKFhVOBo8H+x/ho3DaF2nqMRXdGMMm5W1ZRZkLK2HjZgOuOqaffv9
VoPipFpb1dprEgI9FmKs8vnBvxw8v7im1k1IHcpuQuNiFUyTykxvFVyfDVNQOoEkgXIm67evEBoI
zJUd/AdXiNqrHa3agLZgYh0zA8egM6YdGVv3Fg4c3L//QovVeml/+YnhhbXbxf1Z9+LNPwyvZyhi
iGWIbSxOKa0iITl4wUd0XnWcdo2oPZ+n+qVOsztd/SaHXGC1AyMYSPa/TrAZ6eHaWpGuC/LMhbsl
fIyNKLHIAlAwTdaShsGzTFEn1vuEGrlI2cfHq3VgQ/jWNS9Vf3A8Z1hIjzAQRl+6FXHppyq+nOsg
oDYJ7CJWYKqkmEit+Md/YPU535Pljgri7wz+IapVo8oInTdmBv3V4i1A0ttnvsOfBtQa3CXfRX6w
Cb4kRTtiQgnXz1BF0DeFvzkEyYVYnX5OjnEa5e0HG1I4S9guAR0T37VCpqa7iyj8dw35H1ykmRVz
jF0s2hz/c+ER1qXrZsS0IA+zt+qdpTvbApGCpw7z3ZXPIYsVsh9hlBKnVNM9AQFQA2c5l6YZ6SwZ
908XaAKR6b1bGel1gCyYkQpVGO4bRI8jI1OKPglGoegOVOjhj/fk9Im0GRxIQyUxGzkY/rwjfVN5
bDmP69SGJQYE7obRjKBF5v0tOGUgyWv7Zm3Gf5A/LsN98YmZISnCe/CTnfEB8ILn9b2V5/uh4AP0
BOa5ijPU42c2AogFXUPFmP4/YK4PfrXfq1GW3q3TfhWOvU1XCPrLOvf6Qz2YkIibNlxA8uYidv3Z
fGgnYTh8ubcgqY91izm62crIEAVbhyuKFsJBXFc32b+z7//4tfUGlSes3R1LASBIucZ4zcxuGbOh
p832AlKhPaRPE9LhD9fn9iQwY2DHnbBKZYehe9d2clSjC7im3VYfW4Lb1iXJ7thCxerWmtsDYGgN
lo6siMMEjIUXuLSgUUXnfe0TRJMpeZFbnHFBp1NemZzh70TuuDhKF+gbhQIiZJyphXrxbwd3mDN5
+HNi+oTXPIfhDwpLzd2DW5j6+FyxjDpbkrVv0s7gEwaR4KbKP5SsgyJRbmBNesG28kRr2GXels+g
WAuqFn/nozHRsLNE1XWdREUaW6rgiWZSP4Fzeljwc+8cYHT3QIFGx2mWMb2dZFqvouNUqZCvTvV/
8W7NEyQ2jAIgPhVdR9gaG2+IfElOfQZ0mBQueTJpd4UUUpuoprTkKZodF1Mndo+t+v932TVuf9Ew
hLKuXDq8Ep2I9+5rkGIyX6jl/0syDeAR1ozcWim9MzsOfjdSP8VafzR9RrfGqSjeuVVjkO7BZ4v4
WOkjN9H4n2SaNgOAgKEXAPchL72trzWz5e4aGSr87X9jftTFUQ0P7bQ39WuQGTv6koDdSkqA5Tme
V6Y+++3mC3hEqp+PPmYg2CZyF3Fty/uC2XET0wMV4dxMybE7nxPSkcEmwqX6UmUm3iak0bAQDlUU
dQ4nDvQRw+7twKPKyuwV4or4x1xmmHYiebF1KS8KnqkwJDM/oXf1D6X9DABmeN6a/wotIeEymtTw
LnNkOsULlYWaYF0+V23loSClzMoL/PkAttyY97rvXhgmBU62vFkAhGwEs46lRpXiuEvlYvmmq5Fk
nNEkmHGnM7uq2QzBESZagx3hDpskQ0qxjVDm6M+QCSIEDGlwigTcG78I+NydXyl4QTHwAPaTIhKN
UM0pTQinCKzqqlBjSoOmxvtUx55pOoGaZLZmMRP8B/jjqjM/mnbUFQ1NF9/JV8x7BJF+Op5hIXMk
U6tNaih55Ghm5XaUTw0CDk97MuKXHBKLsOTT1jKvWfoosPSAZuBKCRsynpKbw2OzaHVvp6xui6Ne
mVzvAGnRMyPwCCOnalCStCpHzmwdlzG0J6ST2k/Tl/bjzzaPK2y0mqpWF16NatntvnPFwN6wCZfk
AleuuTxVND4hVXDxjPwQ8hJ6w3CBmNouCXlnv8reM41Q1gEhpMc9/30yvs8Vjgrmib3Dtz4g3so+
GPIaZXdyh5CYJhkIM0V5gjVY3n3Cgeu/SHZOQRJILCBbl83oLm0wBzMYPEL8/zHm+y+xoD/2VFK7
06ZbcqtL//+SVqaJB6ol45PNG7+8sf+p3/2Ymryx2xE8yt0KGLj+sgEtkDA1oNXkwiCY6llrS18K
O96vWYDvNMvmEcS01BFlx7yXIHszIpiwvroh9V7CK3FVQgEJ/H+W8CltAo6dpuLK/oP/Oryc+jED
1UYG6WkzZW22n63pFchuk8iPO9ajY+ApBmrXZcouQP4vp424AFbTxksc+PSQgCVcpoEUVl2bBY8U
sKqCMXpPmlu6n2I49Fh/hrCjMZyUmXpKnuxUqhCRvzqGo3U0xfOFsDIXZQS7VFvF3hXWCEFJ7TjZ
3uz50m6vZUKxE0FF1nH42QWPKKg7v07t7MMrpcvF4Pr00VKhwVMiah5bgx8jGtV1q7GzE/7mHrR+
dKOhtI0K639JXOU8NGZaTxOEwTz+Fg/0lPVklA5VMS5YUjOAidqtZ6a2MuD2ajgN6icOqHQATTO+
mKWcDZy98MmVlGOTsQDr1o+Qi7Zurr8u2/T1FIpsIYUf1KZyyFhSSGQFxgVDi5/uYY0qdwueQW3s
w6zYO/2jKVqXzuDaIP2HSIwfNgGTWkyny0CiZk3MMCE9Ur5d/skyTGZOhKuYLPnpXnvLDRBAnROL
iRsPZJX9WihnxF+DJF6aept/ABvtczAG4fp19AuPPkcy0tWLnbuUKuBWmf/60YD1uC7To6kSXver
BdP0sz6daoQ+s3rIRDNMovFFqxZ1lb3s0UnUl+qXqATw3fFQjb9e3DNigxYwor7qrC6owBPo1Ukx
TepUQ45MdASvj+Hc57C1DEAwbTleUIpZoDXhw4NKoHcXA5xjwMJ6wcOA/8FNLj83B/QJdQvOTEvt
RgJCjrbQYDChIH/0pSjsZ1GWWCfy+iuJXWFwie7ysKppHtdTF21J3zC6+1rdkqfU7Lye14BsgqsH
/VHzJItyGOIbX0az26OzGmOsmYZlBay7TrZimSKeqgqmGMUadRBS1Br3hMs1Iz/zuRlv+1/UvgtE
FM02tuw6yP8QDERBo1uHXOQdF4Uld59McI7FLpHbPIfpQQr/zcPGOMBMNiTgepE+GjXjn22+Zfk7
CmzSohii8JtTGxQO768hJYvNyhHfkcgfXcNgZFu7wnW7VyzJxsXTXhsr4naLmlonWESg/7ADRiOk
VRJsf9yebG4QNUpuTDYH+Jv35odx+YHTywnTKZCHV1thKEjV8RxqKtwhf1TTCNkiajG0ng+HPOoP
IZu1pKOIpdN2yz8Yp9QCOM5nOFjL3p6O9graOJkaU7QaA7gZCn1M+UhKLlapt+GYOYBRrw+GmrTY
tn3W5jW2ofyuqywY/EVmEyCa8DjneX4HBfF1IIITmuf7SdpGrll+QmPLo46EDuCddPUv9Zj+fSwN
9p44A3fNN0WdF/7rAa74m2r+N5gj4zFp7Q1cRSyzKlhlKY79jtbziEQLAwY5asPVBp5CW3U2tHqJ
EoRa6vFi357ato5Be5ikMioBGVUlUqYYV7YyKiV6TWa1oFheEL1SRqKKBMRFpqEvf3MyaWU6xyeL
SIYJkLWWbOk/PvskZiFpaJeMhyOBNzQk9WB238q9ale6nHMiU4ZEIm8X3LykWsgcZDlNQDsJFSJQ
yKOzEyXzjj8m1UmAks6gsceWigo/k2CFCViGsWZ7EWDYJtcIXd4aODrOx2/h4JjHr/Rk4urKBg5J
se1ikCD4NvSOPSFBMZKwCI/RW/UczGgp1/bIQhWNPBAVwfsjhLqK6Gzj54i8LVOOFOuf1ac7sbhE
PEFScwvVWr1YqkiVZK12KhOpI/EbfikU6ooFyvUXK2r/WPP0hOVv4u0WFUZhVidqyt7bqH6iWR0W
1gylDoIo+CXOER/iY2aST6198VhC8mQTRqiTdV8ZnZdVzdhngKDAEn9reZZmpXX9iceS6pXpGQiq
GIzznTbgKNgiNOBzP0wPyLm7AunXSVxVAK3aoVFRBQWU1ilKxG1usMmZfWka6a+yw7cyqvikItcJ
KfrQDxfKSPoAl6WbTuSNMx/dBMxw+g5Fqkqi+QQ1C94yeyrpAaQPD5ZhC6FVHaZdoe3X+idwM6eK
7Vp1qd0QBht3igXqs58ACG6FuveycFiT0SEfg5e2e79TFcUX5ho3RRFX1z0MQvsUXRr8J6m/z4Pw
KoMh06SFeGM7srhfrQjy+TSjMVUZhU8om1uw+mLJz1C2SpRFdPu4N5AHKlv+rjGHtjqmX+q0Q9a+
+JXO1TLTicyYmDdxiPpYjoNArpLuKCjaHlouvBoLpKZFXVu+JiQzbaIZzfj8EnNFTW06dlVYeW1L
UQBGJhIqi+L3rOCIF/e0ig0SP1NYV9giuXrlGuPoI9IJl2uu0D2VZvaEVjxIxG+yMvPCVaiwu0nB
3b/zJ+d7zrYIy866p+YzhKAl/H6thUpDBp7vL4UzhC+0hRE/VUxgDERCQ+2rynHuWEfUpu9uyrDh
X0DJdJLVyLrf09mINnn/RCFkbn3f0j1rspYrsJ+2OlvX1A6W6dZtItcnmUYjINbqLug9XRr8A1Le
apMrF9GCEWRxOM9SSZ957DejfR37yyMdclmBUsRhzXRyV9ytAuRm5MUoKQ8UHO/dL1yKm8R/tcmr
Y+72asCSo/8HU7cD4O1d3FmK+jaLZHh+0Or443D2iAWkMBdO5fCdR4Woy4YPqEir/dGdO7lYNWkL
YrmnBFFDvGdgw4iQr4RbgXDr0BUBxRtWWx2YA4ofCcltg9nXCfYJdIVyc7ByEvfYB3adt47ybOHU
PjaHhpQlYXCpL9Qoh6u3Y1NDNHHhKEQPiQKBfQUqE3YHxhnq+pKewmaRH3s0erB8WPnvRDNiYgZe
hh0b2mAySIQTuDokIZF1+WY6P6ApwyalWBUb1I6tJNHaXKHJ3VlohdbEi9fSJ5dwhZe4YMSlL5WC
xDfyjSf8RkJNBmlqvqbIjaFmBlRhnHt0D604Wj5Ye0CaNZTE3WRutjaATpCYxe94gm4UKi0yBqeF
v1MgWFa4VTdEdee/tuAoL34cCaFnXo0/JRmHfOI7Q4pscI4oZ58QExfG34qTZcfFYkq8Uwl1MLua
i5cL7vQIM5q1kOxeofPeblKeH6kpTD0sY1O+l3tjyxwsr841JV4G2wm6QB2QGN94cqP775IpYR9s
GtOM4TQvYVxaiMCJh9p0D7hFy75vQvcuiwqwwo/mrw7eMigAEaS7lC+AUeOxYWDmNpfsgAYT9dwy
SwsVmSUwm/GLfmXsVZ+PSjXgqvGLlgtKUI63I6qCIyI51jyNZ9BbexhKIkgnXnUuoRQD78lcaiiD
B/aDtPCgOsne1Ewd3v6EbkiH/w4uZVbKmD2da6OwNsoZQAqK/GkkHcyKbPsFlystFob15S3NPZW5
Vwj0mcBWsXNsMSao4ppSO+j/tUmoBXVqsJLTES2CaQbm7YYHpzfmTjERLixEqDRWuD5Auv08CMQm
YtEHlgYbh4DOXtDhUMx7eiMrGSRl8CkglXp8yO4Wdvv+jCzJhyIxkPY5Ble7Nvr1PaHR0ZfPYzir
cn4AC1oKvAIQOn9QRHfUk5omyLU5DSG+z5JXvCuLkQvUXMVxHONoHJdmbVmaGaf/uYt/0m0DBiPC
BbseOIwGDlS0gw5EPGZPu5S+qZMN1QxINAELZ3lEwwOoxDsDThcs0Hi/uQLhmT31crbqoUImnF67
fAN2yWkYIdv4vhYh6Ryjvyd1HtwEHKzZSxytaAxqkGcSuKKtPBEY+xEtlXF2uiUFO/aQMTgaUE8F
m0YDhyX5pHrmM1vOa4wg3O6bFMNOowWk1zel8OqAlrrVp4BKXIAYn+vQw91L8t24vJojLobYzjDL
UBYP8eyCmmtHGLiG9gBgnOmpHKmD2ZOkdV+NABiK7WFBTZAFOYVU1WeFyzQdBAguZxsqug4mnO3l
5hlGkAlik3iI0IVj1toCBrFSZDQ1/EFP3HdCXhlQsxB+voUeytV2uXzMsPoW3zMZgjJVBG7X9e/E
hWIwIB4rOG3NeOzcBIOJdm0UfYeAvF8ifanNGC9kvx/GgTkq6qZoSe5MxGQ1ZgaShYA5/f6V7Vpt
ubxfabKxo6NqTpYfDP6IEFhqGnVa3o1UQ3lq5fwCnRihR1OpvcCN1tSnzyWNd0l28juEPP+1XXOO
3O3ENxYn/SSyiKRoLnwKbWL0xe06OBMEpggDEH0iaPJxEU7tr4+KT9Y4+8TjP4M3JCL7NbyL7oeu
vGpuH2luVEMy+1UzVr9uTzzuJN9ZU6QbgBdyaZgKvVRdjhf//NEGj8Z4RCWuMMQYn/1/4g/h3CZF
tsWbx7qUuFn3avrIdrqFl8/V80YY2B+4tF4Ne/TdGweSfk4LQeeValUokYate5LDudhtR3z/Tcou
BfdzKj/nFrTuo2ah5lCCjFSCn/pWxmGYV/mpl6X6VQRZAjrde07AsacTrkMuZ2xsc6NJ9g+yirdF
Hf4NnAlpQrH+9QdiXssqwLKtJCZa7Zab+CZB/Wci9wFY7r7FDs+ORQlfpwdM4WbNIr+IKrO9Elpk
WF5L9jkzGX/ff+YkxDQkls05mNrzmIWiWkFYUmCd6EBk8spEG3NmL0yhrhC+1qPkNKgk0PvknZug
bpK7iAbr72kPUHF9m/2mkEopaDh0PLvgAzb/B7mzwaNVZG8bHtoIza62k56CulTLeIiRcdeTdJ4j
YZBCkU31nkgqinHVp9l8o5nsnCQrzYG+BJkpkCSOsMBja2d97HgDeds68mPx+Bc2HbyXJKWWjNTW
xcsP1IYnS0I+SklglKCewMDwPySDZVOlDdNXfMV+usKk9XdXLDjG8m6Fe/1koGjhQkLxPsB0WC00
O3SFTFt1jTcsNOjtRKEpgYDRTLTsyye0gFfhIlHwUta3ghfnNU/3LakeyxxKTxELuuUh266QgNdo
a10jfTFj0GOzhiLZwTZyFcrOGVC66RcLv9PvfukR3B/qMdNMogiQ3BP+JU5VI6wQG+rROoZ6bBJO
9PxvFz84coWJOMboCxihl39XL9ax3t+zFMGpuSob2I1peuh0TWUnm3WuyKZ/HvB17R7yfdWoEVRR
mmB6eUa2ncnzlrBP8bfQY01KOgFTJjU1gULanYmCcsLSivOIJu6b8sCy1xIpIoAzj+kHe1INV569
YNfjaAOfKTaShYAM24nLQfcFnUAI9AOotRWWhHIwE+DV00AuuiCMecrEZJ2ZLE0UtlxGKuqWoW4t
5oQStDNHXnVa8URxq4C+hR+tG+LOgFvOHiok4jXsspv+93CufhQ+hoRWkho6s40zOSvKoLMIWXN3
oSaghln/UhZt4xYvtGZoZi3bqkMYOYsGHixDwD7XePx6V9llS5hEWuyvhF4HkC+fdoTs6DBY1PkM
nKLLOOZBFfiLLndz3jc5UUinrxoNqfDFbsgqJ1LW8Qgy1VADwuhGN5Vy/FOdwq/FS5xnyhZe3FHp
GLhWKTUkDoTu55kSidypf3WK57cRl7ssJuzecoYPq3A0+ZqwHl5eTrycJMZoqYAaUgolj+D4YHN3
azNNHON3GuG2/0ksRi80+3SjX4LE/9gtCZsGgjaq5Xb8OIS+RUCx3AdlxWZtVwvTMlXwkIcBdtgn
52TxO360Vtem99mFKo4xKFjTcdJXq+CJ2AWn7EUyc8PC6CVWrm5JJPpLs2l1HiFDYmIRKgTJLqOr
K6y/J8Uc1rwMLYrRpwulV5vL5IHhtIqev7aCq80A0mGmnM335utZw76e7fEY81AQicMe/L3D3XKE
QJwp0FrBEI5pkMEoXg2j+ygrFkc/2aPc3b6waDG9eN+GErnjnVfMFF/Bts/A2/0J77KJoWCnPA/m
6/cSmkcJ0ZJvXUZcNb2Q67Sh1rPG3S7iOsi9LOO4hzkM+68V4H3Dp3f2IQQzTni2yhMWgFbIBjLa
zmV2en+2NYABKpUjT/d9oTgX9EbN+AQNjh6JlhzRljgOztgs1EpRjWU4xsnTG2PkYk/lV5kKcXMR
uBtWyAluttbawTD1sxtDPt+6fcuT84IhPvbI/L8qdzVyZMuyco6Ffq2WvJ+5IlHc2roT6G/ZFi8+
Hn5qgMr2caZrDwO2xJNVrhntpLPI1TeTkbeyygAfNMPVa22QRp1xbbhJIryPCRtWtfaxqqQP3ziM
BUX+K8GhWeCRfqo7zrAlJxMAVe3CJFOytihBW/Dp2U7ymTe1cq+k0VqUnCUhCRSQhY56GMQ0g3gm
johOH/pGD4EPj/t+wQp9/NINpvrFjCUUeBhLq3EQKsp11/2hnLKitWUWy93XHrBVbfKXteFc8Vbe
qN6N9QpxMxVbdE2oYXUQysFQzFfIfRCRT0TUStl3vIjSzvKTL3RxlGlWb0Yz/YmrgvolmivzWKCP
A/KcS8xc+ODkTo+x7TwkluYEkxEgCEOvK/bFA2849An9lyvFZy35iYeV2FfffqJDXGr5C7Jn71jf
i2XBZs8etAWyY6PsL5RDiIZ+Dh4IYrBRCRPRI/z7h6BVkAP/W5H6+WcIANCpOcJLFc41qDoNhZEI
mY4qoX7U/W+C4GFdxYkWS+OKf5sxGWJ9B7OO+sJp7rKd/EPg9LMd4zepdV5XD+ponImZZk+NR9HE
skpkxEASJNhPJMgLYwKsOSs3Aj19KTfOxJ6v12Zm/Hiek9msferqysA8YkeRoqj+pQg99R8BjNh4
oWCNkhmrzxNTJin5HyNaE2IB9Q+YLVXhdRV8u1ZI85a+lpUZKWO5Z/kjwglyYV/175a0XqUyX9zk
p8AmgDk2tgLCZ3DtjfbxJp8Fk7AFQK4Y+idmKwu6+f3lQhaptIFpQY4pzkAFy5vmXoPLpoM3Npls
hNHloSnDpr9hR9p8lXWD/op4pXpaCzOW/kZF7e/VzqGSG2ksvSSSUOMZ+j2wqeYLjdOXiKVanzJ3
aQjRmF+YCRb5CperGXh+WUoU/UFFeJJPBn4amp+rNQFnsqRFElJa2ws9dG2bQ1Ru0NgfK4iDU1LX
Q//9tdrYOZ/r/QPx3jYtHZoQ+b3R/NIlX3QgO3DPMQtqeP7lZqUCtm3KG+YTaD3zO9PkSBMtB4mj
R1jyqDs70H7puo2pS4LDC2KP9wEst5cmeDCkPs45n8OrR/ARzH//wYbdZrPp01ynJP0mQY7aIwg6
kjV5HKbhHQfWN7z32AgnvMaEe+pMebZyx9nBfHwoxr+DgMJjumdcRBM3kgdImicbZqq0Rg+/6zFE
nQMGBBrguYpGMuAuKRpC82z5G2qtRwLs1WtNuDD4/ZIWSbebOmJqFqe1okzHSVGUY5Urklz8bnC+
xKaBA7LEiS6f2jnmQ/TsZIOGfGVKb7Q0D5QrScS3U4wktRBalC2UYWv4Tr1nj0MCkO+fJB69up4R
jrBDEWDLuJ78L8N2zrswOapPqFIGtgrXg3VFlnpYkLTkVeGHlqdcrskKQozJ1FU1GxC9s2JtHUXK
gNBC6z4U/AdU5fVQFUbqiQUDs8a0vUZT6itZdDg6YstTxM+x5c7fxFNzaD9H/GAfGxaT7AFChZBE
iNtt/gD/085LbzWA5+9qIqaStRVZLaNXQjSV/j6Gd/9y52ApgGFgADeHc5c/B9tDy4DJNDFxZm7f
tBVzhs0OYBRG0YY/aTcyyR07cy6+65Bq6NW16XeuSDjgC3rQySx3asyPQPrubqz914rIjv6bypgR
mV5QmdTM4lEgdLCKdG0We37ioS+hu56kWeMbhNmAXgrK2VjHactXK0FcD6nA64zBz5sCkSOXyeJP
klVdPbZAZMbrOa8kl+LMOxjSO92P8clZRX6RdXUSkIKPan8eCGJ+q21g4eSvUHFzZJkDBHy8lK0a
RA2ABlcnCZ+ZLNbUCukLRTOi9rPI+LWtRsBHvFib+cwfYOc8TSO6EQ7MCTRPTqm7dDV46yPGpSVT
I6au5n8BH68707XYLNpZGucFMWMhRhOXoRQwvSJvoXWKnZuoppzBQYQgH6oIIN8ysJuX6FsnoNLf
iNiFnUzMIxDyALbRqMLlmxoPsWHfwdcNn1xHY4U6G7oFmE/W+W0/zBDU9TkitMj4gD59Jm4XXflP
Klkl/TYoy3gn2mtGMf4l7vbWi8Jdf3mTI8rWTB/8SDX82cUh5UBYNNnV2MgDq2P1Rn78m9tBjX0b
Zty0/TvAvR3EDuqvXAYvvQJa+ZASucmW6uzWoILWg1uQ0chbtWFZTK10oj2mf0p9WpMYfDXXelVm
xS5dA8L3rvvN2up8icRE7t87lRJdx5fKYzfqNWXVjmF5Atb6XpGiF8vlIghgLrSAdOd+eo0Co9oC
cZ6BkfsQ8G7Xm+qIxV5CxKZ7Y/Xic5xxj8aGZo4bsL1x2w46E2QMvPNf6me8q2u5BrDBtHS+HcKq
WDVnGGsp5vw6uYyrX/nn7F/hGXQtcUViou8rfrvuJps1KEjQ+Lzl4zH5RW2cBhOMy0yw3yhEqRkw
uFdBDBl2S7XA+iZWLoA9r4CEssucxZz7oQ+hqJ3fDzbz2d8Yb466Ei0nuTohHtBgfFkwFOpeazDT
dU99NUQEfkrCvPVYjoPMujpzy6/NmGAv3skpfx2Lpv0idc3ns3Su4zI3yuxbmiVLmp5Zw5B9+VV5
Q/r2QBPpS16K+mlqaS4gajqL/9YtW/Rd4siMiL1L9M6nbeyf+glzhpMNf3l1mX3u80U5P6Oj8Qhw
C6bBcwzI7Br07NhaSedYY0ex+C+Gzv3bDeOL4qScmnsstO5JeD+aV7Au0U7utd4CzO/Fe/5LVwNg
rU08MIh9qGrc3LPDPuyRyosG2/HndJIdYF14K42YU6BvLBDDAcEMGSG4rh/+bCoRJzltiydZLXKw
DeQROYJkmgeS/eb48kvYdZzzhDVzGtz+w7eHQGag6zZxv/AlZDC92kB5v2Z/yGxM4MXRtF6U6bqX
txPRMcy6WEtWo7QlaRit7ZZ4VIjEUc6+SNIoja1DnYlvir95jJTWEq/W+2YnDTPl4V7tgYd9KMwE
WHCVzoIEFnUqefoyKMJ8e30t8KDCkSLwGPakyxNnvaE07qFgKjNJ4WCDkyoxVpbKoMrb3qF624hg
66KdZYQ+nLnZmR6Bmq6vWlgNYW4jCL/v5Hnci7WFpx3pG0SnQjIL0xJt5P1f9VrHLbBEN7e/n2hw
Fu3dZGQx1Q2YzIpD7Zu+vvFHEPXjW8xcbLxlum6X5vcLwdwtvCe+6Hd1r1639AwHAbRoomLw1QhF
MOiSu/9LlBgQEaw79ncXVQum+S15YSzwwkWgEolaTSQ//yLkQOFDFFlMOVQtU3FJ1X2siy9wPyUw
Vo2ddqKz58iMKrZ+5DjakB5gofqbvB5Q+onhF02rskzMA5bowKI89LNN7tq+ScLBolQNnznJZiFm
sKqX30TcGd2oLO3yXueiQVaecj/q4TkaaiddAtmTA4zt5EOF9QsE1BUiSU0DAw1Y1NTTD1As20Ow
8TCL0dZPfzSn1E6QPRD625OxD23GtI+pd0zl1E6a0A/6PnCHlaUWNqPNxQD/nFIrCtITa5+50yKP
Z40V7GHCmETxAPEdfOFMVhxaKYDtReAN2ESRfoU6q7T7fAd5pTThVGpOXWxKsOWkA5QlHOvFnWsK
ioMmsKT6p6+zJfZxMIwcJ1/nSmdc5VWqzcZDJAaR19+wC9bjwSlubD3KH8szVG7RGdMtM3CgMw4c
Clzx00cFH7Ak3kTn8hDLXZ7Tc4LVnIpqEJg8jZ0Jx+wqQVlE53ARUP3+INYNx2nY/Tn9G+U3Kqle
jhaqycPINuyT7+qGDd73PKW5FUXcMPmhr75btWMDbEeNua4dxBgXJ/Lp2AJYVGejKw2sxMX5JK6J
7Na0Wul19WOedj5ZVOtnFIC8J03db/xFMnf8ayozEQu566lIPLHxyow7W2eLWaSQ+7Yj/i/SQ5gW
aNIC+YsGfkeZK8KVu+gSu7sp2CeMElaiRVF1QOdPJt0vHHcMd9EfcPKn/cFFqA+8/44p0N4ZK+VU
Yykvbb24KizVWpNo/bkrbs1TJn14PlP0VWhgFr9AA/gR5dDEYGOntrnDsBdvKFsEf3bDfq0Y5+H8
c2/VfXVS0SVlx6f8Ymg3qnBlbSYpTD+E/3uljMuS1xftBHksjuTk3Bx3pPDTaAu6xBL9UI5ZuV2j
lhB1Kcfn4qA3dQ5/qfgczfRUr5vSrBH3vxRL9I8nWTYegGoU/qRmQIDIrViad7vpmYpoAGIgrSh2
c51yB+msRA3QrjI8dOu1vEnZDUvF4xWjp8GRJRWiS+rwtKUEdsjPr2s88do582hi/AIWQTWtiLJ+
TXeCUmf5Y4/H6feUYZuWyOaPixd/8f7Gaj6J29o3VgIihDgnc6d0o3xj2olsrbUDXQiSK636BaIW
siZx9aPEjIoUEk+FpHxTHTfszMUWW9op79eA1gC4MLDLku/y+XinNprBuyQ/KX5Hoa3fjrXP498u
AjEfT07uo4jxsVFBx2OyHSQ8OW1jEAhjhg41b6dDsXZLrHEuSq/GLlKYEk9Ht0mxK9KkkdWRQlBe
jvn5lLhzm7k4e7mTI1RNxT8J0+JBxBSVKRL4elbq2Uy0zSLrRSsHSmGlWdcg5aME5QzW+s78y8dr
60T4htN+y1b5SFfbktwWbvI3Ot1u1ozW3SnT8eFTwcc37Rzj07dt80SQK1b+htVD4v8mCLrnSwXC
Lffu5oIta2FM0P+CQhXdtXGAn28RzfljkEU6bX+8vOapRvyu05tgsgAQRuB9SFsIA8K0wu7s+MXg
ruW6RXNR9m0Xwf3lg+JiIXqBpvnC0zKFkAPFz1kvgoEAjUCX8ACHVFjfDKjYqlvwt5vxMDaFyFup
4f9/jyZpWXcVmJeIP1p4SdmfSd4vor6KUkDciXUQSqWtvQyjeGFMaJ8JPrdu88n5zC9HA2symMie
0x66CWouxkmDhWAWiJcBjaQoEbVyr4P5RYq6OBxdY+ysaHWf/cbB9RCJLk+W5dJfNBUc+QpPJKJE
H/GhJH/DOia+dPUJsB7NELYtszLiOZNP1Z4Gb6DLo83pHHiL1J1lQxNVSAJ55UlplknokMs3Qab1
7MQyljFEbzgFWt9vKN/4Q050PgHotusOK0yd0Zc0Fs0I+4awPthxhTWzaTmHzyvIrywwCaOUFxke
j8Jfx3VhPETnFzStNTN5x9WhFukVdnV1J/q7qDBsG+klfzeKofehwRH5lWlbYt2I3xXGmnk1ukHN
yPb6+I4ui/gjL+XdFw01lJTxjRlRkXdFHXYyZpi4vCMUttrahHAys12tUPvqsDzUMyird5EAfTS5
HdK3f7BxX34u6Sr42hTTPNk7jgA67tit2VyZ+JPV225oXidrNHGiXm0qQSnjRpKXbdRPozDYEdyX
bjc0jFyFdK9KHTKfl4QISJm/JjZNTeTGjvn4xV9Nzam2inP0XDCNdtYRhXzq5j97Cs9FVA3s4Xva
zgozgZon5JVrvdpMEHNidZJUkX8oIqLEFrZgDePg6nwBzYiWeDnnQqYNt98j2XiKlzuP9fWw5pVb
9JoBZ/grVyfc0y1VytTZO3rUZkmSFDDkJJYQ88SFn2djYDXpoJWCwCCR1dm6aHxmQQPw++ei/ZpH
pD+SfKQ0Ca3Buesu2kpJa6Tqxk5dcZQ+vijb937NbzH6+gjV1QkHltkb/DqP+MMZgOfXRYqjZNE0
l5JB3BFTyyZz0JW1TQPMJJ8ClnXcuG3PrQ9RQ7LQ2WRij9WeY1l72N5Cjp6rFuBHO8rYnvEzom+E
StLMWa+nH5jvO6P4PnPlLNXBBO1rdW+n+tjNo05EzNHe5ZbipaJYDYARxmE/NvGu9E6PnTGxIHZ8
QtZT1YPqp0+KkdUZJffZwTrx3Op+KB1MWRz+9lHCw7pkX6zjdtG3NOta9QfYok0PlK4ntgcFSfgT
7aOdAtACDgRFdk0CWVbuIw0FkJr3bvQbgEWziGSDmD0AsOGycWISpg1pv38PUwAKpE52b4Tns9OL
MgnLSwqPo82kqSJ1dr6IYesx078ePBWt2/T29Zs7i7czULYXSQwPt1uUcYfVBNYq9dmW9CT3MMQb
xiYdYAOPXdPYTvSLwYqRKeCN4uId7Tbtahe37qHPamGcHeAjS0vViEOBPX0bsynd2qfpUD3QHZRm
tlHOAlc6jo5WnFf3YjyKc/X+DKD/jOAN1YoFeZ2Cmj5JQF4QBpqjkeQ0mtkwHfFZdUfjfeeJHdzr
pFGGHKa9rMk3e9bZagKTgU9Z4u9Hlx/qrXTVnmDZIC3RmXcktcxQG5xli+uvKCL4JhXA7RqRjHIr
FyLK3E/aKGVyG1Ezk9JQ34feIVmVg2CDdrLcWmXH6f0P1Hu/a1DzcRvFeZfWVslJCtk4v06Ugysr
ygAp96qekvexxB1SncYjhDmv122ubmm2qGBZStJ0XTBR9AEe1un+BsqcbpfllW7eX7Fi5Czyf2QB
OgNRPOi+Sqdbca155/c5ENVcC6YkoKTY25irFUpXaVHs+v2qDwdBUadWzT4EX2MLu4ypJv0p/2ao
ReSBTy7BQ/8FEzB0KSQ1iW0N/NTOWsiZz+qwvJOeH72+cOMOgN4/AbCpvDv6WSFDL2WOm6KDIxHH
4yK6h7yXvDibJrivJy9Hhj4cmCQodNHwx5xAmbzCBkkfsdxXdCq7B1dwHtMovcxaOSfr+PlPVyg4
/FsRdtt3qRCNKHwOe/WDAwAhxqNYsocDk1qxxyC8pBDGtgCKdGim1Km1V6OOxVjQr7Nh49yfCYoP
PIPY8kbBGOToPDvqc7fHiBa407K46gPXtp3Z/F5iCaDNqAp9mujClmD3bCpO9ejM/aPmq4DnQo3L
K6N+Cho2CVzZWf07s3r6tnTcILCckUVcFRrV5jlIRV4ekUtJOZG7zHcaGE3q53VVw9/VheuPE6Wk
MAb6nZme/tqWw7FzStl6WfjuTY4M2ingZi27l2I6zor+OvuwYHy2sp1bhEoFA1rMpdfMHXOmB0do
LkyoRldWDR5zbndA8UMCarcxNU1ekd30xFEflkEEcIfKTaL9p80sm95xtdRUMOlgkivD5N+E5Qiq
GlK1wFNJhHCPOrxo18wYUS+aQgcH4EK08rcxHVrODxMRS6FOfDbBO9QOzf46oCIrRCBVqDOT4Pla
hQcob8+jc01o7pdlCCzvk64naS+uSguewXhtIgUqsUj3u8WRKIUtzcuj7Jncnuc64RG/Bk8j0T8X
T/zxhVyiMeHLpW0WFhy7AX7Or79kG2ZvNp2NAdQ49023tHU1upkfkXiRyyW7R2Lr7Q1Zp5vJCfEl
bvXXJ9QOHvoqsEXLUzZS7ZZM2FzPJkdavVbLiCmdXIr6kulrXzR/gxyV+YFefal/oIG4qSwHK/W7
qC0PU+5gc1qm3BDWW2m8QSCjImNa4hv95Vg40imwfvr39fFIGeXiETjMS+DTqyQYk3TC1T2LuroA
oB+YcvE2i2GPSbeohJ5pao/I8MI+D01PZphXDYaFCj+aUdmuZk02ptP6fYLmgbCDL5lrd4/43Bxb
AEdusmJgHtKmzSgJg/vYF9witknzV+DormTrjpCZ/5VPfENHc31BokWXtiHhCmuJdhg3Tg724uzg
hSHL4DGlOyDh9LF6+WcJgoeF6I90e4YpsQHy9J3/GqD+nfauKGRpvGBM53jkt0Z43hfrecWUbyYj
C0RopwqN5lUY6dljpsQvsZq8mUEvSnHz1KXhrVRbu43ZSOR1Rg9m/Mh7mC6qZo2sOPI7MMiRNz5x
rQ8o3uZyc7ghPorqnSwzRWXB7aHws6NYb2F3gWai4OM2So64TP2KxROZeShU7iE06985H8fJGEmG
mThmPX1NL/kT6+ZLXEWdNRAEkiKPW+MVpbYiLbVbk5mG1XXpIHK9nhrs/I19B2u/gs86qVYX9W+b
kt7f8e9w2L0/7Lw2f2NZNt7UM+BzzQGy0uXLLWwCm8a3NOnjGBevnwjT1M2bgaDc0uJjZNAEtNHn
aeqjNV18XahLQ2uYaKbAD5Mz/gC1Z/L4pdU7XsZEnclS2FFBGwxzkukt8Gdejcp1+cQNQxuNcSOd
t5SFse2gM/HzBkUO2A6PKJl+U10VTnaY5xfy6gKQvtBSIa+8ar3+Xgj38VmNX8JliWiPuSF0rHEa
vc8xCtHjfKiKuHKjla2AphtzWGyihjklET5SVpetpdh1Sit9VYzb7PDcY/DNrOnCi43E2HxxDtn/
knCQmdq4RZ/J6eKF7OG485KiChzUIpicmov76/wr1ccE6/FI6+hek5FSThzdalWR4M9H3NNWisV0
s8FazenIbcNEFLD5i+ihoQS8KMzXG4kvk+cuxFR6olmKJIMEWCRqMj79dUoXbbWrQffff17dmRtK
71aFc9OWxD9uRNlK0ohakJozWLgkiJSHsY2IQYBk1tAK96AETG0uAOXra7u9kc8R4Fkos8jyFG+D
7P16g3iF7aUifPM8jxTxZOLTOcOKgaOFqfN8ykJvmSRmfBBQJeGGajTrOdQvLPPdwLSsagB1A6eM
B8ZaNZ8bGUdY3+r2ParLOyE+P/xxm/fi/jbTwYL7nm0wO5RizqnEo2L03CraSHa4xdxuxM6Ijf9h
PH0TI5sSXd4RPoxWlVP4XHNsvcXkQXLCP10Yz/2VnwFHmPuf7m0Cw7xM3SDievmgU/z030cEhdq2
tsNsDOjkxUJJ20Wc6M0J3V5HG41+zYimjFXO3Q8TVn4TASP4KLUCGhs818N/YM1ITv3Km1S3G543
KsVKXpj4J4sq6fL+GTxgtlDWoUh0oKfVYP6QAVf84ny7xSVvE9sPTG956PyWJUpYWKbWf+0Mj58q
kOTuN+ptd6F18S+ViVDAeYxQvmfuWPGho9EmeYtcGVjJBRFLQB3HfWWeAiGw1d1nfvsW/pTdLQpj
arfVux98REliqA0AwOkc8bsuioGFGTlnNYY2JRtLz9Sa1l03ZGgVBuGM09ghXlBDjCJv3cZTq7W6
/uYkd9i0I3/PTpdap94TCRgypuvtWcD5ynv+XcS7G2oE4HDobfZ5SDeq0VLvztSSDY7+fv4Pg4fY
+SOiyrPVMBPwT3c3XkSaqFUyrWqqZlTzGT1a8DOCy7KPSvf+pt9S8T0I2U/8ABvRd4XorPqJinND
CkDAfvyQ6QkIVS1gBYhl+FgdU7F5aAAIsZRqxj2dQs2uQQ9aGc8mqQlRyUv9BdOqAl/70UkTmuj+
pLP5D4uGjNG6yy4NZnIE0hkJ6StBFnEm06HU6q4wArGgkBsQxpHXkZ7P6E7GJ7yCWexxqeKyMDbH
pFDdvCeYD9isVxpXJV7bFHiWzMItXdanwHhasQlqtwRiqxCWleH0rKhTBwK8Xj/7qErpLjqqxxNg
zBH8EeWry1cXCTZoyCM6F+cNCVk1TF656IvojeNXX7iREmegeQj4hiCv8IxwrpGw7KpX+RqPnuCM
Cspz2ueK3aY44EFbJ+05p2mmRB4+WE/eVHFEb5CvVfIS1Xl4fmUzobf/GO64PsG6MXzgCiBJB9mm
PJgWBp47yZuk9WgSLFpT9IfXWU1miO0+Imc7NgohXsiPYpRu7SneqzNTtC+f/5tIHTD1Mh1WvYPv
I07qTOJ7kd5Uk/xUrZUTLDOOgDH/xRHjoG5YDiFS0aDNTGPuVV668B07lGyNf3JIWHx4F/1UC5jc
Vp/vuAQWldCqc+y1qOERbP9g4Qpz/5BQ4uEkHZBlN9qJjyxGSf9G34Nst1keq6fumHPfkvGAJFzY
X7ptOO5llStdIk/U6evDAr2yxVYQ1nVsIizRm6DwfMfRXMn1GetTR9RkrEs8+ZMYHSyXkdoSpTmX
uP03cz9sxV1ejjJ6iiGtqvOrnmFW1KLf/v6hp+UnKuVunkWauGEg/hlbiPdjkXr9L7YXT0JgLQf5
m+YIppvphenHERwezW6idcaMpK0qyeetTMzCxmb7EnFPvvFlOhLhyWorIHRxNg75Elsu4oUNriGQ
Wdf/g6LBoh2T0n7U8GU9bEUyDIrylrIhUrYHYDfJzgzU3u00H8l6I5Vb/oDZxsjacYCk8rXQFn8q
d8ZXuTbFa1cLb20uIadiqKs/OW8H1XJifge/QeYwSOSFbA3DeLb8Z8G8ImaFswAC691vm4cDXuB6
9tLf7iITJYJ0xMyun/QKrAFT95YSEQZCy1+Oxb2vqZEVdg9nqTY0k2aE1WInU9auRtkY2QcAm89y
7vhOYG8/zekaBNstD4iqUZ5A6mXOCOEprnOBIt8QQxQc5v1E6taiWB2wkf6cbgqD1Z83cEzC2frM
zbGZT25PWutxsWeTWS13d0aTArQdiqDN/p67omqJxn+swpS+uwWL6g5LkXBYcUkmtX2GTMUd9jKe
n6A8KFMyh4AQebf176uZE9r6+bDVVyCjrxP7QbAwRL+dDH7LZKf683TnuTo+i8yJ/f7gbZp0gHDL
Szl8QgrH6OmJTChapMvL6z0rbgUJh2CyaYtocJU3m0xTVwL5m+vUXBIWxg89ZGaT3m/N+MhtGOSG
q1txQlNjP5TPIh3WXbPBWIrdXVkp1xFvp2BzoKYONFkibJcCvTbCS2Xsl3zx96I2pDVCItvTAs0s
4FQmtqNE8bpkj/Vt8RaF0wPqgL1J4ZrARd0SnuJPETlN/QFdR4wIVEmLElc9EMviNe64txUpZZ44
xWdTJcq5bX3Pr8VPZrXICj/SYD+b/cgrorcYhCnqfJyaKEfUIyjHS1/jeqoLPJOOftfTS/J3Tr85
omwfSj8PTyETOCI6aOLrmfEcSd2xB9mSPar1DLMgN2MK3TN4H1afFp0QLulto53XqWRFVyO0ZqEE
OMYcaTAhdkhM8K7GWbMI6Y78CvRH0Y9C7nsKEkopo2fRrFwqGwFQ10rC1usqGZN+ifsO3sFuho8T
BHQkZ+eShSUMNDRGosGY17O2/eI9PzV9VC3ZVgrveEQYkmiJy9J5nerzDVxeLSdt0AaKWVzccRUy
C350WaTJL3bchMSumEtq/0fI67bJlePxHJdamgNWmXYssquz3Q3Sd3EgNea7Bg5eqtEZ24KhTtU+
UcT85zD0UE0TT8/HKfAVCZoAlc3BlO9YbnVXIQYsZ5P+TkZ6SJLOZBUXwez0IAWbEd6jIQ3O4OaI
PnUzCjxlivG9BwYdIDpzCR+NXvH/seEb07qFNg6s6hdDQqFhs2LD9ZcVq/GJTY3nWjAFFKPgxaZj
4uli5DL1fPUJkxchotPIH3NgaGsqlsncHdgT+QAHftIt7zMTr5yDpCif8FpjTi//Ywteikjef5Rq
rUGeXwHBzabwneIGIw4qunDfvBmKhFmTwlsrBObkAIk0asRj9DJSlKB+SmRPDWz5He09fAF+qtY1
KU1i0c6z62S3+UnGfZzrJzETuVGZc5MzE8nq/QbkGGec4iNLuddVjxx5wg3+JetTnoAv/vEcNc5v
96r4qzNImmisTb5Y7ix9S+WEVQKpJy4K5JRyInseTCtfqynEyPiQ7o7xgwxLhGMwQ7OxW2fMC6aB
LJBAXRgKh3U12xASbv0yNHJXM9zqdenSvTZh+yu9j1Qdwvj4OrGeJUGUt7XWOzlalm3LrI8ZXJW1
1NxFBZvmuC1cLMnUMJBnImC8Ewtey3iDKPsnJNSEVWKRRdF4SvmuhdVJIgE1PdtmUzIlH9cW4tYD
+4IBC24qXayDDVEcCyfrlr66Bl4q/DfX24VjOSi6+QwzBiYVaQ14bFTCplFuChkloDZwcSpwAFn3
d7xyZflenYRCUrwMvEe5CS90wf9Nsbcz564n4dm8uszUe3r5qw9ijTVUAMTxFvNArk0DVTcgnx/k
Z8fhQ9H2TO33vVKOVyuupvXA1/IQCr8OdFNch7eK4aDzLZYRRbAbWDDIR8EkEv2HjCTgIfWpFhEQ
4SpwmDF0vNOZsWvCSj4WZhrRzIWtHrxKNNKj3Ut3gwjMSD7IDSg5d4XJFxNf7Gt8uqfL9q3e10yw
l34bua4kFx4k67tcerMLArS7LdnEM4on7tCdQj9ckhFPXnt7tNb8hJCWnL7i1EYwuF+v3lGVO3/n
dEX+6pL25WHoQhRVpagnKElC+jkJ4Mz5aa3sM4hjcNDubtFiZBy2sjatfxZL5SK0FXlKQP4AbLM9
MwK/TtklgCpXWRDLKchTrm6JXY6C9NW1+DRB8VHzY10u0/aM6QUccTtVaCajuiCdR4xLjSMNstNS
a5BR2nfgJmf2GQgtFbqDb+3EVDCimTK+aYHbCS3U4D7wyItM5QsGuH1pslJSUZDbkqdx1WkrB+l7
C1bscKcv2BgYEoXsgb+JECSM28TKAxPo7lbpMYZnuxJwPbNaEUiNsuhuKlDa6SxMLZXnD1oT3xNR
Znz3Cws2YzI1MC46CAMEMiiQYqtp/oJbxjoFID/e4f7paXFk/plSDH5wgzZjq87Qy09POALu4y0q
tNxBXqCLM7ydM4944fNX01a/fEhI6XY1um0VG0cQF20tWnHFF4Fkc1sLPRoZjWI8Z0LQwEkFW4g7
JIqwFPhozySufD3bveq+eep3XcC6CWPqD2PcL/CKuOi/URfu+bFKWN8DFXJFraeRnJpw4B1S8Rxf
h+LBfKR51ZQDQy0xuqfn+ZPuv7ViboiSPxoIpd3683gVRJ6CUqQEdRy2laHntLLoGWTZPBC9JJrN
tpsyJsABWAXKPGfqmVombITVELcskHROAnmo3b/1xEeolhADUDUbOGgIqO+464yQhR3a99ciDNOu
MOOxnH+pQpV1OGz9WVNMt8RIgMX0fwaG2CJWkCq55yLFyT07kFX60newqNhWVefOjDh76gVHVTJH
owzcCFe0cgq426snCTj4NBlAu7aVhu0yRnXADcfxwl0iAaSRW5fkcXcr2mowruPd4opQnMDqqUmc
1E7bbKQtf2IGhgVMROwjHpkXE7yqJ7+Joqvit5idDbYJd1UTDnh1uRa6gevZo2CG3pg7ofEXUF4A
cExDFwKTyuhtNE7uPqf3lQXU5rK8/ohhkG6Mw21Xxy/sycCaoiLf5g0UxB30broR8JX4xdKPnOhr
9Yy9a9upBxNmUGALXZSOqfo1j8AMe4IABk7DoStu6Di9CsCf62dn9XI7KEhfmBi4jslmzC7v64sM
5Bc20/Xivdt4QbpswgIZz5MCCKJSq+3Hz+wvQkwUmoJmYBOEaFBe5BHzRmZJ1gmRxzknriEZ0snR
+3IEsSjYUDT59+A+EyivumW7t2sFgCaK3Cnf80SEfeT8r/tr3PVsIH1qRGTgSfjqMTLJva5bOire
SagdjqiZaskI1zfgIs8OBbnUDFWAlGzDwoF0PDLa8x+JJ0BczlivU6YpuWoJi981xdrkkkzuhgwm
1gth534xUmaktT0yE89wOT6h+i8LE5cuSAbPvSl+j1tQQhYIFZ9sE0rFnuDQT3H8rKrUOSrg2Xc3
Z3CaKFhjdtLZeUU8Too+fwdN5VGf6L40XAILXDi2j3pcKkr+CNL+rn28pf7gBkqJZ8J7Wz/9wWve
T/oWAYvWj1l7U4vLOWGFXDPz7un5T8n/E2tFDIH3uLR7JOrhxIfUE4grZrobRiqlCzLKGxY6Iu+4
rbJ+K1/cVQECQyj9B7LdlQYyok0Ef6uDiT6tG3eIQs4K9c8Pm0LMNOW/HPzByWOcIsQtgAn3bahc
1zfoXlFZ5LCjEs8l7DZ10sbzN0dHICR5P8V3H/q5EOb1WYSlUDeUadqvoo+9qEHqS2qAlXTu1Mil
zFjzQir1CYffiY40pQ26ZZdlMLFiiUsodeD6S5lAIAiTSd7yWOmaxn9WFXn2EI8103IWw1ukL7Mj
9ClQNwTgl2VKjb21Bu27H3wL91zd7AofRWwXYD0WYI+yWUyttb7+TqeUMjk5kW+1b//ln+RWj8eu
kUovymL/BCx7aUVyowyPLxpfMB0FdQvN225Xb7OgkRZ4+4BfYOouVffNzidCJbGnSojAoSDaDXam
yGoHmX2ZY3BXjt8p5lh/+yEwRRVHGGumsXIpzkOhmhXSgPsBiqqOR+N1Yhz4CU6zN9S1SV6ACi8W
OLJwy18VTRscfm4Ig7WZcp06QdzYuYrXtXfT2DgRLzBmUVG4rR/Gsgw9iLsHhzOo8kB2bjDEjEQY
vjDV5J5fZKjCZxpX/BkHRpbxKhYsDJQdj9Idci9dvK562Q6YhBmP0AXxMlVLJrjs4PLwws+IU39n
1FySMBjeMS3lKsAwPD6Q8U3gW1xyJsOCW9kDuAVsljSmAPjgaANfGZ9j+A0v+8nnF8j01tsNsJjx
jV2sr4MYNPooUEhDDW3NsN+em/qDJWlCqeXX1PmEvr6MrNNkfabe9EC01qYpYm7fIbTdvIDtcTei
NqZV/a4OfRRSbDyAZ9TQM4CuzceyhhBpFLfgbg13cEP80tP8K0nTg5JOpQZul9BuFGY4qfUAIhm+
wAhqDvdpmf+Zg6lZRPoSgAmHHl3pUUkjl0GV4mjMMngyuBEpamJaeWl7vDrrZ3srJuzVB2A6y21s
8KH5PTL3RkoiF4SuBzkPONXK1r1CT8iNqnlRSi2C7Ntp1PRANTiGFAT8eDLZPDniMxv9odyJ/yuT
1p0fGQbq7Hr2adlbNn1Ry6BJXEmPHgSHHi3mWZubXXelInsVMaZc5R8LmskVTRSwuk2gQxX55FlP
Ortzmc2q9TyVbkcQF+7u5CdvonT9/xCkh/k3VsafK/CoTP2DaPeVBs2Inpl+ji2hSFsuqXdisO2M
a+AqTCzd0Pi/v0gsYTuIBFY2sbOXZiUAhItLL188ZSYO/8O1XAjTN1gJ0QP7FfJiLy+/RoqQo3r8
fCcZ+pVLAIAY+65i8GjTYI4zloVeh+/gjPWgfkaeVyYNGXLcCdDkV/fEMd1H8Jfyfa8gWVHMoW44
se+ni6xQ/4/BGDxuLWc9TBp37JJOeoncEZ34No5qWNNlHt7KFngfVuOC05ZpJidedelf3iH7tib3
wQq2oeJqJ24Vux+r8csDxtn22MPAYtMNm9x9hwvYS5Ds/zMklb2ioKRf36vXy1EwCtfhsysLYdC8
gpxIouBj8L83CfNp83Rf6O3On0RsBcFnKI9NnIBK7dMePetslzngtMQzVFMO6xKmxNyeh+Y5TDeY
xMuCh4BjQZRbB3PEM5Bl6DCqgNGcD97YX4PXqKzFMdX6ejeIgFN1glZNmMEBGqj1+MyInH2vzKNw
A5J8GS/QPQbhyjE9TIK04Ak4e+p+sh8kL9Pw8tpvIX6KluX/h0eNhWnQ9yVTFr7B0LhANPfvVJsR
9qpzwePkVcdVWM7PVQLD5S12c3Ri8+ZLd5XnlLU0dxvtaTisx21to4kdGUV3xuWh98nnJjAAWjyb
RS54YYuZU7KvvBWcbg6woobGT8Fr/phz1o0RPzOAjMvL0sjRzqgDuZLYWkrmKdw6O0nL29EZQzdS
GhU/qGtiv10vgPcfQeTVLC8is5hE15N8WwHlyxBmTdajSnGzusWfIoM+GdaREJCdh9Y9Y8tQii1T
4mCefFtxPdkl7iLRm54KBhNmIgHm3QdNObhDynoU6aaQ+C95E/OFQG7NTDc46+I7hRU9suhcfHUD
hCCFZXza8aZCguTCgA5zMWhREbMn9KGYGjeTnfg3rgRvDhrTtvnHGZUSmMCwfQ6hlhwl2mxUkst9
eULzzUcdv12YZRStzyrN5lUgBzklc2Vtzvk48GIQTZXGFoAv5rRsK57x7T03GkVjcsfdI6gVpOAn
8MHgs2djF3bGQ1/1Zen2GmwinRMzR+QqXLLCRwYTqZHlP+uwFpvLvnM2ewO9oDK7DXMWxoALQd8e
hcigcaBCk223ZebaiU58kS7lBdTnKKOSSnUuWHtCOBxmrTDBspQ0fUs0+vm9/eZL7YmzpqyrZ9g3
c7CYD+vqREgKo3NO880I1LPgkuEpgrAuoSwEo4H28giz/PEd07GGYaIFJLNqbYVF3OpMFGPdbtXQ
PH/pB0qFt3y/1TyApYs8cAruNnuuMIoLao2P+DDcOip4ma1dxY5Bd226dqyil74ttecHbsMhH7ck
nu26O7X4cXAuFnDX+cG24BVFuLevbtAXcyEdBzL3UQSO9D4y2cmR6UfQ4aqJCAGSXAjvLpDVNjwh
Qf7bGOkNtENLNIWg+hQIwSrrPNVzUPM2smMq34mhS94VDUu6D4Ik0VBN3OChHyreVRw3guZlOEOX
fnQqJlH6pWTAICyV2Yjh9YBuro2K8iC2oWAIBqnA+BFivJMrE1QQs0IgIUKWtQ5VEtgn+Rv+IUwX
Ja/MrCgwtzATOxDEL3eoP7sAsmlIrOLfmWwpioVR/4ySrSDE1b0rq8gjP9NbKdmEiHJYL9vV9586
rPec5k9OpyXLEOEqEdfzD96etWcTYU/2xmCdvhtb2GngGhaFaXy1Sl1R9qG65tGUcRgM2BIqtHmm
zXQcg/tjwBmvr3SG63PI4p6f+25AXkBP92YPimy4SD4M4FZ6d6VtkhUUPXm2aVFZ7XMfVya9fLxh
2HZ9IbrZsAm3VlQWLGLd0zjtOmN/rRPwQpGoxDN2iz8Xmu31bxqC5bKxI1zgm1++r6yCkcDi47BC
Y1SyMGiccU2vH2fygl9gV1GDdGN/QxscPTwm1lsFfRNVEKjjp7ZaKUFec1h2GSknfPC4lwdA+P+T
ZNt9YVCSpPAd6Rh+Qgg89heJIZ7UzVp1NZpgyVwoEms+ubryp6LH8cRazXAB1eW8XHKydHYNwQD4
ohej1S3nb2/Hb8dS/ZtD3NQlRlIOOge/i38WF4E3khDpicRR8afJmDUq2eRgCd1lUH56ZhuKtjox
AmVpmvfAa6ExopFHBTAeWnErkPoz+3UoCMhaDX0AB2cllvsTt6qPxQZNeWULwvvoYVKqN2+MgW7y
VWO9x8lI1l7m3XhWD3lBqx4QvpyyvBySYwcrIjVEKXSP5+K6thxH1wSiH/RI4AZwKN5UNpLMznXz
rp2U4ZFOHrYaje9u/PB0eRRRcJ83/18WABDVp+B08eIgwJSH3mnO0+3N3w0ZrTTLZ1ZyssOJTOvi
4rqM/Yvk61YH5BgRwzGwL4/1dyRHNLD/ARS0pHqb8fuCz5eKB4U8r9xReIqiMoZK3lRU8fOGSwSc
bon1j76ClAb/aQ5w/5GauGAK/c76FsNGRmZu5raQE30esHcUdjiY6fJa5DrOexZcE9FvS2+KoNOw
7SwQkl2ZQ5RIZ2uiLCbxoEvBvZhxUJTUaLrXiQOwRjFtZR0zzeggPwMz3DX1iIxBfW193QVoD7ZC
1y0dgfBTnv1MqH/AuQaliqF65eeoC4rdrx9LPp2kj5LtuGcoHUOy8qJixW0AlJ4RNBCMPTjDiH+C
4r/4/ln/MsoaooDxzg3BVjHSLf8enRlwSAEky2iF9We8/Me9uDvHBms1tm6grYn5TbsmEPpCVXuX
HUNYckeQCI9YRNCrEV+sB15Z2bFV1kFHrBVtkpzK6S9tCe5xgK264MbrZltWfDDQ+oMDkxXXoSG9
tpdxF8G454ogNJtip9rjFXth8cq3XqYCtS6dhm8px+UEQ0h4wRYYcd1e2LUttioyoY1dHT188LBy
3zrr67cd4dKpFzd+XX/UoOkmwOEVByVR4sicnGn+ZsMr520jxEiEm1dvyouNHMPH7oHnjuGW4WPq
MphFJ0AZejwXH69Nv2MEZtCJIuV/nff/zfMz+CoeqtkOBZyqXrMheIQ5a8VT+De2bR7pMUFgPQ+2
eySzxl0p3u2eWz1CzoxikzTLAiG3TyV745PjpkB51gJqgpOPF9sIaUpBMuItD+L+XsJ9/b37Uf8k
q621SdpvNjjjYAuOmpnwe2kJQtzl1aKMoRZse8jVS0OeOoR+vao6hZldi/U3MxfIsmoSKSPVpRxp
3Fsbh4GDoZ+USvwnEmTub7iCkteofwWWwcf/AA11pck2sr4bIRUKW9yCG48ZT+D+YUj2/PlYwzFs
5QmYCxwdmJvEglfLkZMwom0kZKFXw4oeJWDhk9SGMBK2dl3APQGiIAmNKjHF0tQH0RnEpNM7eFC5
8H24T5hprh+XzYb5QsaIomsD47vuVV6PTAVmMQ+ZJbsdFTwi5TPn0WW5Tb9UrmIPE+EeZS87bDAV
zWrimV4cFDPS3rljY8A+SM9Ou62Ea77cCoIY+6fjwhCaYs4gYKH3G5R0gF4TwqIBUWgDTAnxaHuP
2qWHzi0qufgOouB5xTi9IK4LmVBLlqF0UKeFLZ47fpes/pTnrGh9carQ55gw4kLu2gOrRtSv639C
MqN/J4gv85nfkcvoyUrlHXH7q3yYhrHJOaySwVMhMYfo+lFs8WXopNqHItXKSy5ZUDqL8Gu7yuIL
nXelxsT5EC8Bt/pCdfDV8T7BIfl1/pBcM3CcCznssDIx9LDMXK7FkV09DDz96YypLshsBXaVIhTe
8+EQXyqEHVSmv0HwQ/0awBBQo5mDNOVEw7iRWFZIZz6X2uM0Ck936GB2GEkQFxiSS+oGSJSYjvoa
8/BB1EYIe/FTSJh75KjXUhfMbCQqAffW73teLCO2YWROFDBpiMpUYcymDIIDY8u1D3vFmSIkkxqL
yt6BrcJYJO+eKLeefDB9gFalf14EcQQKzFtkozePpYSBe1ArDp2vNuZ4w355XGDlZX0guVWcjLEh
3e0tlBb4Jfph++jNyV0+hsWPw6RhU66hF7/ZO09Dgn7WKyh9V3lF3mw80H+JyKnNVJ0zicuoj4FY
rabtwDcmkcD8syGCQPhebRIwXUGQPdX0GRutTRXCkN8gcjZJ3ADzzvXfmAq3LJbxREiHaVAEQEhm
j9v0+Yi+TgPqVJFmbQSWujWWLKsVpBjLN7lcG2qYoU6mmEnxWb57AqwHi24AzBO5d3byUKavCwH2
bKt7jpMmOyW70rIRoy3LVCvMX4M6mSRp/iwItrrFJnjyjCbrtZg1QravH5R9XQBy94WsN0gYl4T8
01diq4mnaDiVlU2w1zUeiyh5OeipeeqhzoqzoTvwGUx/Gy9UjbBtz814C0sDczfGIGuRAkgWCaLi
NJuZKSo0f2z6Rb5328bbniQGeuqBih2lgx6o/XGPF2VltI/l0grPjzPOaGwu0AwXgbb+Qkvd8NK/
oNjSFZkPDxerJrXx2ihiGSAB9cBj/aYfhUUMikuy1iOUNY36CyQPuhK3/3ONmxNTIrcWGoRxNW20
682rCytuU08rSwZnKMbjbRgUQG+R/nZ9NAbjB3OfV/jf3xERxAJ/BOXUuamgzrPhoXrWl2cQtGI+
HEIDUPEQoAfShxufIUJji760iJVEvq3RDYUbC25iq6X8NUf56Dj4lNhohLKyR/iBfSLQLnRboDcU
QcCQj+Bncq7zaq1eosIFatqDUBK5J3z4Qx1+jH6q8nZsCQffHkOibDhwPDHwB16w6wJgLchAa4Rg
mAfi5fCbMXbwm+roS0Hz1pgc6TmQUyqFdpzeMfmKhQ+Fi3yljKUR6AgXCm3dfxRaE5JOfhbPsZLZ
TATDuxAmiFAQnvxpEL8eHDukeCuR8XXyWkYm2KtxTsS2ZIvQQ/oo0uh5BImS8HPqx/nZ6NRo/wyN
j3iOit00YABAyCVLisrpafRJTEKaJXXLxCNeSE0ae12W5uHkgMKgB3hazsij8a+sINcWlP8BaYm0
/6Lpfv8XnX5++OJD9NYx2YKYBt3qCQJJqb1asiBo88XoQHq1nwOF3VeZ3pr88/X10v+qozRm3dkM
MId9PwrxGEe77mPfHCIAEAdhYgw8HjKgSvjBH44JUg0rMgVKhBKx6hlIMi5y58WsXQ4BdKLIirwq
UHyQSL/DULsWBUvsRlk686iBQXZIpWM09qCMAO66QduOuvNRMg9fLE5hKTIRvze4BA+FTMTYY7fD
7/8Bk9ylfDUz2VQGk0OcBG+GWKmp1TmANPId5ZUeflNciHovEAyuzIC7H7rAqmDg8Vay8oKs2th5
Ho3Ym4Tg7XK9ct50dOxIf9FVQ4F5N06rZzwrnNTPBtCs+j7XxlUlKLc3qnnklfz5U6PierQ0+WOC
EoQTiu0ah1RsiQom/g85TvobyxhuMbmBeOTn9nt2ADknPGAYOkWYAm7FYHgpg5BDJ3a3dTNu4iL6
a0UKtrjMvQCXFxK2aT15rRYw6izHy5jXcKLUeZMH/lTLo8oCmLVbTkrZ/iRlCUZ5Z1L+A+S5xf7z
yb3eNYica9QYr9Y2JdQJEeU00U4ZUOdrcwmr6Wsy4a7+yGvn/qGx/CbfHDJu+cjnxGyEoylXiWhb
q7+wuc/m5SC1hLPmPvp5V6DXFc35vBjr0ByEUMg5F6g9qSUMVyDQA2APKIR0bKnXGifuMchxiOES
bHHfHK7Adeai2+MQv/HQSmGdi/ucyMS/lfrLtmqITViIjKAWkRyL1b0xCE6F/j3WNbDWeLk7cZK8
XV88kw7gEa/o1/gLTRcEDKN3RDG3ja2nooMgF9WO+R4Drtr1JhoIlbW+XCX3Af6mqDyyex3beqPW
tnMDqz+Vxdb/lKvt6hVAgfMNNBCYVWyXerrt+vGr6MX+Qpub2bMjgqvgmWDW5mScx9ok5nQrDD1/
/7SAuDygPYOxI/gnBluxi4h7kgcQq6xp7BlAJRWFTk+bt7BQI0Yd8TX0eJnAxAyjKZImxl97YSUU
eIn6ZYHoPp0wL9ItkpEFPwK2efd5qKXBjah22gJxrei0siE3rZ1qqvJ75CNZGgYFeZ+fAthncU5p
0/bsIIiJ3mdg2Xuh36LZeQSsx2/uI2PrxIOOwEp4498V3Erurd6BNDcc/bio69EwMmP/Isul244Z
tG1fntnDOZcDCBamrYsFkidUZwi496W+4C0bW/NHFrD9KJLmR3yRFxbU0avCPTjXSVZ1aH7ukWT3
1Jv/IVWvEUpm3Nrw41YNDNvF2q2zLAl/Jy0u4HraAYL23Hrp+38/fV0HGy545hntHZLgUHUhryq5
+Cbjy3EyzJnMWWbtEdowARfc/QolnXjAjYDhNZ7zj8ErsnV3GPswfVwkCiaPUXD3Kr9jKlMBu419
d3Ql7mpgSaHSZhDFSPexL+TqtPkTto4c6KuKaOcll7c6BVRU+cqW7o6Af9dwzEKzJ06ZOD+KYuRB
SN972fyfwVjuephmzi0o2JhwU//e+x7j8HYr65SIWvaO8A7gqSHuEt3YCIxmh4vD+qcWT8hEgrnw
bY+6hDkv6m4zsq2jJYCJtcyH5pMnNmoH3jVeca4DHLgLiOAoorGfdccQigJ0lSoLPAOqVBm9zvpi
gmMZfqLyEUAX5DVcwyPIYjY5UB+1Ls9BcWzgxABkxh8ZBcsdRU363TujOtfkThpIYfvl4AHMj5FW
MEBgXq9d8b1l40zfgvHKXT4C/ilUuKI8GEQGZqkxq01O/v9DUcIxj5yxoRfOEYHmEMoJz88vEly8
H6m88N754fphb+Kl+nCjkBfhrkP1LUyJehuJ6a8GHAhC3lI5RI9aTgtzZWEAhCmY9vegkY1Qw/Jv
f4kMf7FCWx1jKxwCAf+7v8V+jU/GlHHqE2iV5yntb8lE8y+jIGCD/vG9Om8qYahImRVZ4Bka7xPw
fmMKIf/8FOfFl1uZk99WcIsFWEZm/bVMis9lMgtZjl12DHEvua2JAx28MgI1QSzpnvxoehX38DJB
ylGPxOX1jgKffg3C8YtlPzfA2EygWn6CjCbtGUjNEotF0FcQ/q6gxo6jCPbaHlMC0kmQsk6PcLhf
1pK5TbyJ5U/rqcv/tFNez9Ek0p+i45oOo0ZQ9PBCZ1XV07Pp6z4+SV9JmW150HufIsjkft+LGvia
B9LdxQK5nxX6Nqo51ywcqc8gkU2WgPC6on2xIGH3msTG9yJ5b5cVQt2k4pz3rQGEYhpwnaZnP9nn
6fQL9jTjkPJYvGQ67ng8MpM7d61LKVlm/3gKy2+1vj970TPJVeFszyOSbPVxRx1Mvw2wN4i5cxn2
p3tpw+76B17WsaYEF7psyzqotN51Tk/z159mlN6oR8TvJORSstRwh6G6cgKpnEHYEDzSlnWsnDKU
wp6QbNeLfxJa2jRY1rUy6zBH9Wwkvxra/Yh0rHvhKAGea2iIFMEE5kYD3LJi7DX4CnqJYIsjvqLa
83mfU2DHPLAkiZmPEszGF3zdikVKaTJaJIygecGyEyPCf86ydbFjcXh6suyFC0SJILybcyPQVFNE
8HBKIkl5lEfaNt3rp828ye4T1Z7Wm+GStIKfduhmsxfiD4sYF7P12dpTI1zO91oFA/pyHFucn9zS
FufRtC/3UjyI6hJ33D5sDY3yGUR1DLEsCHbxfbQ2IUhig005uwpcTr2jsJoGZB4BE+HQ0R7fCdcE
dScGt7vcMP9vQS5QSVlvgaNh4xCr0FXimERQv+55pR+SzFzCM6z29b5lbjnn3WYoXinzdBBC14gW
mqNY+vXtSCCzpo+UMwA/gaEkgacdvB9UJ0ggrz1zSDYrhzWv6o5FDPgzYxK9wBGBbqj1W88YguhF
7Da+jCA6OXwsR+r4VrkwXnuCInj6ynJsUg+ydVBwGPsvYHoMUiqf62CgQIxBddVaqjq9k72nJsiT
ezu6iCL8+7DwCWmch6wuJTmMpt7LH60w/fhfABMDc94XT1Y9hV1Y/nIq41sSraOYmBIE9CaxbYdY
IsbiFWILfvfxaaibu2gE2qvlgTl8lFU3wSRdKxIXjeNcvE1byFrQHF/jLq7CrHItAX6jTD+F79fQ
YNRwO/GhGuiUf6p7ZKxSTKNiKT9i8stVlsAgTnMpb6UH8R+bMNTGUWGhNmBlDT71p7ZX3Jca+0om
F2gDtV4GaOgFcrCGgVY4M9iL/B4kI3k6Qkqkel67NIROqU0JRnTtSMPcI0D1cQ7PQQcnRJSntGIc
8lEaOunVc6RuNvH4yHhnUaP/zmfd9jMal9mjIo04l33LmAg0Hxb7cRthXPJt/UOy9NHyocojIOp5
euSNFK2X7ksk+sPrNCGOxbkcnpohlbmDiZSJyYnY60Qb4OvuCN/P8X12ljyRe7t8LihxFnZyw1I+
rnNouCIRK6Kj4GMQz0RJBA92UscPFbYJ2/xabE75aozrJMjCue6J/x8cYEhvsSITinnsAsDJ3MRM
nMJAin+/0x4RwdtZuXUsNTsE/Zxa3xERAD24LfbFsaVNMH6V0VXtsVR9cVXRq6yL7nQJ/WXO6DW+
CWti2qr6kNwchtmN/kLd2WxkLFtNM1YaZpggceGGCaZmNO+GjO9X8YyfDfpb26IoD8eB7JcMgCi0
JK+c+yksSOKthDBkAiKASbHxXy6ahY3EtwsW/X5H4gS+y+du3TN7OpFyG+Mb+DVsy13iUGPKytp8
DDdkn1//qgVUpPHtbmKRPaa1utKEKJa4kjBB2qeU0+hg7pzQ4uNHJXKuH1TNuu++KSGOWfUF54kx
y1JVGQOl/EoYL8jmAENZnBa3ADKrnuPHnzGfpP6m4+enwlV0ljkOP/HTauHlaseP8hVByyqDQbeV
Fa5wHOwyfWc0fJSOQyZo4zXAgk5X7wY3Lvk8dhf/IuROaAG82iTfipIxxGQknJmwRV5kr71o7DZX
k8V/4/z4+bZS4PdQ3OP9We9qke3JwK9sIr85rhsNL3AOnkxhDp4AOGIJizN9rG9SNscmVEtjcBob
hlhhK7kB0enYUaFNCt+/ClpUdhVlqQuPxXxNnnszsafm0kuPDLkVaCp33o9gCIV/h/Sfrp0C3lWY
An2bSjKLsG0y0a/vdj46hNILK4cvrzUFj47dB+M8ZyOYYFWUqUa4InQQHhZlqrddmQ63JlIthys4
ERF4OC7zrP49RjyYos3mS3NCOZ8stfWgIUOcVsdsYRXfzBpH+YYP+4liwObubjCRynapK6jtDr35
SgTGJ49yslz0TU9PaToDSYK06+bhLsBJ9RBrDX7PhEgVgFTDweDEtONv0maaJgsTM6dmmFGqCjZY
ikehbZL+GwBXm4PKkns6+RKi4xITmmR+oIl+G3mQk1H69BjNmeYM8+QeOipQTgHlXysPFvufaoP6
W5XvMZsciqK/zjak73FFpODI0zcvUORgjhZYk6qos511GcTYvkePQ1RGa3DZN90fdT3sj+YPTa4t
Bc8tLbYSoaY5e9JMzaSbkLFhK+cbBtK4qT/S+NQGWwRGRT6Hbsac41y1649wPkbsKZwuneBpe/vz
/ZAgdjFiB1TtKOJEtR3X5/VNVrubbwADJ/HYfe8nhsSqf+NVY3x8K+e4JTNhIN407YaCAhbqk/Q+
YNkpjNMHpxWId+hUK7/NUMaHE439cBs/0L2zhcAgH1Gm0yutAi9Pm009FameNDRoyGeQkwTWYNyb
AB0ktCnF3hVCpbfoNIyqXbLdPBtkL5wdi6ogOZjmn3+GKblPuIW0SH8YlRU9s7EB1enOADGrqBH0
mCRH5KDkFxNAOzxY0oxYvl0+QnbjoO7FcRyx7m1xXQlCQPbTlF5dU1UQLHN5WAVGuiBuzVNEwASK
j2Jx73AFyIalIMgfxo3tAG/dAsrNQYo0xGCB84PBD3k+Z3EfXVLSup8LdaXH8RYh/Z/wK/2Yyfab
PQSrX5QDYjHOiVaitl8PMYGI7ocOsaBZdYSVveUIyYzJKkUzAPbLHC3TUysiBP4hbk389DS8qRfX
PF5I+DPT7MkL9CWEjjTzEDO8KWpf0Qk0AUfjxC6fS9gbTL+orT/7ra+rHefTGwyWbWXvVbuGCxZe
PSRQq0CBEtxf1cq+Ft6wpLGz9gOsomltUj6Xc7/ZW1D9RWw4QOLN45Vdy93lrUoXnWtCxy49+4Mv
Yxw2+4beizeSzhz7wlZVXKOt3OqalQNbZn4kxvLsjIVQUXNCD4ifyEaW9YmoYBIZCX02M7L33s5X
O67azRfSs8QMnQMgCpzQi3rp0z84MUDfxhTg5B7pJmLdzOuR5xFmW8YOJ51X2ZjscvnGibw/mxAs
iMFk/c5iT4ByiThnYzqEF7NBiQoPdw+eb/yS/d8qJeeBtpSedsNblxHwPAd0vhYrzfzyibtBcjTn
6J99KIIpwsO6NBaeAeOcBf7c7HlgLVacnAeimeTK1xjKnweIZzzQtenG5NPgInFIbbxCBXQfZS18
jCnN5TQGtY18Ec2oDoW6KBH8NRCEHxPJ+Tku5wLY6m/alasxDIG1Hj88zU2JtGLJm7f5OERRW7VC
7RyR2B9ssiz4L2S2ivAdpOgY496IvkAGSltXdPDDkTfeTXea/Iw+FciylTBznJxxB9ZFPnIxZFtC
es1jkZq4FPTQ30mZzt38IBLscJW5Mer4d4gWBogT0hKkvXiJoEputpRD8BJBHKBGHr1taNJe2z74
5AEQPM4YE7uEh31HM/BfqdeLhSgzJbjLS4DE40P8zLp25ijmGGbO54RIGBXVrrqSXANfsZjJpfrZ
f5BNUAbMulosEb0eLQGznE/M0CCOPY9Ceqzw4EnbQzWJLATYWz9/Cr9pbhrK8iQdZ6F9Xajb62/v
zwM9SebdIcikl4Fy8Fk/8TwTgb41HNTkPwp7d71STngtw/38HUrI1YimvOLRCf/pbnlKRwmSHxeP
ppVwckoLoWDQmd/YGi1YY03ab12ztF04xKpHXQqW7JTzDqZDxbzxx3NxxAUiPpRxmpzP1ZO/pVkb
4zaWesN8rc8xDwEkheb0Ir0pFtskMVyqemm/M5xRpnVxpa+jMAEuasM7sHkjjR/aL3Nvnu4fI2Ap
SP8ELArQo2kKkADprSt/sWRCXbGBqNPix6MP0u03I2lEZn/IwQoYvXE76x2+j6TT28HPZ83zHpyJ
DTHwIjs9F6TwG5J2rrYbHw8Vass2RxVUIRvM5UL8WTh7rrNPAgHGGhgNbRSLUstKUjxN1BWSNWmU
wx1lVDyOjk94R7p1+UXGUmcVVz9s8YiZ2nKdMa15bzZ6a79DGdFdJUutslvyvWMJ/RFWolaDVwG8
bufltFnnXrha+HCdPxX2T9jQpZivOQFQHMjmcSIBeQ1hZCNF8Hk46nM23gBXivITKbTKMCtfa/8X
uhC86Z7NxOn29sCt2tGNGn62Mshx5c1XQWYmfA3ZJeoxqfn9GKF904IOgJnf9RPf5QG7AnzMkn2f
YvuZuRc7iLc/TjjqH9bHuRXtE76W89rUADmK+3OFOL4ajyXWc8VhCseS8rBVr7p/N9McvTBc2C3X
dz1BkD3m52zCTG4ncs7U5Oyic6KaVtJ7PpLN4AurO8ZULVuhwHzgEIKyJ2BNXUOTagRuBUYkzsrr
CYTjqry9f0YlxtfGTx96Hrxjh2Y61Dqk8+1iyXNae+shS4Cuh1ex3BS7feIQNG17WuUbpnKNEutG
m0eApaI2aNUtYGX3iDJEs7D6L6rbkluhIUDHlaukcYt0Eg85iFlpI41AHFXtNtXArK8ilMeGkouE
z6XHKJyETwzCWEJXS/1T7S1QoMTMsDH9rdsWc0Qvv26tmNTSPFu+MI77AnNdTIJwrQLRCnQ9KOUD
Jqvot56ANfMj8Ov2greI5StiB8ePuefap3gGntAuGfJ8YaNLafsAgwdw/TTbGCZJtQrBhmHYU4Q7
ZDAdB/9FjUuVs8POjL4dbuPgEEAGE7WIQ87WON9LyWFEP+7tzjpyDMQ1rUzrSm7Sbmy28trmS5gR
9MYLm51bAXQWI0brcAAw3ZxctsaddHSPsHqxxu2M6s4XzCMYnyH3TjuWwhmjh3L6aPNnbiF88DeE
qSZxrdshxpbux911vcDE4knNJR7tXMQSBycdirX7E8l8wqwaGqXWgucgsZheUciLUhokxoGSCaqb
8nFs7RxIh77Dv1cMB9+WBywQ3aGcEB0H+jjeRVfJUNpw2VBnQcm9sRlTPlcRkhWmTPY+ju9W9KXw
rLdtCN0quOYHjGwgofQkfoBvKru3RPYIw5DqZbtmpNlc3IIGz+kIsPkJZ0Q8ZoBTv26ja+ZMzwcf
YgEiDWdxVTs2/Jt1pOB+bv2cpEmjJA9iS2bC91XmREyqTH7/R6HZElRHWcLZ8Znel4DhfRVckG4h
rG1agK0eu/4T8QC408FMx6IyMBh2Ow/W37R6Ix7ghftyC0T4d5uPXweJjw+etXlKEN7X79/+xpOV
FYAvwnEAeG3XKktIdSelhdcREf2b1Prj0yXXAboYR7Vohv/1VfSXVVgSQf1Uv9c1VDPKRkdswtwt
JmEBKUycLBviBUrxay9gYDpJuwcZj0I7MC5A15GdQvld6pT+to6q4514rDic8SGuySLKhQQZTzVk
eS+Y/ICHpewwAhPuu/bSIhvCr2o0c7FvWLliGUKNmI30SXvoYmq5Nel9ahj4Ht95G+vl/1jYDnWU
L02AHqbFEWdgbAqFwmXLsg40lsiGT/o89qPF2dLViexqtBoU8niAF9U3z9KaEjdMqq6IME9H3+sB
ajO2AB7K7pXmUE0/ePnpj03OQYgaDTc9nvJ/WHEy06e0lzc6QDTk/lNqgwziVOrVmSrkHP9Q17Qe
C964mI1UmOhGEsuDdd2wyUWYXVmrjQcHzbYiBbOhi5Ytb6Gre/9zXxXMNFoEgYS+u6/usdkY2uoh
RgI5KLjQImbsBOknh3GXeZWkVHBs+5XLWZChaDlQ8vszr96/n1iqeKqNneD8EhR1illLueMnX2Bv
K0G7coY6QRkjz+I4F6OgPbfGWrjaCuXIUhdA6tpzHNsrbMyIXrD5iqdjvFfiRt42Pm/nZT3ZmBeJ
2dhH6BFsdBJM9iqApcI7W1I4cW445iiMLixsWekZnih76YfvnnqHeIQcfgJemxx0clRGtaoRDfyf
JKDvlp3je6Z7d3dY5Sf5XXWxayM5/2XhYXsTTz37dKf/d5mZAtDYFkAa3s2jcZwNdWyfN5lLEeUl
3ZJI7CWsj40Diwraq4+cVluCPKVYc9AR9yRCBSWWfMcJd/G2LEEz1+EjQY3fHI5bvKe3bIE6Vbqi
VsoWUPfib69ZjgzdfUr+ti/lZf4jmF4deRqBHHtGrcn8y/xz20NYUq65CKeCCePYf4DlQG37RReS
6tNnn4RMwnOXHRYK4h8U0apvrgonlx8KEJPS9mfpoaDT7dzV0wfR4+teahYTesX7Bt21xmBEHRgX
0p1V3DhTXWaGBUQMgkHGFmRicJCSGfDX+8MA5PGRAQv2JiFUSeTw5dzd+xJnrEJjfvtIyQSY1wHW
eKvbA6ZRtdP1pLbM700pYZMI3rnnpWCHmO/04pV0DxLmjC2scjtTGS8Iher9bNxC8nQTjQyLSUQh
mlI0XEN/cWnik7T7Gpa6sOlTQ+grXqKx5Rj7TlnYkZ+c1ettIzJ/tObz4wo62UbwkNi1VlqpyIHz
R2xOY1RX/E9YinKpuYpFpu93JtUElLK6tHz9e+rD4kSCiRAJ0jEGg6ixS0GQ8zYn25+o1wEDSv03
MwY77wclpcWkz9sAh7uK7GwRP20idxPij10DIJ/uyXosncawlJfzhERPy0twLiXPcmyUjOt8DG3n
g9kDjiYwuEKtu5Qd3a/YfBKTDYqVh1dqes0T/OJhSbjWbfSEfNWPRT1c3aTfdusV6fwKf+LfnbqL
KWFzJoqgOAWp/iLE23fwvjEf24YjR46t0ks9hedYUy8r9fel3Tx1+V4HxnOmxCcaE3sjukYqaX7P
2CHkKWxEUS6/NJiwiKVasOnID7G0kf7k6s41YfQjlbAItLDnA10l44CWyc6fy9QHXESNBOusDG90
+3vqKfeIEiegXWnIDevGBrI+OjbhAu22eqMSCFM+n6OTj8lHsIQu2pNqFafWn5ouB6L5bGJVfmH/
PPN7cGFnfFwjjZR7QH5Ip5vX1h6bc4Auji2sWs4BKFryBo4VxZnew4l7/34bpw40wCci8GN83Pk6
hYSiExSoFPt3RmOeV70TuUoIc5P03bOMoiaFfbX+5vnnlWiOqbH7yt76Zilw7BwqxNNpv717eJ8B
hhUCIK6QX9eKmh4vQrZzRWftcEMmx7VRpkhaVgp9199QnC+Y9frygynV5rxKrtQ8t4mdkAchhE/w
gGaFgbDt2M/fAM7gEUnw0+aEzMNeTkzraBYKRJISyMBY0TLZS5W9pY+oCzFygNXilD6BpS9cg6uB
TA550qrsZaWQQlH19LBnYvLYTPU1VQVpfb5cii8o9pYzyFFzx2oaT1JsSj/5tVBoJVP2ZSJNE5DA
tQF1jZQfmKRE6gPabeklQ9QSUcq9J6sb8CwgzBZzkBIF3MGpZegS4n1cA+KDpuNR/ONmSRz9J2bZ
BEC+BSkFQ8ekiI9+pUfESMpZluCA6BJxjSdXH2aE6qnrrv2WtK2eiy4/b4rSFsA3VFfeq61Kwfa1
xt6E3GjwukYetKReCQ7Gz9ZEfez7kuMFBm8witQFQ2Atj7R/ozmlo2ix5v+L8KwGV+GGdL8XyqeX
I+IEc+sNWTiKmZiyafcKOmB/oivDfXVdIKwWKnL/L2nPMqwr5dwLea+3A1s9Y/Zd8KNxGPJJlvPa
QsVpw8o/IRKvH8Nz7EKCEXXxX/veY4FQJJYXIheaxGRHQ5Gzpe/XLZk6RlYHijH9uirUiF65nK1x
qEHEvgVnHZY2hnLnDx3XeYXXOVJcfVPBhOOcMI2/G0T0CU4gIofOkZiI8RaY/oazcAEJsVQhsjJO
bEJLkjzXoJvhC0muvU6p+eHzKnXFlwsFW2u7sZjK0xttAzkgzo41pQD068enfK2iv9hWy4TRX2+B
16BzcTvJi55BHeNS0EHkk1jcqcZ6xYbmAgdghgil0f1Yyw/n5qQVoR/33pjZvGtMEfzkjCz2tubK
R460SfTMnvLHqZbcBI/3ga+cMbRbM/NoG4I/HQtu1yRRb+aKvbnW2SEZN13iSqnTuURgOcyYskpK
UkxZp4goHK/0RNjANl+WgNqgahu2WyS4QrIzmq4ONAOKb7k+FGEKsqzOH+tJDXJSH0v4ojimdSx9
vvlQzMR2xdNsSOVV/+UtSBrhLIp1sTmlArp8ntk5wQSPxri9leC7QZ1z/ckB+7DCuTnCi/l2KfLL
/v+X2iIQweOVx+yDAfygQU0nc7UDiJe4B1T3iiyETd1nWITaEDBifZ2YKkVSEFm1q5mbmux2ImbJ
mqlc0I1BKtOQ0mL5oCIxi+GxVEewG+D29tQ24/ejMd0wsXYgjb+Nshet2LYUQzfNMqqNTyGpUQoO
NPMrUW09N1Gq6XUMe3X+v3hZn5g6IN88wOui61eDJHqTf8hwzHTceKTf3WXdf/wWH/OPTzKTRhcb
391IIt7LfnJ6IAZ4/xizVYZZeG8Aun76H0F3Ga3IHFv/ueWpQZrCpR0h1cDPVciFgln1vGzm0jxu
V1l0y+pWpeIzRrGkWIj+0F7zsfg5dzqVL69u5najTpmeh+dBaWIF1Lpe3NcjqkTzb7GUzWVI1YT5
5UspG1pAcVfI/dllQO7Fi8KYpMqUKtx5BqCuT7OIqlHKaJYq0lYWg/XP/2fJkYxM2T/d94tfufDG
fq+L7TaKdOYnOum/cyduwgTBhXmbsdxWUEI+1NRHHIM1ha7Wh9SwB7YmBWpAIU1XVJNjUrt1mSy4
Mx7AECE8oisWYL66jPk/gqcuKQ1LSHq0QwMisItpe3oyh48B+wo21+HfmmRIXWzz34gzNR7KBVsO
aDrmWl/yXEV3cmn8ULBdVE1KzsYI6Tf0rMuoRPtZHK7C6yBNUDIk/m4OtzEXlAE0mqNpjbzjeEYq
GAilW/jQeMOGZObY/qV1cC/M3Twc0cC45UMh3QSUc+qWic4zCzJU1XiIDqZdwgBZ+fuvbJar8J8y
hKeRI1OO/M0pAtCcq35cTjIfDwvyUM4DxHmyPmEAp3NWELHmqStcsD5pmAGaS4Iq6Mf4M+odZwY+
p9LO0onR8R1I3vfS+R0z5qRU/irPwl3qz/YIWReBlmr7/O9I3zcJKf7CVWLEqNTfJwybJSoCOuXZ
8woWicR6HsWZ6dePPUF2e2B5eb/OXa0QcuCT7gWvbMQL/xCvMGajmgrzVc+XrwV5AZT9IvLJO1Sz
JD1/DINa05LqzUjcfXHfBcTYmPVeUbtRHGt5rbLZj98N8NEzt7dKDT6DneaqHkADlmik0e6iqupJ
8jELpN9rozjF6mTzieQj6U0mzP2dKYhVOwJGtc6zsE2TkB/ELsxk5ECtivbcBBTv63bQ3VR5+RB1
k6bEnDxBxQAF7wxhU+myCxXjyjdtEZyswtlBr+njwy4asEFO3mAPXBFPLLW+0B/K4fqw3XJLw4WV
9hwLYb+/U2g0P5pUMyKyAo0xkQITW4h0JyFL26yfhOEJcExf3L+dJgU6vUOoGSpld2jboyQT4IYw
+8VTVubK0Q4QlK8l8Oryic9JVJypf/GYv3aV7M0l6t1JspK+f8L94cbzaxbwe+neJ7GSeekVGsS3
tEZKLME/OGe+bGfWFDrJrRnhx3Uz97bKmxuYrNBZQ9q+MvzStrCmret8xb9t2SixPH9jXuThEH5P
OgbXdwsPYgoH0ELkj4RCbUoI8HLcajUR9GiaTNWzTMWaTHdzRS5q19uYiTMjlvufX0YYRWScG20X
X29/hgjxzIqjEvOWxchuOZIuZwEEj4PxthSk/V7nSuwmBn8buvB0ZpEy+ziptHNsOSRHyNuumJcK
Q43To78RJE40mY9D+JnUmtETPpcErN/GsvXuJNY0/EZHkjitOmge1bucX4ou9pGFQILki96OZ5K6
HGtpLngut/rG3DdKwO831t4lyHv2VNf+ap87iwT0IOl0SxDuXmbPZdXinLQ5w8Ip4z9oMtkmWKKu
QePDA7JrW5+EjYJ5yi+Q9bkKTv4s4acFvqgLQEI//Krwu10CwDIfCTHC16PejxYTiQTn1Kn1gT7u
7x885uH5qZSlrHtJg3RCG/l8VsJyyv0fzktnz+2wYg9U0+kagEZPyIVZmicD3jZWHtyWCujletZ5
BkWY2/pul2Niqw8D6yx/4abXt3I8rIOcAsxn4beXwe06RyyQ61Kp0oXd6GuidgdiY9cDmUCkyJ5S
e3M7pMUzybZgv26xYyNRuWoWetapkd2eQHWnmT+7jTYjN8vpS7x3ybtpT4sWcncGvQiNHiofrBHw
U6SdrUnNx4vBHRp9vu9SIeANa0cGEw2+ALVAUyWi3DcJC9MrbjiTwwX57E5rCDEZ6MGVqkZM5cUu
1YxyjRzlOq9LmJhAk1sxGGJPjh4EC1AmMeJGNKR9TuRYItyJQenCCVA5oCWWVQNw10LAWvIv3IMW
ap/M5lqIGm5J31Nx1ZsUnvN9fxwbztSJwz7EBwzljjCeV/Zru2IN3+oXZxIeQf6WzshtCjq90whY
CJTkmtMG/Js0hbLsR/aYb30UPM5CHvenwW51fDyFFsoguJJXtCBf6rsWSCnl0qc7MV3kDirxXm/L
B/a8JPtlesqIruVUrc33fTg2bJz0QkGqPrXWxEYzVW0gErcj5igkr35qtsFBjP+pqt7VRXtxiafV
kY3/TqAyj/VZmtxNnqLvFsFKYssh+XfaxEXAPic1K+Brf3jkXWdfXIGuRRHU9+rKnAWl+635XsoM
k6ffiKOEQNpMBJvOo3oinc3gLU/F59z0jUGIo2hyb7OaGTqjRm3LyE+gMtQk0PGPjnsCmC5v1MML
QWPW8nWO9mvjetxoPNeDAGJkFhhjKWVTs63Fi41Ec2syTG7Eoykhzfd5qM1+b7xwpxSWySi2WbvQ
SAsj+l/OOZvle29aVIgZ2YYQBp49z1tl5jv80VHZ9m6su+bqki15Iyu1HHh+xBuVUqvyjLwGmij3
Lp5v+6MK+QHVD9l9f61rVINuKuLhUuYWRg5x8x/N2QeEG6KB9Ay8gVzEOJxK7olHJe2mOlFjzJxz
NZdPFDAqO8a2ka+avx7FzZ+2+6yEDj5ylbaj8SqgZnro4Bq0fEdxXkxVxEQJrzTQslQXm8ST4Sgn
ewN/cPiLplwMS7bxIq61QpZ+sAojuNKvHSHW+cKzCOEjwz3MsRcB6Gwp1AQQ4M4lfMVjQqxteJZO
wqX6iFonDcvE/QEt+AxUgUvwJqTcLnxQEJo52gTXqkorkfx0y0kbFr8mEN7Q+Ri0CllF0zvKXoKF
KBKVQ9kpkw+d5F/2Z9KrteqDe18hUELadxHHTdkZ3hzFzGXVKe0v47u7aOtDpGjXfNWkS0Kvzzil
DK9DbnhSceuUL5lXTd2mmSmNErkJQS7nj1Dzi7oHUfu6IrwWxC333vjf9HnKZN2lzyk8pvR2ub+t
phaH3vzT81WPsT36hTx3gFDepU2GBI7MtYezswX+osZJRufLJcWwvKbLBZ/ItSU/tHLtsrVUSBZp
OZCGWWCI7D9dK2ZrKMvyxTtXZ/f+zXZuIbMLi4p9QsDXOW3JV8K4f9lEc613tJCmQ/Uxv4aE/2PM
hVzCz1fimk588uopHiWD21cGcEb8xx+cki+49UNlaWPBdlPorvNvP1eRKh8FevVQrz81/wfvAkFr
XEVEzqaA8PVIa9AwqiFiFHsct+a1Ls/dQAo7Jz+MRJOiYy3xBMPuwiz0hWJ6z90r0Kom2lyatXqC
HFSbnLOaHvDrNnq3EfH1jzL9J4fC/09cYMuKqg6Ha6BfDbo6IaKisGgXpiz2xeZozXaMAGFvsCY/
ZafhMKegp65BBqzSJ9qdVo+Qa67PZjG8EKqlMIOe+UF5vMzKFaSNI+vbu6xwWbDTR9q5ewmYsmou
+2CeYwKBvF2uFMUDb6rS7xWSsyx12N1n/peyT81dIpmLx3jz5c7p/vAN3FvdG9zLLXJf75u3BwyE
BOCZBY5RV8M4fd1HnEfURW7ojpBDD3T+CLZHVbpkrEd2HnTimXVwDP+nYPaqtNXF/qc39V4T7NEg
U753m8gXxCfh2kw/6ThKPgp34Ef87/M7sQHgoJVLadQEEbKUjSBSd/WBTcmiZyIYwB3Cpwjw4kMF
LJ9IT2oxhCOF9CgYi3j6iVe8bkPYt8oBjV6eqoWgDjbzLY/YnF9IC0juQp5hi3KqIf0wJP1Se1ZK
8YsOl0XF+0pxvmNtaI1krGOgAKtPFHk8WdQNzzTjUvVjFOtgePdtqn6xxNjoDSOh28j3KPWtjAOn
ASuLrv/PTmNeKzi31qpBNUB823g8Dkof00jKYFt5oDfSCINncm3lIu9hgiQgeUAz51P8IDTYwjoY
NzSqBFIZ9fxVwvi80g3wDpT/rRP31iewjPxYKbWGCTe+PkaFWxUapEeSbGarPW/NOJnZzt1hAQQD
YFnez2Lp8l4+6MyohipEgtkhw/8BoVseJo0pj4YlaPUgmMTbAUXq2m+Y2nKuWzZSgoFI/tQjBKD+
3WHDGnnPO+9m3vLghsujHl8sHhieDfDiwVKHNQqDH+vANnEzNFkHM+9RyHAqF3JURUZWiKQvK5QW
W//1tWRIgdtt1dv4cVAcn7CUOsvrrwhn43jhTyvWjwRmVfm4LrrkAxc8P/6o8mCXa2XLT+Y0dKaX
ZQ/OrCDsoyIn+sHuqi3CiqjaNGwo0AHkGY3u2P4/mF7bXRobgYzSyI6KKkJ3m6kCtPhdwcQ5+URe
ZNxmC6j+OvkvB3H4uRrvRXCZxCIycRO6jIcE5f8fawM0vaN8dghoF2/Hepp+/zxTRjrwbFSROD1m
WGmCv4kYJ5iR/Gj8ovAV+MTKEQPE4Iev/QRBv0FgvB4fUL3jEPI6CaJO2jwQy8vEkCqbhPo1miTA
pt3M8FhNjxSP2lyiQX+4smZ5Gk6ALaOCFQfkQKUj7lXSflsm4slDux4y/e/KZ7YQ4BdNVh/dNOgj
mr7CehKnJIhq7JaIn+pZry490xYbiG8BmFSee/6ywc0ko2J4NfUq4qFyUcLJtaDPG000CjVybGi9
l+yOt7p6qyRaUUjtO4+8uFRd4zkLiNnrLP1zhN5A8K/gOWfKMsjnH6jxJTLXEP4YZcYjONsXWP5K
8VJc1QYyl2ysYwAuw0HMwbKIiISjFlR1As4PhSjNsI/WeXkosqizCUeIzMQvMGWK1ACgYcGJAcWc
+nTVbmoLPb6jqe5jK+3sw0+h/DzdCXqgSPp7bF3E9gowMRVnnow8c5Z7P1wsDkSvFVdF2l+SbNko
wsm19nbBuW/dWwYF10LoKoO+4nd1EbcjNSz2jyggkorPr0Akcp+ZngQYw7IvTmJoNM/t74C+c8yc
syT4NJNvj1CMnUYgZ987lh6xE9zVcU708UGeDnlxkxzvB8/WGMIqEWOJDqNYD1DHW0JK2DIjFbbs
wBlOyj1UxYI6pozJOPjY0T3WN5aBMGhp8Kt+D8GaAX/dJJYYotFw/J8W0JZKl0HnusWrQJ2enKUx
8wiB+RVUXAjk+yDSPBwQHNkRJANq/dOyiwRAQ1NVVB8r5GKs6Clet5rK+1TPkjA52zMPAHyVc2Gz
omOZMctxnK7vgnT/MvaXUyPKWpCESegWJja4bY7r272eaWZqQDZ9I0a+EN4DGzvfd4j2Tgc7FUYP
o7JB/OlHRclMOH8p4Y9Iw4sKvQUCmp2gbvN+6uwwKBy0EdExtuC70a119PHO2BqPFJA6AOmMGdbM
IiDHcLr0SrOs5MkhltrY2AfO/HdIU72Kq8GGjvY7ZuHfnBtz0gWOq8bqUcED35ACpYHhjuzHeVBt
dptUVhWwUx3k3ulJs7K66MeVeSUWpiaefvY/D5oZ1e4hJ/Rfo65ZunoXoOHRjSenU6ngi37j5ram
TWNocZm2yMJ+priZfR0NX3qcAA8R6V5PmEHflQQHtV4mfrDXe88eMTx1ExVHag6ENP3iKh81ZwUC
ZFjMS9fOum4g2rQ2zi5ZQgIjzqYiCoUZBOFV6DGoKETKrAGVCSoprB1+BucE5/DlVJdRANb9f/db
/5jnzYhP8wKbDtqspQ2WDH0TzRzbtqs336/uD+fJBeaeAv22SgQARbjsLsLQnoMhvqJfwOMbVCcN
DMhY5SUmb7wIbNHGDfUbCWBVrfR+3C3zdEYGVts/ES/I77WLUxKrgrUPfXouDFMZu+b7MOpHuQKk
94l61XRYX3q6UtK5Tt2o+4C030LRPBzDnQ2h4IddmDV8igKg33zEsqXUZ7fPQkXFBmvCIgi6heO3
S4Cn1eicBNKHA5FcskhUwcKhmwBq1GaeRM0o1UcEi4HaoLzwYU1SCi6xWbWyX5xMqJd8C+6a2cjw
Oy0vVDbWEps/7bzqiGAgAf6Ppw5fdLp1y5cD2qZi9lIzwShOBVJexi+dBnfh3dWCJCesP68v2Kvs
X97FECUucBd8JUJ0CPpPMAnqPAaSRLa7XNtRpfDcoMLlxmkaf773a0/3FQvjYoz+wuowL9oPJMkj
oOEQu3+O9fleeVkeFjw2inJyukArhR+xNbfJahsYkdnCV9mkThecvcylXqRf0/jxbQBk6LaDZCpm
I8b/wt2Now7S4r4z0K0J0cSRfO8G7DwsQnmWbqe7TF04c1D4CBZrVQjRW8EyTezK7fpoRPDBR8nA
jvNOQX2m/t7dY5d1rY9+/U5R8BSXTC+96qBFhAcP9mMOk8BuVmJbdo3rRjrywSSvaYRiQsjfBaiQ
+vbbPLb7V+S+pJ49moepvJno2pU0apXmKAJVLFwBeC3tJ1gAj8PlHyEuqSmfBv1f/V5sAldRF1Fi
u8C16eYAxifs635U0Sj9ftoCYOOIN4nBTpMnoLb+1YkBAOOEqjTk3lFiQq33a/GCPRBuNWf1+aW+
OO4FTBMHWCPKs+BWGJ7EV6V5crrRPYrr6F0Fr7OUKLAmV8SyoCWlxVGxQf9kF4gbp9n8hHGnRTnQ
yYYyhY2j6sCKnIN7JBI4yyjLy3SKyymHraTiwjDvHhLiUldbPUpDpMabvOpvg85evIyMnV/r88cG
y3u/7eFS78KrjkYzS5/rI5xc2n+oRLw4KShMZLpf/BWmZiuYsoHXB+yvlcUitfsE5s0xrVb98G8g
daNh2asZ8KrjzCWXhayNtf93hotKbqlqWe8mhZsYhVZGAQG1kl2sGT50J3CaB3iaAaGxF703jckm
b126bE8qSDwIFlN4UP5ZwD5JkLs5xonzaRzmKQVV7aL9UVj8jbWw6sfFxLQsWDN39AwcjwSHLQcS
9CnJzijbaNcDEoMa7rdBq1tD3WiyNULcZn6kJVKMjvHa2RrOjQBJWr2ypGiF//KRSd17Jt/pX75b
WmmmdABofCvnguFYoC6Viao/2VL00J9K8rJcbPtqkMuwtI2uNBVXBAaQhZdWGnq+M8T4DniAeJ7d
s0VZc8foYaKt5GQjH/jQHfDmj4OHZM5I2qUEZ8NiF9G7u+hWjXqHoPDhObaDVGq2BWiRsktAjwcR
OCXO0WKDSdTpZcwn0VxPxMcuV3Ziuq78AMVBoNvmtusWtn+DaZ4QxNCpwF4BDjqgKn0AZCdUo88W
jpHNMSLeEv091vtK0ttsifyp1ddFc5z5XOhaYJ/uJmE+WP41LFJ/WU1W6TQ8Q9wZoOM5faodLXhH
5hDAvUfzFz19eUhctUvgCy/YVFpSKfhDmg+neKnEtcM2j7uhAzapV6mb7pGufwr6ALvHZ0Jrg52E
WoVGRwwAafwpT0IOA5fmKgaMEMUTfO9cSJZqSd1gCrkCE+y6hUhet9F5EMLUpCSe3YfKQpmJWE5H
c1ELPGO8e15cwoE/N7wC1r7oJpDXYt4FVdsubCAN29bnCgwuP5f57RHhoezEnKYF0lT73poyKUxq
8gR5m+mYtccnB7PFVbnEVMD9GUeZzuri71FJxfMWt7EVnlopb/1+nQDocMg/2PJT/c1Z5zueOeX8
KKaH0LbiqD/5qau+C2ima7ASoZVI9PGwyKFxd6eaFAMqV/Q3aXeyfnANEUg2WxSdROUvTorjzCgE
/rbXOG/PjOo93mEIJ34T3TthrxmLNwUl3o8BMjgFiqeeT++Jr8xjtByKA9wC/OekXLl1Ybi9rkX2
e0M//iv4xoH3+OeYoroKEsz0OomBXe/OWV+iij6bqd1d5aYlTIZUEJPrVruCqP9qlyplGv1X84Zz
MMUXWaMW5T+dzxXlUEwMMxM3bcujKBq81VapsAMbc3WvrYHciT3tL0Eq7NrSDuokhEcF4wnHxUgD
G+N+kQdGJDwywKup0nL9v846e7pEr+H4vueW2B6Yo5Z1bEru2QRIabSzULI4Tf9Jl624kqekjU1h
dCJ6U9jw2Rvvgd15kgWv6r+X1rP9xZqDRRt4Hr6zfWWgdBlWkMsBGkSUWR0bUy67dyz4pPDPZ0SE
XhiHv6VXnAAH26pFl3EjRF1f2kXjWpbi2EbpmM6jtAlx1lOWVLLzYUtFDv6RB/2YO58coOmtC+/T
HnCR8SCR37Wzs3shNiVZG8DgsGS/ersa/y+4LfQ0kdLOcVPNIRcfZ6o9/Acw1Mpns9VA2HNwuujp
fdde7WvwRmUKCcVWcepSz5zH3AkUH0sbUgngKoTWCeNmok2rP08it/fkDDljjekDBjj83mLmb0WP
O3PwH92GTRp76Bduw9cC6O8PYrk/paf5CY4yI/jNETbyDBtdgxzuUWkc1SCWQXD+TTP5yvn1a3Nr
Xmxh8c3EJN44dZdIKt7aJGV9BUlAlagda+Kpnk/kC803CUSu4klnwDVGzoqqkwsSmB9Rz5eQPqK1
n+ddIlJwakrrnKBpD7/Z7t2JoKf56niC++gBgn11UrEgay0FSCHBFrbxcAufA5khMVay/y1UqZ/V
lCIAKJXIC/KFxHvuvHOJkAuWGXECZrFmu43NTaoScNz7gGNG2Yu+5Y0Se112+xaIHXy4mdj2eKXe
MYMWqmUB2HBMuSUc+qSksV0LBpG2E6EiXknKZQf9LJW6VFlsjNBll3zmgyKry9v5KKJ+h3lNMMzr
UUFAPSPYFqkuD0NAP15yH3bL7O2lXut59PPXZWxzFzWXOap7pY+G5Vz3pLqHdX4p5WS/BpRRwTKz
dnlLZR4uuEqxSWyqR4Iw086KFsmqMLt+LYpDJdbjz9Aoe6JbO3Sku8kjK8Tyz2J6y/r2m1n/+JbJ
0crufSDFnD70nn2IsZx89z1Ni2wXgsvZ5ExP7SYl840vpjbyN23Owo7hLun4SYJHOtdnxYnx9qT9
Zs6yj6Bm3chYEg/tWN9pSqKBfH6rYNazhotvprsb+ARYaNHrBj/gRpJil+Yi9VMETzlvy7blbQ3K
Bd1QkG+d+CQFfcMn/wFe0Q7rh89Y4HTiXJR7hv1ZUGA9hzQt5/Zkwwb/lOeHB759Cq/kzAM0xjtG
K74cl6cCpXXzeYunZDVdJCAIbtPgxDbC6KU6//ZQvZTKA0hde6a1N7DWA2kWK81JixAcNRfCGGvl
iDMrOAV8mwogzPAR1R5kXBmhQ9b0cy/wElH1HL994PRH2kHWCuZujgHPKfi8TgM8LtDcdlKG1thd
4npUqxpwTX8nDl3n9dTVa6rbtmpzopSoOdkITwy9dKT6kQ3PSkrN6qxvFJ2icjOZcjJsNLzstAsf
zHLO3fN+uBlUH1vY7u1df4q3g1dqiDkf4WoLeNGSu0AR3cC+/n2uhTBGgG/LBtDd0mK4ArD56eoF
T/obPl8Dyj0JhlKBcGHvQCcvhQx+wsOV1YMN0peBzijPK3f5frWwH8RO3WNtVRth9Kwe7TfxUycW
dn2SK6Xr5tcV88FFIutYSs7TWw3wGFtsiLjb+xAbi+JMDiT0mtWejdt28+wQtDCzus78iUJVrP7D
WfO26uBId2CN8REAr2b1IsuIBlX9KzpG8Y/8+LBQJQvXLHR5enXg8sZulVORDe0hVdyheqyNVVbz
njO05HzHkjk/2+oJUQXgNLnEFHzHjqFCd8QFSSYfFUWtMCwpIFlC1W936LAQmh7Ei7zx/cdDvHSX
+l6gR6RFndNxobU6bD2R8dcE4eS2lPAVdyFqQPJWVwkShJpMyZ14r4L/Fpr4Z7FhNCxExe2eCOKV
I9XSttuJXU4PtLS5ShOfgGWPSVE53n8iAy9tTrt4CLMdtECu1/Rvam9zzayf89GGiN4cUDRhSIT8
xHdasDuD8ZIFb0KV2Th2H6XP+DEeONnYlgNHBHHRIjoXei5MoRf4xpu02BwkVu9rqm5JHgPIY31b
MEK/tZW4Qf5GirqKCpEcyUXGKqIOsOnxUlpnLrOWUWPF8hxz6+u6ERWt+w8VVQayaSs68cwzZk7h
sFXpOrqfcqdGyawLfdTUxE3epeYbpqVNydttJqV6SED/VG7iSnHLCNaqU6zzpx6KJOozo52jnPSn
zzXjeVB8WD/NUC3WiBq6w7/ApBDJjewyR8gRdvl4RA5sBRfGMGWnnHWopGlP47xamJQHfqW+iXtE
t6mRr+/HP6IFEcYVY+mvOwNJ9f9igbkWvgM0fHl6Y0mV6yDoHB/qWwOEbmhVlziILdmK60aLOd5i
4evTvH05cbNUzmcF1jRZDS7I778rCcTpwZdA8yjOJznqB+qD15rPORdQ4hyFm22mZua951Phq6lm
kCoS9TV2ORQWaNuLCMhNYTNUhSXFjOv9ykfKzdcfYP21q7Mhx5BulOUQLhLiaMrlg+PhBiwV+/5+
C9R6zrV1836ErmVPmOrg1OO/qFZJnDl/4W75ZPUZ4sEzOH89xACevTaR9dFuqAyycEtovyS8CnDa
LFmiqJCbVEw43MvAeMvN7Rl8k8tx7sIIta3cpKCi6qKl9VdO6vM3iq7UiL7mBEFk+Vm1YXZPmdmr
Hwk6izgICRc4rPrDu/oNoKWLFcmDcwaJ0BthG7taxA3/8YzrkrbY2aP26DqTK+evJEKdi3W/R50g
CdbIuE0Nny5r32ZmTiAD9wJk1eo6Zds/rd2yLTW3odS3bqogNb+f62rECZ1L+td5c0W95G2dmJ3M
jfGSBqaEQsvli7Qc05Z+nzvMgnC66+BSQe+P1LRvnm4MM9HFXLYPtSpnktsZZtT36z90dkR88Y1o
DJ46ESPMRB5Fe8X8xP3c78rDe8+VMgrAN+3VyOaNHhB+gRIMesFhzyjGEf91QHHHORYeIJmftOyf
X9LQQEG+/qT01oO2D1KYzyWVNFXg22Rt+kGlw0TiOY5JGIEe9Fl5RjZFtYhnu2l2rpm2ieGhkqJc
Md/b2kVgtPcImD3THYFqAKZTQsXdD7CL2cZT+Mff9yFfuu8JXL/oftWpXolb6a1KSD1i0JUAnQ4Y
R8rEDKm9vNEivTEgy14hQ8I/AOtvJJ/xJX1gtq8CGKLN0LibquQxavi5xmIugrRiUlL8XBnvNUlg
E+Vlv2j9/D4RZ+uyMUdUUOXPCV8+30zdf2jlPAFCJAQzNjpNKye1syekRMGQhjzWjoTZIcd5WkzK
nAekFEu79kBcm8WTMvGMU9PHvsKwdlQFOZ6tkI42Qllk+ACcosigtg0b5rppoo6NlhZ1MSBcavHg
EMRjBmmt4lMr5vznAmcWUH5dK9U2cIiFiKtJpkwnj8JzyAVFGWR+k2BN1Dg3b2+NVBr7enh8GaBG
G9OaUc9j8Kva9Q7TD659ppIhYXZLnnCO30bsh5ckQNj6hIkDHGvGQ8ORgmNt9GbtsnRNr74s5qs/
79NPf+OtignCgmPEbBPON7s6yW0Jrr+CwhidTmkeuEsbAQ/qZO2sQ6Y9Btq8b6Xtud7aZTKPsFiH
jdap1wtxU5uV6tT7K9wyEJA9STHFwKPDkpd0rg9nLVqRTi66uqeHHXz7NWtAt2qugGeTtG47SO9c
BqKUxN69b4Tf95+Jo6kz9rkH4xvX5fDmh8vnfAJ9vk4Hx702HpifjY5cwDOjI1w1FIhOcIMA+AX4
g8RUuquxGRmWgJZ1jSik0WvLcfYhCgV/QkKxf5du8fjzvBBz8fctqWMoAzeUpjsVBeKQPgKoavix
bn8jpjMpI2x6oG+ezyJ7zSiDQ1GsUH9U9V4F05/edwQ6Ik7Y6edzxyG1s3vwiGrY8qgSInLSfj7L
P32aANB43B2fuIeJGfHxuBwufxEDBIyDVrRffrVQSrLtsUCbulje5zPkW8jAaaAb0Cj44kSne2FG
gJcyNGzBGn7lAQ7o+JT4UmNQNVFjAoenv8JYWP7HQ+JLuvA4yMjyNseJqgPEGuBEXfn9qBaSZ0Xf
jnUvOzvufLuGq4yrSk0rsAutKnSZu6MCVAYydUFXUWqGM88sHLCtuFipJ+FLslsfQPnyeDJUiIqa
iFRvKsbqClMYcut8Iq27SS/yBntGUKfg/lBCc3cqR9einohfhClylMQB1B99J3W11CRPgkITwa1s
ssMD0GmcgzolqpnMO0c82tt3UMI0s4kbxsf8FqZMOvEhgsZZJUFPyYr5kOQMUxAxueVTCsbs0aKf
V8BFojVYhZ+yX0aqtMnsO3VVZJsvXlHEeDDZr2jpyPc8isYzqyBSUJSH8QZljtOSP43rSPyEsI0w
M5xnnk35/QaKNpedfvOreDBo+fnawvSevDKztWadCU4TcRqc8KRVwX/1I25lCkftOI2vtLYlnLA4
JcSyQVYeHjrv15QOZbCnjbh9KNLHC1LUnnhkx2S6Fpi21kH0Tkv/DPG7MpDPVPwIlEjw9BSPdlIm
fJd/Wo1ezTxVYhvR8uageSChvWbNSZRYbvq3cLmlseomfdFK9kyBCabDMrp77D4zKIDRT4xUxoQZ
+TMPhW9HI18iu7l6ddEHTYKmlhKCOI+i6SnAjtHa8jKkIXJTaa1Q0PYw/k9lWkxIrkPzo2EizsuC
DxjLqV+lVunN+4Fdp4qKcmzPtno9amZA+L3IsHvev+hGrNKRjHDRHKp3g+4WKPtIzcu32AevFYCY
AuSH0jJyPka+IV2nGRG7xKy3M9Q6JRArCApq7y2mAFO/CYM8euAfhbPi6W87A/YwE5o6unI6pPkf
n4p+S2jOvJ0eW0+CYjlOFsczIgRF99l/H3nj/8laDjvZ8aFg4xsKlC0/KksN/uO352fkkvxS6F5J
6Nhc5xhrY284hyQ47dB7y0qwfdp0hmUWtfpooct5L4o884A5HGNBWXfw0+4mT8qTWpFUEiw/Y4Dq
uChvFlXec/k8kjJfGoqYkx3qGEB1fIHwu71WIqMLR1IUuxVMcaNIzhPRmVMk6HvPnhCAmvSTX+V0
aeHxyWYWn9KvfV6i6Bfr1L3Kxwtf4rmSIz4VFiPbkBLc9HQx4ZOhoBJPRkr7XDANhMqahN7n1fuS
QeQGB9dCoAv6x+Njivps9q0sb3iYbGhN9uk38q0RyQ7VEZWKC/hlv2O+sMh4fh6tTAWtVp5t1duT
PH1kclnKupSPmK0vkIQBrnUK1NMWLrnzJOyfoyQYyqqjMVeCP+1Yj55OG1sHOKKufQcsiDo/xG0n
Ehz3xqr7EbA7OQ2lqliNE+r+j+BS/JeEJ9UwI1oYfLV6LvISnKrxk1/aeKFdTxJGIzWUESh0p/J6
qmIoixDCiAm9z35DbaLqT6n+bS0FBbwMKEG5U8qctCigDw6zSEX+PgmZjmNS+UIGxqhaGJeopEID
Qh0PdRtL7r35l8VVZxqJ0XFCWrXCnGphsAXpzTXdEoxGz5AFh8fmhhZhYp/6SpuAtRvIa+aN/XBN
y+chcKxHm0muIec/2kZUZypyS6w/KO2PdTwOSSs+SfVGQtTQsp/TLNXP5qeSC4POBWpOJ+JKjuEV
QBCPQcyZp76+utoiWISrobnAkY9rIyDnqI9hPFfst6vs/uHz4gdz/rLNmPhZ9mqWHucRbswVvref
/2YGbNIzHIKWl/tteOF81ARRBIDAiG6MTdIRSRAMJyyckF9OyfFOOtHthUYDqWcLMfdwyW5HYzch
TKN6BQenBt7E1dQA5tgfGhtSkmvrM4JYRKtWBWB9DMdjZXht1jixq8RLPerIPrmgm1nklSZfVuec
1UxnUsvdEEMCVBwKi2J+V917z2i7VDYcGXvNy3aumcqw+nuWTubDwW1i8tC/vWJKj8s5XrnvWf1S
i0B/zsY4aIwzsCbizgKvFleX4wQUmq4i44mF6WFBThhQeQucA76ZOvxWgMzauoJBbIgdebJIt6al
FnAqfSHxEFCjcW+l196rNWtojjtigfva32WSZuFjlhrku09XcE82EuU588yHdN6tq3IgdCWwnWtU
e5WHqIoxip1sOyq4zeH1ZCI1xA1m0MaRAx1+pqcws07V7Vn2cbWSjQ8wFaTkWfJAk9fz1U1BufvN
9M4SW2qSFoTcDbz1x5TeXgXYIWKMwlhHJwNdTnv0ypTVcGWzbGIye/s8xgLO/dfrh73DflHzDTWC
w3tIYpKTyffxjWEw5m/bFYXa/pGi/00Z3yERWKF/XKtad5V617CF+Mss+H8wEBu1jggiZbvsrtG8
8SNAKhEK0KH5E2KT8j+VBKhAML+A9tUBZBlILVPJHZwLQRuhIowm1T7inFxmg9AETc/JQ+fUJEJc
yghPDhDhG55goH7dOA5KLLHRoOaybiEv3FgqGAJZ/p569pr6M91WyqnpBj3SAHIUh5tBZdBModjv
6f9C9liMIEzniTpGSQ8eUr0RXUS5liZhaBcmLE10+/s0RqxZModL+7I3GtBD0uH7lgC3zB8FxgKa
GH+dye3bpUrbO8kR/5ieWi794NA0NgmxKQCigq8xkIeUQsxoyrrQOEJtiNnlk+JHHjNEKZnULCTc
M3U3rZGJmFVhQaaJqeKXQANlC+U1oYx/rgwfASCxavcgH4ZHsCKZWKwBivLjM5v7/O3TMm1Eki9g
vkqWiOtQY/UynWD4Da7n/gMicXybaDsravhQuIDTHh9Ay6ZaSTfiuVSLmgiL9LPbQP+E8mVCxc1k
Wm1OWhsD8APIRG41KvHtL09K7Zx9Ceke8j4cEazBzOBWB/ZCKi/4hiWR42aNHITGVWKnGzGRic0d
61NC6q26Q5CYGz7L2+cvdo7bufjfdbekJ3WDSd/8VOnakvVxA8gG/Ro5ARLX98PBfkN/Q2L5vb9/
OUFOUIqWWmZ+Z2fcrDWniKVa0b58CCMiKTe5tq6G2idR96zPaQJzC/0l1GXgPHeH9CDuZv6vxak+
N6ft/CvjJszVoCjkkuijAbLApu8OGP2BhM0fvnFRme/GPEG4x7BWSVNt02FdTDdYIpsg1RMhOcNl
D5qXRm44cPfPjNuEkeDVEZE8m9iF4xTiykT3hK0mTFDfyvf1nG+gYFKffny3YDfql/B39E/Ld8v4
9jPlgtC535/w5M66b9qSDsigspd3jMhdcqWgTQiEEu9BSuft4SUyPmtJdVq45RG66ByaemgALCnK
3kTdclIIl8yHc4zIytqTo/H+mYJstPLOr3Y5OJroWMQSElULzpzJ5tbcnyNa+X8HjnQC/jZeZSLX
mrDiInMxsWhVRL6k7nvHbf8M9CJ+FLAtWf3GuYJgXTm+wBvQVwYvusFXzGWoXegE2tF0IKJ7L7m5
2VUVSfELVuiNSK8bg8qvyqPZkw6Xx4im+5GTd2BNt9TYvrUs9GjD+nKg0SAdoWYSJjKtkeYro11h
CqKaN+hQ3GRBetJ3OUD5VgAxPbC5cy0nEc3OUz4UmMuWIa4f79HbHLHKb5xBGQivDN9XS2Ro7wMl
gl0QPD5h3e+N4mRPSrX45eI6GNZcl/ewobSr4ApiRqjaQle4hsFwrNJ8aYArxYRqUwo6jo0QgN3h
9fDkdtlTJudBw+ltrM6IyNcnjjg6D20UX9aWDQ9w7u0hMmR7b1E9bXPxu7mbmvFsOBdlCawcuR5K
bLP5PnLK+Bpiav7TwVF0dHIjE396d1nh9zF/P7EKe2IaPk7n6UDwWdDS7XsBcH1CGWMX3+xOSaN7
f/qBEi4eEwyox1NIT+6TMHFlM2//uJ9yBlVcdRH+JIufT07KWFc8yhnRUBNtsgWA/wq69D1BVbkh
S17cVrRG2sQAcAjb++9C4avcFiRo+9++LCmLBWKLktRD/6UJBXSIKrfJ6fb1gx1z7LH6IzKKLabJ
ypnxKT2OTujBlTyyZSmpE/BzQ/3W4vUl4o5hGxZ3My3pDPdWE8UHWPf1lSa6pMKwCTExgslaTT6R
FUruVnfVGKU8b/dFsTAwlGfTSeMl4jSKIH/xXPN2anT2yyW/EVHN0jxh7pbWz8E2wsurrubKXszs
9GhN4Hq1SDDKd1y2UrF3d6PXOcNyHC8Us0adGqC+IROWfOkOV4j+w+Czq7SuOdTKvHOlLHdsmFXc
V6oT/BvjdjnagXPERs7FSAkCz2TCrLnzyDGCiWuFcYb3O1lq+uafP0KmkIUp+CRu93vqD39jeYE1
u0e+Kl5Yp3sOXL1d8ldwCGiegBQHggTFDfxUfUx1+EVTq51AGpIzEYdDQdrxIvGx49aACegiACCr
fnwhlA69RcN3pt0xkeAaQecTnupN4MDIUbCNbA+nTOHuwOYPR1gQSaVfg7GHNKZbvxvtAWv8e6Qn
S+bf109EBSoXpIIXSE0GJn5+kJ+p785qeH2FCVYGzl0HaM/6fiQjzAdGMKctqtZFxaOJz8znWfYs
FdAr8pDdoLhVUFh7R++1wB0moBniFPU8HLGGw0bBHUiHJT9FHOKU4JCS65p8XR7TFD85a9emkuqn
OT9QtzP/Y9MqbLeMoBXWzOGX/w/Y+L4twAzs4sgl10DbE2kX3iAvKTL/l+g8SSEr245k2VKws/5q
qSJa86gUby02CBYuTk12PBalELbRLVUzhSrn/sI/4fX63rg8qDghOJT8cukzynPSw1hqgLzCplj8
JrUS2P08UR5m9kLIPqbDLN+A4D+6EBzaPS+k3+tVtlI3d1loLaa30rqJmYETIapBzKT6/7nC7wCp
JZSSXGxKOqKM6LHsR/EiazIxXl7Q068NHDFMMI9fBY+eOhrs4aR5zodjSpUdvQg18Fv3MEdnTic4
YeG69eZxkrzvxTWDNA+7+8dqjIVQBvkQ+CB8zoXfKJs2yw5pTfIYnm3gM9NLGRshnVbORIqu9rfG
GNBaJwdg8lVIKif6BDk/IVy7yyMmZVp1Ei/KHR3wDJ0rzPfcUHgqJFhm+v/OfdRV8IuAkqMdxYIg
iOGdK+RCA+OWv61fL3+qJtDnGilokJjj9JebCQuXxnDbXhDBJ24z63MP9upv4TIEKojpf5sKEGq1
yf8C2ZBStKGoDlPh32Es/x+2iarj4hXjIEPLVUfRPMl81KKLM7nyIZbhE0tIer2koRgOxyxiujOJ
FgRDYXSViCmrIJA5h4YWZcmsIW2cC3bR/3ydKI7z/Rc7AUjXfq7NInTtrJyZWZLTXitozVrCO8Ok
z0Z7dm/PgTCTeYsgEjW6eoXldfZDRnDpWvuKQujM3zH4NosW/WbB+fuvMrNo4t37RMacnKKXUncl
636nLceL2vPt/OqlnerflP8gjgxtTPel8DyvjpiZAeXil29fvz/+1QHvtQVpyFjqSi3lIsp+lW6p
Sp2vcZIK93yp2ASAs3P8AlEDqQcHQgrqnSaboGzdPEjnRBrNjLkV2TEr6fcaCOERdYG9Kt35xIob
NYMe/4exhzTUy8t2tQrtbW1/QCldqqjPJ9ipb9ej1ZiUf4DQPzdPyIWzzKI1DBvEe4XohIHf0PpY
V3nGqyfPelGrfrr2uyq0CUHmzUz0XXuSiRTXhY+yHOzNamnra9oAp6waExAhC54rHj17/nlVQ7+0
2Gdw2heYP66FvFMRq65O3PeJjH/22SxvJi+cx65HxmDAGtm/8UvWEV9UIvBJRd3EfYx04ad0RBNJ
ADt6CNHWR/1tQqCOXIeE0voyeKGnqYTNIq5EPHUn4LSAnTVZn3qz46ZLfK3cHNDNdoMdo0xTZlsW
2ZL5U2doHu1zl0HCP920mP0XQ0QuDO1R75t0NAyNKh/H1ZUiW2IBqvb3t1OvugbwpaioATAMzzbd
rURyhW7tuGT5Lh9HwnSfSBweHzEQSPS8M9xMnzGuUbf6KE3V96LyKG/Hg6RYMo75AmbrRnDdKwoA
xPU+TlRVskYpGqeOCHNPFJUmPNVOVIL5naBOIx1/s6DOhus+l5h31elE5IrtAgxjkCil3T84ZMod
1kB0daphdHeTlNtQHTd+xpH9RqM9gPyPKx5i+Dgz+Tx/LaPb9Mxy0Iz4ETOv9TpfgeF2iNIdgEBb
la3oNIkVU+dyA3mNdbvidibf7MFfj2XDAo2jFJQ30nLBOhq20whT9wwpLccG5lwnVxDU2VQq6NwU
AUHTRdsre92ESY4x3YSjGBi/HZH/IflLlh5FzVG+tdpwTaCapiWg23Z3M9zTAgW6zuVLWlP0NhAa
istDq7dwm2qrPOBMW6QZmba0UHrV3Qd61emqBy1zjwXu8o2M3evJLZuA11S/DjlH30wTcb4BMvZj
3ZopAsp2ug1+SKKdZCcc7N+z+Dt8NuZcfaq+rCWY6YQB6izZYmMP6+799ppBQZsNghwpT5vd9lld
a6C7xZab3PGb18nnBRVGDEIcAuKV8cgreLlXEjyT+vNgXifW54Gj32slh2VzOL8cwuF1I/jMJtPw
nTYwWuFjAjHl4XutlKl3UC4bsyPAvkuW0dvRtw2qGRkpgmNKMLH2wia2W5EuaV5DCCaTfSFBDrQN
36GbwqoOehuYD8m0KYLM5fx6iTCibHlIHU6tmlCrrapppHGHEX2HYl3SztuKstdxd7Q0V/uyaTE2
7DlP4L5jepnW4YYKsIH1P6uVp61baxBJUymrmyZNSZi086P5m5SH/i0YZZQgSv6sAly8vBIZ5pRC
oKXjcIT1qDgKHJA9VCgZocKHPhviQnpWDwAAWUAdba4DsygOOWDmeDJJ4MBzXD6afFxQaXJCOuPA
b+srTEFD8aJ+Z6nhiuik7wToNuVs7oCzrXy4N+tyj/AcFftuZosd+MYB7FzfyTnJya47d0J6TyWQ
2X+u09BBEY2ukvE0/YyKOYybrJab/tCRZ8W0dMJ3GpHU5kBFyq583BWHRH9UFvE1DkZguUXE8Bd+
3o0ExXEyH1ftVCRq2qJEm5v/tdwGg3sWY7mAS8CTk+wDsn50zjMZMg2lfVbGxYGo+Kwo5+q052j6
lzAxC/AoBXIuKVI8WGugb30guFIxyCS7uWchII2Slh0meZIyRt5YLKYdyE9bdEuZ9Zf120eML37d
n7+byzz6WAyhXgRHgdUa5DIFfnhtRpJLve+HCzywGfZAPW3BKbS6gW01uLrN8ZPQ/UTN/cJDfMvH
O6aw/INomZeP/k8JCcfS72IOTviy2nI3JXI6edb7PObNaBdOLLGV23x82XuXa2hsq7mfHJECArK7
AH/2FZNRKXI9duzCnM4vkwHoJQ+atPu3Bq7pn1UrGRjKXEPQe6oMteamUBXCDYzZdYucmtKE2jEB
fZjbuNmtw7dwUQZizmnnhIksulQxCC1fA29Dgww8thHIYfvkbNUuDUMqWpDD7kLxslvJXc99t2RC
PEZg4L1Eab9TD2qX0hOOgssY5KLeUiWJ7ZRJLRHOFl5YhVESu5RaGc0O8fIcTvLq9asBPMai5/5y
zvUkqcWs+8bmEo0CQoSynH1h8KssCWaetFsct6O4oFiGIcVtsUJow2U/L5TYZzA75IhQ7PytCQ7l
s1Z3jqbHaEno+FMvF20y8jyJbqpkKmjzPqXq0dQ5UxugUlVjSEGSP/he0aATnahN/yeOL8Cnuzp7
oXhyxFJFn6svC2SHEc48nlouqrKjnEM93QUSb4ASR9Z7MmRo7s/WePZfjjKySvE27RA3x5PvSAPO
UF8/UbxeDfuNWc4+qJu/BTQHU2Hv43pEVqQ7Laxn8WRD3+D7YdqurjoZzSnEw9KGGTF4M6R9Vx6h
NKkc8Rgo/AxbHHIG4dBKsbGN/QoFMGHCcQBz620/cgW5DZf//k/LcaIizEJLmwbP5HETEPE7qvz/
tSSqDMniylPJtnZGOQEQFTKe5ELotIXvFk4vR4qWNViT/oo2RFWqEzhYfS7tgAw5pLHuGny94xZ7
fynDdrUI+sKU+RGivEU6CV3d7i81dIsldyk+/hGFuf1SKTm4yCp3RlO3mY8qIwJWCrMhXCX1TdcR
Ztb2BIPGTG8Z/CFDRpfReEHwxM5z92IwCu9u+gYgBmf5TsHVARC4VnKW4bhD4pgVSB1CULuVlheZ
BxwhSkdkDirXqj1FURSDiWiRcjSzmTGeJQWb2IUTO4ueESw9IH9lDNXwaT4Kyc/bnHP+2DQe+Ic1
IhX8/Bg4nQIcx8GQ9YnCO9VD0FV8KIvIe5ImqADNyOKFRdOa5WV8KJy9H1NsX71XYpIodf+mKc5S
+ImMyGsVUXw++GpY7Njm2Pu44Sz5urAjQE9kDqdEXj9/QJvyqKlckgX02Hf6U+ZbV1Q2/W+/w6/2
uZ05WbR+Env/KxegcqaJKTqHv/X5/a7aLqJH4cKoZIfaGq8xP9u/Af/O6PdvzYJHCxatTdBjdFK1
Lws6PZ5lzoB5JjFQXAP2vDliFhlwuP+chf5Ai2IV741cdsXh+tTyMK3zjT8WE5BhV8fr5taIIKPH
ojrDvvpnVhKPyQMLAOgmSJy0nIhLGDtqiOZwXXSilmiJYaLb8E23lWz0nt98nxYAAxPHfGeAF3OL
GUkcISstPJj7/moY1Yi1FM+m+r27v2sOJcsy13s3sQBhEMtPc0iVE6MHXOABqwxfQ/CwfYtYMBhE
C/UQ7ZZOgzFzhv2NzmJvYMc6fg5Y85uIj1zetY9Jqm5FoH2YPq19lEa3EW09UBih8cfZ1uQcB2ex
UQ+v1mBVjStR0XQ7Hn2nxx26+bu0+HuXy25Y2lG7D/oP4BjMHp0rwRBJsSS3I2POuaQ/3PcVyg7P
EygzIIjNjFxAFRlaWcCHmrfpOPu/+7txuDNHZmgB6ykkevzifMzjR8bRwBwmEBR8TOZu7eZC/f2a
myHrIilEnxLr3GYkqqi7WJprya7ediVXAPpvOykdOt8JywRjOj4/D5y/Nqffh8JRKccHfx4l22P2
XIh/5nIQNf2PgZrT/s8SLwV0Kt187OTmkJxeYU/ZbdXDGMe2vMKDz9qk2S9ccz+uPl52njC9lIx3
7JLpgc27rl1iH1p7PvplZ5MSW9lfi+5BaMwsJ4t0v9FTFYe3x9pudRrOZ2C+XSY8oRqeUKh8Cxvr
T+JGRKJOomxD/lInKMJfjBZOrjDl0154J1vwHnV5wJnYx7bsY3ph3YQxbNk13ME1xHozMZCyxG3b
G/Kl9Y1VtOTXntXknessf+iYJ6pA5kHepwq0vIPOaB35soA9/EPOd7xBNajLM0p/RoccwCFa657h
qouqAaixjBDsnV705LJsRbsgSgO2noqOqp4gHMMg3c3tYJfkkzTHacAJqQ4yZglIq4z8lGo5d0UG
jmc2zsM4B0JjEIe5n8uwF5cgiJjXi069X+3j8CY+tCkAtfQyBsvzfUUeHcQkhF+fh1IVIu31Rn8O
r6FVc31A9uFmNn81PpANUcbZN3GiwqXRZM9+cpWsyjVv9Ebs5TS+vKHMJmC8kCtRAsXytUWeRZY0
XRtFodGe4Usnb5ixsmMfBCq5kc4WpMHUczGw4D5m8dhQQgjBhUnmn8vFHono+KokxDImkVIm25we
ToxfOt4WLxV1Fz+2+TodJoE6W6ZvMHjfYzx+DxamM74DPIjZqODqdERG5wTkrfjkzQ1h8FdO3cak
x4WHAAwvtqGN/EQXHkKZzUQI/FwHYOd+AZTzL4gvU7J0LpbCPI7qU0YJobaq9CbueWesX+d+b6z+
XRsLmrx9EeLVkKIt5fUenNOR4y/YxUxBVd7jBRRdE4PK3Pqo1uWYgJBYGs5BwN3+0BKyuIrIMeX9
WMEnbTxX1gbZU4NCllOOanpb2f/tOBMcPX81mOM5zRa+zs83DynLL+SsQT/d8Nj7AsAK7Y9572SA
fKy33peg6R9Wi9RgWEts7yUmpCXTcSSUkbhFFtB7AFKUD4BLeqTMlQEsIQSURxi5K6SAzrx0MX5Q
MOMoRsvHo8xeZlSJPUeZcIknQOR2ayFjsmnWbt5nJu+6Wij5Y/emt+0Y/xav+NHbTbaWBmm5Rpnm
IIm3flIwIw6feW0FVgeEXn2khlKmkzJ4TZetTPrexXlJC/+piNSz2ILwZy1vh11lhChIQWbupR20
xXzH9jI3I5psbdDQHLvcbZBWeozzQG/KswUwqOLmoQm8NFjRpWwGfDmCsXoQw1RkbImdTpyM43SX
G8uyQjcRPOYR19x881BDoxVImdMpLpnNQR8DYUBVPatJ9yS33SD12UTOxryGw0PIiEK875ztMbk0
SW6TMoH4Sw4/Ohm6KwZfF43P2H461+mnE6LbMup1gDKe3/yNVsNN2ISBVx2YRXSefkaxQ+bcLTo8
BmY/uYP2ygkdCfpfIZ1OFyxon7CxBVvT66hUbOBzldmkJ2oUD1P8mUmQKXWkVLSVoJAU0TUS/TyP
vVPtzDGF9oGtD2Qf3VBr3zdHRM1IbNP2zr0IN0JU+gqtBjpnCUKMn9HcaYtS8fcwgbqB/jiZTkOk
Kp14n9pmDpQAZwjmlJlfTCnw6VzjbUt5OtEj+WQoJA343QzokzDj7KW0LT73GMauC34x4Qx51kcE
Hy2SXYPjuVWpFMswZ0JMZgnlT2kEviFleQiu61NIN273bc18ehREOMOQJMGCDbIypi3LNRo5tkxh
cpGiYGs6ZAwfp6ZbMG73l0wVvwJUfujIfwddUYIc5k2IJTN6Qo38lrmpg9oFzLhyTNP1ZekkMgza
qfooIKxvSiGFh5ADsiqt+9bLt+bgaJOh9FsxGn2qQki1uf0q4fcO7eJ0+fxShi7xRxKENTPYg3fY
O5aUQ5ybbP9UwxyZpLYIG/VD8LPlwfjOv2QQH7WeuXB1ZqPRUycncVffHC9dsvVXv1ZCE/U35Szn
/tHaNJ5dKVbgE5H8alw1H52nN+/zaMqLjnKEo0YiUpnxQ9zgRr6Gm/DqzooKbZayGxz1JGx2YeFa
ju0dwBOR68loVjSDW9i/0LlVirU736CKONd5lqC3YMIuVVBUhEfL9O4pnghYTn4hCfxr7y1/7p9T
XURTmZ1wLR+yxUmrWzJ5IwPuPnEys8t2Z4KBU/mehoDjoHwfqaOUj8ZQS/5lzUkKkrdOfW98dEfg
UsUVwe2qerJi2bdBIl0K/gyf36F4cKpr8wu4mFmcXj/ItV9fpSi83HvrnAT+5RJoVSzB3UXqIYlF
xT6FB6Cbhmad3o3diyV0w1bvWXv4QyMviEispxgi5TRw8KREO4u+Kpoub6d7MmQ3IhqJ2BXsv4qw
ATPfvgHQPyqZn1BGs/0t9EoZYlyJvH/R5RVsbFm2P00qMCmb5LLod3D0yAOwpyyzCTpFlE++UtOj
ZxsaXoGTW4fJbHISjWo++38Q4uPTB9nl4S8FSpN1d06TG6wpjAmLEbqCpmnn1Pc/owyD1CExAuw3
SeZqhzI55OqJnyCiNexfXDb5+K52NAMu2RT4MuDV7Y57SMCuW4IEm/wAdOnSJ6ZXrq1K07eNThP6
jFaE4QvNauoAGCNk9EhP7kmQpoVIaoBYF4sbHeEfAe5oybBLRAeraipKmg4zItEbjBLnN5a/4wk6
ZIZEX6zQ/0A37OEhVrAHlWvRexN2SgjyG86qW3n95WR6nhtqGi1Wk2ItwcnzQV7m69Xlm7N8Zomp
oJEhk6mNWmIKAkTHlSmih+VJilbFiKpQJM3HyKrIM47jOK0SsUqoG24mkmKKHJm9HR/cR0VtcC8K
rrEVieHJrSDNDielz1B2jWcEEx4owuXPGdWoV8H//OA64cLREcnpe/3KiBMlKv0jL5lq4myBJFL8
aLO4eEigZJkbHuY6PuBNZ70xJRnR0OTQVtNYrllIFA9twra1Q/6ieNKN5Wu6jgHr/KNoJEwRS8j7
S/m9hAyBarg16RgAZCaBMvmAO/UgVAJD+NFl0TOpjYJyySzVY1ugEdedQRaHWMOEwdT254IZEuUx
KbXPUZaam8gSSDEUIGxtXmeGOzqrWPK5+sgXTO3CMFtpJdkBoIX/Gk9b77hCF2FUUTv4osW8IG/E
ox/U4d3kKUUB4s7r01zD08MOqqyBSu6h/GXcIrywN2VpZNtvfUhcbu1AXq7OEL6u9eNLLW1PcKKd
S00Kd8jcM0D0NDSuMognJdVNrwhsHJr2Ak2sXgUYeHMbt9iOHVDudX+iUx50Ot5Gs1J0x/8aTXDi
8YnG2gCRD0JWY85sa0ImBW6jZAJcslZ2Eexj9+tlTxf4BwlF9xMFqBnW4DqGxNJTxBHWca253ZK+
fPZTG9akg9AJOOj5XBa/I0JoblGi1SInIqzxhskTRdcGYGeXvjH2IB/v9wTZ0OSY0+GGGVwOF4F9
NIkDBlAeyPvIHDcDWxm25fYBW8bt5uW1hYAZlzyFTs64iE5C8c22KUX5GcCM3KmC8BRlVESwviqq
/aOqXikpGGar81ZjHFr9Lm240tlBVlnMwXMxzIv2UROHMWGCCwrfNzxlTgTK0XwoqRcTtWopZ834
Hl6SD5Yam1WWYDXJmbRZSHOKCmbzOt73BOzXZldzc7nPbqno61ezbBygsSv6uax0/U1dxG1XSGYr
Nl+m1DWl6BBIuvprgToOaTwVUTuunLqnKzFebWC/On28RtfZNroz++2zj572LH8o7kF89ku9hX2B
IsqW3q++PGj51fC4X7MJIsbrHF9iLZzFW8X7PqmnWu99WTSg/w4Zfvo3DeW3HEkGg33prli5Y+hH
bIMHwkdfcV9wRossnZeMTgKuWryKS7nKJg4fy8oGLLHJNnxi8iVbW9lObf0AK4jKXhwg3sbjYCN3
vRtIs8ARO8v5FzcqyY2r7QLNDbAV8di2U5oNV/4/3WUtkXRXfkJrAC60HzSmuD39vsfWxhDpokKU
pEX8hH1QgDmr5O1PZEN1oN55LLNpuDwbYrL2o7ebOSklRCam075GCdVmaY23WeZR3aj++V8gLCVG
qeanOa64axYRmT4f8k42MU0tURry2mtbftdhVlFi4xanopv1F2G4LgdNO0pvk6glc3XYJzHOBEiX
aeF1zuoTQJ/53JAdaYd+e+Dx4UierFSMMWqaXRR/K/wPOn58KuAz9WSh+xE7wwkkYjJDwys+BaUa
fpcbwr43HZh6FKYxP8pjRKio4EsmVijAtLfk6YZ+ZQeHwbkw3ER+Bulk3zNoRBjootqi41CL0xtB
wyoanEg4FLsjon2LeLdv7OtXWecvlghbEyKFGYy/MSdA/2Ho5bxDpWE1gONJiE1jYBJrlpoxq5aY
XdSSOr0lVKaUQxdNmpqXnRwZ2dQDw1OBByPvzeynuMER4TNoKPv19rPIc9jfTB2HoeM/QaZTemNe
Mo1m5bgv5KN7v1nHCeeMpdMQHiLhLClYqSIlst8gd5/6IpMMRR0u4AjSKwwUiJXJDl6Ay/XcHkUp
VlSFZZilWAN7g+lmfpUKVrEmxin+7TGVJBUaY4YG5lucrUByr1UnyQlmKB56q7fpWs2EWSdibjqu
ylAP8VTjBccwrHx2FUZHFaJryr9Zecurvkmmb5g5NpU70/7YslgKTa7x65pvC+RSM3ZDoBO/ILzf
isqKDjqCvSnzNsoaNltsiTPtlSYY4D1DW79bPHqDSkmLPhe7ZUXHKLiAar5/KAuzehxibuttUM7L
FeVOUhcveDIbADfXnevTe016sy+zUyRnKRQk6jTY4MRx3xZLGCWE9VmV+IAx2TYkFqAxPtpmzCkt
D4YAkcvllEevJe7khmCiGCfzoN0FupQRPlJuba8KhvAQWYL+xv29PeLLbIr1un7puirtbX4j2UrM
Y3bnwq4c36FITk0X1ZqMF4BudJI3Qj+Y9wC98yuUtaGceMfhI0V9TbYvY7OXySawvrg3pI3bDkul
02wuesHCjyHdu9TYFOtsBUcz5peeC9M4vXNLj/9ElaIEezYV2GrpkHl74dfKx7cEmjGVoyihg3YX
2r9qu1SEDlozTY/1wBH3xUU7VnIHVQGQmLdQOVOQqZx4ZFQ9tHqHry7ZzT+R16Slxcu/x94DUCnR
CDwaoDGPdYn3KA+TbdC57cez55GpKI1YLuRJjfXTNYosJdtZJzMnc3YzqGjcwbr/0kK3qz4qIJLs
g3XJ7uLFg/nDqRsHqWdtz0XZ9LzoMCwjA+2swtPHrUsq5day1yU1+8Qw3qyTuJRyLS1VJl5Hz3lF
FDG+hwt2z6API92Mu9kZTATsmS/pZuJQOC9C8r+X8nIkAtiahOqMH+j+/5xqMrutH7JXPrsPUQ8E
aW4OVEYbDHmm/jPDCxSU8lzy/MiSsioEmTLIWOLtdsn3IRP0Ht5bReJlvEb/q31L0Go1trLNgb7x
yCLjhe78eoMy50D4JyI6Emt8FSjQoFJ6PjINyGeSHQg2y0HCgkrKPdhHnWB2cFz+oCxE/75cq3RG
u/MBiWXnTFSoXUS8Xd6Y3nkhQgqRblaIGsankZpZmAxMpiGxWkQ8TT9i40D84ZbrmKN0EWeSTUN8
86AghHE8X53Sgzf2lQQez7iSmFIQhHCv3OwjvI22ru8iLJgychsr6uMJOsFGUCgU6GNIZZ7YZhDR
Q9ZMSfh0xJjCSZaNufbOyecszQM60RL7/IV3FK2R5VUW+hXRRfQ7iLK6Q5FaoqEs0sn6vSXItVWL
iK+oCICSeGTdQ2LG8aao6xJpoQDDConJMExV0K7JH8U6NtzpwDu5CL4KUgQcMDmRBScvn9gSS1rb
euWkHhy0CqTN0p3dlZFa9+m2z6mpX/TGUQs7OsfZVNoCWAAMacFzTcOOQrpGo3AF9Zt0hxl9ckLm
fbtut2G/UtJJ6gSAj5IuipM1xVVckZYomyf6crYNsTAFIRPttsNrsWC+t3dgjAqK4180WOMLPM9K
t7Ve7SlytfDQ7SfyQI5yLX4B9S2mqs9JvpIncJCzexcInx5UoM94rFmqIwTItwEvHOgvl0l2xi1y
ld9foFx6sA4jQbU01TLnT6dPl/0ScDwuhwSZGEEHiNY4BOxZqyTXT3n+S8XsoGePshcihObFdZF2
p3n7QRK6XXZxfCcr7WT7wBgr4o8+IiL2UV9+QDB+5NAQWf1IwLrc7Ojcadjha8Pk1goWt3v8o36F
xSqvEiTkKuKv7EbTHaJMYiyFghoCtkQrQ1N25dEA3bYnCPJc4+EXoKKqnXITGIoytZ4hiH8or/H3
SjD10/z6H/PGdsxY4DTZeYf+sWgm4zFWb71cYkrrv0GiLnEMqwcLU7q9eemxwtOevbMSxFMuwjTG
h49mcLY5oCj9h83amDXyQAn+7Gux33sB2q1vmI5CaqaFooMNk12od6jOtVaNfZHk6cQBcVAGIbhx
CGca1zsY5tDSgpn5tO/1MWS/8ffTCXC2d/33dpmJK0xZMjgE7ANVYTPOo1Ec5v8m/OBcwzKy3n0M
8GjA6DcOPm9D+HvUn3EgqxAAEPiS9XL2G/aOe3EGwZPL22SDrrDoPYCTDRANq/a1eZPtar3Ho5Hq
UqMMAQYfQ/XKIGY6JvDcXrSLvgI53uSZnchbi48RpJsaHSkkDMicKOn30qGMVic0BXMMJn5Biyc3
hhqGJ7CPyC4aSQXdInejTU4WYmJM/o4x6XLzGSbQ3n2H27l8RfI++fXRcSqlBeLkgzpqLp+fAIBK
LnHZjr9qVYPjp0Lq4Q5gotCYz142a03dUf1bOXaX5DxWXrEYJs+MiuOu24yqzvXAThc84g/L0Xwx
ZpNglO0IiLzkMdyP5Fy9/bRu6LOreKwJJTvanR7JbfzE9MpWkls91KWI9+xODYx8PmhFE8R+NQmR
FuP/hdOcowmlXDrjQa12wi/UKel5noe/ZjSDLZXnivUu6nLOFacJdorhqIgByi/4rx+stMUb0IrJ
yWCJ6viaz6h6qeHrAUqqOo7PoaCAItqKpu7i+kCv4ExCXYzILLBAL1eFcvw+PE4x8dFVEgOMs4Rh
5oWr/CFZHwh0cmX3rv0vq0L2mQquf8ny4bGRv6wuea1MfQ2Tyycx7y0LzbvUprUG2IgFluULzepg
2yu7ITROGqZN94CpSsXrStw0bMZ5nVgxIR5f7fz3umgXyULZiq6PWFm+AzLpis7FexvyXTasx13V
1CTozrbRLzQqzSq+/NesyMzsNfrGoYiqN6cIrBmja6apa2ewW1q+Yl0ugE7FCgjVMkR/6EyiAjPZ
4KULtVoh/afTRrwZih+ScZb21nfcs1m2A5Sk/uZ/yMnsZdCEctoOFd1F4vvQQU5BhhH7QOPWlMbt
JwFdVNQ5ayzto4DD27HRL76yVEe0qhs1LPVKJFDXor72jrSStiCkw6ME2O3NgD/OhnYSLMTNa4G1
hl5FxsBnvlXVoW5pJ7k1BxT1iU1SFKlLO4T7sAEB4eTn0r18SB6QqWVqRWEjR9HWfeRlRueOioqL
jjyS89F3F6q/sUIqaPIQcGUFc+TOUt7i0TEFoGMgwgssnhcsk4TM7gs4FWH04PitxocubyjBkLkB
LuJZqIr8J+qw5s+uF9lX1IPtEuvz94w29/plHMhL6xJzw6LQLs2vdWxEF42GrMfXlu9ZatXQ2rmw
PjkcqjkR0E3yx7f9dEYpXlnHrRDzIokuztrXmJ7XV8euC4mPH8DAqfOsrgEFFjvJQkGUGy7hnvrL
5JT3E1fplt5HZhrd7oDQxj3kM+ziGLUtx7iFIITS40sWiZKlT0ozPY778QM6K6+LBDu7lZxRFriN
uAM8YHp4/fFPAeKc99q0NBhSQjd1iDHjAW3fqkXS6ehdszFtdW5En6RItSPsRtxkvwdks145o/ka
1O1/rw+gv9T2XuHuyTfbCnu5JjRIlvC7+6TP5OUpK3przOkyOCJVuVo1CIkEmTBhLiyz8CbQvmXo
Yvu8OCnSI14NBZDVaCJdTrW7NIKNuoukeUTpaHaf08B9dqoSEgUDjfXHRSe/tX8k11NzbucO55Vv
eYa0SlAyqOuJ3nSh06ZyRSArUwTyrOVtVRsSAsaVCY6mZci8Ph72S5tvIWxiskztXTPseDSno4yl
QG1Y/dUOKulapefNgfVVWGwf+NVmnEpOYIGBmVYpMg923GY3kaBldpEaaxhoJEqtrN7KX6UERxxb
BBr9rBhDkreJQC7V/hl1i/ePZuuM6anX6NIjBU8We8id3x+vD9cqherw06DhE5zw8EFn5ij5slas
PsW7+aFfD073cmRSt2WwG0ytVghD5UAqmGGLlzA2kaHA9v81d8t/mrI2UrQu6GPpd7nJxJPy8DSw
I0gt7uZlkMzUzYUSsmMNQ2flxbLnJxn+LRunlK0ewVCHlcPPzMEoUJ/Rg0NP0bAeuhywiTZY5vbm
d0xXOvMYo6JzCqIK4NUxyZhhGo/urixR1jrxJF9rhL1IrHSQSWqib7yaheR/bdi0YNyWOYswJqH/
nAJpa3FjwP2ie7siwdrZ8oZ+r1cj9sfA9KDJt8Vr8Ic6jRCFyvsjcd27MjilegGgM1FwEID6P7k/
8cf87slXYZRwPhYZVkHaJ0FoGakAugqyAcn8gPiBDd7fIC5cRShlXFgVtlcD+SsvKoFwphQSRkTP
Dn4BWiLCNUPLr8gSE0sZvjtreJX0XT7l7B7bUVSyhUf7c54qwE8raVck7h2DEoHZm6XeGqjwPseB
58nRs/2V+tCxu3VWImoYEBmB9WAMF/SSNdCRM2yQcrHrm7a9TJu2F3QU/u3U8+tnTeVC0jgioEN6
gC/8+oSVCEsRuoX0wa97TYEtgy9GnWz0P8uhHQhqS+JYM8Mbh1rPn828Aif5btMU6A9iLzZdsqxP
koFhkr+Zu1MO7OqvgEJKWEWdEi8yV2sIqWObl1zJnGcl23fVQFFC5hT2Q7mf/VBeoHAUop+L47/C
PCS/YE3ottnGtI5TYo/LkbD1tuxBBN1kidQIx4iyNsN51RiI66rPVkn9YZv9YKEe3eB58JFJKKP3
nmtg+1V2m4UK0vuSBuXW1p1oc/LXpYQ1INrSCkUVOc8FyujMmZnpNz/Sq66qKswXVn+xZIa+eW6q
adi7ejiAbiVlQxZlUCARxDnROos6m8jcJhQRW8rSGiF+aAf4MZ4OjqwaUlhw58L4jg+BwI58jMVt
LM6W8G5AEfr9BK+lP6eJFgNlOimRj2MGn13pOb0Xdtr3LkJW1Hj6etiDzyPJRGQdB5M8UXjgnsaJ
S4kGFsofpM4NBHoOF5v5Hm/+E9pcOaOAUYk6muerpw4FEwdve7zF8z8vP3EP251VIt4FWD1kInQK
C2MQZjtfXGUG2+NmM8rRz0Ry3fJVPH48XcBstzSQbXwFnupAEWxeI643gDHrRt9E+xRBpPIBSJx4
j1KeF4hfwBE95qLvlqYUwFNoaUQmkxZrqHpf4wh5L+Nr/e4Ax9vbFgPFN9lOjsQ/oiySU+oiqPtK
SyiHrllbHsolUXU7Lw75vJU2/AiNOX/jvFXJKdOMac0dXcUYDDKI8kII+fz6AzMzImTnsLZucIC/
vm31+UsgL3pqeuIQTPQehONkjx283U1A3JPlkfqiuz/s2ZpBAumdeZRoR/4IbqQO3D2Vy7qK4/8B
rGmRQjdeyXGeFHecMzGDfyGgqcPDNBNEax/1EXo2gmpRagmPCDyHbTgQ4c2SdfI6wDNtvwTxrnDx
2OOZANA8jtJsUWu8PEjRa1YL8nxsIzpQG/Wqwwzswi51rPR/L+vqJtE3MZjeqFiyXawQT7gUKf4+
uyII/fDfeGt7kC4PbwH6BZMHphUYEIizcEorfxyDsoIaz93JyrDeK2eHJkQLBHsz5+CqjYBz9COZ
vz1apNFruywXYzRmWUoF2FQURCV7YqZgiw4Q4ndxoY3soo4PQwS7h2ibh5zVSJ1o2BPx5rD0udl8
suEt7z805m9tyiQH1rIwYq3bdQ3Jzx/ixYTenuE+xIweOxjVsu5c5VDltmjdQP4c+d7E0ut8ifIF
sDHmK9DwpRzi9nYs3PKRDaz49GsFU3dqtfKclMhdOFr/ZwcBVH5T5num/BDY/6JwPnJ0w7RcSIlS
ANb2bI20M5xyUIaS0r/TiGhmCp3Qq89nN/JYqNGxnfGtpJ6LH9ZwdSeI1TgDsIrRsv2lM5+8CJdZ
0yV6GYGzsbjH49dZFSj7bDe4AfEppyHwiqft8HFRffWDNuqQeUlNnVSQPa/5ez34bWQ0QcuwQ8fc
iqR8octL4B3eefMMRUpr+GatBSQQCudNthPFF7vnIbXqgENg3E8lTn2TvbJH1vdztCk93aDGKLFw
An5p+oDS35IBHMLc5osCtS7W6FQfNDoFNEKOz70aw2PTkBHrQc03RbAyHW7FLxcFe+a3kyBxQlEJ
5KFK0UPVZSzdCZSyj7YzPSEp3itTRBuEOzsm4rVuwdTEkL17rftfEhejz9IH8H0CHK/9G/4fgVoH
55SX2hx7ARH1xwY5IWvxQHpFZqkpVg0/z2NT8M0TtT1urZ5grJwINL4atkPOdLX36dPOstqfLigh
zrr0x1gL0sILwK6+ruKWFf/7W3uDADprPxUAtqR8Hz+KUOBL7IVOe+SpRM5XkezaADY1b4pgYL86
Vv/WKCYlm41Co84xBUR0v/KXI0U3OBktNOPUc8iOydXHN4Cmvhso6C9HvNad4sgoZ0IEr+S3OeUO
KVVHtQ/0vj+1kxytASn9M2arZfQdlhkicvyJ8FlR/AEcM2920Rd8ewfiD50fYzmtVQi8mtVjACqz
n3c4xurG2jvvHftm+3UM9GftVE1TfFYjzuhMfSHECXauE+/pe6mI7h2oB/PalBwWc/hN7hj/v+zy
gCqXBoII0jWSjcjc981m98yq18H2yiEh8/3wpkrmLr9AM0YB6jIsJ7DcmzEsgfbkVW4ufElN5eMy
OqOm1HUt5d4jY7CCpHDyWKKvX49JPCzpmVYxCMXVavNwvORnsaR2oDKJdoREC/JyaaOBPzIQxP7p
k7dtfMAdp0MPV4u43ePrRTIDNPZdGqddwLDfRQgjPZ+AhXRZzL+WCN5bKIJbW0NQgCwmToIdSqqm
4DjcVX20rmdG2XMcmNT2aiNxZy7RFkB9LbRjLbe5OR3KJEx5U8DPZMP3leGxPHz67ULOhpkW1jzI
EQaYPvBr/lW1MuSO224VZOduKjT8uOsrI3mVlAPZxLaHIolIB1/IpAIvXXW6M8cxjWsfpeX/VPw/
fd2t1CHitCqTFm3vIlz+wPiUeKHA+rIFVZ+a7MZbIoG9lOoqCGltM4AbZ0wQCcegdaTbwBD9QBU3
vx51+Ak8phIxo6mV/1Gzu2METngwOlJsGlEnZECp3YVtQyPwCLP/VJCNsnqOPaDZo8L07mgei49g
CktOJXLlcYdC8pnQgh5JZLUXlVTdZ1Ca72TuEtzLtF0/SQawPjHqNL+gHst7EYaYgieIGHOFrn8l
HZfSgFW8aCZYvYO68huzvMoNKm9Bkpltg94fq6Xlgx51/uqvmcdmpufgd/l9M2utwvZmBId+0bMw
gBIDKGEIvpa/Ed2y0Ek35SNsjqaJcv8dfeL2O20hibHUv6O9V+iB6KQj7UMVc7qFEVYHgONJkoWo
Lcp6JYo9Fvib7deKrv+/mjlowI/z8ksa9XeLT18Ek5rnA0KzlEpjyzIs2lcvaeXQ4YCAuxCYbHD6
mAZj+QG17YwpzJX9tUASPDNsfksZZaegbuuWaP1LDK4HXxJ/GlFn2N1htL4Zko13qLrZuvSgpgk1
49oG0Ssq1iQB5JOGtLK8LzBcUkrGIVSXAUFJsyjifObTXeGP1RyMezvDYJaLef2aWUemjZvK38o1
kc8UiwMo2aKoHlpJRnztiiAtFcc5E8boACNLjsP2Be4EoF8cJOKrVcsAz20YAxIyvgV4Y+NUjaZQ
Ddzn60vlJ9v+e2KL16GJDiHhMDvLCbdVgiu9H4fmRAYk2l4HX1AZyKdhfKpMFHbRZtHR8MwMtYXa
cieQlhuur6LCRbmOGTqrOhjT+HMD7XKKAEvF5iBiRiwJ0B4j+SF2lw3D1Y9h+NAblIKxb+iHwm2L
vsmLfavIpJS2fAP5ep+QBiQL7vTkgi8vVCSxhRNbspZBSVxZrB7W4XIS1MTBrN1eUFlXgYhEtArx
RFDE4qZmSEQH4X+j+0MjBLt3F+WP5yh4fIsqhhk7PXacodJcKqh0o1y4pQO0HiMiYwCti5Q56+uu
SDBPEsRx180A2reusE9nXk5GKWiyqhqip42Fnq8ovrK2XPuh1HOG4fwuJJ07awY70isOvilXEJJL
lKpC1oiDbBP7HVFN1aTlcVof33Pm6dQhLAbnfhzyBCEFbmUX6F8EI5Uq3QUMaBIPVh2KQf2uBT1J
QYXIOywceGohFbTyeludyCc7uPOpb286mktTDwmM1H17MQxJddqLhD5o2EbfHKW+GjPzi+tDd/Lt
WNdCGkd2/SudjPHrUl1APYykYAHY8OLrskxOicmtbocQEbfJ1IIrqS1tt80e4B/KXe+nvqn2wq/T
QSRpgN7ZAzu8zXt5w0YoGPOaWS0h7ThN1Vb1oalpmYk5E2Yde+xd2wWNpfk3/w8eAqAKyE6MY5dt
FKMAGTTEH02HloK1n9c4DUcD+QeBCDSNgUA1QpoZ6FpmRHB3oEjn3q/9yErfYFeXIrp3QLl2vn5U
uiw2amoRRLcFLBTJlRzcTaLy4Nxh0tynG8kv1aJCbhKkdcYtLjrb2Vu4mKfEbmWA3yg/3g3AABD2
+lN0Skn1shxvSquSZqlgdo1csUkvdlreGX4DH0O8cbhg8tGwVHEqjq10DSaOVCZikIOv7H/UwB1P
AFwpV2dT6MfXvCcROxhgM6r002KgJvrigISQbPlDu4zGmB7Jocee6m94Aj1gnVeaEQMiA3H5tufM
fZv+0dSjEeJxOIV3OpiucxmyBIF9P8/uMZdrxAeI5KJ0HfP4TXDLxMGpeENTGV+lvIIpxq4p/C08
Lwjq4eGtglsaUTFRQjMm5Pc+kXqhSTsQKdwIIINB+9WgixSb/6o3tdiOOjGqy06LL9pu+9un6C91
U7EPlYPlAEq/UBHSodpBaB/opJACfooDKrWdfYyLDx8if7wdeVSlAZBCcSb6ZSghA4Ux9ym2tV6i
uqjRWEfJ/uXAAobDD9Kh6TrZB4MiF0nQXWjidtB0J9DXtzWr1in501zUjZpIjwT2SEQ91ColwjvD
9Rs6LaJah8TRq57etLFUBagCNvZKy3kY0dOLnAdJQnfV6Ff+Sl7IcmIRKb1UffPAnP0oGSrZd51m
7GcOrYcEPepve8geW1B7VgHyvT2xWp59iydYf4YnIuRNHZtRDPNAD0bRe53bl87RkfVyAHv5aPyk
sB8nFcn2dx2g9nNe7zK8hbd1S7SXmlJCB3e1AjCnyFrcCPirmHSqnh3pcnqLtM5KwWRLO+x3GdiR
kZQUPcKpApFpoDtjcQsO3/+mRy4Fl6UPpWWMpQodM7QFjhVgHvAGmdiTFWz7K3fDX57OHkrzfT6O
tz8P31jtnOULXC6j6yoCgV7tmB2Dv3KQy+rPIMLL9UzytDqYjxkYLkNcOWwrAnslhA5SzOq2urrH
8pq+X7uNfH4RcekzBizGv+mjcN/bbssk1CWD1NJvQ5Oi1Uz3z/RPOgX360XGN9rDe+47DIluKYkf
JFHdIKOVa/6oZ9kNTuqocay5/a+N0eWve+pBBuXpYm1280CZBQ4EbBhMmnK3ZIN9VYTyahLcaqri
h8ip994uiJW1jnI10Vjm3A/DqszYUpScbO/hE3bzoWGVFHd5rp1nHgNvZjVa9M5Hr1mCF7yWrge6
BCBHb+U5+WOR23zVp+t8zosGUBEU+x2Xepswx4rTq30/TkEnrQ5+yiDQ/oxo0Y9GBfkvJuLUfFMP
ng1kvQFbw0ZwwjKt7teLrWTf9/Qg7NXWQfDW4S6FLjk6gCpwHru/ux37UJFyU5Zuy+eSvq1Vi44e
ngF93l2787fVvEcnkuHEVi2R0lj/e7LIV3E4Qhzoq+73kpZWI8Qa+VKTDwKv0UMZgdfjzh34PRM8
TmJcM+dtMXPLfgkW50LQNbChV2KYZTioOITWwLURKVOBNV5WPFj6+oFa+aT32EAschBhxnhwZ2dn
QiXEOBZZ3aWrsBTUswyrgLakvZTmuKVQp5dyHabWX5pU7kgSkHO727Va4Nr1+56TOMtG33tRg+v+
IBWBuwjt5/F6E/yUmRaSO+37oWyUMbrLPCeKeMLWOLKvRa946MxrGHQlntei+jVlScnr52+LdyYb
aJo1Q0zWn1YPNNOSsnRBxwfYkcy/IGuzhbS8wm2V8gp08gjMuZqFLUYDxjfjOwv4scWHQG6kuurc
Q7tmB2HppiKUvXme9nM3EIBpEKg2JDmmfs0rH/BiJDXF9epRUI6oMki3F3YQBXMp3fctIZO2K4te
IInTG/42BEhdseJOwqsH5Bn8Xxz0TdSLi6wEV3o5Mk/J8+6F3zcECXL8dN7qoba70SK9rFSMHQIn
Iolf7k4tkLQW903eUNScuQR38Dr/uc1F0Oq0Q3BFbdgvAkqTc+c7FtooRdJ++HwmQ9LhkX+prQg5
3FcE32S2xBerfQzJQX3GN/2Yl0kVJrVEedW/pMlpYED3sVLgtnOZhsVb2o2FHbiRDOi3jF7Uv+gK
aA973lrSNgMcvS8Lwk30zqi8WerTZeGJ8VgXyEe5cZA2gAk8yf8bqmJ0QgXDw3b3awYUTIiKc5pZ
PCByYgxoufVFnFPQvZ3d+jqeb8Kk9tmGacH4i6PGYPPvRwWf1PW38QBzR5+dBsr8YodVKYNNCs5G
1i1+TgsaJxRpUSULsQ7HKycSNFtr0cKXOSFkCvM3FaEbJPzgmf9IgyP17E0v9nX545fjaG2Enwro
TGr2eW/Bms0wi8Vq1DEF/op9sg7oNpaR23/aMWFJMB6MBFJLniuA8HM1Sn7q+ggd26aPUG+QccuY
FlFj8/j1UQeU5Sh/qcURKyECOMHsjuhIqULG4BdLd2PurefzzFC0yD7v/9V17H15F/Sb1ayVWOES
p14Ikuyd323NJNXIVRkTKdoE9y0iN9V3/kDSs+wXg+VkLM2BJPIcK39Y8nV3mVE/CrypKWfbojw8
6fJNAYxHlSAuzDg9VydBZZGLMMrEQ9RVeaUG4tzwWzRq2MlktS2rXryfdGr2ZmSH/n/N8HVPcTHU
+zjSgxTKtuWuGAC+S0pLgi6ep7lVplAwZGW/2Sst6naAW3y//+WScqTW7yN+nPzboyvy7aGkrhL5
+5SlhHTOI3zspGS+sbrIBP6nWiyUv7wCiQsqN1OWdlYw4gdo8GW2aacJuY5ogsDE7jsBk9ahsFQC
XYIQzWa+YdRre1fuSjEUIK7IhziDmZKD4Lh44Hdhy0d2qWSW7bztGXj5AENv+O99LE9aJ0xzkD08
IElNL69lphoeEkpMsL137NEB9fxnse7bw68gQGezFIKxiPHE7N0HPAp9lYjlj7pL2o0I8YyCBM53
su4Mb5crrZmWGSJpvFMPb8xb4O89eXgryRayGrzdYhx541jFqiGAcAcz/TfY1yZVEv33k4LaaqqF
f3DQtUll67jXPG+v3Wzs2PfejJly2WqqrYS+/J8KJHrve6O4yuTS6aNFeMQpadURP4k3TWiwB7Kt
tx+U9KL6h0G1L2AY+flZACU3TG2LkyDwtJuBCtu+Gd1Z+7KDrBtJIm/S513luB5SagNFWy1b2AeV
AV057uy+Qe5xoywQ01vVfBu9Y47fUyLOwRCKSRmPwLW+T2DhRxIO4S5Zrd4me02Kg6KEO7bQsFeU
ZCWmQncI7G/RYDR9NMo7AtNHMzkD93Ffy4vnh/YXUmOfXA45ocL7FncOdY9ZAkeBrW7C8hnc5/14
K//sMAqbF4OIEVqgpeOF0lflcru94xszfyE5XxnbaRvpcR1G7b4idrfZgybE0fhYDVhdmyBURx5S
j4koxBY0FcQzFcEmu6aT5LJii5YpOk7X1FGH+Zs+2OwtAwFXeFNSsqopcp2iZu5qJ3lfLK9Y4THV
T99WuVdKiWI0EHhT9GsVtD89hLRY1OEc6vYFxduQn0IOEtINMYyyMWuEQwusOkubbaVDgLpMFrKq
MC18SQL5sSvHZUK3uzMtenaOWRy4d+auvDA0jno061XU7fpC+JZ/XPebrfNoZ2IrJRiQvW4cHhFY
R2SMpWSPF/QSyu5BgCt2eEarv9nA71CiDJAKkWdBuv4/v1b5eJrFL/sLjujZ9VPVtNZE38ndRm+Z
24t/+ljkrhW7Kexd97kqIB4JA2jAy6YEY5YXsa/OtFQYsTxVUnS3iCVYphXFE2foGC4FuDowez00
DXpqEUYIrzPekSHXJ6HH5pfdUtOKUShTCszvxOxoO4h/wvch2b7ghkaxPgzFvEHCUPXVrUcpT1cS
ygEFnJSt4Xk8TL/44WzUkbODv8afzlBoZXSeL2CbkRe8CPNTvB7F7wMlkfnI9BytqNC3Y1BK2+F9
HFZ1OVYmi8r8KHsHWzZR9UII1aS3n2h8GJoemBIEOL9n0MFDeYMXFviN2S9Q8xIKVBXZL6LS8jBb
G/YFmjDu/ACy+dkEhPlkG7+si7z07iHwZzhTWlfyfDcWenlIOZGZIPBlc55ymzW7lN7dS1jSd2cM
QpvV+4h357aOGcIZsCMFzjizSGdy2PRcWWTI58zSIYOP/TWDonDbh42pVT21sd9SQYrqFkn8wZqY
xfQRh77cB8BNAdEwr+3mFGDl8m2vvvUdst0Lj5y15ZrM8OAnHo929dYo8PDQ87Nj+BRdboJoylrC
0FY0HRfez3ij7LMaWkF3ckt6Z8F2GG+ny/lbkmuYos9lpZmbCezuHTQvI0mLqcOp0E8jQsug/3D6
NN5crNOW2k6UYYIF0FK7qkDHmOwi+mg67a1tLA5sKVJo1oP1xM282k1ffek/dx/3CkP9Q/OFtnC3
7tH5rt6bqbyLwoJwxjg8/eq7wWZ5KrNSWV4qAJuQ0FFZcwid2EXefEjQtmqDFh9N27SQrLYOw6RQ
shKtNu6ntSa4Mtd1AOtJRHA2GbKPS1oAUBf7ZI6TCTlh/8Oz/zL31UJR+bzM7pYsMV0kxfm7ZbkO
LjkFiUmU4whJKOFWFhuhrbuLIDmYzPqfMUGATtGzfkrvWltyOz6PJlvdgGhpWaWok43Z4792wa6I
YC7/w6g6Ms9494rnb7AeCki0iN1NhNyWLzsgdek4FDk0SeLARh3uml8LPQJvJcaKPKahESHozMlc
V+Ad2+kEGe4x119IG6CTutEuucU0d10x6Bi0HP4FNSn5DWRC1tv75R0eRiaDJLKM6WCsyiivzJgh
LIXXofL1//qWdEqp0rwJIdptOrccoUhGH8CNc36hn+LA8EleMf+rt66FAX/tPFykA/vo5u1RNVgf
UgGfO29PFI6+XUf9BlHkaJRGMzzzq6aPkwsVuiy54UEy5+PUDVpJzU1eWxhyicBq5ayK3+z3iesx
AeobRJsPmReC0S4MhglKDMuOL6h8YIgpEj0hBw13GbqiE2AaEBpfB7yqt2l0gwh6XuWtPNvXbKdU
3thxCKTiqUBqhBN4cWzypQo0QnL1TcX+NWI0q0gdAs4Ij+6Z568DLFcAhFc8GjoNyQgOXqJo+4N/
jtWX3Zu+or1XOfw2AwA4aQ96/9wIwgrzds7sPnM5lcotTlJKzlvmd9hVUlG3IPzVRRweqwR0PzL+
ATZRa6pumkYgnksP65veYgpO/eW672Q7x+YNJyX0f0NAuiMD62cjxVDD+4BUZC4YiZkzOKOuvjr4
ALjkrB8YJ/AwFe+PUpS5QTwoQz38EY/B46L7E1mxio3Y9NnbAagLST7c4kZYc06wsnVYiErCEfYh
MSxxOkqHccXFHcO9UinJUte5dgqO9/9Emjx8NRxH+w7LO9QWefBF2sfmVov+fawcA7cMP0LZPSTW
uuFEcQfqQXGUCIqyuKS3bycxjzpHLK1uXpyrTYMH0N3SSLvO3AJuYWMT2ql6DVZHYzNNWUJFokFy
ykLmXhvqN8Ne/y6ho0ryvIHf1209fgHIhCc220JgF0jVfx4TByBF35w1WC+WHcMfvHtFULffj/e2
w5jHKLu3RIuvM2aDzW/j918G8hwhcvH3uZytcp8H10z6WftHgE++bAGUmlLD+w3RrVjXAa95YJzg
J63PxNnHAj87EaSPvFKw/jqaup69l0A1TabwnCYMkexw4lUiNAqAFpKGN2xn5ikeYEh2of46jqIi
anu+p++lS4iukZxzXXXozsh86OXhpSXEbK+u1GvyaLoMx2wOyJYdIeUtQ3WMEBgHatNPENPhWien
+XDFJrypLvL09A9bqSaN7b3OKsimWNDfxjx9a340DVEt6EqTMBmIqGyYkkkqy9FSjGly0sV2TD3+
3AtAVXoBPAN3vNF/9gOXbknrYkM8NH8cL4MfwP0c1OIXc80YA47ubs6fR9dDo2HJ7gTf7uNAMXoP
5zxkZaT4uYKkyeSTKIEpa9TAI8/xWWyQ0kSzGecJYSJ1VXgZO9O1eIV485oxAJ9urR/w3g0r/jUp
DHGeklJwgB6uRpBnNBhN+w/JTQYkd+pmMTUm32b0u4L8pq6RalQTPnvvEVgwG4y4F+I0NdmnP0YQ
WbzGA4wzH4MgKT3TWJOt7n9YjnSwm1bzWSYYlu8gJeVr136cSTyVSXPhNmJyDuKe9noe5ht9e0zG
EmRYt1TlNo2BLrjoDt7b7Mgse6ODaQCR8cRyLSqGTM9E3qKtwJdx0/QfyKuhmpf1fJyEMXnEQGfS
Uefj8F1tMPYywOdfM/GAoJftbsrXSN8d/nUa3DdYrFKmiwIOrtSx4sEqjv14nodHv1xurX7G0Geo
M+XVrc8WtOpnZkOVWsoVxfK8hxDz16g/N6laf2fAntURVVgTNCOpBHuJzQPRFkzukB0BtE7C1k17
+fMaDum5aXJayPz6zuStjGGBAQxkMKHN470ZsbM/53hriXGYwABcHNaZ3WAC9wDBhDVVXsnCSfdA
xabSwtZ18y2fMB0kZjzStS9hQ+oK1e3yFbQZnUkHB4KmeK35UQtZf0YM+XrI71KM1bvoklNcMYj3
pzUQlE0Q2uwbG/IaeAZNdF19SQ13IJ++LFK7sTqEyGpKQ4uPpGeQ5kVWRy6YU1YRMyCKwUikSHiA
HA10Jn9KB0x5/FYaxu8KO9zw11I6C1tA46+O/AMKFcrA4OBGVHO0ws/ecWo3x+EJter43j86Fl4K
t4uZlQfp4mC0UtTle3Q3l5q3djl0AcYjYcrp6p+XkzHmzO9R10u8v3CnTHyq2RB7Gz8IsXLxswT0
l8Slyl4hjeGAxkRVYCcqzL734k35hrSJqYdrFQuthKW5fU2Mqi/w5fitIABjac6jmRTm/Gr+67T+
acuRaAEuaRT5m6jltfQwWRyPKgdeZcOZIZx1eCJ+ZkPTbnCWjRLRge/e8iSA80VwQZYTeWh4Q0jk
9QPOYevXEzKnnXVPp/ZPvwCNOIKAvWHBoh/EHOv+FmLoGGw4dqKCTz8bD66PIle4Rtfro/ueHi0/
YDaCK83ajon7rONXLq2rQPVpb/zAIVEUeuHn+xwjIr7+R2LLqL1t51JpK9cI8JN5DxwgEkbde1RE
VCQRLoh+KeJ/c2p4bGi+edGASVBf3RxFl1jt5r2x+YsItbDOU27EhKirbEzI7nwHZV0KO3288rlp
GAnqvgUHYwaGG8i37iPWKg3CuMZ45s8fq0i338dSXf1CpYbUjbf2u/sCwZadS5iVUKBb1WVAejux
Z7IcTFk66CSHn/44i8eKtYJT2Ss+T0yTczzgyk7r9oKGDRZW+e9oMoD6eGqQYIb40JxOc5HbRDJH
sUAYviyDYJsMYbSCgUY3mjVEk+pbcyC6hzh04mUOf52VK/bkdDmvqxBDKZ/Qiz9YEbVQm7Tok+rv
gYoGFRmwPZWWRArhzmKez24FhRNVL0xbo04lfN8offsj9ZRcfISuu1Obl5tDk0d19GiLeKmOuO9Z
4oO+CwpwKowWHlWO8FjSCfvHXz8Keh56A0AD5jpV8jSENi+hLH/SsSAoM6GPzYUcjzwL8IgHhZeq
DyR9UPnbUy7VR6xjHjQNgM3Gy0B2Q182f7I+WSMyzipzbRD0NyBLbqfTISQ3ND67rAJZ+jUO1bmM
9Vtjw696+Sc5ZIPZfsdzxQyFDxLv6zcrFW6l9y+f3aU59V9ziHLKXw53duhia0nEfbfc4WNYRn+u
fWMbdM4pxaOPh9p4NinEN2sBRc4ZJp22DomDoLoZ1xNT6Vz69gEduF25iUaH92ZQOAKJS4XQ1Cyq
/O4rZOTsYimfr4d8319PGtlY9pmU3rKxHcp0ORD4vZV8nEQddmduQH7emft1W9sgIWYhMTz1eLeu
BiB9+X+sY3G3ly5/DBBq8DoTfF2CbcgotYlN7llKOG6BYT7kEeqWo2oihzXc6qnnZsAwI2tBm+8/
Cwz2zV7yuIwPhN5fDPkupO0RoZLmI+vZBE1tmii8Sgf2jycJl5u3kUWEJohOAQemAnXmy19LraQL
8NLr3DcO7//CXYQQQ2Ht8nS4j50fCZSUygRJiY0Ppb65BlAdZj7UGFCkoYDdVIzuinabddhb/Pdz
DH3KWlnNwiJ9FjGxH7EAIS7JYvQltqbvm8sECaExhrKuxcXbKQuBQ7kFim1QUIDr/MPaTyMEl8vk
/Qv0K883U0RxmKbcPCVrVQoEAl2CYReaPOi65rGjxPGYpc98id9YZXqdIX0Lv7F6x88za+UZ9seI
3FZfX0zwYfWqEfF1nNVGJq95wt1qKF7WJZd2+RoixTFmo8JeUAktzytGsUQk6tbF9KhFLpuChBe2
ZSQnRfNeqIQdxW/vJe5A7NLZ6z/BuDYrhCT7TiH2JfujADc/WKMgvoSUE5ZyurszUiuRVQtfPlpD
7cQrN0Sz5+qGCkBefak4sAzgVuSXSI1VqCyzIc4TzuGUbgRD0eSzu4x3lEok/oAULz97Dntl/7st
2QT+wIfJk8EYmTXqshF6iO1pG6XwqkXp0nx/x2OWKBe1XD5zT457I/rizPklVR58Sa+cdOSPhIul
ih94xrf35DOffq3/R7cOH1QSPELPj4s6S20rj/i2h4ewcvsCQ8+gOEL7+suSLMw0Vebb6auNxEJ5
7MqqQrstMauiWOeQjr34PASs6EFSt8eGuSCf+Tfc8DNmgaAvCMJPN6bo3tx29QMdoDEkyY/jENoZ
XJ6WM+OFfGshn2fVSJoRa3AyiTlVotxknyxgjTWcV7RdMEoVh4Y3m2MAfgW4lk8w6Rs3f/AQPl2Z
BgD7bysNYe4BkCESoG1tBo46LhJ8dwgQyuQ5nkircHVG2/+6ir5W9qC1S6VfLIBiDwzUK3Oecm89
IDoqRaYNM/TTeFW1QCPdu1EH96kPJDkue7KzPPshgI7Pal4PQGJ9bjpGJcA2mBTYDXWQT+XTWDKC
pkgas95jV1L0jwAyxpARbfIXR5PIVMxj/Abbv7jLelSqEcxqp64N60qBrz78PsAX6uALMwq93+Cd
9X6gE0vGXn4jH6R1pkeIWHQszwQti8C8LIOh8JusqYZ9B1BdYE5KK4y7AxemneW9jSO9iDbtuFMy
IY87nlVgglGgsaolyEghkJQWoUKl4GT68L9hlP20p2aPJ00z+aRNCXumYqmtZuTyHpuRrYgOL0SM
xm2JdjqHAbZJkvY1wEI0lcqskAi8m3GZeiJaaaSqv+aOfLgx6r0c7TZTMngeMpEMBdwWyEORePvM
GJCNDD53GiDSBSm7tN4beDocEl2rGRwG8bJo07LV0G6eprjrx6L9Ssal49VDRbsloJX9aNTCig4E
UOqJQ7TxXoM6og6XDvrbgbRWJCO+W6azC9HrM8TZmUC/p9y6sWZOe7uSThpVA3TLH+mJIFuX2P54
OEx+ZSKuBCN0Wx7y0eyBWmBKw2BZGvKWd8R+mzhYebbsCXpsQ/CSSbqlulpfdjn1m7l8IK4NljDp
+/IJSaTSOEATF3XSo4kwTABrNG3cUOh17hXsdIO/RcGHyoqOma/hB4UhiBzGWegfOdD3JADIQdZv
c05Zu32mC7PWLwxmMti6mxNZnjWCCyleN95xlgR6osZYqRuihcf3vo14OEn+GdYEsQ/tzKPpO9Sg
5GUsiKUeY1RG+EsKvwmbmR3BfzWWKJMLPh4oPC2R3JhrOpJcvpf7+3T0fx4JwtaPJvjahr2JjB29
HDE7GOSOvxwKE4tyvltIf+mr1Bp1Dbv7udzECOUTqTpfSl5fDUFhBD9MgvTbmN7vtXOrSiOGU8FG
IwRkVajm52dNRegj01UJDNQ6zACCaoBjIuuSzA71PbtFtur2OxUNwomtAxEz7ad1d1Xg5AoHyXzW
yWulZXNi1ueFVFua1Tr3umoFLPmnCyfBbp804RVgMnRa3ZSuHUXJgzZy8pR2g5TThr2cWqpONfGc
6lfJFyOxU72zSMBazLA8RqeAN3gH3o7xgRmsS3xNKYkF8IRkWaRfU/gZpkv9GmVG01gqdB8LwZo/
hDLvn9ZaL5JEKHxl6sdnew2tAa+U79nsnGOEXyl1mFXGUzg5uRM3QcNSmxm7m/iRSHqO8Xze3sVj
2FbetzScMUge4VFxnndR1cPlZnAIiIzRjffjZUEAzTV+bruqWHUSBQcbW7V1qBqMSQmjf0fa8zzu
zppGf+WE2bt1N/G+a5krhBtOPz3TDL/Auiusm2e2jbvZSElz6uYIEmvt6dukIVoBlpwX/ADsNJiX
j5WMADPVye4dtYQ5V3b0yTUX990Ys2RRIdKdq4oVxefvCV3FNOJcz2rKb18zDPGTGp7l/RKMmqeU
mT8GIiB6uG27n7F02GQ2R1bkh9WA5Dk0K268YYWsFPK+hc05EG4J7e+4p2l3G2fK0tqjXR+aQ2Cq
P04jEuRgCHqLLNLHzQ96jQNFcaKgZ7pR7fupDtXy694riM5L7Gk8X4HeKK4raDnNBOdv23hUcTVi
94ATVVISuvNN/jc3SAUxfzuyVH668BGg7Z6IG/5PcsGSqUj5JUhXB1uO9FyFVjevtoot2FdKU6Ee
Lh1EdrV/9eZ+rTh5m9FwbUT6/WkaeykCkRsgZ66ndu9D7nIKjXxAKtnLXY0iACD0AINusKoTHEVI
T3uffvkxo41B2Q07rLQR7Oby46Rq1oGE+D14A6rqudD4NlLTLyvct4wzwx+NjKTyiWWNIwzPx9H5
y0fGS90n+Hibqmnc/snao3HhclsFPLb+bYYGiX85OGrs6cz4tA8aAEOJbssfVE6SFrPf2wblJuJ5
C9tAQkO/0GwQTPMTxkIirtPYFQhzRjUGnZ5WkdPtEzJPlVm1HFDegOViu1HIKh/RVFIC5br/UMn+
QF5EVue21DIaQ8v6vtlpR+EdLTHTl93eUmSHNRm7+S70tvrSW3JXxlNG5KGy0o7E3ZGC9wm1nQLU
MNUxDcSy3WcvUQvn/JJrWCoC+xq5Nzs//FT5XckRpaVoBAt2H70EGBp8gYzCDMDs3g/mrM9eH7iN
ejLJYk4uGfPoeJ6n+R+R2+vAkERLUE4WrfvdkZdqbflB5E10lFobMjqlX8kvsBviJrq/JreOU4iP
OBDcnM2a6wtR/EaTdZaB65sD3BYJFvpktr4siGFD7kMig1OKpFdkLfUl0yxJvwgoBt6tIZ6UdtWW
7txk/pNwCSSgIxv0ebZjw+pplGZ6hLpLONyjyrwyk7tIJnUPBNlpya7MOuEjtf/VPWq+39J+q2tG
wDBEaSz0OGlEnnbWxDf8EhAnbimQiIzP2fsuaaM5I0LuZDP2UfgUTOOqGkbF0bKA9nW70m5iOnaM
jxmMzD0zhqgLDI+L3ALwiu4zMmZFrx81pbcN9DKBX0G/FGV0jbejYDI5hxFVlsEU9Wu+5k9sbhj1
/2okHhj2IbdkEqVvKWKNYjXnXv1TsvgQnJrtKJrI3US7EOrcK5bsKWgN20jSMKkZJytK1JP055oA
MsoreVaUGNNKP+poeiXlNF56XbGq3qn02870BhQz9yYyZLXv4NKuk+kgZGvc43UuNqiYqvJEZ3nA
/29ZZDl5XzC/N68jvZ8aqs5HEbOqZo1y0J2wV7Edy0Esy5OPa9qHmNQCS64OXnVhPAjEEZwrDfuP
Y7+bMz5mE58/f5+hKy4ZC4T2okMhdkiR2q2bKbAZmYvwBVQ0UFHugLkiMF3c99Ht3QuAPV0HTMcT
jUOiqpz30nrCpBG5TOQgbMDCec9deRjg/Ahk3Jh7PCjkEnoSQyaDh515xVUedaqtdhm/r8l3PaSw
vcCJSKmt3Ny8YI4SleiQ3da13MswkMCxXJpTAkFX8G++N60wTdGe9iFYj+zf9FjBZRPAhaZk+yB0
ccfVFn6K+1W7V33Gf5MS0K/teD7FGijJBybloxmyuDtR5E2F9aIUF99c6XIfGmx+LGvrqHvFku4P
FzgcHefe6478Cf+hU2DcY77bglgHF4kKDA5jxcZvJXCju+GPOwesAqm3B983q3kpnhpAgmlDegMF
Bb/Mb7HKmpZoi+1V5uFj4nzzFDExr8vRZZ1Wp5xT0GkuA1H4GutYWFy4r/5UsSFr89FW9bJWKSk7
pKnzTJ35iHvggPMzcTYj8hQlTz5DtaOXQ2VKBXYcBvWvsjiIbXoUBmprTA7mfhEIGpLO9lwdL50t
taYIrnTYeKkrTH1oS+9i2oUfqXOGMxTeXX2jxPYPk8dDRJDyFKK9SW32vz+AAXjBefudwVP+1QXQ
pymEYTiqANurZ6P+w6jdehORZ53sUTRfQPfP4PYutRmslICAzTTtGwKlxql6eXsCJAjYUrbaCFEE
+ZnlbL46/UgcONhR5BzUDfnlm5P7vyI08WC0F4HU0H/0pNh+I1T+GK+c4UfPxNhgNCcxW3Va5b4W
vrGVyVBmv+KyJ2YtfqUW/orZcPpK8my/lX+W/E+cv0zEMndnM2oBrz47XZ/LG+LNSgxEhP+TGa7J
OKQZ48hAybsOn7Z7vDC702f3j/6ZPjhTpMTO8sLUB37YlTgfJSEQCCjMDg5YVYcZ/cOiIW57eSPS
eFz1d8EKthAzNPMTn+onPyY4HsW00BQgQ4X3PxsIbT3PtooUNywfcrfXaNpKVgqRknJ+RrIUSto1
38zm0GtqQ546C1s2RG1udv5zXB8vPuHUrsSJtxS2GWBIFNn+We4sQ0MZYWgLKt4J/tWceYrcas7l
5cjNGTIMikcAlzS7momji6UeOWMb8vRaZ/f8LjwDqmMto6j6pWKKwN0A/jHfkclztmsBYsz1/Rdy
62NjqJmJjeckSP8QvkXC5Y6CNkcey6wXiZ1v/7lheR1b6AHenStAPwXPz+yeluGBV46JwNLfKfnV
TOxaO4JqHkX6/t4gB4xyuo5qcEHhgpP8VGNsfny5O2WOdny7++KWm59ty1tqYo1XX8NirVD0PFkQ
OYChvBZXOPNVn0AooLW6wY576rRQLk5o2wUM3gDdKQaWK9yIyGGGKaOH0xF/dVgSB3tNhoBnk2LS
xhey16twfw4YYAa7LoVfzqEcX7fi6RxlRVsslMiWsmotHtTGMtMr2bNuRVd5mITajCrttbTkC2n1
UMA6KhuvEI/1Oohp91vOzAmY4W0ylp6LFnhY/DnEoQkyXO4Mn3n23qXVHFh/g3P8WUmrD4/tvVJg
HpTX+F1K2L5iBWIGRMH0X9U5jY92+VOOC70cpvy3jHvgAeMxSODLuj0a+66wiqIap7we1P4+1Tfb
rP4r31h0mvPfulO2Et5RGbNiXEDu2ln9nd35kPQsnlF7AVp91va6HcUBeWLdTfOlJe8+KvzxBQ6g
rnrVvwodBk2k8C0m8i24lKOGiDlPIWUj740TizxQsg8WP9iDDlsWxrytAj9SiYxMO91em4B/m5WY
IH7urvJytWq9omkRLGgucd20fS0j0uxkV+rNzh2EXw+lLEA0EwSZdTlBn4jnPaCdnIoMQsHNxh93
gGO9HtzeLF6MjaGbaQ/hdgWbSsQReJArCR5kCizbRhyI9F8SEPI+woUDLpO9ed21RUR6XUqEA/Eu
CgUM0qoXAtzEejrv6H6LI07bgJ8iVr6/Z/6uYEq4xbWynqDD+Tb5DMVOEGyPL6OqxcmsltyI1Tkh
8CZ2dtNfBwv0e/T9yiTGmyqHxJIAY2eue1DKPxpwc0kvnwio/ZpOjkCqBoxbXwnjqYKvmb4Hj2j1
s09pKRFAhfy00oHWNKImGuG5xs+5J3FhFV+U5K11Ay4zvOzJElwgK9fiSeUlYaEaDVdAj+iAeL4F
sEMfuCLNuRvXFj5E6z43udMGYmBx01gBQ+zB8lAtv1mdusr45t48I29ja2wMHhbjnhpjWtZO+Wmn
EXslVGOglAq/ZiD7X5+sI6MCf7SsqirACawB3WaB9HjRebcC8wZbMFZSUOCrY5kOUdmlr9m7cP87
6XDi1+BoqsEHITLxGRQg96c7JNqO948sbt+UNofYthSPa8TTgkf3vWKbhtWfDC2KTl6phmoXAs58
11lTYwC9NqPXpqBik0e1WZv2cuV/akIukfSShED2FzHwww2d6pPi8KLq7Lhzzer0A7AiCAcANcXA
lfqVSr+6WRfme5B8YxSjUmcYFWrVwRFsK1gg0x8bL9cRQrH2Z3KZGGBLRycADQ3YjsOru8/g7J4B
5+dJxIVHdHY6D9vUJRrik3gPky+kjSXDBd/mW8j3xuL0q5z7bE5WXlPy6aDXYKVPU/UiQDWPg7UE
2qlV6m//DDPPlAD9SDIoeXKKjy8lGyG7WJnOLQzWD2Ii4cPUrj6DtbDdgRF6tQPh83RbmJzuePal
DVMm7T64jK3B/0pIX4qwCcaVC3imkIBJOnPHsTNUy3+kU4znSKalKfD9cYsfrwaGrBt3xED605Yw
YSs2JJW22vDpnTZ8mxF5FDJQlsH1KYRdpOha0+KatMusatuE465w2I3T9cmWu9zzgZnQzwFIMgO/
n7ju3+trXh+8MawyepDyIqcKqOm5reXVPh4GhwTPPsGconoKWu/3l6S6SISo2+FCBcMA2VChtmpv
oNMOBml8iBWEzE9vaheeF+vAFHoL4l4Df1CSSq6EaRPomnyN99WWzORANXJqVPDXUPNeHckODMmR
WbJ2M513jxslURjHaQ6LaKawJCx52Ro0wn5ZDT6wYRvxyz5n/HovzmMQPYWLPYXCBg6u0hzyaMY+
dDPkpx5CEV95au/hpceH42B+LB7El65qbYAGQKbdNkuMApb8JnW7mwznX9JJHCgu+4b199K5znSY
T64dq0JPQZknWfn8Iv4rG8WkmpYaPPxcBu7+pYQgK7qzruJZ9dNOeylfeOZjVMz2lUd0UEVw9xTk
siA60YvOynLccwfLZ+za1j7HlMc2HldJV+HbeiZgJVCreDrGot5vyupvY5ddKD+1fCC+QYvNOpYe
SKVh9p1PheZP5zzVu9Yem+zGer4ubQsIcR50lMS1wvVbOGcPr7g1E+aGEVi1QbDQKarQxWsHxyd0
vUYuG7kgW+sXRwNo3Vu8NqdKn4jDem9BHVLxmJUNHRarHQXQ02xPWpERzgmJHa54ibm3I073xAvP
JkIZ95qNEJkf6+NMIEH5g7X2X7yYEVQyXWFYLLJeV0nEtre/b2uMd8ozvLhaJIKY4l70nwWUM2on
HHQ8LWv5OjHxfMgbXKjDViiYa0mxCuu4dMEByZb8I+1rcPHaCw5lKE73knllYI0fuTvC+OB10n3Z
X0/wx52wY0RfKop9NF+heF3Jfip1duHJDhFfDh5VSbla+1R/i/1VpZgMYS8Ywzq6IqBqsXM3Nu6R
jvfVDaof3LncaX2oXwRDYBxpIiX0NTCQVVPujERGZ2QF3yYvsYhLeC6S5YY+1mNEe3EmLajbgcCe
9m70lyWwxKUmN0Cpkahv0cWJoNs0OHMw7SaTSi+hfC9XTNu4TLP0yf3PWAKvB4rAOzRa+4Mm26W7
ap8QlyjJ51+/M8dzUYRujrFKcJeWNo8jneXCfQbglnhX2PE12EaIRlPvJfhF+k08b/CIiMXwv2gQ
CPpUN93XWBNNPEQQEps/VOmOog/Fe1P3IwDYHMHqbR1V6Fxr4mMp4km/sFxPmj7OaQeiSyq6yCha
Q/RoW+IWbFPeIkhYFDffqQhDse6fe1EQIxLy5ha0svhKh21kjec3zeJEw3el2VDSrEGs26VPslXh
AEUTlhJSYW9XmQspAD94ocPu341S1OZi0b+ln/G8V/CHtrEg+OhWP0eD0+R0pQNlUM3WX2s+D8vI
N9tTuRJfcmdggUVYTWjCyTM/P8VEpj9kD62RziD/57ZAV0ZBt8fcQzBwfvNCqcuBdtM8v+sx/ckM
OIkWKlEiDoV1w02mLeCblWTDGh+74UxDx7vsMV7u9UUtRpwJl2snSU8hBeVkZnOwt9o523V3bJ6M
AGwRMD5G16Lpmet0F0hsoFJ5+dHBB+bkXfmkaewwc5dTD2rGSipi3b+c4+9bEEh/mgEynTQeyWqe
R13s5hPxcLDsZuw8Md1AMbJlvwjzYKvvVCOQd9QL3QXLPih0hJqosqgUgNbCHRTiTUmUEWZvhHko
O2oz6oaPFoUa4upvzaOD5Bs7XqU8zodZn2IbTILo+dPpqn050PrwvDDZMYVdEqmDXCEx1L7VeBMV
ZA0VZuYI4OpJ/LzdlTS+5PPyBrrTfvIrJgFhs8ZNyvpikQVwuvKbErx8r4555YzOGDSTmMByOCrJ
cEb9V1Dx9UY/rj6uTQQBgzj125XKbxlavnJi4S4dNk/GWM3rpD2u7foEwLdLDWRNcm9OyNJttEfB
gZ6ntJupwEC7dZ3w9Yd2+9n7Tdpj0d0NX+5uSmkR31JWS0BoXe2KjpO3V5Oe/CFhFVZnqmnRzJdO
Pl4w80e4w41pHwkVRoOB9jp4Z7IOZ3vhCoJN8lnIhgatl9DlUaTIrAUPi0rvC/x6ACLDQvsvqNVx
RIzU8Y5cg49E5BWYUR99uO/+xzJWx8/Cmx+NqhTvD4bT1j6yFfUtncsyXNKIS4HXiwTBsOy1n9hY
1uTQDbDyt+GITGPgsxHZqiDaUHoMLWrv6CzEnxAVKYdWZ85lV/dmAB6b+jIDsM+2ZKSPtbpM5de7
KwlkRuHMtKAJHs5O5TLaQPv35I3Oi1ptwDE4DTmU4v7MWTM614y1BS8bJkhBVrFGdqEexJnm7qRb
JyDvnQYZHnxbikr64/4AiWYhSYbdchhtI9KZtCtjUQJWkSBpxYZu9PbXJOybx1OIrz0JAyIncUa/
pcPwO/GuOs+fYyk6WobtyZtXd/nQxDbqF8aZHfWI/9gFZsOPTHIsYlRMu5TBAhB7HE9Vc6S5qfA8
LLlkx8Iheb5B+1cRoI6bSh/f/SinYYswq24revPtmXmY2R327svVfn7pQNVPP8xpiWIkokvflNy7
0k6XtO8equXuhgSCXRU7ynMScbtsER3eK/ZfwcB/KhcNGm9kseaG/9JWT9zB1PCwlYFjLkJdbmBY
+D0+SsYZh68iSgEgWx4VQPYjeV0kc1bAw6AEnvEc4N+jeefI8gbHsYdrdLUywl8iBatZ2LmFZvz4
+JPGXgKYs/xSgP4KzJgqvOMrPZgpsszvzrozCvhMIzzx6NwjsSjHEOxmP6r6ZnK91+qI2RIGPLzH
TL8Jgwizk1BbcK35Hg3p6DI3QoqwSa7C+xpOlaUfAwuKuihTW0Ie4xXMNuj5CLjDK1PGOVpTHNMM
rAdhJOpZNd/4CPwlTcUpXXBQgPoPh05j1hQOL3RB3Ft2yDjLnKj1fHx75GwKkaaMgvKA20gTZF9b
MkuX8bIam1eJzQ5Z9vTe2eNdMhFFIlGk3J/PMSy2tmhswLHYeRRgtX5gPd3iwbSMcuI7Ads+zaXC
DGHQsK3WhltxxgukWo1CmAZwGgRRac9NXRsGRXV04wcvUAxZ2r7UgVE6vbTd0RAeaCt8KDBKY94a
QaT14N8JGcoPHR24otpT6J563hdv8KiyH3uL5jB5ARqGtmivpvynp/JaGrIv5vGqMhQYQyTGqLu+
3Uw0dx839oj83IUq50gJPeoqCgppc0m1XwL++J4wNburaFyVlzs9nXqqX5WPf7zaZvDSWIWd+KZ3
JlUcZkelHBr3SyPDiKdS2Y12OsRSFsysbzxZYC5rdRO5apTu6zhfLrokqHkKw/rh38UGZvBlU2cj
l5Tt5TgbYaNqMu9Z7S415e33H0c85UmGjmVfqVeO28vInLWDotStT9zxrPvnovB0oT0snQerYSVi
N5y4ZxlcGvq6uHun48Vd9DsRIWBYOr9jGgagTkXvJucFp6A3OfNgVTb06dZG/WsMyKqxvJvwTe77
+mH7hW+kl4R80i3XrAkJDY1B/WSF2S1KeYSn7KcZNjwqaxcO3gpblNX1Up1YDiMw3KVXLPA7z/RO
5yknnF10lQzi+Han4Pt62a+lC8eoG6WswX/Wn1EwR+5gOfk7NQjSZlkLty1+gCR2gWsMI1OAdu1V
N1Fx5tsckloaA3HlXSN1zjy7A3REBJdhcLdMUnwYr0P6hkWlj3mOwM8yPZ6UymCjbeSSxxLHxglA
IPBWamuSDEnsuU+v5rh8nJjTa1SB35jTCqWS9j7ueLGRvG/yS0T9qDQObW8OWCV020Zy6Agljlwt
aZM5g6oGPph7ZLSb0zN7Ex/9A/KQwtphbGUJH+6AvdMb0qxDAI6vuXyIST+uknBY7JpI5zHuTn6s
lyt0qwuwJPMcLzmx2w8045rw6I4Pc4i8DVZECWPR4GsjsKiIAlOw7WHGBAM7YG+ftvRB2QT3jbUN
W1vLMt643z7rlysGu4LcFZ8vEYDUynPUIeFmsKWscortAhqQd3VEZC4JjYp67Tkd7x9eThOndsif
qtRdZj4gdeP9jWT/KeuPwCMM92RuGx6BL5FZXRfYJqOg2kd4V8N4NmqYZfuRL+tjQJsWV4GN3qMh
KGT8ulSmmyRwOAos8Rn9UekFgimfsYFgYe+NMu5zAMgVSC0R4Ct/lWDI2ONZ85X3IPu/5eZ7RMTb
fbLkELy/6nOx9e2OrD3BrCcfHYG5bpKhAKYeUVFHnz3DG+uCIsaVPcbWz8AfsEcbrK3ZFF7oIYTx
Jyzfj0gbmFXLlDHmhd1sKl9RTK5rebfS5fbowQMyC1nQjJeh2tF8bz/6OwGVP450k2lELv7+DCOg
YMRGnSuso4Outaa08aI9p0pOC34fL83JZSsnG+KnbWHxB716nhiASywm30Gn6k8BnfOqOfvXSjro
Ly+fSLu4VZPpMhJrQCjXodQPoXTcWXgG4olL1Mu1nNUnI91VYcApFOoFNRKLb65Mt5Pnj31sPhPW
kJrit9Li+n5d3WCa2hTmjIlTWVRKKy4d9ytiGczclqT7XhgRZIlT+ktbaQpVoBX3w9h8YwVgG0vK
6Fv3e2p1WRyqBtB85XIqGFIFUdZQjxj9be6IxxjXZTPb0Lij5/k55JCKEJiZWIL8hkZAJVv4ADpk
0Rx0B7edWoqs9Ic5zC9iNcGFwXwuRw/tq8aOAR7veMndFy1mAf4BK2TJ5Z6WV8YORxcIen0qnNvw
WRiWj8g2BcbjuzmsQLCRis92+qUS8siZy/in74KfMG9eIoi5cF5fHypHjqxm+MaXXOi5CzufAe+0
zjgzmQDZp2OF5+rzJ31eeMoLsfQCTEhl3EzKia0urhaQPkJvA/m96h1pkaiQ4TsLva2814qzaTkC
NOyZZ3CwVB76VPo7CpDJE7OIk6Tz9zUyd7+75iDryF10zs+J4nevq7TvGhUOlA7n3wBeESMoSIvj
PeQ7kb/eltuwJglpsFj8TaOMIUjbFcadnhkqAsk286mvvFwAE0ZkvoGMaDI4wRKFefptOMugC/aR
u4AsX1kH263+RviZ51DwUByj+1Kf7ulO62lwf3umxK7R4luyG+At2DRY803pN3VHX8n7mo1cfPIC
7Lw7+Iig/fUjI9KuewsNXZkijYXJIchCBdLYTdyE3W3gFfH9BcdzG2R2bLlVo8RTfNmG9HShk3A2
ewKzJ8EU7JDL14b+IRDAvo2uJ3OBIdaNG2DcLfHtN2lqPwsRcH8AjGGxia9kAMHatgDBcx+HbJqf
3Tq6VYyme/LbLCRbpNU0j14aOH1fLdq0+Vhw+CREF97pWT7wrD6p9yXvKo7XAwwl3oeTvR1OadiR
VrIIowxCIzA5sQQS3zp87MdcPOQtJ2Rto3np5QIg07+Ayd4dbCv3DaMj5oqc2RamSy9gkhHwGUV3
OMk29ryjqQy7c4vIbirtPzNJc8WTA3WY7tVs484L4PuogQAgaQIhRGn/ZOTHFHIV56e5qXXgbZGp
o9yun/ODwc6P6Cbo2jrCPcrX8TLg49meUX8j8DEHzES2eMh7bT+p9TcxxOJlx3tTMjKSv4ElzGOA
sbuCDED5YFofTOayLbPXtKOaJRVF4M/5cdMN0xIq8VTyNue7EQzeWQNZ4y9yWYaDy2dYWZLXKcg/
jfSYkcnN5shxbRc55o346rlO0Iv2ZW7cZ18dhDsbMDsQjEvzKnSbm5g10goEwXVAAwJ90KOzr3JC
fxA2uZqMXCRz7shJoXrslBTMiFG57xmDExLo5VnULznTPqb9DIvIkTgn683w+WM0c4NZ8Nzn6TqX
7pPtnjJQJ75Jn7HgkeqTeiVLRZv2HI37GBew3/tl4z0ICoxx41L2V2z7sGykQSnEh5rcyPfHKIQA
cfzxCf1Rtbw98muZM9m1dF2qYpndlsiZRt1Tf84aPrKB9MNrD8dYvVX8uOPlIpvX5XUnoHcDBi4p
NWRLbmoXZhxWluq00AsNxLdGo64OgDbDbkaVAsGf9jgT0k0U69gaVkEv8bhK/rlncPD+84BU0n9O
2ObK/QrJEkh884IOfLcSCmiQu5CiP8auVCBRpwJ1YcKUtAzGr0ObaGU3T+awOVi2JLSkXZS0XK3V
RarslGhuRU8IwiMDJ9znOn7IxcKP1I7X629Ew4ZL5YRgWESMkVuTBUW3yyHxk54e3UbFgX6+RICv
ZoZgiDKm+KPEKgri9ItSfaAHqXiNnGqVWa7rYdz4YeDtwU+YKUvTlvu7TjzY9saSE3lOupze3iDW
gjXGJ2MJ/ue++fknt0AYrKFwDTiRDRqsf8s7XltKCFtOhh8YqF/FJ91/PzSbFvuDZwey54Kpgi9W
S8bmtxaKsyiYQ3sE64dfZORoox7MKDH4cy/UwS9ULPZV8wwilogGQbBgET2jVZ1X0Fq+3PgihIwQ
UTsPFJeMCpIONuJZA3yXtbYrxG52xZb9hX9Ma252omIc9iTdNTgs+gKfGwT1xH7ZZL04spxLtThr
L1WqhmnTrptHtvZqtYKsHkVxeiVKSiWKEAeGcbmGQn6v46iHCUIsTyDDcaKGXOrpHOc0quSch2uF
4IE2ztiY5kJZXDPcB/8jDrU7ASJMGL881bc5Mdqsvb5GfYDFcwFohgPmaj0wCkGoi+66KyVvvhZV
gC3hmfsr5CeuU2YGvzSSMg5SEP9oPU/2mqOdBkyrvoFFQibe++slVSN/L0cw56f8KlJ2Kn8C2Q6j
X+G+TF4x/ta0LEYl/ZSAxlNerhTYi7aubr7Uyg2wBgvrKzyHlKXsZzb+agMVuH1vQvZWcuCIPf16
lbrwfvitOinTBaKYqjCbugW7uo1FNaizpFd437H1gNkjiQlHCl17aPO2PlnVCQI/hCKlgN/vvZvP
lE1/4fw74UckFSyUsc/+/qUfCDOT1LCyLg6QpR3+312xxhQLPP5xrbXV0/R+0oOFXOTeEle2FeMw
2IbrsdQuunG+0TxW9ntduu7Gyhuhi4agRli4QHJsmESREm6sT0X+GHfr6eeAOpDMJ8BwX1LuoPJV
G0Zl6hdj6pzf/D6wo6ClGqXEb9Jx6GcSJphEKM4gQFhiBzcVTzE1FAcCa+kGOvSqfXstiiLcxSjr
Y70IyuJC0EwjakOL1quTGGhfzcC2n/jbQ26D8x6pL8zkCQOvU7AwOmXD+R1DhCWu9vdbjiET+rtH
Xn88J+RH/k/N26dWzpAyvDvY4Mmx8gpkEJP3tW9McRGEDIVx2OoGcrGdRkx/lkKE2SLE2bXoBo+N
rrrgRmC9G+z+Duo1hazqSq8uHOLX2xgcnvqeWNVWuYMcfUN0uvtbYx+c09ky20fM2Qcr9rlAIsH1
tJKUZz9EPxO0vtboF+1DTe1dSQO+a1sJtDf8DC28zjHoCqI2kUVAqkmHVjJUaEzc/XZc8ikvGH7i
792+zTg+KJFLkLgIDlS3h7DE9HpUWdsrOh5Pwaimk7/hlILQeSUWrJ3MHQ8zKwltkj3+rc00o6fi
PafNhKd/F/Lm2CGLPvpqSuSMOLczCk1PtKN3tgAP+J9GSIgcv0IQ/PuNLaiXIv1GgvZEUzPBnH7C
4cvRZWPoLWIcSppvAJPOum6v0uv2si44VgzJk0wvPyVw0qyBz9DhgkdWxGJZZlVxLL4npmUKZSmZ
JrdHlhqIMr3ivh/sCHmgVfONNpbEhLfRN5alggoEEfHz1lv1TguXarqIduqLL0F16maMPE/QAvad
ArxYYnHm/7HQvZZfoRIWvIEgI/6M6ojndcZQNZj6CeYvVty9O+hOYSaqNhzJJ6snOr3BXM/Vv7zn
9b3gVLam3mYNmPCmw76Rlcq1Pxmpa1dfw2NdFu+CgTzkCNl3x9CNt8RUj/VCctHlYD7VEAvAIuf/
7tkj88hLqNjMdR973E3nVftABEkROA8taPRrf+ZRFmE8pVuc6smDbxgp2gjr8c8bQ/07oG9eSNkd
YF1GzeMfDvcaTay8o1h9LvOlvSyOkD3tVt+p4FztZGiyzb1TtMr02FaJ+KIvm5IaQbHk5dbQksnq
Dflx2U5Vu2F/Ig4tTZwiX1hHYndTma+7wPyNqaPVl1PdEjhLSImaQoM55EFFxd1WbHdgyH7Rz1yR
3XBevJjQkxj4Wp8wXCjN9/46gMbzj6i7TgUnpTQkYm0RhEXAcSykJcBznS+syFydlk4EfV8jOkDl
tgOLOEyi60mOtksXAsVkHzQy9r2j8939tLCaRpl4Z6r5bp73dxBuvMwWpkciLTKftcWicd3AWx/X
d2CEUsQtfbBkF0Afwx5f8cqzaZ6w6f3mlkVxDhwxwlSO+h/6jFWWUnnHsuHpXmeQ5iw/7u/65vpm
Q1SYH23pMy0ArwfidlCjHBijakDC5JS91/XzV+pQrtPhX9Kr+rum4UVDc3MMueao9Vjdk9PF24tY
k5Dc+ZPDb6ag9iCV+eEix41G/7jnwVaCnB7ZVZiKJJaos5sgMZlllECnzBeNxyQ38eKrypsHBKXJ
sg/Zkm/AYjW3182ny16ZcBixsu3AbH1aGNtyyERuco3Z/Bt8CLR71o6LxKnplUaCQZryX3SKQExB
TxnqhM6uhxdIm9V2ehiP8MX4g9wuce5MidVzdZyYUlHrHly+kuQsCmQ3XLPYFyd2lumTojPhSupU
ty5FDH7WbPv0Yu0n/E2+D8LcJ5yob7UAJD96+gOg2AdC9AWGg++dAhEivWuU7nqv2tY3dyk2RrkT
0FQmwPBl/8vBnrS87KYL/vW80l9ozqVX7f/OY91H8EdHDMgu/nqBDRzJWxWCugGTuBxB09M5cUC8
Q9897Wb+gCkrlbOl/nF1oWF8osp5N9zmQx9DJXJqiDqJkelyNLqJIWhlzY81bA9Psj0qg0OG6lbQ
e0scXAwd0B74JNi6HqocEkaq8nSD3E3pfWUfPWTC593Fk8j/YhhZpgQ3K+7Img9tOixTyNsyK9Nn
sDjcZCgKceFX0v4LrIe+Ein8MjIcEW3ldKEmycmbslwAQs0ZIb/yCHNXqos3+RDJM5QWDSB35dPM
IzkmVM6EV+R/VcwiyepX1JjjW42Q9lvyo7xhzNXE7zGIWF0oYwJ8EbkN32k6hvg3t3ytdEQTF5+v
0EL+a9vEsFGt2Rw8fL3asSeOC9Un+wzMymIqMCeK2nhqSPVXkowldhw5loZf5la+MOZRJmiNe7xT
CkFzpVP7NfzV4uoyhtJs5mel38cXZzwlW0dCDJquGxWku79DUZmSMSRFZF/xiULu7kGKyzTL0a3o
SpXMfiia/Gqn8zRbqCyfkJF7/2f8xBOkdjnqv4Yy3JwVqn1RkssjNcYSrcJ/ywpK4dIaYQ92+gWg
A/3G4OtgnMkZqpdoSOW5BC5vupOxvsPQjHXlSYlFeIOV2peQHSDjLf8LVCaeiuWV1t4kWQUfjVEX
sWatvkpFnrSvdzkyp1BF+DcmTrFEZeUE8ib3GfR2Iv3NazgohyeQUFPxie97GLcWh9zsPiLvUwJg
vSBY7XyzfDsWR6tDvt4yGhzfpG6iqBgKHInnsm5vYJVPawKQIrW+jAvNkbyaYICDODwDEG89nDsb
rLJDFDuMnAo0EMX1yOP0MrOFwPn/ckYAJvdfX4gYFi0d+wW2wYHHnQNimeTJ7fQQXtaDtz7tElxV
7Hu1XJtn3l5V8gR/hNvcQrZFUeFL48JJfU+v10123zH1s3t7kYXSOidw47EFgkOH07jJoIe+gGEt
6wrDV6GeGSY2nu0JXjuqZxsOq2Oy/IitX8hYS5IIEivKREhL0Zk7NnM1aRIh0cZOz+3icg43uk+J
iyOgR1TNglxSmYb7vCm9pMKXvFhDsRyVNwHoD9qc+eL0+O9FZ6Ko9C79iLW4belkPqFcKfiUgkPt
RXutLxlh1m7iuH6/BPcHUADCssp9mwogGKv7HjDE6yTnNuJGzlm5QjH4Z2hj/mjk0YYdYFViw38o
oNytnS+bRN2io33YUS6CiH1g/bSDvnbXrQX3R23NU9q36i9wcGrHG1e9t93+tuIjQbgd7FcBl/nM
Y/Kex/quAFmcPlBUji+atu+GR8blXxkp0mQwQs2fjuqo4nTmGc5caJjhHalg+AZN1LqP51cCChIm
CfX8QN52Vo5NscCOkKa9BDlyGou4t66McsPebEbdSqBwlemBATPiA92ttCp0lg4MA7ZZHhg9hxIJ
iDwDHLGHOAG9sSngNbxeEf0XKuuf82Q2g4gPe8xJJMHgGhQNf/6M6pInW4IgDMoIJKZlZxGKpFn1
LqS45W+d+oAxdz5NQd0TWRsWxsfw4SEKeeyRkJrbdanDfa8ZzU6f8riAxAMKLepdKXOhJGRKyjEl
Fmpt0lZoKG1rM0TKegvBt9afEwzBLI0FtDeuZySmJ1U4MsHQcj+S2xUKRMlsTqpfWfyW2iIyFj+r
GmMy+rDicxfo3+FSOv52S+kITbJbUc7V+a1XWOgXK+m90tr8eiBGhBDTsMvZht0wgUMYyFDN30Wk
iM2pMU7ZuXEy3sbcGtGvG+2LneQJCEeqZN9HXDsSEsqncsKJpsBKziwxn4uRdhETvRO+h+NZypLq
pcnECXP4gkBO7q4CkAJvB4a0xyPPJw8dOhHVnLmXVkvS8BSeJg9OoIrBDNFDsJGbWnRl0jvnmk/1
ntyCpo8cAULq7pHkSwBfm1q8NkIRi5ZfVrm3FmonPzViQW94hst7CpuSitonK4dfvYctxAgeDS2b
ysH8eY9qH2JMvNN+NnhLuIravKMsp2V9erxDAsgrHY0QIcL6Gb+T1PtT+jdHn+KWkx/PG7Lpc/jf
Txj4tbU9aQgVWf/M/gDZCb3fIEGo7xBSmwlw8f9y65/u0QnabpcluIAMVeUck7+P5+eam9mK40fK
4xRh3FSujPfxdzO9jKFb4WxP5A2Z0f5BYttIT0o0ZF22amW431rD0AAh0OmPMSVt4tlb9ZUdEx7K
ICrYHT7/OU7D52JzmfHot3Y2wOjdtxB0ekhY49YJYoXeps9A6PGQTWB4Fmq1vbnQiPDWjRwcxp8M
FyPXlKDhnXPubyqE80mOXK2NLASneqfx7k7g8t3LBRD8U/sNbQz94QDQQ4em7QLXgM5tqv4HMzE5
8ggobQwkS77vmRCOiTjMwJQjdzsA7bOc6Oz6cTzGXvJVU7DJyYSkDvM0Br8FMc7e9pveCJUDdW0E
GbNpMjfMl836mJkdUEHCIgceC3nXTdLEOYDYBgzIhRPq/YhBrtFELW7o5wWbSLsArRlBgSkuRdfi
1t6RHhdmds9A+zNoCR/4M7IdycHuHhjTwdfioyj8HduNe0lwQj6EOxy/mnjrEvVBftVupa3KDyno
627dwd3RjdZsgqdZZ/gNKu9oTRysZAEXQEP8/zMHltIf9wLUm6vn2ztXbqmt1Y6Qv8RWD4JatkgY
wej64DWMAZQRalba7C8KEIBbVXaF/80NSHlKzeS2WFx0XOhdHhbnGKqu3Pv1582P4VqRCizjooch
0Mr6VaUXnSwo5BA4aXi9fHrHqWTa5fmn1kIO0gQs3VR0VhVi9chOOaGXzBU2hYqeskTl3AYS7NoY
wy3qw7HYjkjy+3L1wf8jbZJc4WymhYAauaUtMk2Y8ds4SsBfuCFq0yR9bU4xxXi4LPpHDFd11If/
tqzaenU0SqGS3WM5QJ16+84kw6CROur1JR9bSlKrECMTAXCgMGJ93vAiJaDJ/gubwL7EnJK0j5xX
CrIxrW8ijNC/iPUy3FKttStaBjiJ1EvccL8klR19c4g2os4RToUJLCJ11hkcPEfgNSOR5h/SqsPF
Gx2Gk2IXflvbpviFXp8i0bV2OPROXz5kG1ND2ieAp87yHOgJa5SsnoZgrqRWFRr2Uv7porjyIbU0
RtiOLmnuuPs0O99ReXxrS7hiNzAeUjckcJg6PEDZoY9Xal7it/yzorSvQkDGyNuP6LCvTgx/nCeP
Z6A2LF//E55VQgb3Y8qWgC6qweRgz7z+haLYug/lXXYq89Clfg7AOjLYhYoc/v1AOV1sO5bMmuun
yG6ho6lFbCEo9zVOV2JPkGcXMTEEchhEIoEONhKzvFWqgAV5YpgIponu6qYdAmvXKVR2L+MAsDXr
ttDYnC3i978sSUKeYZ7hm58k8ylq+RaFz7ExK6y5lOmF6DwyHW/FemXxQHtRFc7swt7KjVqp90PP
WGMcYvRzkrk9pbZoZtAsQvWDda3UskaRyC+BtewKVfJ4U5yLb7OpInGBjdy1UUCOp356+LlM9BSA
8zdsNbdL+uG71yFMWVqA3mtJBzz/l12bcS0+jr6RYpVWzo0MDGdWsojFYldyuUYB358xac5N6GQj
zK2ebaN2HT8hzLuIzP8JtH/pMMac/P/7aAoEcJhGEAoVFSdby8H9FMXefG30/63QekM5wkPSRIf5
MDhmCaRzfw0+jGrhlIUFFROukYMIQyY8RGciSpjcbgkSYmhEbd+LQfpzyMJgc6PuGEZgAkF4ZNuh
IuDHfdXQnaKk0m5YQbxVSQfBWWwvDN9kdLKAneOuXhvnKDgdYp9yTJJwFc7xam79OelEKc4DibMb
ZazqKPRjPPJ6IBp8kid1JwqUvEglG06b9oqC3KRLDguytMHvzfVXMSJpYq/s+fgq6BAgTN4pAs9K
tZ6kEfqsppHoP5VD3Y/X43EPc3f6VLfQ/RHLOjG2APGbXVxt3IcxsspGa1YCv+W7rfIyN6GxNUOL
jqJDOZHNHP17HkQ69JacqpoEVX4LN/duHHe1OjKBpEyGemDxEBQAR3rHiGk/OaA3AY9oIhzsZ+Ob
uKzGRF0FGY++ob18Pk2XmFOLVWzYR3CJ/lhYvdj63bFWBZAhwHmm8/nImlPJiVvu68wZbDQRHGlr
BmdJRcKr7JCcMzTgEuU9SNK16LEo3KgsFqPIOjlX2kjb4p3S5Nkc7Bu4fD5J2zB3/CaFe3Wy7DtD
xMH48TNJ8EMlCUADFrZtyk0TqGSvzquIK5SyUA8p0f70o7zEXjxnCnN4g4rJ8rfGeXccSTYh9w8P
7yzDSBAV2/wGh/JEKwjBquasbIBGge4BuH27rZbfApI7Kz8c4APj7VC8ZyBDGsTG1Yi4n9/3SS6t
aFmjt+lQao5vbmYLQddCuwBBXH2f0LjBeV0IEmT/q/B2AWh9ezWd8VURBWbJ/0Qcxw5n/sbQb1+V
mlIOobs0pFhfdT6fQaVnyRnqcw3vWksf55MF8fYQfTiQb8k+wLTp2GuSVcfvjEa2KXIC1Xzi5ud1
2KhRQDrLCout9UyVNBWwCNnP63Zn0ceM20KEM823si7PRQ9j3GkWyC/hQPNm9nwiPw5usuiV72HK
OTAzR4i3XmUkHXh0uUce6N15MM9yNehvElgto1vPrAz5iWcYuOs9GGzy+FP66eE4p/R3UbFq4cYb
F7Sm1G3MwNNV1OAMa3cRbr3vC87Sl57nmpSO9woMI0Ia5e4uXbJkalmZHiqM1Pz3b+0EhpehPlgl
5S9tDjKPaOmy0RsAkeBZtV4UZbNm8blR/rOXpF5b52jsnFRb7ItZESXlMup6TDppg0jYXTNZPOQw
HsF1JUFsdpSXZ1l4sf6jsK0plxW6y7ojVdlJJs1h1dPuiSeh6vi3Mr73Htu3C7rm+dAk3X3oCL1k
nlAjTDrMB4R5DgEX0N/tOGTC97DVDKqVM2S6zeNY3NF/v/LCvzj91NpQTXHNjPewO8HDGp8AUoQA
40WOBYn+fA3DEPTjfWikBaCv/gmv5IM+7N7Za4sVLAOo/3gdnad78A9ibYmatnkHqS5/4UjVFah1
Pt4bxUiB7Mcx8zkARXD587tDEbwPZZMFVJzKSDi6vX+T+1Etm1DABMiWsgp7sX+9ueB6Lh2EJriy
+eAuO8P5Ic7QPiEF5fno6GhFkrXZRtBKwFmPlWsfSogoNTzOVfZXKyGJowNqm7PuAbiL/DSTIBXE
v/v5KzFucq5OlcSDa/ABl1Mh2vZ2bM3grYRfmG2iOFTgWuMgY9oUsb84V5+i7ZV24clMyMf/S8Br
nCSv3VkMuUdzY2KL4AeDjeMoJUpE/jFwQmiIoyK/rd5U6u5Okitm4FYTvYdLxPZ4Bg4ljrXPHX5P
jiFttf1E4Y1hhKm7fM9W3LdP1i7TVOXSr0S+ViU7/UQylQpH3VZJRV+TRsmg6hdQflXaxF2PutO/
WtzkJMJhDODyfgR8vafjzdUtaJGBKIVs584S4h2AnfgWytW8qDfX9TT4+IIdVosDePTwLfBu58Ta
mUflnTG9yGh9i7YWHV5VD++VPVpn2s+/lMq3WrCLDwz/0JbYccshN1R6dNrtSV07zZjIQg9jEOkM
os3cuA+Qz5QmaYEE1PoDZSIYvBT6ChflKns+q7upuXCdPC4BDx9f0Mcc93PamUX8hWm1PO1er63w
dmfX0LAceX7/SXWXzwQexUaMrYazSaGJKssrlWSOqh5P/QzClSNemRvgrkG/CEvIUuTGfG9vLjiP
FDqkOwVUs3cEYe35oemxiRqBZAm+v6FtQsfuZQ4JCSqlf8oIm7fATvGbX7ZiiKJNPfeLTp9cQtGc
B42KUkvrPM94RoF+ba3QoTc3RyiRUfaAtshgSIsuF6E0qHWGWG+8d9k5Tb7ScumsNG2i6Ri42QXt
GZ3HSoyyrIRSUBAzB4t/qkJpflaUXEXQtm95QMPamzvD+vFWZXVu2dwgwWQGLxSgVt8MxIzuOdtZ
pV/rC22DE1XNBCVmZTEFieNB81EVhOCZ789s+kSy/gdXESmD2mJ9rdyCpItFcZkBoo7EkuagWwm2
7nYFTHwldPwpDzpsDdOnXoMPYmsAH72Vm4wOjxjm3zzbxxvCAOPSkdoCW2BmAXFhWRZ2CS6GDeGF
9UrWtdWkD1oFGN31SuENzIE1/6GzcdrvHrf6XEAMuaINPn9uAol3kdhHt4sfaznVorlzAlQpFQYr
0p7m3Bsx5lIYeJJbmXemG0NO25WZmnDPYGax1Fqv8gvXCeAkj4TcohGW4gFYZMoV2fOa+ldJPyZC
PnzSwcEijVYhBtloyy6YOm8/WBWrsBZmVmXabbnWEyNixkUF+DtT1s8KrHK+paotZPCndfIhQPU7
o89ZCIUVo5jL4x/ROp4TGymdqYbSYgt3a7vLt5t9FAoEDBkd2Gp+92ntrcj1REbb2CpD7lliHssK
SbZnRHftlqIllhxp0v2o6a1ikkPyIypXJHuAI05FEm/nJOM/v3T0ZV0FXuCO0eJ9pQ5tYtPzpRZY
Z7K6Px327C09vrqHnVsk2esqPk7uxImn+GOMWz9azFSFCIhw5WFyx5S+oyGblLN+JuTH7wGsrcVC
YG5gswKDCObO0fZ9XgCudU77iTJ7kpbNnrvHRsGj6cpwJQajlxmn7lBUN6CbbuDxpEoouJ5A+Z62
Rl1pE3n99mYMISYca4IJqv/a0wtMF860ilnrBtKtYMtCKqMusIH0b/XmiLTrTvcsIx9Fv+eSjNzf
31rgB7NFG+oGxcMrf506JtjUJajPfwuQaq2vwgEnxYkoynIExUV3YbfGLk8wyN3Z2Nv0B3fBhWT0
LVcnviiQprrcaWN8gpHI3MfEspI2jJud2RDO9I2W8r7zd5LH/EvO/Db5ylgdEPB+dJVTNgfUVgKr
oodeAbtT3OH8CF5QQoIKOKiRoEfGYj/mY1Jc381MDy95kI8O8xY0ZlKDkuCQ0VX2pwW8Jk7HoykC
zRUg0PNTxocCfLDOPo1/S0BnTefqVpp0DW8QZ3g+69k5/nedC1nr4Po6ltkBxybdB3xJA9eELBB8
LhAQXRmYd9wfPtduru8bw1rCtt0KNhawhIC4Mrc/0h4dwz6L2YN0b7Gj1jPsR6FNwr+XRn3rarrL
WNkUAfdGKhblJDIQ6LiWjj8g4UcKvcU+tH8rC8F1xzKZ46818mcPWjVbbIHxYj7H8S8i+z2lkyQt
fMHDi3sQEsn/J56obpkSI9oCgm+XGw/37UL+xF91kxmp4VWH4Q/KuiMsYYVIfIffTPmC+IK5y0L+
lmAvNT54NC5FYP1vwrwoFFW6WazJIpZztActkHwqC6mP0xBx1AIzj7bCXoX8wYvYdIv1EZGeW4Do
TMuZ4V3yYGpfIDhXLwmcubn9K/a/9o9IJ6wHE0kqWppva+ANg65bTTLlGZ0HVxdRcs9n3Pqlc38d
388UwQX/PI1HJp95ClSBMnrwUFpIOnsEWXogOCsjwoLI52EfdEwg47dRWb+9rKFQAh0uZn6sRlv+
9DGDzDfU0RgfK5AKQrssxL1BpDYRQUp2yMTvbwoBhXjr01Z4F3FecxPKDk7GCwl4uAPb+ApejjT8
XSdWd1FoQYXZQgZ0z/3DPUse7OJCufhAxlekmm9A0p82kKz+bYFKL3Q8wEiQE3pImnNQbbVtK1wF
86gQmO7Y9YgLwdLrP8beUgq7ibGwo8Dug/avfPJm92hKAjUVDFMKh0Vs2JHMyWplQ4vKeIsHzvYp
jh6XzDil8G0XNp7J+8pXYnclklqKUh+8K73yaCwwJ69oExlxVWECEa236aR3nmJ8rkNkNbBYWfkX
8A0vFTp95sERpOD7Ly8BDnS/AveR+B7W3UYufvdKZ2EiucreLylKF3MZCp37c2GH5pauDyq0wBLY
9AViWHwJup3FCH6kYTq5M1nEgpaIzPZkmLSA+cfvKYoaxK4VM8zD9ZqzW2xhCxp6YhaM/rUlgpc+
QMXYgWkUUXrQcu5JVSx2C1idiAxxqOkhEdn/Q2YZqMYilCTTdfOZ0Oa8blSegeCipZy+ZX+0GD5i
zm+BO9JuRrCX2igPXdOG1wrtgztydC1Um1pKlQIGx9sH5xpEdDfmLC9+8j4r9bkQserp6iu2afP/
dzET8maJoisIiOIPo2seagAFLCSwUytOEKvZSsMoHJINxTnQeXhgpcDXt5wgKtws3+MYCeRKwcZe
5LvMD9aIe52iVPiG6FodeJH9Y7tktdqZDinCzIQO5inQrSPgK9RdrF84i4jJo6WS/hk+y7gFFX7B
cOywk9R3iDQpRFs7OHNDlDstIU4ptRg7mM9nXmBCnXqVcbX6mGS0gfOkoe1/uka0/Y4SumEy8eRi
yszWV/2rHlIRiloR7bdEIqLEf80CnJ5z5hvgqyXr7NkGkLUFXNsOymxbUBQgDWP5CG+6y7c+KNB2
GavJKaaaF+bMEw2bHf5homtoc1houhzaq506vYLiyOloU9A96zcM8uBly4GyY8gq3Y8VP9l7f9+J
VlYeQkFR7lfn8xV1EhEuf2/N+NBhxkEPOFK4hZrVzSRHHaPikC/HeqayEp1NqK2GRdDQWPdEulR/
eh+qg1ArgzMtCK46hznQLHF9Viesb8LEX+iOd3SAnlImIwjHvoUDp5lphGmIVJKQaHb51Oa1dwcq
E9J7mLqikRwB4rdwxZhc3AVcR5ow59pTp0SXeS4yD6Mg3rywMqFwODQugAqFwZEFzINStN7JrMtC
EnyCR92Rk4PP+zor9ybfrovlA+6e4rLax8lWBLD3bM25oTjtemvTHRu4SHR1jsXfeqilPoighc0F
Co7ZWPNmL6zJaDfekBNpq9kDP5ofW2SW5kmPEB2WIaLPPHcwbeRFVp29YKfBY5FP8gVdDBGUnDED
3leDiePRDpKJFpa/jOdx+KBsbm+vP2R5H1IoNRUy45m6Mfbaw4L5/KdeelF/PK8JmkvoLt+KV58X
Z++RhkFKzgvDuCgmN8phfM61iwdLYndYkttBqFawJjxZ6GLlG5CfQS0Svm9P/s+acnVeKXtl60d3
9pfkM48umb5SOS0fYzIT3/S8jHDKwy2/MGo8932ezi6GrR4N3fZYGJSq/6xdp9Pjw4+BpdlhW4m+
b/ycNH0AUGuvk2lN5Lf2/7jzq3qiojdiitbqP8/Qh4lxPWEeL7tFM6CXxqV3wOso9cGScuet6R1h
HicVi338YLFuJWs9pLRDi3tdFPKgZ87plijFykC9KLL+lhMWX6ObSkduCpCImeDu+oj+JjqogMHA
1HVFgkUkn1lwfF/H3sRnM/awDgGonv0O/afJOl9EaZTcSo9DH+0uZsl3Yga28rsvE4l/L4dgIm/m
9twxb73eTrgRRYXB3kQ7c0UrZSf6jboT2+pOTKaqPn7raKqSnrD9YvapLfDbuqFY8h0cnmxEm7Yk
C8l7XAFJzYLELy9zCGE1pxsrIemgpoqI89iZhASBvjV5d3lP/N7OjWvPoC5Vq7SnzxKhr2L5eBOk
N94g2xRlSZ5Cjqi4mD/Cy/utHq5Cx+FqkXUqNJD4G3gBvL+SdXpHGXRgbiWP+ZZzWQ9PZPJ6PDxb
21khIaPfuo9d4cwrB/XneNU8cH993bHJIkiKTzlMBHzk/6WuNuLp2/Mi7w8kCmN2uldPJZdkZA4i
fVSzlALMVSrzjoFQWx4ZkepVmvQE+c0cOJTgJGNd2dmolXe/rw+Ja3wO/e+koi3Kg693tEBNbHxn
qoTVTs7GzW+/8JJqN2YI8WLA+snYVbsC+FKu9hA6g/HQj9EHnBwpHl6GvDUZdXIXzP7v8QPBBauI
JRsVKps4Ypx8DC3T/BIIdjJYW8DFLPdihvUCGFxgtOCLu9tQxUD1JJK+FFZc5ij/9EZeEIcuyVUG
x8z47m9OB/M+zG1xdcXaXEjy/G0W6z74HFifWJB/ig21m6gh3y25iG3yXhIq43KRKz9QMCAdfH9M
6glw1cxAYhoFaie7O4xYhA7CN5hS695BuWp+m+kQ7cx7FzIDv+qcm8Pzd4dkgeYK43Tvq7HrZAdq
0INZ6tXMT05FK2kgsJO1k/T7m2eoZzqHvI4Irr6Jb6lvvvtIqUk/c4xxzs595YaNwM+n4FjAsx+r
teTyg8XOUMd8j8HSQEo9NgPHm6RinRJguu8eMFD4CMFdk41NCfNWA2ZTGT9hA3W6iAf2O/nEs9EE
NaYepOjcqbfvYLY5BlNIy6blkAz7h+/pPRV9wKG7q/fNhusjBSdIJP3Z4+2E1B+wl00MfnoZt19K
yq4nZTWqm3ZLoqYbMIZDPGmbyofU9oCM3BpufV6gJfGJ6KCt+ucKt8qByPAP4R1FKpfE49N5vEf+
FpFBJr/kJ1eOaYrZP+XlWoWg6XTPLJze4RqOr7R5jGuW2NjvoFO6WxO9dCEZuKWrE6a2uFSHaCBz
uaQoTlDJKv39OLkgmAZoRosJlEe2dnsmm6feMDwlW+SeSeEAnUtX7r9xF9ifLLyZEAbkXdqXlxYW
xFuDKgkU8qWlCqqHeJVKbSP1U7QdYcMXBecMGZ7wLG9b5IWXWi3XZvnH3nZH5Timp9PJQbINYaKb
BBuFVyTWXFsuVenRI0ivviMVAeRWFInZ2fMgyVlX7booemeDIVFkE6lO6nDlRN2JjGmKnk4sNLM5
Q2dyFGuCfPHle1+H9y2n8JQcLTl2ArO2veJfc7jGFR+wUpwSNmsCNPeF8abGrRWypfx2gZ+lrs1V
ZVg7lZlDJFYQSwWK+07TsWpAzA7+rSy5tlOdAjwngUAT/5fSmRsN808XEC4rTXZkwcI5h0dcQfLq
wHcCMTefVqFJTwE+EsgFlfexiTT42SiyJWL7VzWrcrwDLewfQ/Tld7qc8Jnq1TT3CZGpq5zPsi4j
jTUEyLHXulTJyxMtu/T8khG4hZw2cDATTmowuwm5LtWwMjcc3zyUv+eC50qNZKUPvhZewq2aZGVP
SrvOamgFYHFVN83SyoSNIVhoQ2pbOTyjpftMeC2gWFMgUL7j0KsH9AyPZjBbTeulOokzquoOCZYm
ul0xuN47njjgwdkkHC7x10zpHICC5em0KTdi1FATP5Aw3FSyEHYEL+gBhF7QPJ7r3wmgyPq0aAjV
8CH1Tp1hEP5J08YcJbMFZODAECPj42igGXm6SAD2t8+CRxqdaFLN4ZVvUYOdlZYtMDuLW5STKmqS
3U+icy8qtTaYYx5XR5nNpomZuYDHmMH8JJijrrQEJcJGw/+Jnmb1vh1YcXEVQEaXO6fSmrV4c/jM
MJDzhr6tABImg1Fug8+0RsBQyqhnZmgol17jAndDocY4AesFQHMLG8pdBtdaXpzTqDnBgWRJQTL8
VauX5hbUy1wIeZQqIgJBOa6sQWGyRBM/9qJIiw6WP8qAQcBRaPzwrBA9nfrSH6rStBKDAfM/F3x8
aCxb/UY38tKPiZlS7RSkRPczHI8BguyAvVDrfbTcc43WCwsERKWHb9y99qbqCtGHQH7GRlex0Pvh
Abb5TA/zQ0JrZjJNeJ+kYgcJreuA7DR+8lbWpDEyofeG1nfbPowXxtzpmHhW4CL0EffirjclB26s
8TqpFJJcuS60z5xvmyjG8x4FzQ6LIxLMBTt352njo21q6S+13YmFlCw8x+wuwzDZJpZFsxztlJ/x
osnyyTKRkJ8NtajoBO6nn30Y66HXc3mWOCcocSujlzZDL6MZUfoa7Q2kyzk9x+RV/vtuXa6lzaGz
VrK4bWIWYuvHhcuJZe65snDYmr6XA7WG03z4hxa/zoZ7p7oc1qZRiaBIAultdkJbYkGCjNSWGyYl
gbjGlcSiyRMcHrDF7/00mLASBsQucbNSEsQMyH+8ryAGV6fKkYAgTYiZNRkrgPfmvacaMbdO6vq2
UbVMvDcyHpYN9909Wstp9uVsnz06YIIix5aZAu9Rm2urCtEVswNgFBwNHIWTDWKQs6vTYvieaZoy
/TU+wCr2tFI3u591ns1gjn+xncN2+kN3QThK2B7qaHAYCmFA64PvfTloUpJWjy68j1Wpobw0m56b
tTycW9GVnzHuTH85QhCYIiiTq/HXMm2jk5pckVZu5HG9iqtS8FItk92vSurtb+2P4yExaJUrCFK9
Tm5BE82k6V6nCtDCOGLyyz8L1JdTlfyYEwRR1Zt/rBv7KJtMFM6Oen1EreisIA9xOl8z9zFWBFL3
gohfMS2fsGNHbFopbNZTLg3XnjbgaYki6YX9TN8iLY3v0MhiLcAfQSyaVr+7hoh1oXvut3nCeHpY
mDCNJaVNojqEdnMRV+Kex710VrBHCoz8tFHsKOuiNPiyDXaqNcbD48OhGClSB8L+CdhthASedAlE
sDuOqYr3dAszPVKnudCcP4OfMai0YeDrkOPP6XmtRstZnejeDf/T25bLWZ8VAJXipcKJp+0+yrIi
I37/ksTIqH7h99UBPisgJVS7uBM17e3rtWV723HDQkCRlKUOVGYmHtNvfNc5bl1hE4e83l8cbk6p
jkiwzDT7QJQLyr1wAngaIj+9uqGeLyN41E0IaH/vFoNjSKnsFMtxE7rURORy2MkLK50xGuM0pcfv
DIeqeTS5QDhbGO27Xe7FMk1BWHkh6oLjKdmCMRWsl2SbG4UEDV1DYW1u1VW6UJxfwr13szyV27XQ
3/eN6RgHmCVaGFcW+GLLXlDcOKv/Yr9qRToc/JWYNCsPd/1+PHbuE15V4qdvtDkydqsW1nRe+JW/
7StAgVMpjWu3DKIDzupNbD6JumSFZIasShXYlQGk3VCAYlv5a/tZoKXvNLWUE1V3HHMwyhlXPSxA
MvN9m58eSRHrZoR45QTT0PXJklNyCVyfO8iSy9e6lKyEfbLtBAYS9x8uBqBDPHoOhmjAQTMvGSkp
akiPF5ZHFlBV6UmThYantZLFGqbNeJOWzCNk3xShAdeq7GcgQUyjggXjfOtxq+9Z2mOrHxKDJ46+
ME/62X9qOCf88ZIQ0Kb8ciEjH3VV8PxCnGN8GZ5rK30XslmQ133Ll2ytAdkMgKQ0oorWlD1FRFl1
QHRoZfFYdUbm142DrN/oQJok0jYbv2CgHVA3gHA8pYpPBmxKJk9/tumfunwn9by6M5lLyub5I+Uu
eREVOYibJp+sG2OLiTKs1bD4Z3HwkEOo+MrRoR0VbIkoH1IVsVspWx5Krv0AUnCsmLrZOzPKVl7a
+w4DbJEf3hfR88XuLYPIKjJr5VyPdRoesfbYufqXFVRWzW944uZUQw3ySE95GP6h9NCMltXaSvhx
6jAbW7SgFoAOj5Kp4nKpaVnC1Czb5QTQfxqPasT7lFDKdGSRCiuRLuAD/CZel01a02T1Pp9+7VnI
SdLx0n1IxePcVuTutplkgY3eMd5Tipa6DYwJIftY1G2nlvd7Julue4zyjZkzGWVowiWoMPZCe6bq
oLWQ2sbXwQADryOXNSr1zwTXzHclbpcBmAsAQLZL7LWOf2FvOboIm4iA9PtS19pMIyIbrkaQ0m7Z
Qd23HFij4Dxlpcv/u+BMf1bNyvUOuNDGrLA7yHEmfah9/aYCKO77MeIYMDnW4U+9xXO3C6Qd+qnX
1Ybux2VUFouf748vDiwrDk2OJixYsnl5+SnXmelwYWf7twkmA9ccij2sXPnr+ZNGatqUc/RtouOe
cugF/b/npFEUzayzsCdZySghmEiS/KvMsoptuLiS1yOvTnD33REApWRbDMNTFAHpt4Xe1oOdQK4b
QdTUuE+qNAvjV44N5B88EudbY8g9MaVxcF3J/DAJasJXc3hwT7Dc87FEAAZwd2rQ68JPSC7gWxID
vTr4YwluLQjgNA1vRdR7ZVijdKf/qQ2L5LOlIF6Q7D1wx0HX1hq1jjFxEKDBvU/umoPWO0b80kwo
UCe8Zu9pRHYJan8ZcSUyzXYDr907vaTyBvAIMkvGehBPxupP1xJtwsJVMHvD6vADeXtlsJbBFNTz
+XohQtUWRRmTUKBP8RO+wtqc0Onvs8hlMuEmR1DIxQWqLkrpK+HEtCJqks1h04xI18VRCPqvV6Fm
4PqYU43XRGyi31UOhwUfw3b4ZQpiDaxVJ+wAm9FVVIoLDykSQ2n9Vo2i/jST+84bsU8x8JCOUJrf
LctsFr0vJEleikn6eCG4m32piJJeycJ7r5NhGtqWiP/Mgd/oU4jUjbfqWifw3PBZSaN3t83SP1yq
NJUdafIisw8Z8U0lOhYe/BXbcl+tipHfb0Jrce/s0XVxHSPUYxtQKLLS8NxAAvq5YArW5XczVvCW
RpoPFnZdqSsCg5750SmODHdvxQvk/DyJnoxduq7QM4I4ZDrvn9nAi6ohtfwTUVUxHFm30OPcSsfv
4lEonBLjtbs47HIxoRRj70FicqrEVTJxFss++nf3edVVSd7M7AoUT70w6wewDQQaRUlBRScSTY9P
rquXpbQr3j1pKJPBbuiDyYba70OhVTe9wi+uDn6Rje/5S94stdQUqyree/y3NheFbs11ZoxnUYBk
gFOr6g1CkUQgR1HqiyMVl0DP8Kk4n1fOD1UdmT5Lr8+/5D6F7uyuhWYz5+hNekb06lFF3H2bQ+Vh
4BHh+Zawc2o3FK/dTxfSdlaqBOlX+cTT3h6oIYad2qb/UE74k88+FbO9XzkYoPPO4IA23lCL6i03
wKUHK8kg5ufp/RcoBukiioPCJyeo5clGtUEH+RB/PMoiRNTAuIcK6pBBmDJPbUdXf7a0WPaHZnHM
Va5cGwXQ9UimG+t2P+rjW5nRAAaokJQmkXQ30uEvat1ulRSWP0VKy0yy7CJyy57Eic3Z1dV3ybRR
4nqtvKOtTjWsYLV4gFMD3eEyOD+/ET6MJUMcgs3ehKENjFVuHKt/25etNhiJOqaCntmCMYYGPuWr
fMX6AV54KH2FZZe82Z1VmUopffFFAC/zL5VL/qfE5corixCVC6qiLmoITn9a+e8vUoXrNisTGCw2
eaiUz1Cb93NM3kJOowBEe+SyqmmwNRB46RvMFKr+9sjzgKFOjSngAW3SzuTxAMzUoJDCuU5l9wHk
gRG5qn23R3xu6O1ZdWvT3WslgHUdAX1UMnW2nZKPdl03/l62+QF1oYKkY1YQrjA72VxB+LCD9TiA
jyiqlvq8cVOFv8qWHNv7cJHibII7NlFprkFpOFziQ+H15BKuNqWwz4vZEvSsqGIiEySKRchwzzni
1JvwnxFvayParhtGsK1VoMaaG0dsVN/TB2n+kOoDrl3ILCZcAsonIDuWr7tf5w2OCDKK5d7/Lgw9
5Mr1Dv+XZ6hOMuD7F51ABlEQ5vMYqKy2zf/OFpbfbk4JOdJN0jzeqHh1AV56sXsD0SQ4yA1Parss
ZrVORuPN6ikmjiLAh05W6z83rKBxPQ41K0oXS57TtNqy9giwal9p4GgCrm3FuJk+h7U4nsEW5Wko
lVWlkaokBFLwbfHNP31Ym4jhu5lw44zMEQDJgdTPVIwAzLnt4UnuNCB9Ej0joXu77v/1xy6KjkGN
gkqlAeORwwPF33evAeRGxH8e/8aYaKHJ7xVZDTSeUjhD70BPyNV49MZMo/dT0OtvD18uyU8s98tA
mLG4BhOWV+BG7VdAluYt+4i2n7zYVBZx6ek9CNAaMyVbQ6F/4AWPDlkm8+voY9sXDFzAJBCsuEqL
Xo/eC4EMnyt++Kv0CAOA6SJcG2tlXGiC6+N+8PmKip2Fr73b1aRo/whKDV4Vo3ROK3Oplkj0B6jU
uHXH+zMAhIkXtWezrzJrD4PL/OqX0xlx25GJsoaKEv+xBIFd4/BCqGEk5ZZIuBgWcw2L8ePyQccd
oJfF3kNsYx3Ostw0vx5UeJoRh9bJ4zCoudVhDWB1y/gqfFb1Fm7KuqrnwEHP1SzvrPpp2qnTaKZE
j+u8es1rRAIn7xdNssA9P14uMUSZm5TV1kLu5bRp39jnxhOMsEPimXYrif2xAHtKe2UpyZQqG76K
jqgzR+r/MGLecf0twcrvTl3eKMXy9VHnu1Fqn8vz6mLjJPrYWSkHONlfcYMrV6LlEiCgLIgIL5i2
T5zygvpGuB+8aJVERrCX/FilHD7MgCJgjKlw/Cxd2b5gHcyYiQKYl6inCwCNjxVDCZq0eqkyWNVU
OgREXL0YzweRE68QMJP7P2H1y4qmC8Gda0TtxMqJwDfbVRRvjIgI9+lArYSRj/rWeQ/UH5BkhIAv
VHrqOoW37PY6OlhQ84d5VwjBzNldCIm/A0sFFmn0H8zjjWfJQByfR8pOLTwCdehLJZCLSBQCbLwP
2tietByKsS1wVs2XXuw6t/dtb2mo7QgSJ+mDR4SzcM7XBVRnKwDqV1MDxsVYEpHZ3FLQxkP7B7eS
sSs+XqJ6HKlWPZX+xZDlgja/TBzCtLvDs5lk29vZFlGQSgVgAaYlLAYG/V9LksODSw3YJ4u4pDFm
yNOmsJ0rmPHGpwuulykKoXsvI8p/A0x56GvpG51i0UlMvBHYMiytTgtiRhisx0xI1J+JPuPVi1HN
j2VrVZx4Qd9xmRze+ZhUSm1nzdO3Y6LeYCpXsGIn9fZDuxm9avu5pwUKbO+fj8unT6J0fBo6LDyE
wy3lrzsI7oDoIt7xav4gbc0U/j5+nEKRwp1y/ecqarR8b5kXmERsOYEGE7kztwU6p84iCBvAQ7Kx
x0LLiVkOr0CBXcIG3X92gX0NYstawAUO+Wx2Fwo6guUt01YDhYpPR6XuAu4tgu/TXMQufsiW9AkV
C2aNy/zt71Wb7bu8FdV7vS0+oPugFxW2xvZT+RXRc9mHpWhSoIXCg/B1fj0CBwYUfgKBMJ/l2/gG
zIP4ERGh1QWl5rdND8PVXpPrshieHy0M3RYr18BclnxvkX3Iwz79kaejfwiuwLI5TvXRLHFuhXZr
HMdVgS6AL7QhsBxyM/GUb1MQBThwfVXii1aeZ1ksQNCh2sYmCQx+6hvftjBTZrKbOyHuvPsu6r86
CCox9cIK9galhsILXWHnKkPAWxGiwuxaNPr2W0sAj+YivcwEuQcib4m525aRJ5LZyQg7SQe6e6jL
R39/f5sl4V1B7PwzaZ5X4c8VdbPIsqB096kxAY0hPvmS93835jw1n0RafQ7KO18wFAOjScGKDgtW
KGqCjzk+Zaxb5eIZIIumbME+zaXPPJSzFST7TIWRPRb3ttfXpEK8UUspfVfi1QuEKYLeeJfTXVTV
LKIMxLirvo8bvW6ZmIxMwfnsO+CpEz3to3PY0NO5tJATtXb/tmFRmqhAvaDRtihxLRi7swkckUz/
1vdxD5Gntx409qmsJ28zElZPfYJ3YGdOsoQsaMwwhtqyClNod21vunToB2v38swQVkzEPbhMfoPT
lP0PBi4Y0dv7DH5aR6uVZ5DFuc9Ru0poqtuxOXsB04BOvHrF5jb9RVv8MHHkI7tRc4rvwRZCGpdD
Y4d2wGNb45xGrWC41RuhcW7PhysNKDnZdPj/2ggGCKNd3lzX8LVHAhazdl+xvk4tycm/bJ5KgGDq
9r8T/6vE2OB7yS5INWjf8Gqu3gY4kBJAq+BUlF+JInJeK38r4zFkNDttF1mR9Q+ZdHdkrFBeziZy
kRgK+wKCl9xNk43fO5VCY5DELK28ZuQ3kY9otBLP1IwBgmOv5rdefiIdNn55VYC6+wxvLmAQYCON
pzLkAQzmaXV5oA6NfjiSZfg17qYb6DMBLfHGdiPZeq+eFuRABNWhIprK0g5BR4ZJrFyPoE2GiLyO
3IrdzYYTXPjDYmcdWt73wpFpHHIadcDnulOReFBW4VXibDQzAIVscsDRtnTiIl9rE6+N0bwGcIXD
KPVPmOPmIYkWg1PpOhaXbaQ+2j9SlAd4kLLFJGf1JXZ8pA1gxhvrQ9fHWvzM5JJiWJ/R8W9donda
R0sy5wWklMTgpMT87/q2yfoC3cw2frDKve8J/OoLNttP7euQyKWB9wErCSghUoL1Xd3TZxGOzIgW
ulXmpwdXIKIwzvPCxvc66SIrUhSK9BxMaeBLCbs/Y4ZLwXt+qlU10lR9PcaJRi5r0oADslz92D4R
EZodLlUsQNR8BEhrWnXWSMnWM85C0d1E0pfNvGjN9TkKEv4ll526tim0CkHZafGbxwWyBFC2QBk9
765sEe8Be73hgBBf8L3lMi5qbfjXCXTINBq9KOXPgu166ffU65MFpq91ECCKP8nC83cOb0Kkh+xB
p8zJfn3qZDKMZPGdWGV9AEtYqYBQQd/OAmQchIBoY6c1Q+sXh9LWaNeLzv4aY0iEP/e5THP7DVcQ
JYkP1Bpc92c/yqebKZ8htFzHIPbFPrNmZkfB/KzyHKpRy4yqJLIS7PW0dEYxKVx9c5w8Z5AFZC6F
qyn09zv3ZZI0DfU70p9HMB5wX4NT2csdPdlQ02HPm+s6byyLWPtVXqkxYQ5Ewj3rabVx4OuJudNZ
VeR89GOfKhJ8sbca2IG+WDJyYnebuGY+mM/b0BBFdzCe6zUyJT+950iPkDimTODk5XqBwKau59+f
5RkUNR4HM4G1+oF4gjx7bATYUpltK/xf7REpGesiN5PAjdt/3rtHDR3zGf7T4D3l5zGE+1URFCqp
LQE9tTpYzG4CHtPaem0apHMsKw7BjfORwAcxudOmN4FbzyyTqv5q67xwQQtM5u5947GyyIVoagln
rRipTyE+2yOVnObcfcnR7Hjh7OJTrxakLCK32oM4JVPI0DW+iwqs3yvToXmvpaMg37URfF62tFhj
LLabi7g2wFFvVI8ZIc6OsgpCooXUwQSg38cqq5ofI1VG6kFlg8jFoItENpszAtWNGqs0N1bz4Fx0
GmDVmS2jmWjj+J/uk2jileKRIk1XHw3CxqFl9Gh+BqUpZFaDf9ZJ9Y5/1jS5gFoAQjBPi+jmBcud
uhZXRx1DF+mGiGDgsgPMroKSOYdHgqjcrYAkqfwFPkqYg/kuTWmtlIK2gF7xjAzGdsJ3pwBo4ACX
Cj5hRbdm5plZ0Fqs2mbUYhH5eUQt0jLEEQqC0N2ddXmLxyCF900aIRs91SvebX5LkdFR7rQaBdLw
Mm0ZojCFi4S1DhLUX7BQLfgVzg2xwShczUHG223CncgR/teYbLnovdY+o6RlxP8a0toa7oCP7y91
tnSfKRjb9BLQq8mX9oS2aAmRRMHra1ecFSNP9FxDwWrTnZ5IHpa74zNeCCKqgoSw4CZkz8F4MknO
sc/wZNyKk8x729d1+bWrD1C1HlBr6bjYi4eqwjI/ocSFhpEwc5edNh99Wcz+/4BHVujeRVDIRKxy
ZzOiMFIGkH8Zb8ciqpaLWv+zj3wDvADB2lGZEUzu9+tDd5WbCTR4ZygM0BLxn1IgaeyBC3jErIuH
FxidaeDDcrfrNv6wxDemwcg8TGZtAIfRCf71E064dE/zpquGsJSo+EI9Fmz/TOgx+1Zh+YfKkNt9
7l8jJujsHgrQqa2xWS39WgasvcMM5NRElvhaFRmMBlCTgccQCdppNm/fJwOnFvTPm9yUiX9FUTz1
4dcVvmZjUxgsoD4dI2/3EAI3vZF+UHkkpUqLeMkeEWMB0p2Z46eVvNXsBk6KUUTSSjop+SBP4qyB
l93U5FlKU/NYpbGrBeX9UCfMt5qEW/+4IKxnJUhXbbYHxLnHVM1bSS+ISki+qSljzG0D7TFkyAon
gSTFEBJQFBRof9zYQVDwzCggGsW+wtomPeTB0QsuEgTghe1Mg7VYwMb4/uHeejN0a4phEx9JG6lk
vWMxaUo43iEtFddaTz/rvM+h3UO1OOOOJhXhPmpska2ALSvFduecX2qv8YHGLW0H3oFKvb4cB0Nb
OBX9N3Ctp0p3BzBGLewFYKVN+hS1D4LMbHTL1vQZ6ksCqyPbEmTgboPjWUwIVkBbt2DDIFIHuc/4
+kjeMqGTn+24fPxl9JDaM1Tp+1RHJFri3seizqg2Ku1RGu4UhCisgb4238Y67GIOYb6OsVtKR1P/
tHWPYZPl3iGsGUiWyR7gAnqqaCDJUE+PDKzpAUt3YR/bnsu8RXWhe8oyViJRPTKJyT0MxHwrHoAT
96202TXmoEjDlpnKe/AJQlxLrQbsbrjl6YzmSspsUQR3y2QEPhpiPftrZIYT2H2NU9aZdJAWGVNq
CSJjP2C8Ain63Stvm7icgmonhccTcnKPZtiqepAJG79WyArVpC8B9H6aqm2z18pR4wrQ63CzERnV
DS3hEFeZ1wv1Ck94jqrt2gt5IJVV1iwg/JmVGP3uPl8I5cMCfLK6gkehE50w4KrrK6VaeD9LVKfu
hqzk4VAhmd6LIzlrhUPlHFBxRVEGFDzTxtfiJ975jgoFazMwDA6gty9vLiBeFFl0Ldrmv+gKkB4t
mXFdQrxXXJUAHoXQ96xZ6Y8BULI0HgsPGmeAKhiJOFepcjd3CdZEYi/KV7glIfgmVUlbbZoKS9We
IvHy4IGri/5qqDzJ8h/FHecRbvZtTRemT9qqlH6srQZzRWqXeIg3cCrdqb2dk+fFb3hrLkAsomoY
G3/pMlb9YpuX/RP56BLFbzY7V+3qiuuI/RbsjSVFEnCFCCthF4npDkjwfo8G+P3QpFDq92Y2dN6T
pnk/WX/GWoR/fXD9FUu3gJxa3aZKdpvw5TQj3/3PWU2bRMqKxddAdA88U/yeEcSKRGru3wHPCbK7
HIGY8WtGkqPcjepxXlp5T3rsD591j1NQ9kSjavmBwf3g58PPt8L0IQ59mUf16daFsqRombqPyFnq
nD782CTN3pOCRod+8lILOajdmecrYoikiOMNY76FhFlqttEe8PlBvJCiULPMlWT9QI1mNGTjtYMG
Kc66ENXgDMAyP+huWHA4XXAA2B89V4Y0PbwWDiVV2jWopSqQ2JjJSlcCrciL1ETWdXRMVQyCbteo
VMuQHMxGezJ6LozNWlePAGq7J3LVSLGkgoHeBUgc/wcJAUWJJ2DpRUS+3kp+pvv86bUEp3SRNXV8
q3nRSDD2OhY+I1STb08GBulud5+LEq3JCCSLAE78MwggaIQCM/BZQ7K9Rt6CV2qIwUJUI+3cEOkl
yoMQtFqp2mdODbi6SiigPTSNq37czoWCXEZEC1g1xfqtyeDzjI4q+bkR5zGm5UElIG6XNnVyyxy6
XSmrgkmk1UYSr3QADHoMBxJA773APBFsn3okxHbCgtY4wNjgaaErirrAeQuXk6fgdebJ3y4pzqCu
BiG9NNJlCB4JPek0ymzodwYpDXCuAzJifief1PUVTv55ys5+r3d0rBQV7X233hfOgfzoIIzhsCIT
bBs+O8T9tNduChHxpLKp0fGhDo7DOEW5NHUh9jo3BDCoZQpaH1HXrLl39FBjpVCbhGcCHD2mMM9T
tUrf65pcEFdkjs1p6aB52DiCVOcg7hZkPmRcrQ2SLRScsWSXPc6SDJ5SLAg2kKHZrIFQ1Cei/E67
vsvC629PzP6wDILqMzYDFTaTMAi24U1gO+vwAJhgUsIWK63NJWJC4xJJAbThMHmknldu68s8PRWu
yLs+me/eF+C1NpG+NoGgtmdOAod0Sa9Bf/BcerO0mDXDURGSwGVRnyNIsKfWckGP8ScyNY+zuMBj
tMsPSQj0Ks3mSfhg3N5f6ZOYLAiAzd48TZ03hMo2W7O1s1lIjnlnsLzkOUo+ms/7XBbhkgcAn4Hz
lf6xIMGLogUY0YvitjRqqN/zUM0u0Aj9ygpuwWgea9HRbOaABSzNjltD3mYRYojy0OD2+7uuLv34
QQTPiuDrgAj+L6F55wXn01hLaY/KEwzoGjcGgmZLxGDfCr/L2zia1CvfHHfeskWUYnoahmjwsrGX
RVk/+eG8IuaSB5/E4psn8wPE1O921hbVTw3ZTXiQ/kCshHxrUN7gHhpAbZXmTI1WqKtjv/E7xXb6
Ws+Y8Vvx7jYoiaPOPDiaoINZE+I0JReWE8u7nxgnYfnU+U6deT7tVA81e4pLii3A2aTfXf5+sPsL
xdHV6jJnOkTlBK2y148pQoTm31qWgJ8vkVdrNkaa5/wSup9Pp0jEVS6cr/tWe38jkeatEEP/MCcG
CtWS+dDMNsgjhTKpLXXvwEiI+g07qgwhXJexm2vspDyibG8un/jNRDUQfGr4BNSxJ6nNy7pqFA36
Eu6PV8/83wY2ScPddlQGFEjXWIvc6CecnY2zilFBUZXVxyy0Lq0XBCwAdn6y8qqFCWGxVvPiYrD5
U4DlbJpjArRAWggzWd2QeGpG0oi6eryLwG7k09gTwHOwPOOjQfblYoZbdOEB4XU0UORhLhdPX2e/
STFpWQdNZv0+xxAGeahbpZgFeRQs6v0k0QGomeyyIGoWSchhquvwOq6Fu4KQggpvqSatJAYmtzep
VlHgcoBTsuT7RJPskesramKehq2A54Z3+ktGoh61KLr9aM4CHas3IUagzOajViE6Fd2WPcsWlBE+
sHl86FyLf15zioQ97Ha3U826ZcHjgJ9yH1DENMbf5sby6AtwPQ9HM91CWJi2BAqLFJaz0yiUc/07
5dkCmecy8wSKN+EZuh/+cVGMlrnL6vmBOuP2acdf7mASXseEKN1kGcqVTNk7iLKOhYDCY1ohxZxF
AVMiiIfQr8v1BxUPMYVQlGH2nE7pzPYcW4lTAHt05xAGufy9AeeMiDpFLnd6K+Vx2VH6+bqoUfwi
5XHQyIN0ZoO37NAWGx++DbwRWGL+xFhA52YXnWpFKz0jmEpnNpx/sIoUJ65d0XXKwMZZdmDwjkzD
FP+vbbnEmAjKJZcE7uQdhS97BHD4GSmBeJ5H6qIHfoPLpQZU+QVdCwIUld9v8AZfCTwxxTP8Sguw
VLK8IPKKTtQGA/2UY6q8Y+oVKJ+S/BmrrUdM4ZPf7WC5F3xkkJZjM7Kil9svP0hCmqd6Fr5zKfjL
LFrBB71T3oeXt0GwxDUlRoc22xgr4TCJFqdSTh18Kp6OhVzteJwu0nOZJd4xkZyjzSqIALgUStZX
RGxXT1bgXAdfU7/bRGW1wznhpeZGc0znv4Z226rwKwXbHrJcl1lXoW8zYGyLDa9510rJp6+M8XNC
v80P/DUUrjDCO1/AR7ZTiwWt44n7AyXDy19nnaCCo7mEQNYlGYfpv1NTl3AaXrGkE5HpUsIZlAD/
GNNQXK2Im+xj+kYNeRqgpcPsTfjRby7ooTzgqPwyvHFv8cm+slWHU/4bPZjWG23ReuprxPho04B7
lCjXF0xjhRh6csBiFzPO2C5+84OnvK8L3Nl/EJywutkEfdugrl7M8+D5OXfh7g7UPFWJBemynmFM
u8M5w5EeBN3TMZIcKYcFLRLZN0LEHUZge2FL8ZbhmBvPtPkpfJfz2Arq/wOkwNF25VEcMcW2Hk5e
vHrWuEBNMXoDJPHyn8hwr0SxhCg450/FNsrghv69UiiJKBFLvWsBJSPPGuNqOq3Ef5DotBwAL9kk
ekZAr8/BzXi3RhpWD7aL6+vIsAvfZ9eynoi4+kxzHrr7+Ge8obAkv3aIGWM+VdLrvSIsMIVzBWfA
y3UKSjMsnHnFScEUa3eXJYFDwpBGU5fc0RO7KBzmH+GsOPiNMucT6hOowjSSZOwaZZsIR4gshjzK
t6w5Pi2Y4Xfsrn3FFarmRGSET5Dewnlf4heHOMex45+i+kY9439bjCoBnLV3eqYDTOMS7CvYWAq7
Eirq55FUtrbG48qqTTTDXbuLhwJGn2MXxqj+w0Zg8dIIleLl+kVBlAOsnhZAvD++4oygejnerRst
iNPOb3/ImFjZDPm57OthjqUEQesNuVtoDBtRhAEkH7IuduE8jwyDT4r3tFkm/CQhtCQ5iLQd7qyB
xNNrekKs0bL0qrjt9NhlKmaUp2ELkmSA0WzJZxZmTb+63aDRj3l5o8GEN580sruZfhHtvY6hZqL+
LTVp5Sao1g+PkvLrOSDioOMUQBuujTQJxayHAyQ1CA3VVaWBdCbVSWTCn0qE0pBXBh1Qx0oRhN0O
k1E+sKc48Xo84bZoPysuc0hpA9rl0xgpYkHjr/VkkQ4nGRJcLqdtZeufuWIeGbXNK/OGiH62CfrQ
u02Y48Qj4309CkWKNMkqaJf3oEZ9SQBFlLsrCYdMvjMYPNM11NgZ+ZDZX4/lv1OYbx5mzbW8ubg9
iBkIWw5d2tzRRaX3GwORdnOBp0YubZrRlw/ejuDW+KRdoeafXhrSYSL4ClkVXeqkQphjcJgDvTUA
JHIWNx25IL2pFQtEw7U6vsGqwhF6BSGuxMDMXPBk6NmXQNn+vo782UiFKH531BE8dGjM6lqGPj65
X29TWwMnD+FBOG8l0JaAqgeWK2LkK767/Fq5beazfyZpbQsVKBDOMzgqn0D3ZEeruwvlVMZ5++3w
hx4hPRZE2yEND9h/YdXTK1JAdK18kDbSLJnze5O9pq6ygUdPzCWO4ox5o8psxWTPgAD07Rz2tMxL
biQknqW4Bp3zpgjk6EmFH6Hi4Q+R/tyIxJ61HDL06xMAWez6t9kW39DJiE05LcOGsCId+HEe2JtF
c/QXG4C2Aq60VQ3ONa68tiBe7DBGCdauIoxmYSoYlho6Qez8MnLswGc79pEmd1QDZVx1u9TJm0tJ
KT9wt7YienrfJAXcCrJCtd8wv4A6IQkCr6N73lmTGiRFMYWLNRsQvUH2anwzYnG9WhnWeWp8Pjoe
rRDPWDUZjuPzISrL5HpviMgQpyxpbDk4E0yvxrVx35O4eaqPh5A72hB1klRoDc7w00O5OirzOEBo
Bh1A2XEsev6GdFWlXAZBAsN2So/CgJG7g5ib+aU3u59LBDxwMfWa/Afa28X1TQSlg7vDQp/dRIds
4fXA2cAWWORB6j5IpKyNtQjXQo9lchW/fDD2tAT8fs2VpdJNawwe6G4EyuJNi1xBVWLN27aYMKqN
ButXmBpW70xfI5F1RG3H/QEwv9eLb/wlFtgavVmTsyAp+/fOeOKy/m7Fejak3JU4yN49VxdLmjzq
Sckuge1tZdeHgP4xPK/Qa54x3VY0kDNE1iZIqXdifPXDQFKtIA+ILXQXTSfe+9Bm2oibo+au4+AE
6TvNVhdRoUmhI+vhWDOWrpYunt9Mnh7ytNGk1lBvaF49NU2ygJ3rxLFtTD9EDQfgTN1AzKBqLwQU
1y7+9+9FaK+y4aEAg34R1P3+Q2yDh6Rl10tjYGoKlR/N8tpPgopDn1ifeR3Xjae+4n65iO2sFson
HsP4KyX0nBrO55fzFm48APY+OY06DHRGuj8x96xxzNtEafrBlQOGgoEdImWI4mcffnxIA/EzinxM
1deTd02lHC4ys6biatOhARzoWE3NOLGsAOuR9F2DTRkyj7RgC58YaVT/vELLnJLHK1jGwlzBsgZn
gKuUNSgz6b0nyLUL1gJiQUkcgp3zg25rXpHX0BpB7QWfhaefRRUH1+20iM8Sn4acdzztUKbbi25T
0O4ZCiPIojfbKrSpjQsMkSRyuI4afwC64nMI94HZkQfuCcVJF+HiCrGMSVa/YqIGZOl/wwJO8Ii3
e4CKWlFY0Hk2WmhT4RWTBLqjKEvE13ZZ05jBKitBJKjHgcNTnHIlX0n5bcMf2AjASmzZWX6OUMh/
q9eUJJlUudLiuARvZ9G8psVxgGoameFMkAd7g69I/5rMRN9NnV9I9E0WdZthI9POThbD9BangHlG
bWRvZFEHACieBAdxF7kiMOfsiktSCXGVcZxkC7u3G4yzJV5azeP5QJL1mE20hxXjzxx8xpdxMx0T
zGRD0EmCHlOzE9YaPrSW69HHjJUGbQJBBNnVZXtyBs2Lwaaa+POOIXO04RmR2BmCLLKHKF0ZGmuC
0gWakrXr68fCsogEqzHk1D6gDcUozl3xctd0jTc5iQY0tuNYmEmQzgZyBCW9Suk9749YVAwBpEoW
Cae2ZW2//bAstufcaQJ+a8T/LG3bZQJNZOyzxPp7Buivvo3TUOm9NOSRvdTtHPxDt3Dyeudpi/si
OZHvIr2UYEmwbSDtHYyl9zAY6jQ3MwuuC7HA2s6RSvvBC4E0zX/xBPdPDHMCXfqW/hbCjQnOHrkc
Z6Ct4slp0iWaGtlNZhaqL0mK285D/fZ6iK/AC179Gxm02DeeYafuH0gKRJZDvjB5tVMs9ciAGvqp
OiIEhseeH/VJTmK5Bf7j0dI0SNT6WpHcXwdBZfn5nzwY56olQlsxr4PCw7EnG7VuCJORgEsBtrQC
GEGafNnu4BureGQiY2B6X9IXspiTGDDr5IZtJ/YJ4MwVT+pN4W9vU/poZndsJ5wZL7NzvavFFOFY
cKlJ4RyWXO8FTALb8ZuKt/uLMa7Lc5ZMzBzxBSKP+zI0Ai+Q0PoZASm1mzWqI7BdIp9zfeRIbVdM
1ONRTEIYJO7luAPRjZae0xSJuepngn7z/kOBcO9hQ7uE7bARdBanPyr/WI/BuwDXmj8GGLqJZ5Md
Du0GxSBUH4AapIePQtDL/QHnPAgyqQPOLkZulaVhGeTi01M11HG7qaKB5g+IiYofZYbV/aEwWbo4
G37DIc4LRIl6a0t7Uf5Zw/JIrLiPNwmIIyD4Lw9+YB1JkCA+lMF18pR0Mpj67oQuMk6s9dzGVbb4
I9SDq7CXwuVF0ShEV8ucaGBjajqWtXJV9yI46Bo+jeUa1nqfYusoRqSfO5A4zLPv4hg3JfuihnJN
4ulmM6eITTFc4A7nvWgzvKgevpf/NPCzJlnSzbE15iJU+cTR13pB9TSuhw28UMiGkeini6RgEGOm
oIlCyyHG51TDcvsNkNxBWQgZop5XSNOXSN0Q04+q9GfPYu13Qo+fATwfgyicGrXKeUIw1tYp/Q9l
c2ZRcefZi7zbn+3USSMwmd4ODpaQNqyqJdnWpj6qSoJyZzebJRc22x8uzQL85AFqJTinhNEVyYug
Wdu/sYRFqRE8zrGV48Ov65Jw3jsSmP9ZzX6dtwUioNr7cBymGWmRsio3AY1V5U95tjYNm7qAQt2l
4cj2ImWwESyqo44f8Lkt3f7zZLzB80Pxm74UCJ/gGLU6zgUBX76snW17mFe71KQvZ4rLMr3ATC+k
16/TMAdtSR4zT9J2WXURCpld4EPmMMIy+fvFXVHkNaGhBNrhQbAsz72F30GAQmwR1OmNvT1fees+
hq/UM7bdkt+krmyxoAVaYNBJZn7vENG0YNyvK4N+CT3fGnTRMMuzwDcO4Tq/QgiajwcNdlgAS37y
11vAaSuVAYoc7o+2GxhcfZUsJ0qsD/CAaTJdYEdUFKohpJsMmf1XLb1RKYBcb/s8fiTL2lKveVAX
UyuJ1/1PbmCm04PWid0cJlOoSXW8cGUYIugA3U1QfVqIyAvGIA1KDaJeUEK5R7mfJZS/D7FXWKM/
50o351WpdFOBRxUeqyarBxS2CWufJ+2rOB7vFf3V9usCcbp9f6RZXvn01IQi0ve3mxSdHexBHWK+
rDIzBMJuo7CTneZIkfIefTY88f3J4212CJrnifPmCZZpx0MUjpyDGDd6EuZAn4B9wijZJ7BsM4Ic
wdoq3Gxx3NLL1kRwCu82A2zZTzNo/D5jhQ/BEJberh1vmIaCHA4/3AtJOTI0bnL0vVjS8qw2tkt/
BV3ixrnCjP5RYbQdlU6ldE4Rp04Kv9AtJSe5J8URY6kI0K2BSJo8SUlypaXq4QwBT2R6cjYIxNYe
ank7YB221uByVHZ+mML6bs0iSv/BGf5XqlgAP7Id0Vb47exfCISnAwCNLKJJklHY1sOHZm0TB35m
Is5bDg7eipQ+Ij6APROZ9JRMWMgcL+a2YawbVuSYO/2FD6Cd0DwaT9o8hmWfE5id0zJ7YL+7e0JR
sCig7C1pobNAlHtvmUiQBS0uhp9GoAJIbEIoFzc9jlVONxs59Y/Qj5mjZXek87f2IxjBTGUgY7QK
SR7rTRoHEJKYQFMDV67dyLeWXlZhvO79TpeVw2OQHct4gW6+1hKRZ3qq7KnxSe5lp58Xgqq21uzl
90BsqwNEpi36D8VV/tdCwCfP3LVJ4vhlymQrU80KXnLeKjyhL/k/CR0Lmd6ZY5WfpFYgXoYD32HJ
qZR8QzAl4EvVWKPx+HRGlNh7t0WSMSVTFLuNEaGgA3DhQXaAZTPOrTB6FqapPROXDFoVV0R1qWeE
6DDlD2+QlQ67BYI2ggoaJ8mQpXEpDsy1cgTipE6IpkRLEwUNJ173Yi8cv2g/wPSByNG48wl696c3
2sqidM7mcMdCUemlPv6nqr3XKJEK7nWZsCeWZ4G3yCyURzypxuKeYNQWKPC6xQ+3wZ+HUgovlI7r
Mk3kj2Vma+zEWe5Ly3SLeNsvB8cNxz9WltRX/YW1Aa/VEyNvw8Iy9SSDvDANjCjUBFwTXZzpN5da
XkVL0eXWwFszLyadmjqPlRuR0/aiM96l0KxKKJ8nUtBspNKKRRjX9EXNr5Y2xxZACdJHWnF0hItn
6R9FZ52AbojPAjGyWaKz7lthDSxyZXO2b2yJYxmFytW1s7ElgRRe+sHs3j3ecMhjjVUmVjOXTW4N
p34c4TEsX4WLBcghG85/uTkzIcj7aOcdJYqv/NCETKrwcc5JN2OQrsaww4GrM74MGshMbLgZHHwO
QpDPYHpJlVpBmFcpsfOohxYtuiypWksqCw7kuCsh3aPq6lozDwwiZrdiZCMhoErRK2GCCzyn4ekC
YYYlkux+bOSSxSSljHTO9JKQ5g+U4F2SM6PKtDQAITbEn7a22+PgLa4qIhHEqAzs8wHMegu6FCru
gRkfjyGe/3LyvDTG9tTM51maR28XUPiElgA7niJZXnbmd6qqFo+/nzRCOPdfXtsmlgzUUkZKq5OP
CBJEZlkOYLxHJNNvjfZ0SuMr/eQeZYlsROORtLuO+KFvzCCBtEJrM+JGUwgWDBEiYFNHueShMgQU
+BeMl96lt2KnAUAvu6SOCsJkG9wuB2+rViPBTkn8ReUWpYK+xwNqRLW9UzrhSD8eTWJKQKmymuE0
R7UTYN7pPnNOWbD4aTxmOCavlEhxl9HZNxdtiLOcAkHcjZHNVnjyINrYQK07FoI51JtaDGcL7Q8m
kjSBV6ZuYPeOwFRPCh022PLeOnEOl9NNPG2eboeuesO60IjggJEi0a1fpw6R7sFZ5WqtzSKPWAIz
IEHN9pwR/jYNsAWQQm0HaTa6QUVj94dR+jS8vTMOnwaCdh4EXTyXt9kPSHqSLouh8HtJMu+PBKKt
ohaUmeIdc4GfPnZhQdX0uEjxYlAllp2Msq1JsMhEiWdf8i9m56ocI6AkFBNB9vNwWqLK7cB10maD
KJ/EJ/2BypJ5NjIIm6Ef7CSwNTl948D2+NEi3lDJHyNIkrH0PzrYZgF0/1Uc0gYBJceIhDq4mM11
ntyq+r4RigQ8ijU3rxZ9DQVHG7N6w5veiJ3vKIg5OPd2WdjtUSwzRr1R4iQKamtm613PpiUF8oyA
7gJgsHXaht9NYGGYtaawq74VSdh5XIaRtuotEKR3F/HDzds8EyMcnGKsH6ZwzZ4W8ILh+sWTKYsJ
UtdN5dEfup4dwUmGJYiUmmTz8Qq/eSdE8TWkTBYhISbuESM4s3flkDBlp3QmnazDXgxEVrpO2MeC
O7Y0U0DeDOw5hBgIzT9z/1YmJpBk/Da3NghV+ZD3LPwHrcAAqcZEQZOYpr2gKHZtjmUd4ShKDl5N
Jp6y/N2KoZq9V+jBit3Cywl0sGo5YwcaOyqu+lf0r5aXDL5Ouo4CxJdq1yyjSY1+5Tb+3nBkmJrL
M9ztrH9DHjBaXOtQuvnQLP17MpU0M5/wD86S6qU755tBJx6AE52K0DdCs5oTfLK+1o2xgIkUDF3+
MmQ8M9Fnmdr+W9pdmLo5yX16fkqdUOmd14hFU3U7vBog8c2nBfqZxy9y/KaS/BbGPFGuEKpPTW8z
H+uBYVabmFEvbcNINjLy+j4wWI1ziz5hqyTtdq5dTiWjMDL3CjRNV+Sgzsxo/dw8gRdi3kPRUT36
ZxIAOXrCiMoeUcWypB7omGulCiJ9BBbrrUxc54K24ZzZ4bKsU3zJk6/Lzv2bLLmOfVxJ+egDn/e2
gvuN+1UToA+nughTJWHhrKe08e0Cu53b6PEThJiYGxcBJTTkwTVZY1amVtfMS3lOktiMaQuAKd6W
aHicp6mX3FJSsAueDNAO+xoedyPbOUgwuAz4reQMDR+w8WkhypKzRkG+hqKBOg8X3rReqzw1hjmh
9c1QkLXMebgtP/QTKV+6oIGvkwqrlILevwbtxklynAqW8Oc6lq4taeXGxMnvjbaBaM0rS+2Va3ZL
pJmAI4tzg5vk+GLEe33PxCfYrbMWAYVAvvz3Bdq9GLJJ+RK2t1M6YunZBL+l/X2w5qO0Vz+vWbQy
qkzK7fSjbLdg9gMqlTo16LI5lN486RlXoYK4n/qnDKTGq4yHrdRMDAs/ZHxVIFisIOO3CMM571HD
+TPGoCAItAH/1os8tMuddiWTvJhlCrkkrPNIphDKe5qgy8z4UD6kfNQjEeFgVHY+3Ce5JVbrag/8
Bf6wAXIsHU14fJGEOOaiz3Be12n4cePg3F5jrrqd+bvF7YG8gnvTasGKHqYcfiKB1llNIJi1jgpb
YAZPcekcU9eyB+lW7aqVBcpUo/3wqZXYbJMFcHvqZsedyyct/FiSfxkdUJduwj1Hh0/tMKGcyQM5
8wEEmVR1QUZvJ43qPgH218risJMBOSMGqsm+b5Thb9v9eDUD04R8F73CcDQd9oll4q/TbO5kWzyx
UBH12Zorzk//f9B/Wyvd7XWOdkquwP6/VFf2BdYPWTjP8TZOFSqgdfUwCP16cbtduUsVRQoj3QsJ
GSfVebeiAFCV84ZccDuD5w0OIF97GAXrinMoX3sdJ8zaa10GCwGpwdqitoEen2gB3+aGVcohLoOm
EYA0EujPTw0d6ysgTqQ6x5GGt2Zjmes3+v6gL2720PtGV3HlTTqt4RVe54eIFxtC/ZyXzxHc6cvn
mplVw/aq3a4R28wFDaVdN1HvBProCO+2DACaJ2tE6qbQ4QrVhPZzPUgJ04I7lsOq53YAzyrm0X3O
aYQiYlfPv7bxad/cBDMmm/zaF0062WEdUSJMtkryTEZzxSiZ+g0dRhVfcyTxXzCHT/rvdoeQ68pn
fO3vDc/o6C1eTUxn+B5zx9h3AwgCcdI0hWsDi1J/CoXOi3Nq2mNB+zyB3EpMIWbXBMYWdPFKHz3a
SMRfNUCggN05aUAJG2nLAPqPmKRFNrVLG4x1O5k+i7TxM3QJMc9YmMeTUlNtVD+zePt7sPptUJFe
r/9jRQHt4Y5KkIeggy6I6qHPWskbtKtMlIPgLSjZGpjtIS8MdugM6XDNhidOfDWmw05MjpKP5j59
gg5ZO4fUUX1TDEzBjRKZxbiEb5a2HLLN0Q3+iOTtKQ3zdVzFpMfS3scD1eCr4qvTu6FLDl4L4x44
MvdYAWMUJG8ODiiXn9/fZ4S/qsdXEZYX6Ng8CRp6w8GpZTCYXJ9E+TsOoOsl999XN1h+3uMLgFO7
/DPmZUAF/vMMipkFFqEMkMg8dP0S74Mn9ZvUdI/uLG6pUCto8NMvPw1T9zYroCZQgt0rHfdWNnct
y54FdI8gZ6nALvW727TtqmAfDrPfYGJXkam+An5nmAZaycgC3izg0KB1/0IVU+dZl0XF3ZMXFeE1
GW0/dREQbNgmzF3XgbU6KIwhDHF/2uX/S5K8HvaEegKNzst95xaAMZ2gT5rIdGIo3FiXgvY+912f
vNzvi7ZcksmPRihzX8epamRFJUS9lHhMwcKJ+zhSBtfmVrEPg3/n4M7Q/EegIWwdBJd5hFmybUsX
EV+n1k2AgplYuQxkxwaYWVO+pU6UYRFFicaa2u2gM4qBjRuoDbeOQAoANMyq8sDlP/lDEd1s5nI7
QhGuawsusIan7+kB5Ma02Iuqyi/0W2JGBgGxx8mtXLAAvmDHd16NYLlCVLtTu/Tpabmf6mas5sCT
xJ8G7fiE8WXVU80nkxeSxQMF0dRGkQLjHPKkUfIgSGsHYj6n+RqQDX1i+NN0z8cOGYWRIGzqShFX
i6ok5ZBbLwFPK1OwFC4h6GlfCLo/u3bEWxdOgc0rBDuIy+w6pVvVUJZndhJbFQjtIIt8LSX2cuQX
lNYUqPIBTOjj4s4QixoBjeOcTcTW8EaXICqAyco/0c6cRDsR9VJOXSndxycygVuV5RIonDT9nj4F
GaL5j8NFyQFsFlMWunr9B4Gv353u/H/CSj0ai4IzXeanWfRYEnjs7TsSG90DLOArDkrDrlp6v/Hg
arlAtxy4HuixGKpbST3SBjCU28LhnQ5JU2Yz9vqpHrU+o06VHo6Qe8jBK4z+qkNMGV59dtOMlARr
dv0RjKjjcUiwcEpt5ObH+BYoStXmx8uRcuQkMlRwENbuu/v/xbBqufOxqTK1W6Uf+RDVgLReuUrE
4v4gtCHEzn1rR7HviG9qrWlpssV1lfWUYj+jhadbx7Qssylri9qtVkvTA6NMLlMmDBs8DnuUAPkZ
ncQri4NQyqCukflTd6IPiyV6UcueGsLidMHttJJP7eRTi+3OgoIS/TO8wUAxMHPTlHmc6HkUAVCI
Vl6xKIxuuW9KN8U/DDat3sLczGplQh15tg63nGLwx2+V5egfxOOO4z++wxlibkIDxSmbiFBbylIe
9WXQOdqVk35/SrAdi7bYoYjrj8DvcSsUZ+El8L4BeGNG0sNREyHWZMSyDZOGD6d4qdK7p2NJnz7O
yYJxu3WDCiOssIp/aBEWt6JRM/OdeaJ7+lZXyW20fJ4U5eLmusrf5au30UK4E4X8u9vAoFsG+8+u
WG2eGHTRQBJmNvBu7AcpMaRSTrg940hwWnlX8n6d7Uttrg+EDmndcWHdK8g/kMNcL9AdwwW1Ph/R
rEHklI2lnYZt2OHPIwnAgxuu2NvfSpbJWw5bVaFcPoTwXIHHepoW7FJDWNCG9lOtO/Rt1YKBcI9c
mbR0IEdOfGMDaG3Dmygp00g0h/WtkPQh9HZwYz8jt+vEWyigI5oWeruX+tBxyUh/1uhYdVUnEUVh
neC/+Yyn8bYAgmLDkBYEMrOHePBqJBt+eLdbHekM28YxoClRS4iilx22R4/nsf+qQ0cP+gWGxr3O
7/fNVAYpSOkWNWs9KME6z0A34nWZ0OLfr3z8qrsmCG6FmZhB2RXdN945Yr+W9/2h4AkvW1LHh4x+
0EpyCg0/ATEl2ndxmrWL0IeY7nV+Q8XC0BOuYW3rY/zOW43s8rJUqT7NzUM9MXmUcgvxayZNwndc
Pac7ybjGa25McumgGhfCML2NCqxGQI6kqmJeB8CwrG/t9NDOXGIqk8QkRy9xKzzJ5TDtH2BgQqxo
SziJMoqOx8vyx4W4K57kciHbN6iARbn3HjCBHeT8SHBqDjyjrMRO9UAOEifDnI555jGNSk+L5H7/
RzzDBryjyU2jjS3tJ8yGJK9yvZwfYNrNaF4x2EqAno58QlrBm16YHXdj7h3LtTuUjDzmi26Os/vk
2MZB+qeAniiPxvHpoE6G5og6XApes4sHVdp4/JNqQCuU6s92WyNPuX3GSdfd1T1OzjnApBjzme+v
+DfOCi9TEFjDZY7T8QX8igRUowPg0TWZeBSWa7frUjk0d6eV4SNaS92iiu4cbTdVAOn/wcXMBdfa
O9uzCS6R9kCgl1qxSuRYRhftQFfrAyiGevY/8PhfWmyMRbfX94CXmrZnnUXeCN1GXCvUfAWylQdc
15M8Kpdw7SHlPPXxayWam76rR2S7nFTsFjXy8KK8SrgIzeO8/XhDJ25obpKurN71mu/EIKdNaIem
Jy4giUZ5BrebuTfhwzrPMmEuTghu8cl7ASPUpIf7jPUmtrQLbKxhOPwwbbLLLe90fI/OYTDkzL/m
W+/1bnlHk09bk8yjm/z19ZqzcBcZWeZzJ4N4be0vgzkL6cN6oAzWYw/MWVIAd0F4fQ9LFu1ZeHLw
hgkTt9iPYtqyN/ggdB2pV7QxlHieqcWSG6ONmNqFnCkkqDXo0JFtlge5sv1NeBuPhp3Loy7ogJ5A
atq6TZWIkYJIqS4WLSI7t1bmwfgVTp3eOPCobEatQ5bHULqwQMGhDBNYnJglIdTKQEwzuGKu8xOI
9pbA1b8QT+X2qF8XNpJJKCECUALvdDaGVrhVHOKQ2jP7iXZF0tgnyE856jqBPYlMwZ8GO7oVBaou
IRbH6bCtFygYzU4zL9pSYhBAnbSbNWHHzA7hq2/Yi/aR2is8jcACGQslxOTE/njkDA69EEIDRIwv
EAW83NloJLZJtaicVaPu0+/CdUopdLlB7VztskryY/Dv6Ue3BH/bd6l6OshCdTmGV3uP4IKvs2i/
vmDRVZfpwDyrl1rQ4pVqy781HjisGARwZd5Kqpkzyjmok459eO0BdyWtm1DTmp1HIWwpKeptEPuo
ghAlXadEfB5sqKkDkOpCCsSU+FDVa+iWZMxvtW/oM8rKOyltOWCo1SlMx2pDZ6GDTCcyAbsAAkX7
DtMr+y158fhxroigaffF6HVpkGbxci+RauxVzBNOTRLOuZSms9nEaN+/ttTrKHqG4Ly3nLkurF1U
gHadASZaVBkZEuqK7wPvE355IfbH9z2UeZo98TGwrh9BTgtKSSSla8bsukeiIvunecaOj70Gd4gK
fH+oH0uYDBrp/AwPUzHIPbJKrFamq6Rh8TT+dWy2PcZF0e4sTkMybqKn/qFDhOfqGNmYK1snbjxK
1sX48njpR9MDAi/b4Pd8LxTeMt3o+k3h2U43LhjmxMvh/5SuL54ZfCuvAI9RxFkkaAfpch2XGSm3
vYsM4BeoR6CdjFLeiFJNxnu+C5W+nChnwc1WuRdTObEoulEwhuDqHXJoPnnFlxXGe8WasKEdbX1F
odyJGtxg4tXo7tlvEUsnjMI3XS1Z3XvT1guDfv4ENJhLQInD5JCxNWHOR0gO1So3fA2WW8pFizLy
6CISMvmmQUg8b5t5bisW95WBqlngq28JQkHK3LrlN5feKtpB9oj3LjzDBWa3ecs9+NwGdHPKZhPy
wVGWauHyAZYToc/ZeKwVLdv9uz7jcv0fcddT4AQosJNYAnSZDFdyc6Lo/UP52CoS4utXbNS/XbDJ
AdVvScvXfRdsBkekRp6tHOdkBJgLwJ5eNVMAAnIDH7LaK4I7zJ4ZJULoYVqGXvHyJI3W2CP478Pt
dgOXaRIxhNfx7u6W19glcWkSQOKjUQSrmxhodjjo+w9AdpJeWVLKPXpknDRPZyQaY0MYbXrLqA6x
2RAEDA76sDTqmgi4AEZ3cJrVoYIAaTe7UCLc5+OBXHJfuygJUaK5GFr2K9uuZJuEM5EQprGYYSXO
DwRffqEUVyUXwr1mYborhdzQ7isSeaOSiogsBwxlDbGEkoF0dun3K95aAQAJYIefXkKecK4WXXF8
KdZ9OLyqzoQDAIpHjvUisRu4gDLugivJ2vnwgGCCPv7TD0ZnwtXg2d9Ahd2qR5cUtBplVUbd9r2L
uv7UecLPRoimUGWJmyGwmnIgjWBxSDn+EPSnFMEqEaSsfjQbK2ijwYqMFuz9cvb2gCeK4kAeQoPt
nv/b2FeLUGoEO7IS8vCX2uHCUfzsiPQ41NPIF32a0DxU+RxpBsYtiZWvxSVOzIInijhmaQ6NXHSo
FxPsssgX40UtN2HFyhbYJxMKFNtBfLX15FG/0tZfS8/QoJmFS/AU3mODPAUeiXtayBssL+gHh9gd
OsY3CBXmgzA38mMWPz9xIGiNdWOkFB+/WFO4jCelRe7ZP8Qvp0wfo5LFJROCxwNerShCaMYf29h0
ner+HFCMgViqjVGEwMF/HpHlw48AG7tkgkFB235Y/ox6dZ4Lxm/rMFybBS2LrLH9zWMNR8ocNZDf
hKR+PBTxA9Ritn0VAbFHfAVUsMn4fkrk1jobcqdoCwG0D2HRl0mBs/Bf7kab4b8TlMFZjJBlT1Mw
rarxsS/8WMcg3LiPI+NtJBkVgCguRrvM8MTHQznLBlmcEZZ1+RouIry14zBkZY6nXeB8SH3i8wTD
DBWE7G5gAf5SiCjZQaewT0rNxeBSgqZ63Nz6hRA2N+titJlrsbM1NePx6mZ/fZOEAIUujMjsnhY8
+V2tVKjGbFkYuxyYU32rk9nLE4aIxnxijUAMczsw/cd8Or/PnujiiaS/tcxst4hYrO2dRpG5bmhB
s398/ZJSreCXSMAkmLWG/6Sx88GIcXQrkTRx/66unGhVjxosFyxhKO4gS3GdQjDVqhecIxSnSn9e
KxrcvLu39SSwIxr1xKOuccPvrgtbw6t/TaDIlavZFne4hjWRE3FZBquhkstKOXMcgCh49B6XOpOq
Aw5OzWyIt/Av3O2BsoVEHTHJyZF3zl7IgtdGdQgBsmzUppp6j2t+r3p4s5VShfIziGCUo1ZClALW
SuUsu7iGRjHQ8CIG+R8Nf3Nq9GLLC62EJfEHHZhMiQQVrD6EYY9r1nR8bwU16zJn9TbGLXxBG68Z
bW1uy9Qmj4qcXImt9T7sWbm8AxFr8tB0vRcpbbCuldGHR2JY+bYWvY1dZQ/2pVJSmuMDX5pUSgpc
vK8dWOFW4T6MGHivW8AxpE5749+u0pDj9Clb4a1CZroF4n1ZRsSVIPv3eQykQhshGonJT2yxw9a7
Ap6GfU8aGz/+KOpdMVZ6CxczvR6sZXejB9AO7axWCIsnLC4ktg8rd95b6odxJmnOpWrQEVoKNtZD
BV6hU9GytfaYNDgF//7LtFTUaZfh+m8JJb0/T0hbeBzwMZ0L5tMFe3UuVTS7HGwkDGFrgd6KCYyM
8r7eLHS+n93Gyua9zG+DrGIqdyP2pcQfz2c0xsoVHTd1eYsuYzFVWA1BhPsuSIOgMhmirafJLGL9
B0ofZjikBuC82n9UtecMcyQTKvfpH8uU9CZzosbvf1eOXv2f/lai0+6WVSd8ucggiEEwJhW6P03W
hgVmjsaCSiuuFMi+4m7L2YIT67WM+Dg+gIkVBVZF3Wd56IjXgLycAl+iRk7JsW2839lm/uwO5f3V
BJxytjjn9UB29j+4ER5j4aAAwOtRAxQAqH9aeqyDEZKF6Blzd+LRVFy4985/+Mle0V2oFf13MKrP
busvg0G76I1gtLeYGZ17N3tq49GIw0FZEkygTApg/t2SZQjoyn3T+xHlG+zzq3dCMwuI8AFKijIB
W1sT0DMuAWBBVQodzl1ELmSXSWlqhDjhqWXfYlmSn3Zq6y2MYou4SDWfMkNxQSMZLLzLTr1nkSn8
ubgVuTSqvRcpXUjc3A0gQlAj0xqW2gBywwDdYBrpBYvKcpmeU0y1hnSiaio322wxZxZhdflb3cbk
TPh1Z4iIkRWkAVOWKy4WozXxQQCvXj1idhdfty/I9KEB7QyaO9DCA53pzTebDj3AyJb3MmeyomFd
h77cXsW9VLj8ywprxXe+crzJx5yf9tc4EDhHdptfg++gocW7tbO5X+fxGJF/zDb32ZauZHpzsbzO
rMaAYvnymNDqKHJKuh2yO5zsf5CGTGkxmi2W8pnsADiLLMIT1wmQpJpkUeanQaZ0q2Ys8Bsi7WOK
m54TPHy3+iT7JtFkKlvXM+3MNWpYizXYN1oTGqGucxDI6XxCR/12YAYMUt+/8HsoQg+qTqqPTIjf
usgr7VdFiEjtNHjSNgVGoN6ww4Av9Jy6CC9sd7WhTbGIHq+BoxymYNxRDuaZayttgcIHZtxXx7/S
50vAl1SDEQ2G3lvHW6e1KwdkMvVJgUkV9S2Fu9e+r6ViaMjVQl2Scmb1lVnaGiGIO3631PQm4vtM
vtCZ4pvcRUAyBNSDWhsX9xPHRgyXozskqXNXq69xe45jnQM9onCqvL3PiAZfPBetZDCBe6ntbCLU
jlGWeKTIWpEtPYLuj+V5AUlXev4jMzb38o4dM8+syp00GO/iL273v8Vgyl1e2ds/2xr6DqWyV0N4
ug52Ir3bqIT5fVmk/DSZ3sdoMgKAB8yjQNCHbVU9S9PahRsBog297ubDEKriisIp8tiMDuC0vjcT
D5wFogFYS6knvVofbtpUlFSNjtwbyBxeNIjClSYBvBYgpe8xwVQgA1iyM1lhL8rl3685fN6Obxhg
qJY0BFeqeID8SFAf5mvqCqUaa5bGc3VnGdvudewccdIXjcJivv054AjJh+oNFEQPjrxRCMd1zLGY
l1pj8UWItzH0vWJXd+dTeIR+aJb0nxAaVqIEFFDwUAt8j65qNuz2xnhPyq7HPqDwGUeKNsxSWkrG
LCnUflLe3deNeyE52OnHFXtHooMU/h4xJ4/tKNjhIZaqi7ChDpKRIC+8XHtUV1UHG9V+hXler3fR
3mXCjSU/JUpa4dnlU+fZZzcuoFIs9hTxbdLRqA+CCINi1Tnod3otlQM+WJyllAgVmsv5RsjETnae
NLyciyMZ0a20hyS6a0Rfi23HKSVVZFy9qYAmVrSfvIR0T+9ywFTT7b41rMFPFPXvrXvSPJQugSzY
vX4G6tDmaGcmoSMtgKT3kf/7r9mutXOKLV80kRJgc1mfQvYfXYEDM7kn8/Dw2slIT2Q3AIvoP6/8
I44BBb6W4ua+ZUx4jYcJuYnzfQHAg7FiF8FX+GDSjuKgyGlvnNQCbii1RVm+EocptKsJzVNQAEDM
h9BISO+qI4+47COlwO6xlI5rBGh7A/hQk2Ye5xSFohSkg+L3aWgupFefs8pvbRaN6h+8ZAkjgheQ
OV0pV1fLuQf44AfSzf2pzBY7gshsSJG/q5FZN3km4nyPdkDKHhXPDOQwlNgy1co1eFlgUO/XDa/j
rEXzS3Bbsoo3OHTMY57tok8kGzNvjVjw6mi24keq0iwPsRTWj8qWg2C3qh5FdQWQLAg5xDY1q7PW
EvcCLXS5JdSAlb6KtHdXz20p4KsRxEaOnhrCfK2T2+qV7j1tN7+tDXtZDfgGPggcw9lXBlGXh5kL
zrjnLoXgDIWNWrLA/ZHbWKmsAkAJMmvwwYOv5Hg5fgXs0Fj6Jf3rPi4IuZFzrbyDnFXV5X41DGCb
4wE9lS7qJHhbA94DZpPz9bDM81ZLEHvKIetcbniM0D7nHjdIpGdYnj4ZDbIb9IjVBhL+rCaBvnr/
TD7fz6vEbyxHf512U/gtWN+Kx/YGiMYOUMlaxEuOUMv+fYLteB3OlHsfsHX9dc3v+84S6VDKWVbo
gLH2uHVfMQDjJXrzFVPtQAOvMGDR3daK+PMQYu1rfv70slHvi8h1f/Xu2iG+C2zk86ie7dPmKwKp
KPpnYBtDmNuO8uIhM3RRbTJPsVfJv1EQb+5PP7mYR4RKfs6Ap/V2q55FYfBJ2Bmo0nfwcipEGhiY
QsyHfLT49cpfwjuUNjAV/H7IEfyEfHeh2jyIAUOE1f9GYrUS2E/v0CZ8Ofn4+txeOL+6uulWfTGG
/sUBoNL6CdVOSH3Qh9SmQo0MaF3i8WzZ14rqBwRQX28huzyOMLudyzmTID5ZH1nY4ktj3PWBGvyl
YH3Y6earMBhJpkpmIQeE3Zp4Xjo0dO/L7PrjqTFZQYsWZ0iTHSioEBZzapyLdOWmyXstcA4yWIgN
Dkns3qKlYcqBwDJ4FqURG7GBXKTQQpTURz2eHOmFV1PAwPpSq0J90i6fOGT+ZW8u2drYaGlGLd2k
h5aJ0c2Gfi4zKn0NLay3hyBgKklsHjMDkupxXJVs33hrWtVeLzhb0dFkmQ72y7UjgsgpDxMT+d2W
DyecZoyHGvl85C5NYEYBYMyDaM70B1JgDBsW8SveKz0pSk1I7EmmM+K9rhd26Bh7QVjiCC0Q6A1l
ttKzYRDAWhYmKdcrgT087wg+Yi4g3Se/yQaqQMTGTACwYPURtIDEzqqgP4Oi88hiRHHHJDyC00uL
oDipuCriRoeCJEQfG2Y86Z2BZCSh8l0W8OxIF2olaTiSisARQoVL/7Icco3wVkkmSoxN9Pq9mbuc
2Fgj795h/ptWMwY8CDZta1sLtXNEIJx5ve2MbPKaxRk7k/6Rg7cJeEmmtWwYK4hmD+gOcWrQpbtl
nw512qb/F+3xH3EShXHpVQEWQQBz0QJjXMlQ+aWju9TYHSvobhA+ZjacCeFJl4RWYy0mI4t50Q5S
ztQ7/2yKoqZjCPY31Q/p/cb5xda3d9Ihh2zospUQO1j5BWvTKoE5vogEd/JUHvZ8Jc9LwKMKL6Z8
iRaDuev09aJPubcP5dq7ir/Xma7HCKe9EM3AFdrjXieqeygcCSu7qD4F4zjipFbl1BGSgPDb/Bj4
n0gOwhbzzdNZQ0L84Fy9VsHVFBngN4VWmaNeQyz1gf+r+9Cl1K+5gZckWnwwrhLqGefZ2Z4lUGM7
phazLwU+15FL9+800Vqyw+/CbYGENzNlb6AtiH9PQZV7/JF+7uBM4glvcGkwQbtCvSfcQF2IY5rK
0V8MPhDhPdtevU9vBTaNLjZsNgp8ROOrDbt1n9UC7001mDpEtcWgKsMX0wk5+44fU+4M99FOPScc
0IYQZWEOODO5V3r704LXxTkXuMQI0LHHTMnaAjq5GghfvbxFVP/WS40tKriAjt/Y+l2vLltzQPK6
DIwhz92Yfj7vfKA/+3OXo9oVoBBHAowS6P8KepZGLsywijZN2EbzIK4DNb3LuMuK5RbLxuj/EOqU
tTkqyKZq/FxJuSjC1Ra2hl9AHQKTArBNXOMVbiB0YPskGc4RVjzVbTFlyB3EzXhsJr2KSm4dNQTC
78wx/Mc5fPsOZME/olV3zAKko+GiDLetlLzRAjdkbt7OtPvsaphO+kO5Go0wv4vU4s0C6AVxTrQj
SnQKe/bSWaJNmU91sV9uH/xlHR2AjvV8if+2qdDMLZUEk14pAMXVm46wakYe6MFTfAAJ4+NFDD+E
tR0F53h+fqk9+aTYzJMWmNTmL773vkxj9FOSApyQPmdJbxT2cLq8LOEcDS+fmE5j8hm0AcsoxXsE
SvhHEi0wXN3c6/ehqEGe77JUhU+htl1xelQRYShSyJlcoGtfUIvMq8B0+6YMhJpj7wpApPgyQ5YO
BMTb1odyMFU3e/uWhN/xuu4dzKJjkcroWezqz5aIQgxV5JtETQpHXkLgs+o3IN3yNnYy8aViNVTV
OHuVqhb7wXPRQ1/ePC6vRcTW6M7DFzwd1k5fy1N2KXQb49WNazEfwGKXR9mMho+y8NQRKttmK3bY
pmTDtxgg6RBzRaKfIdgmzGy9w8drBDOfgyMRIsmXG9JyyxFzfq/NMAPKWXs4LZ/5JwM8koKQVPCO
6aylrwGtBPY3KWRWjeiy5gxeVJsAQyenFHY7+EAT5Kp7C5gpV9DsKfizFhiIBeTpStSgG//6ZLkU
UVH03YpFWCD9Mmxi04QUJ/lr/1v2Z66qEZ7oEp7EuArLWEYGKSlQzd59czuEbzW3MbOsu0Cw93Rk
0b2LMfJuTDEg+LfVgjanwO8YDojV4s2lWGLihiRhkdr4vLIGJBrPZbx7ftWTVm3AkJSdkr5jZeNw
dubV1gIDlUWow4v25BBs85wbOtwXouUkxnxLkXi3auRoeM+YZ7Vfo7wv+HqP5VV4THKRZT4IB9/V
Qo8+KrZhzNoJg7NWe0Sc3+BKh9aXBTLZbXCp4UH857wWy4oH+De4P8MXWaJOMyiWd/CDQyvMWmLi
Cv7y5A0oE/tEbXCONiCHAKN20oWP8OqJ7xyy7ZeevS3kvihfJxBC+EaDigwmrRXYM3EMRf8RODxp
cS6k5HVBtNXUtvD3Ji3LDmXWOvYPOEzC97x962nUBab3kdVC7DpQBBzvulRdS3k1dQPZX77E1aD/
s3ZO3os/z9GYgAry8smPbmOQI1Kc+el9bsrwvoPIAGs55eicCBynuC4mS0/SIYkX/LNuxiHoRW8z
evcM1wqR6CWNCycIfBdpzA4kFF8GCrDM6S4NjAiKA/74xzIGfpQYVzPmE24JlVEo1N3PhOdOhzao
7uuErGSKKmcpDyxUSNkw9vMqdUttPbxEWSJ7qNYbM5PHOs5cUIDRThWOSlUZamuP5Y1gDO/47Jji
lVfzWXvv8LXivGV9z+nXVkqNM2nTG0KuzwhuQZkdthVkJbcjrq42LnsfmnhoOki9w8rexbZyn2ZH
2GCRM4qA2Zm5V34pEpTCQsU0GGFvy60POCQ4SM1ru9KGeMQNHZjGtqUOiC5xszlDUNhWO2s0LAhS
twjfRJdLrzoj958l9ZuWbNlVMOjhLjfWbWqvjwyBeQcSIHz3IburhxeZv8O8ieoA8uf1O3bI2Z2n
1VI2fQPXaQsprUiVuKUvVECrc8m/XQYARKG5FQYCjEmmuAcQ0qmYT3BCnx4JOIgwbeG1hmjX188G
WiPKR4bC8biyexAA1suEpBQRTec/HNjeVamdYxyRS8UYdsRSNcnpfJNMUbFsjQ8IUjpreOBdr1ly
L4khP5wjvlQGyFOLFy6Xnnza4zbTY/6HofLuBc2QS0vSBUD38fKDK0oK1JU2paPe6hAjviL3qsFN
5pCS3QaXusIN4vmmfzkVQ10T33CT+Aa+nPvzNmlMNjMNAHFp/6Twa8tygOqiFaErns1j4p3me+8j
bZvS/qpJcmJTudITMiyXpG03ZhMKVZ23xXizWJP2ibFRZ9iC84soimoaVsup4UKZUwV2PkjGFU26
wy6NcMCnlKGP7FFcY/7OtimdG0mSy8mJVqLvdcICTA+cqMpb5TFTRPqxnex4oCnbsVer58LCJ+Pd
dKLrYp2SfbWJ0R+MeVWaSXLAS5Ribglx2C3qh4017pKWMoKmSZAqnMYIhGFlGSuOugRdMdONZnXu
1OSAzTNFGTHMiVVWshNnVEIGFknDF8nKp4jvfnxCuzKGhF1/UDY0LE1su3FCak6pnit2pZOfZ+BX
n4DJ2kYnHU9A18TWI0J26cZAqntKWsgkAdaGtOuyH+Lv47YzJ0ypYO8khti2QRqW3bWU1uhyu7fd
EFSnfTyxvRUOtbTFd4mimrg+9uZrfrXb40lgvTEogy49zOL6ZtNKk5X76+5Xm7zNk3iqCGz3Ct7E
16bZBGVTMsO0MOzD0uQmqL934CHOm/z43xqHg3QjlMJBXHjVcJo/7WPoJfxDIlLJYWp7b6uv6dPL
mDNWJfxcE4UAx3fmE6wi2dx95gPvIToaSvuYo80nb5fbbn3Jbeou+WBNLn40CF9oQIFFDOdoiQq9
Q+7+YIqCejy6aK+nCB0MxIShA+tiWNSQibc8isJrROgmzVjDqt7yXN2vKYDYqzZMghtWP59gEVaA
2nvuru0UaVq4pdT3GWx1xKvNI6PcfDuNruQq5uyXK1SPZ7iDp2qzckLKMV+qmWSibg1hQchPh/gL
JdELmrxJ+MZdhWQsNK+7Qh5Pt0vNIaPmmNmPoUMcJTA5+yJB7JHXX9oAwB3nW0EsIgUkOUYD+nq4
2LJqjsF0hLR1EUf9acXNNqgyHKlnn0vCPVBeZ3FZPYHxUMrOWV6USkqhO5OYKijvPCIEt3NiqKq+
QTYNGmJRcoDisdAey++scZK2hv1x4Y6sd4At954MxleMDJSF5oSaVzYTzLxjKf329wYblF3bEP1O
ufFChf0+bQTHeehTbT8ItBRXCvlmGU/iT8ZPgXgVxatUTvwzB/QZvXtmBVT94f4CyHZmHV+df6KA
oRgnKnA5mSWQUZccaDwc4w72IepOVYPdYOrKSlvqKkFW/gnXM7eBDH+Zn4NBV6ElkLIUm9lKv58W
XFThHEXoIDSUHs+YR6KNcTM3lEQmJXdGPZJDW7u8PIPF8WYn4nbNLyjYrR1WoFP0uB1532Q746ZZ
Vm8jWSoTjLqiIf2LD+0qo5gYzkKMclqxf5dUARWDE4rvQuLjCt8J8nVVOelacE4czcK/FA/SmSzn
SXrjhbmtIeNxmn0ftplHVPCHZxgy1jgFCCordKg11OTSxW0uSXP8EFTKjmKJiwlTPkBmskR7nYBY
cjvvS9pAcg3TV5D1zWOlhx3JMWr4wRkhDovGRrTx2D7wnpqhNNb1GQigXd9g1ReTcNg0kM6r8Tsy
33oPGk4NCWAKuznUAyxKjzgL/f8NiHWccgVym9CBn69NXDWVCtJVqyB3mpVUexVtQ2JvreE/jrav
cw4sRcWAnNJGtKyAr9Pz6nfGtalcV4AGNvrxxl5lQSZpV/38rOkgXi2+BuePTsvncXyWVRRUsSlR
eU6bS9W7pyKa2JByLA78235t03fNskWZyoG+An4Ia25finv7NPSTAgCQXmVKcjWIZgnsEtbdJdo6
ZirIFagS20rDcZo4fjtrpOZzBdGkvwHvJLSIiwBcUjuPwYN6G2qpMkgtSeNexIt0zwsZLwW5bTZf
+4E7tSaYmaOLsK4r8VOuno+XnyKbiViEy7VQ0mG7JrvfU0pCMaVkDe7qpFMRP14aWm2Algpibbdt
DTehPYq9GAZFQeEjZonWe5qgRYCLSuM3Q9OSfa+X8tej7C7PRLkfaEgWQb1O//Xn+MRJGl1SB+xw
Hp2UJ5uG0els7m95TgAWOekP58JBcrmUYgKOjhXsd/sd8/LbBxKaZ2OQ9JFhBVH0YViyYEWydnng
BSRVqebm5If+qngfKurRgPHb0JiCipuoO3YVyQbaLCDb+GOxOJIPdwzHa5XKW4VKKg4V8Uf32fJW
a2assrYu62fjNJ45e6w+vc0QE6ApmEGgb1nHbclK3o5qeiAUKGIRqTRxTT7PeGSdaAENt5n/qzCm
Bfv0WQ4pvBEIo1zpZtFL0ncOpw0ojp1z8KBuUb6pHAC8Xr9wAX/QMSm09/2dQauztNqEYlmYpJVV
25Yi69Gcc0VipKB8ZtKUZpvhjzEDFUZOeQvuzNpWNy2mcv91Cfej+osU2h4JiQNUlEnWu+VA6b05
RP4sN8ujJg/PxVP7mwUTh/UU3yXAqrLelaTAA3rAFNgIBYWmTe/HDpaYdYxOVBeNw6S3B9qzLD2e
wbjykziPTn+/o7GvQupCz5Jo7jjmhmsq0MnNdBp3UKS7kwRCUhcNeHBc3CYSWSbeKNSuJ/8OUfgK
TmVGDrpmv3J848JiEKPebZmreR53EDs9ut/crlCgrQipRTL2b694hb4DVYkU3hsgY9zj5KtcER0i
2JFIBz3fsOBXth8S7D2aRM5MHJqGQ6dahMD0OXlYTMkOPA1W2tNZRgPqP/KOfar9fdVUn7oTkeNo
DaAfBBh55nnp3cYW8avMEJQQwwQUZDqQUXJEZpnHlgTttSHrNa3a7XtYIjojRfFWMxhxkKaraec4
1JGl51sUEn70fcSfJSilucp0rx7mY+Ehm7iUvqesSqjWoAu/g5HMn7wUYv2+6OfzJLND5q0apivo
mAraFTtOfNokKBBykni0Yl8n66oTBr9zxpTU1kGJemDXYHap5yzQQBCEKAi1X4oF24lPIHwDZeIY
lSOWklMegxYUEiCZkcTSl5LyUSVnPYCgS2/oQk+t9TaRa+echHDmHntOLbq6n2nU5ibZdE5A+PYF
Cqsi7YbYI5bRiAkI2e2o3lU0iBSyyNO/2teqYdIZqqbxbVTJoRmLmNBrmy1ne7xp+c7uvFbkzjwm
kyrWnb3bZ+5S6C3BJdJeb2ysLzbqVj6r6m+lI0dHyvFZxRL/e3sqlq3AsiZ0EyA/+2wd4SosVthB
xWm3SLnI2loLzh6BMizbOMO5U4c1IFQy9JhgPayaqyLWvM96nR2AHR8heyuHeAvY1XVgTTShzMIh
nqJx7AImQtUXtZx1SKtqleK/JKuZ5YPSwZiVtlk+d9VwTVp+c6dwzkZe+rwbtcS2uJo5lHPe0Tw2
2LHBXN8/TRB1V7hlDqyEXP3QEkPg9u+ZQkxzggZvEPl0l0owa11xvpBLGuJWyAJZlersrUFvHMeb
S+s3khRrOKDT8SMSd3vqA3eQ3iqo6W8JmBzED373pjXpCNXqIQISw9j32mOEgYp0Q0IvHLJjwEgV
ij2Qka8mhmPsIhc/AYHlknqRcmTu36cab+RXpx2swE0ed2/eeHSd9J4bRQCqmoq+tlAGmNAXrYVk
y6vVeXgCNZ2In6/SoKY7dgMPRuSMRHDrdKO+bRlLYdLivT61PAA4qFt29iOfN4PLDXCHoeGzvSUq
fekXEszh78gylnJ4M1ernRgkX0+nNaEW0BCmqRYe20gI1JdPKdj2E2hpQPyOU/NRZYnoVJoH0WFH
xlXJ3MxL0ZxagsMV+fWPEc0Z3Ure9VxiXGtr78gBIy9jtyEP3HHt/8gJ8nDPFHHW1c1TeIWSkI/n
sBtXbGM5FwyqJ+q3aI4hpNohCTNShktgNuPjgPkBv98dWw8ano3pQX6YUVp+w12ktIoK71i9pSeL
l+6qLdQtGoRCROU7lo7cFqXskHRNB72SV5mHrnSDXs4xnhaJh3z75Fo9RxbM9DKYmUh/Q0Zt+PmK
oqrhLcb/6UUBC6wFmesPOKOD78Kl02A97ecz8b1MeBeIwfu7YFHCr2lnF4OO0BSvulNbEJzgNuZ7
+O/s+sb0/V+2UQYCmX9rgNnA5bZNXVrNgQE6QmpASzUz9wrugICRP7xoNSS5fM/bFkHEeCI3oCTq
arvsLv7l1LgwiUjg19jx75jNheZmdOnaeWc5Gi2FrTsCh/BqvZdB/sATtPuVESb1ny7cZG8ZMdwl
vfl6/4KtzngXNPeSGa/PI40qaawASeJ3r3aFOUpyZQ8Xm0oEiDOVVWK6Ni76jvH3QMS0BvGgTCt4
w1iI7MFdjJY9PlBDz36qOIIIRLdKOqSXAo0jbvgh4c+LR5Py5c/o0YSdm3BkuNSevcZvIlSYBiqX
yRBgvB/OmSSdWWzZCroUw1IK34iuPrCwsT0NxAKM+eemHBMMj9bK4kNkPk9nQ76bf5u3Xy4C9c+I
5HNmXCFjaFeTGIH651IOFCmXsyJ4q3d27NrTjqDg14t1bJ42Hh+l7EmvRZ8DQFQO20kfLChtcsu4
T5l6i09ZI7iuzINuYU5JpuJYjlw6T1lURiojQWi7+h+9XI5P9zF2vaKhgbSIF2+bEqFc2dztjxz2
gL0ZuzWM85jsXdck719Hyfol78MdekzLyyPULTGM3Bqa46qpCZtgWK9TUWkedvNAUijoSZoKXhNn
M9xn1kuqQW2SgazqoPvhpcpK0eEqw3TJ+g0XU6jupOyScfdBFb/PsP1a3rgfy1GFgezlAnjnlk+C
F5GWEWvrXjzWvc0zquS6dMDGUQRYf1SSbmlJl4q5hcOuYGtGNb9YoUwfaB505hEHMQSkJqfsnMBH
hyUzSEOGnUhFLt2ZLlsrqbPN7htmRdIPx0Uz9xCyMl3nI4A3PSymtRMvyZM8sYZTGLrybrLLxJil
SWINvo2xYpTrAzXYekzJ5J19bJEyDGwTk/IoKF3UMPYw4l1DKKNGIeGYosk10bgnw7QWtDSisu+2
xJv3UdGCk25MfYiCbX9Gv/L6Lb9EnvziIXpdd01OIfYCZm03ZnS8aV2yg8KU/07e0hCaX16nlPXH
+ENlfmrzEnIQo85/4R+tG838vKt/DpjcKKjjZjW6GTnGozx6eyyELblMLYC2hyJOHk/YQFtr9v/A
ReCzbvPGga3CiRbCU/wyxiTv6hIp4IOYlXA0z9W9I373YOYWddd11rOKgZ8c6kiGBx2Dilul+bs0
xN42Srp2Ywn5oqGhQfdPSOYR2FcjVEOY7iYk+6oJY5wWxll10CflFd3+iIANYDdklXJFfLj6ihAL
BsExgEnE3vKXgVqZCGYlRE8QkhU4CWg799mBDa6cWnIsFtxcAxMK6n/BIm+Sa7ngqll+elJi9mSR
ORMhE1+Ikxu+ijjLe0qXP47Q1s87b2L6wpt3hgXkZbPBZsNIsnM8DZTMFyN3OcQ3WTIRzhWhghy4
7s+IddMoG+aJzlA4BGoZu+Pjqco6XWOk9ECKwN2AXfi3zPiWGgmoXfSH2CZC4sMfEgbAme0DpL11
tq8uvwOuKMZDgjJegwy2FaC84TmBrbMn3EHirGodCqh4SKXR9Jvby8vd+c04TgEh10nrwijiEni+
076aNpsWk2xhlFYaQF2kIXFvD/oPWDhWfV+U2T+6fF2q2Ohqp3juecU0OCM4RbpbT/chGtBEp7Bw
Xw3NQO1XG1ZT8+UGIA8bWUewvd97djUFqdmt9ygWLqa7U4LMyJVmpOKfdLoxqmLaNrgj1p0/vQuI
Xl8Nzd+MxlLxFpW0kDsl6vDkjd2PYPx5Foi5VIFkHCC0kIbkzVJLLMTT6ruCYTVqEaTqXCO7omiI
PeCjm9Wsomg1Omf2nhhVLq1X17KB7PjQ/3rSn1tIaFdJSWxCEbNZZFXLLI3WyslerBSLokeF1S5f
NC5wA3cWTx8gGMCL03+kZnrYLg8ttN4zLtJfH2+XyxzKofCeeBa9Iov2ZdeWlGzI5dZd5uFEYgeI
ro6leVua3idiAw0e8GW1EiPGIsaThV1nNJQIZgUTDlp5XTn9BIlW5dFyUdi5qzu90bYRDLB3ZaxV
d9xgrg3llWpS7jvq7ivw93P5cVCzKHWaCvCHLWev5oGppL6NMqXid4hPWGyMv81xrr88f6r9WFs+
hwL1bqSfKt6rS6kqnilQF52aeCAJlZvm8CsSq81Adw7cSSbCI/yrLjlC+H7fVJLxJK7WGD8H3znL
zhWQF/UKx5Vlq1fYdTolMjGWhFlA04f/ty23O5PoR74mAd7ep5LlA0BclR8puK2Do61TV6R7SPNy
P575a5v9DjAWN4xWGWIpereOFcNy2aR51I+FX5rAEuVgrj6BWJy7e3uIGk7EFXYKV7G4sCHYg73S
teS4cJtJ71i28bLI4S43I88pLk1gxJPcnaI/Vx/sjclvgxtXgolFu2qi3hWIziUq/0ZQCoO8zmfG
SNWV1vilTvJ8x2vrgCoNkQOWr2PBJh/mSH2bdxVP6Zfhc6V0vL2QBU1uXvBKR6LfiNPZEmQ+5Thr
deFgBFEj6XKwfUXyTJXR2WJ9Ncbi+GUaEo8XUKRdQnamjStKeqj8ZqWdDUVC676jXbnDBzzybaaG
InCiKpweRcMF+RekRrZcKSXOd6Rlavwc4KM2P6DN0xnYSzZ8z45eX2bNtAKmxnMu0M2noQ5AtoxZ
t3M/XC67VQi7HOcU1Oda13Vm/P1jGLy1ERuKT7LPP+P2dIjITEqU7rQESt9nHCZyhkBHZ1vilMPh
ewTJXDV7Ji4iS0TA2+8YhjRCePeMzeuuku8cXlSt4u5UTL7++WQMEjjYzDgD/d68uLhdbiTxYVXE
Pckn/+cGbCi7ZAOvkIdm2NdLpVyL+T96beH0IdIyXj8iwQNNqJQYEzMCEUZHFORkOwu0xZbswFLE
i0QBeindsJ5TPYwUguya8pXS+C0yas3BlFUGWf/CGNeQllHZVZ7829pG7GG42f+jngCs0TsNLGFU
Y7gmY1Sfun1EuvSAt5+2u/RIWWLSELmjzIOSLsn1Mq5Hndgop/bIUP71Dya85D5BLyZOJPuMjgda
OJbQhjnruqqnKHrpK+TTndvtRsb62561Z790ITfEYNroNjti1NkrvHGnauwdkX04GGgeGLXuhhwx
lWLc4nWlqo2OZYmf8W4kCuRtT3atydwVC7hhzxwA/ZMzqmxO8/XvkJJoU/r+4GpzlRqGn0kKaHx9
3SJK1B8SXKH7070SmgwYSu5FCiCy+znYwqwGIrBM7AZp1DhzBU9CYOsVihFL/g81FEXN/RcLDCwr
EaT1e29yNZGY+zqu18ms0lJQEGULDn5MniDDRa31ObqBD3bu+95rdM1WZozmM11/8L13wa6zCt/j
zjOVJqySyGWuPgKN5QvG2vV9835vX58dSHi49Oz7GGnL8lKi5Dx9e6CaE0EAPYibNCcXjGo9kI35
JZf3D/rkAEfzlVVXqVORcW7HqcA3gY6xIpuaGMBlCWfeSTyKuv/x1SSROp3bTg4mBwlokUXfaytq
CNOCPhP3Sj7CLG2U5wl1c2hA1U+olG7iFikGOUg7kxbdq/wgk0r8Xt9q1HZFJlMxE31X4NGKACLn
B7VvTkq07nCL8etMHLoWE00VtI8fqis6aDKRl6Gme4JOVSjeAT+TzNbbCHMAU2HAgiFs3KeXcj8o
cPuyFrszrTJEcDSrNpAzqiAY5B3eWxuOayEnrIcjy9G6Qf/CorAsx5mZs0kz4AZM0cXNoq+BN+wa
U5TewnSnRM3PcpfaMr/8IDOvyPvbDFQpE+uBc70x/PEIk8p2lJJn0y0z8y72UwaXbWn79nvaVpMW
oId02M2+w9AbeGgqq4y1Bbt/CPl+qRUJg1Qw3mzVPMyE1mMVGv/jDBQC7MtNEgymqp0q67kCfs7B
oEXnYoMIX/Qml1Sd4hfUvspGH8vGnEogNVE15500eSynUPcWwJQWME0uCqPSrT0Tf9nDcCX6GqKw
iGwpOb2Gr2fFzs1IoVftuytTs1WAyoX/paJVe16AbZWRn9whwW8ql7xUPrroqzIyUdGx0+b1HMuO
b98azu9KT7ctlnXVx3yAJHchOW72L/KvDIgSgwuxwvcVk6CCobkRAx3d6d80aYUsJoGzt+cbQl5k
0+bb4SIH50XS7UXP23eEIiBRNLTHtVAGGbSfBHoyud92RB0ODPDQI26EjMcDd2fa5tIn/d9mIt2y
t++AhPXMsLjsL9LM00bo+D2sS2YvthUo4+zA7Y1hoknokmWBYgQwK6n9G4NjovMve94v8z53qbUT
kB4abdbVaFxR0V6GB1bXQ65Wna//Ia8seTGLfgENdRwYu8IvuE2/fV1a2drO1Y4gyt39bXETEWXY
5VA78ubdV15h2FPwES1EU/RIf2B2p8+FVsuSD9B9kPIq3d2/uS2jnHBvO1/8G6XCWYHwEELS3McG
J/yubMfUi2rN/thmWzrHShDtXq2rDhsDdC4ydM84ZaWw11WJQakiBwm5dKPZaYQJuHgdoZ00bpVF
vhggn4VqSoy1s+c4DMrpkZ1uCGgZhHa/m/rxSl0TpJDDYuY+2PUZBiLeYkuYVEconDcfPIxKj2K9
jrchhodm/uFTzvGCITEgmfnDIvBVMjXMsFyfpl9vcgd4U8Rp7SPnzjngM1gTXPaPIQsY1Plc7CHD
+PhjWqDZjBPQ1H7+q2tdHnlDkPiBWUFPVZokCAs66qlSMmXvPX6cWbJa7B9z+XKlzUEcAFwJznbz
HMKLvucROVOnLYcOM6g69JAPMQ8OMLxAR8+CBmVrB8e1DxeZYfIbXUF950TBjTjio6xOreUaCkZR
nu5TowZfmgh/dPYnom34/MD2iDkANb4xgiUIW7kRDkweA0U3yGukrHvL0GSF1bIO6wGXiVYjCSsU
uoaPCPHM5U/7JGFP2vmFsqKhN3Vk56pquLPjSEYXUTck6SPHTldaqjufFkVMbjhXMBkyzoPDFOLu
c6goO8laQopnr2g1Bp2N4m21/FpXmjg+CWX50sbCb1XFlmWCfzYogQMypX8wBsWdH3J+ySFm8F8n
/uaswWTs4kj8/pUscsYZ93NRqjLKdvckjNbalh1uYuRaYCsde7pO0b0grwcW/qy2s/7wxIPy7ivY
JFR8eMQgCtO0ampTPthMys7vyJAcIaTo3TBWkXcjb5BDJWRqEPYely/AIsQmA46hcQfOBkTFWGRr
vu8XxcpPDiigd+WwQhWfsyJUsD8iwnZGqYPCSdvYHqpMMClzr/POMDvb7mIqkA7TREaK6501g/tU
4540+YM/MZ/KKxnrNtNr9gOfTzcHPxmfZtKkTrivSLpS/IunLWYhOaOfNQTqChcisRTWGXIwS3k9
K36afZ30gOcD9mkjincNoIGUMd5KwC3iHVNaJDFUZjDlImg+IoGrlT2G94xesQDzZeSVIaRcOV66
JqIvXZVAxYri6KKok99naXC5l6q4T7oMdzIMEjMySm/RlwWMPtoY6xSvliqJVBZnJ3L6aQ5TEF5/
hod8T5/rOtD4WTZMkE3og9K5temm1D98eEmSwKQZll3aRmFo/oLLYfWjLy+aTrt5aPz3D3u7d6B4
J9YVSzXWXXyxdTDaE2uK/FFfhNODKrv50+JQAhUvbZM/4PrhjuhjwvZhSKRcjuy6b6mDlGEb91bF
zJR4eeB9rTtqQDfGWM+1GJ1h0/ia05SaEPN+GnoWeGowl2cGbhsQaplf8oGeOg5wDgQBGLnSvYaM
9bkY27ZAx9U204QDGECJ1gxuz1yRUVGE4O8NSLl7asnSBpdzniiUYkSYbSyBka6vpAd00uxYomV+
sJTGZK/AqPcK52McsziIYkHR1l7dfBRswbNZe9mxeOKCCX151ylhYNDbOQrFSIZp7tgkPCwR0B64
agZrifT73sLlJWWcZNJxcHQVoPkPzLqyW91slJx9txp74nk8+9qfRsukJHu/+XWS77NcFYziYjxf
k6FBRnahf4rwJt+rjmPMFdvRwXOEsn1NXLfoxUt4QKqt05oBNpHg5W5jKDL+fGN/PA5yt7B9bRf2
hcEqmYH6mO0dxeyWp5lwI3hOdf619pUK/97NUbeZflU3bxf2gbELGH9zFshSSm2/8EA5N757si1f
tIA0RSSsNSgSlAaBv9m4fDk0CkWc28hSUbLg81I+hvv3owMywB04mjvLCNNgx9ykSDNROjCF0xw+
hOXzn7hD5Ed79YAc5Z0I37BOYqKynzq1EAQngyHzNovlsgsowsB92y63QKv4uGBQqz1y0DZTIR87
AK5+wfAF75TQnvqlNKXWi9ZaY9Qa3TSVQVEehWVleOh4C7Nx6mSUkzdSvXbVbnEv8BxdT6doNpnx
sIzfs9KstnIXicVoQp2OPCqPakXUtm72o4tr76NeRqT3YkSJ2XjGotVN+rr54lPA9N7UCG3HOfKj
QQwNFMF8EHHVwnezzZG82vwizACFdTm8R/sgZfSwzrAhVeL4L0H6XjIQ0VxPV0hINhOjfr4U1Pcw
Jy8iD8POMF2nHongjmkLzg6xjNg1AeYXRg/cvEpj0YCKN5OCCVn1zZ/4G/bsSDyvHbcuWLPNYCNE
uLlmbZwj0qLqvVY2G1UXlDd/HlkBa18JGH7C5R/CpF9rHmgaVn0zcO723ArV9+lLDd+MUCXNMxAq
EQbwbqTZXsSbnQ/zJmG1mcFhXsfRPqfV2p4BpOi+74dPC5pGlEiGX7eQqR5+eNZhUh+nWfre+Jgy
mF0E+sF/k8SietMIeiY0653yXZnF1Z1bqhDUCnXad0uj4Puy2BAtC0ucWL+gFfJM6SVkG9hBK8uM
R9ZAPYf3EawNLV8dzDzcFQLAucA14ma60OgfKrhXbfCV0LABA7yOKU/4UusyHa2pdqJbcJF1wvpa
AbEIPoPNi6BDV15RRwo+/J/39VZNZZkNeVRyvAmsi08I7xK8YRKaoU0IQauuEBSXj9vJr0KRpvrh
HDz9u2eabY4TtojvjTso6RgkVi1owTVl/B661+5li4i06RHIMeNHIgVB9tPXXiIh1OxNBWonkwUR
N1HiWs9sEfR8cd+5lt4aDKp2Gf6xLWy0AF9dnz23cmvBm9ImraD1i9x5xwI1PMZZaXuOsj2myklB
dQNMS1Cmkp+ypapQHGaytSqmVku1Un8oe044ovKJ0Pl+ZuvMUG8IDxDgbwpNBUMCKoPhLxRQmgu2
PKBoOJMCDfcxwMAZUcAh3eMmxeGHsYGZ7qMbhpNCHaIvdz3tsTD+iXKFDK9fThnSK0j/bAJa1L0O
f7exMv7KGncVbN9tJjExw/SrtpUVixuHveQ6VwfUOLB4ujVhRu/C5l/FIZbHrSCFcPXicY0rdD+i
lMx+RH4tnnhvC74zinExuOnfljPwltXjsIBXEO+uSxH2uuniJpVAoXerokZpwiuHcS+7r9Shooxj
eE2T9Azhta3DI+t0syxm2YeAwbZvuwSmTuzQ6V40KvhbxpGUPcKnAzCCf2DxDAkFhrLNF8AHbB/7
zo27dGEzIcS5LdUVvZdgXxUHR4lvdJtAdCDY61dy/XEu8ll4xT2qTvLGq5JoqUPuQ5EzNGcddWIf
wirOBYi4WxD5K220m1MonL6hWQ8urs+yMEvSkNQorNdDrcZSXcNhrXSnCmW4/46J20e4516xKpVw
pALxKd6XdbY3WwMA05zuqRAdL6Wkg14DhY2u8jOr5k4+GfaYBiRQvvlSljToGblXaJNVhoXMHqZE
quTMY9QZSF/ndPO6gNjBJToTZq0oGT3nIG3OQGvkuWpoO7/V8DQ0Fu8a5VjZ5G1S2cTR6kSB4izg
FWdXNZcbEB4c2T6HhA/h60TledBXinWwfnUper5+wcNbvsTYDO3Lc2RrZrjZSuLdEjN8JTtZPzWU
/uPgn8PB+mjiqZkWHE+AmGEC2+oIOdA5bXSHRoM94lbiiXS3wb6VBIn2Bj5TJQP1dzYc5n//jo24
uqxovl2FExP5ZbqGYGT43F4q/DF3i37t0YubSANXHPMk5W3/NcerkC74I7swy2NvYlAjWtVvh0nZ
Rqq+XyzrCk24atzoTnIjJSLN0JFKY9MjhaOKN60DGSjPBjhMx+f2ixQkHMyP7UzKI770R6OWY0O2
UmPWYX87Fyn2XeHMMOQZKK43M+3d24Jk/zbO62w5tGM06jGkV8ofrbeDyecn1XCe/e7oahbBFdeF
rufJ0lm3q+zJtZCgTRRl/a4FVK0aSm2fvheeAYGlL6rbcUP2zzT9w31n3Qhe8t9tDq5mN7YpIBvS
Ql8+51PslsWo3C7quKbAJivnzaQi16aRCA9c38jHomQDUgCZxGx5QmmYAjY6XADlqFIK5RSx2nbW
I4wk2zuu12shrDoIt9YmhtvOzfKYJ/RzmcK5ZWrMOrItWNTRpRcFa4nZdpo6fQkJJzmz927pa9PN
E0GibLIqsRML36stg8dLW7d3wjlxKPmm0BjvdMoI1jjxqSYGzXIfToryfoOm549XrNdNWl7bF+4b
qefIBVPh/iFtWf3luADcOw2H7IqWKLkA7qrFpOGwm7P95RMNz6Gn33St28YgIiBbpVNMxW/zxMPA
XQWeviEFSq3YibpzylVFz1z5JjuJ5+BLH1AZ5cmRQ1pGJjK0VY30p6LRsn3vNxuuchbqUvWLnJ/Z
uL994DqXqHxhRaVvY0+XeGWiuP6aC4D8s1dPTNOPRRpkZ9F3e35wZiFUwzHg+5K7luuCDrWs2xwF
A3zkeVHUjjt7MnaiMgmYiD7mbPuAOI4Mlww8PGKxSARBYt/4H3lWYpLi3r6DERhJSTAfO0kAv4Mz
OoH9+O5lzGNgJoRR3AF+aQHjGYsyet9sPctB+mfM0QvkJhLXCnkX9ed+QsNgAtPMtzYCgKNoDgF2
0QtRWFRvmA2lmxzggRG4XrGqhcRpLJNp/cMm3n2gYZ6TfdTOHFN3dTVHIJl3EzGtVDryX86I+QQY
jKhq+S56jBjzh8AXEIhglCh9SaGCnlRFE5Gqzd99FqGBr95Hv4hu5lyHV1egkAmrbiQtfCjw0TIX
A6fNUSd4Aegg7Rxv6/WuWhv7JlrNKs8KhhvQO6oI0AYnbLIe4uhN7zFeLMIWeVXHbTSKfngD6VsA
+XabBibP4KiJcjPZK+jhICg4ipLaTnpM+R/xFUdsFTQd+WtmYy8xPLt6QgH7YtSgHn3896Yyk5ZI
ymFyop2wXL2v+7ThFsE+789s259feTlrmcYep1hwVXXpwlJHm12Q6mrPSMolQCSTMUMFkCGyRmH6
GSlv12yKYqecfHM9TJiBs6lIUlTC6WCDo4Q9+rcDexAK46jHp3iPE8dS16orpiVuu0KE15Nqm4Lt
nRzXUzK88V5s0sPSULWr5y+yKVomThpQB+qVWONO1cdIebJxFArRrh5QOHjvDmiMhJ5yK/v8Gcc5
mcEhhissHY1VaZR6EgE1v5v2ilQPeUjJWY8Q5UrEIF6yoUdOJ/No7dhaGmNoqPprkCUvtKlCN48H
qMZZCbigh7cxmJ7bhk/2bNdwFMOPgMJd6oQRQgQKYGW4zkCCOp5MGgVhd+GKXCpUOXzPE0VPojPL
hkFvk9XlaoX9LcQJm8cUCV24YlDU1M2mhwj4qPwQGq942aowP0yXxmBaPnL0rDCMS3JRv0t1YONL
IzAorAcDxeQg1uLy42hSfbPCWE6G3Zwy95CWEDRtfEJhnnXFG1/PRQ7Y/7Z4pfS7USlbgb7mtjYl
XAQpJ8Jbx9/qLMtXtG+x4ApeQKDWAStk4VL6ikT/gMYLLfp/bFEqzexxQIKAydmLQHXpGFH3WRn7
ZUkqP+G9YkhrtQGld+i5tf4+CTMmYkqysENkU/pFeg03NkVzd3MuU5LMH78RULlhIdiWlC7DwlH6
ghVjNicepoDg1AaaVmxvHGOWFtk3O8HMKHtXMVhzr2XtFQ52kTyGFxcrk/N2xz9W0nzeLweCsPmd
aHOvluUgbQLHJkiYJQOMeylY28oDLZZNjPeFPsx6PRtMs+n5LVWOUj+1D+06rFyHf0dxjVkeP6d1
zvRStqoQQMG5XJHg5Mnr1mn/lDImir9hGdZIvgJ6l31lgcS7pvu3elI1L5JRAijc0A+xxkKv21jm
QsUya0dRv7arHd8G0POt9SRFUN9uUiUdTSG9bVEPm2s7pU3rgCwhR22fdHN2HB1qBBoZn75wXnUh
bMS1hvBJlo5Zd4IUDB6CjOugzad6YUfJQh76EFAtguKUxBimY6JS0fOgbvlSzWFnNs+T4Zl0HB/F
KeIQyopOd+foxqyW9sg+h50Z1jkkPT27denl7wmZvmz5YRuLpOnu72d+fnutYDgMKroHYmIIs8fm
Dr0uRYi5BBPqulTLY8gZSZxMsuRBahB+c38H0yw4sFKSLp9s27G1wwu5uEMmIhHZlmDn6Xhkot/h
1zySnXYxNhT6+5sgLNNGk/7MTkGrOxNXORlgXEXkT41la6JSjBJyUDfXh5SyjagRAC0ue+hQBPNe
ndidr1blbxmImslIZ6iJ9gDwt2dCEmfG54lXFp10Sp68Zl1Av5SNtljn0ItkRi4TpL97qc6zQb2r
pWK5B0q9hZV06RrXfxUOb7sOhtafg9z8ji6ljd+Le4zMeY2+SLq8ilf+/8c/JJbWhNC2YDl61BLa
dOU9WXbxQeraCnFCx8a0tcZv6MJ/V9v/eVCgRxLobYyRYxzpqO/JuKwJm66FKbYXOXEykXFwFQWI
wUY7rpmE4BxwS9hRJg++pw6qm7PK7IxgUN78Gft48cG2izIKKCLf1/ztZUJAoZzhmfy0ppABZE2M
3awvAvJCi6uNWObXLfqqWONva3wh4IwYgBdyOi8J4Buc1W0xNrf1xfWprqRkWltdjK0O7/vCMQji
vSlR3LGVsFf1HyJj0h1v2utWaiwhzFaEUBnuZDkTMmGg381OpRZULJHjuOkgJJEzpW/79E3OodV0
Qy5zwJGsPuO69B7BbJaCfmptTbZdV3NV/4xjNn08XdkVrJF5Y6cJnf8Mf6XngZnWebQeNAJNQrrr
RUJqrJEDktPfIFpOfEqvUT0y5y9CvFgIlMbmCQhp3r6G7LtF7/d7p7xvhSf/1fx6NFyEENHDthnq
4tjWYLSqD0UdwwKOmjU77a0FqAH5FR4BJrSimNGPNZ75Kn8kYL01tCkdJEZ9IVSTNwxEMHXylkp5
qHMiJgZc4nVmxY9X0R7IG3mcJ3IoOkwMjuq5krC8r/ojMP3BT40Wpfmi1PSqnYouvRkLWhHmCYPS
jSVye5rfHtCZt0C7doam/Zna4XwFwDZ9NgCZJI8ya4YexmowapQKn9aCZCe+HZ4S67j4T2TfnHm8
FDpp90euSz+gRTeXjDH/zLCN8lyI5iUSqZwnGDTPknlgcgFpehlP96UBOfKAYynYNg8pOO/CoM3V
s8bJEO2WEc3lx63wlOhsDMMdGa274viRLDjhfoQOI1BqGiq/10c0NaEYem8NdArvGrMQjVbztuv4
GbGtKBwwLvRds21KjRNVpLc2VxvXrN57ly+HsxHSL4HYcRWbFL1ldO00SJc/ktGC/PF2M6E6Cl0G
+RimfIBvoJamKS6SNRGcum0vCiVAs5mCg67WdLq6eHx2LYTepIHNeYXRDb6tBxXkQBWC7KStvYlq
xyqKd9z/fk8SbmhGadEqaXVSRSgbDkvkioi6RVI0VdeDGHCZvg1hXDyPj471s6rveNlWM2mrbcwj
Gyv2Em9VZd5MAVrbVn4AXXDQJ9swVE1yZ8rDip1HKmxtv8VJUZ+UZqxq1/9fHxZySwyAgCGBSM3u
0T1oUoGgenVDn5SAuJfSRlIeBZ9GAjOTbj1LOcyAQvWYubswmepqKQpWW9r6LTK1Vf3W5yR7Hzig
HUe5qTmOSYyOiT10D7CZXb26ynmJXnIGXceIAKBGNfj8wqMNxhOLykhBPKGTIn+N5pB0Jh7cdg8w
xYKFiXf4+LErp7LnXotG8oZ0kAyeTwIjQMs0VwG4V+gpRUkRN4U04wkMht1KVGvd0qOfjaPaPmHO
CoJA0FugdmHYR6TZL1lDrGUOrV2/uYA221NV4wZAD60t0sBidqH6RgQHe+4gNYeCwYDLhBlKNEED
NyWQ/DXBp9U4gf6rQpvoH36wn8MHgf4iQUyTFLQfDKo6d3brX7jv6U4hwVGAXQsybh3+ZOcm6XOO
dlUDfp9xZb8X1os0oPUKDVMq9MXn3iCxllztjJf53jJryG6o5f8j0VogmBECA4NY875yEK2FSJ94
jxIAqFx3F4chxlgyHkvYcXg71fN1VRaYHyOVaq90DNRE3aMNuWNIHjNVpMTjKfCUJLqDsoqFLC/w
/40EzA48CA7xzX4ICIqDA+nNcdfHmUt85RTloiWpKgjyYqTesjzP3GsnFypyWx7oe3ag6xIdlPcc
aV0DQqvfxmbU7SBk20uE/dnTJ3KT1Zh5iZlG1CTBpD2Gx8zv4bNuqYINpOLuAT1d8P83koCIVIIm
r9o32YFXdY0Bsjrrm1zlUcsube86veX5tGDAnqtSVciLBFr9A0TVULJ+JAVUZ38HBicIEgORjOZx
sPFdquVtK9OBwMVR3IHunlVCUA8B3mwHk0eH7CciAQtcSGYt2uPE/ZsqgXyyLiXmJ2DyGFJaW3W7
N2U8WoYwWcFXI30P6DZazpwNkLufJiqO8TInptYTIafauPkCkvpZzW6py4zDjWu/bxt6G6kxTRqU
PeQwv5X7BoYOKGY1Y18q/BaDcZnlUqJoNr8SBLidre8dIT9xOzimGBQ+I1PavL8LqzEVBmkLyU3h
wTruo6LxD9NnUitP81x08TYe5j8w3XPe6BdsJVFNQLetrUdZYFGcn7GTXw77uKcHK6Mgh+FmGf1L
8SZfM61gS1+YCqImrEHVs6iM7rwaAub6qZL5IWRFY7JR7LRAcCnjRh2YT/0PE1t19BQdFYe2Gp30
vkD7RdMnQvzZutKK/k3b/174mnjqRrGgM9vfwVEEdWDgwYoLtWEyOf4blbeQ7B+F04Q4QO7pb42O
ARayxJOJgxUSNbTSumNBHMR3qDuXqimYsI/x+GV7voxze6PbUCWexh5IaZeZmCA15odzwTvGGkw5
L+ZWutLoTbtzZYGKUXibOtl+wvWbWPopb0atGudcSSEQWCmZ1ylYjKCPP+usafK1TeakZYqagnt9
MjxH1KsMkvBIygEMebBlFLp2SokUy8RrDaO0cT601aZzKvXoODm0NKnCL6tWcwlxj34g7oT6hspS
uS3zRNHpr+3UGWHKPJ2avo/iWKN19R5r1FwB41nziV8PpMdJKm/CmLgUG5RZCKhBb86szImedfA8
oDOkE3wjMOeUjv+kYOJ5x7GKCy2NzAHLgNafJxkEuwRzahEc5Z91QsyCNGa3q9SRHIImOPS4BEqX
hPsHWXM96KoVtauo/RDlDuDp8gclebUxwG94bpuvtgi27x/I/ABPagcmamotLGIkgCzkre0nIn5D
ZNIF9xuy5Ki9qegsEd47ZLRQqqu2iOJX8lJND/E7mwhuJIv2V6qr5+W3P3piq300cBoGgjQxTA12
HQulfCxY+1dcNV7kLQhhd24edp6KhX1ZErwQ02hRrqVHWM4ezQxtfkKVyGnCVpu2L5XNQ4RQf38B
TVW3c1QvU47LmgwwdgfZcFQuqbtvNdli4FfJrNEuR+jTuQlgX0FF+S1F8Wci8JpbP0aIJRI8b5gE
16PAVr7ykv5g5xU9pz4AHC1oB0KbaHrGDdtsjF1xosOy38ZPeqGW6lmxqayHbnZ0UVUmBTbJQB27
0XDCMe3gBP8k7nBpOHsIB9WeZY8VODQZnnsmJq4seaIXRQiBCWnxaF5bgMbIze+5neEt3vWWczzt
H93yIiALT4zVVYkpfMeCWcHpM/Ok2rjJ2cf8pCpNo/P62Y/ub+aT0OA5wQ02AvqlTsVWos+Guiid
d/r8a9RBSQhvI7r0lLFCWCeIj4eo/Fr3KW19QO9Efyv5aCfdat3BTMSmqiv7OGCacDSDoKchegUU
tf/RXZESOVh6Lr7Sw0ODAg/gjvg9AadsFQrMNmi9FCVYxuP+2HpM/Upqn4Ns6BIRkPTlFBcCg+su
kknPKnnKe6thie340q5zzqTGMPWn35BlggJIHlkOC/hQgPCrkafSXTPv4YlNrmSjks6hgNbX/4AU
b3fdGPs2UnPj3+N9QSVkp+wQ0CxBOoEVuUrYBK6ZjZmN2LyXNYu164BqCENlY2E08joKKxitBrQH
y6oIVKHc3j+OCX2Gntx0za/HgEQuAcGRYCnKv26iXIK2/MnuIHxNeKiDVCJzKAarglLtF65wyCvY
hoqGDyAyA7QU4NukvEnikyvUIcpFFnWG/FI83/BLxOwlni0KX2002/XA3XJ5tvCmYiW9m4mqmh9D
lyWngKujn/YpLg9ASXhz4AysF/4eXSxZi+YN7iXzgNw94lEMoe0dHV89jdbXTPW5gC3djaUpasax
/H/BR+ga8KnkkpCM8ytENai/UlH2ZqJ7rHMwltfVIT+7ISKvz32Zt4W2Vsa0jVbcicYK/dEuo6OB
C5BrHEbFuoMeTe+my2/d7Do622z6Ral3b0O1Qe/D/hesd+lSqki1JviKmAlOGJbkS2sIbL74OmWH
X5K/f1lBCiK7ruA1AJJXzUPTJenQTBJ+VjdGtf3lDyPB8M8vXu2pq96DQFtfbFdMefo+Q9yip4Sb
TG/gPk5Z1UbukpLKq4y10Rm8vH3rfI6QJbbpyq9IsZhUmZgOn+xrPEfOmseG6NgJANXmn2LJzCO3
k2x6KLQldBlOzEm9sMbDj1U3L2AZ56Dv4TBeV33BEbhOfBZVxS6xcb/Korrbc+uEW8+/etorisvc
6Mp07DGVr2iH3EADrJPAjbWWTdyBBg0xZrlxUeRlpy9i3xWH1AXNmVacWGwUd4hbBsyTmuwgXfHI
jL0oWBAZ+cqPemubnLC72m4DjHwIbMdbkzp2zL22psosTsTSeJyaVMC9/4M+AbvlPWBTd8O7LSON
v4lLdEyedILQGiyNdgKiwFR5B/mziR1PUvZxJU50dAPxdCSJXhs9KtBt8ZeeN6GO9koO8db7Do9K
fLVhIGj7m0RYu7JPn7/TbYZS7sMIS0uYNtzL17OypcIw7YuMeQUGbbEIIOI/2wFeeCXGsvf1MC7I
k/QNVpp9BWigApZelkzOdt9IfNzUPvA6Pw0lnZR9NRzoD+qmZY1CBZVYKgDvCC2rzpVQZOH9WQVV
Y6++31vKeXwpEfiIX+7JKk/fOkM8lDavV46mb9h1f2z0mpW5ESceKxZpJzjD+XyF/UBTsJmoCWYs
a/FXZl/ZSSOGjKul6VxgNRSqYkO1oQgyPMwJUXRaL8oSfuxtqPjv2MqBfIAwM0Jutiy9+AvqSCPB
S7Jmz+JMDRRyxkw+u/2K3FS7mFF5ol87RQVWHjjrknj7zhI8Vuq9NJ5dqifb5FFvgEGArA85Qkv0
qo9lLngRd0mlHZk6Z1tKGKGRFbg/wBxuJmCWWkjWZ2kQ2v7vIhGusUGosnPF/0ZvTvwh35sAAl4B
E1hsDuQjubhuwUnxgDUE69+hPC8zkmdCmwJoLU1yR4KFWhZc8YUi1Z1nDRPLMmPMXppXE0WhssUO
u6PzGajlxwXWne7Ge3E4mqt5aVlq5Zojt9EWxS858VkV3fGGAbCtZS+svsom26D54zd0W2DbvK7O
uFO47I5UktG1rR1iZaCIAD/BWhkhlylMX8+v0EZJl8wrx6/yiwaBm6nQ2xmXA92vkPpgfra+x/WK
qoj+qpHA+YBI1haZX6GxOUUFHAVo/sLj3eGY2FTPZQsWT27rFPsYqSZJwQpTOjnEprMJDSnPAsez
q0NnDpezyPUUndEgzJbIkvJqZVJ1rukrbEc85uKzczSTTQ+V7bXjhDdyTZ7d7/TgJGr4oMPOeFTZ
JTxMGE9CkfacofkPn+hZ6ZfxXjOstg8Kwzs8WQyKXn3Jvh+YPe4JzFsFuDA5JUQLmA/y1/xFbnMP
M5vs861wt4hLsi6gxXuxR3MUmmdHkydZCiOUZVq2Z5ucNiga/nCJE9iLnKwyY72NUvhQ4wbuCAd3
pqxPhCytzeIGE6QaqT77m1Yq+JiGAXVpZFy/DC8n2zitKQnWp4Bsvs/aQT+y/7cfzOnOw/FoaPKr
GAgw7o9SsLeSEd6SBfWrxxZX5swP3fSlxqdeoUJ09eo7864+EiU+ScbckT0q2DAPhj+iSwVjY74c
+tcWwqehldWvbXvRdNxQIcJwu6YbBQuFLd9ERvyw7g1IPHxyXZ/GMl1bXGRNg6N52I9fCy4fervW
4L181EyZFMb41x7inPODHv0jLx2U80peBTzLUktpS7IsSY7EvGhNkMrb4zkLYzaUWpiGN7NKlyi1
ZHNOh7gJgw8carW9w090Y82rWing/d/qXYUfGCJSn4V5ur6z0sKxsMdW8m6Ids8Ia7hYpuklCJ6g
QlOj5pfk9DTP/XP9nztSmo2+UjRjrDQ4HHHSy7FTKr0whj2SCI2VcpZx295IXmzU8AH2ybXVBOxs
klr0ZfJGlsK5QJWDyzX+dq2NBlqGlCocdqZpsUJ+k8OzWf+SFmdlA0O3CLnUy+bSh5J/75ey6g7A
jktzHIKYSuxpqISFLIQHs3pjrZun2mUZ55EhAZs7Iyp8cD6SWw0U9o1U/RQHx+bRED/ObDhOd4N9
hKR8hyVATUAX20ANc5NZK3yLwOfZz3r/GrBRZfMp3vC42KPcoJdVeBHlM6F8gluak9B8DpA86ddG
uNw/IpbjryCW3Qjl9qyqYBRxgtWB8Jl5ckPObDjEoHzGqOzqT/+mw84Edz3T0da3JtNmunRerU9Q
XIimXgfU4gplZEDUN2ss+EeRMNS9gThhleD9TNMdfhP1xF3ZsF0SdSJdNhozLyu/lzcI6Fq4GYUA
uwFQExW4m23M8tK+dZrRnk9ACQfnuDOE4QgLKpsPayLftikZ2o4c9DfFmE02E4BcrNyZ8E3RMOO7
Y9/Zh0tYv1gFkUD3HWDt66IKTHVGXBeBdDalVHvfN+uUNyrxi8lF8BLqVonT+XTImOdjOvosSiNd
iYREH8tWFgrw45yIGh5nARfjrcgWWPKDiv9oSMuar9CSLWSMtPe6zfmrU8676gXe1ESBbvio/NwX
G92SkWnAD2Wr01sfmo0rhGcu+k3wT2fAsvgjqXMLAenUWMa8ZilDVFv1h/JLvtJyH1fSD7f2gO8y
vRY3PFLHLfLE4Dtu4ee6r178KGcH/jgh4pghZMcaNLQM8xpM+xf8vL39ude21NKCgn97eDGpqQrQ
rdmuz+/bn000Ag7kEvo87NKzAi3EkUlsatwJTcbr1SKLSKpLOxTEcMex1wjd5gpem6Uw54sFPDcz
cUiRhY5f19vU8+hEgDJfYoXg696a0y5x6N5/f91g0if1nTQGPllYHkjRASkVBBMhF/1BKg+hzC5m
csnB9n2LO28DbF85ho6NzqGYpgoGW8n19nfporG8zxfCnnYuw2i/PboqJ0DNvAKZ5nkLGD+n/0Bu
sQ3DZl6fhUC8SVtInHHXO5SKKvlWLf+/BjIb1Fm19yMZRjbfdb2z/XtrPM+5bJDfKsJDUXxegXoG
JxxCIgx+XduxeNZFAWlwQjymz+YA+kfarWpYb7J6eaWyIGwGB6zaiQOI4EoEIofgYjDzhtscprNf
g+kOP8mXBsYD81XrImVgZR47cDx+kjN/SJAT4Nn7xDU+OZ1R9ZMtgIG13/jZz6cHgByXgqbh7eQO
fBN5Rqp6GUOBJo0uuQj2JTEzg6/XfBrTagULJtTTfV4ie8rAn66CTk+co48e2wKVM3w7DdMh3I3B
jus/vwhQ2jkt+MOiR/kHknr7Gnl4wFUFcyMaGM/XZ19Zyp8t/P+9rcaPDbZXrQMtIlOKgOjNLGpS
B6q97I5IIgG4o9t3sgW5+QX5T7yxt0lHOcDEt1mr2+VqSRo+YZmtbalBySnNll0X4wfJUmVVTDPl
ZFwRzj110H5Hnb6puV5SxyhTK7trtBKMubhGE7s/YfxQcJOSYYE1C7JpGLl8mgO8+FgrqR2eW1iw
G7jwnVWO46rRa0dHUEAnx9LaqG1Deg16WJ6n0dgOysgWDOLZ2HVrL4dhS2w7CF2JZmuiCqg5daY3
ScHXDoOw8oJV+NIyGrzk8rAcgfjShB/4AgCkYSqqOjl9kjb0oTSUomI5asn1cMA24ZjyeU8fI7IP
RR06ojtwuD9jwm+Fua/4YdRonBCtqpPY5ugJbNpR3aRkFKnRyZH4OtP3392dSv4xyeCIC7lf96qB
MJD6MHr1KoP0oAf98SsgTGKzgYnZlrtw7uOYA92uwT2p3q94VHg0TDpPLTV8zUlHQ0npuQXkgUoK
0dadSySo6Y8NcsfvwZ9JF7jn1azHwcB8Sef5jmBiWznGWSW3cPlKDESI8u/ygCXKOIZW0fAWfJGy
GfnaEMRcxbJuI6xMYCh35YiD6FSEo7Gy20KgXnoxdOWhb5u6kSE3u6lIbZS2n3MMqZj9sAVT5CnP
sdkuAvUd6fEKPKc64SxBDz2LkxY3N7U9Q67/Bk6w+y2lAzvffjuxT7r9cgghKNXaO7NIwnVVknZS
usNlr01R5FRN5ztWUz7JO4qtmgW2Z7LpZorevxd8Vqir5BdcCoYXexox7voTCLjeKrLUh02X35Sh
eSwXexVQaB2rC47WuOJAj1eAKLEP0OOqestyMi84oGcvVOewIl3BxuD+cWqsUiFQMMqLnhH7iQsT
PLBge/UE8zj4oOpG5XEKLGkBOmD/Jhgok/adKBTQKPtJlHyXfwOXGiCYiO6cKqwvdRp4u7mFEeTL
DF493QpNZI6cJY7uUZoy5QJ9TkspBhEUSsoyPRW4bEFwdfYSn/RGgJyJUpO/j9QsG12vqyMoeNLI
dfRfbQuth1emArIk2aYrwDNnBLXKi6Wso0TrOI/cBTX/q8vKcAQcaU3LqdM+nqKlLfp2P8HZ4zLC
xm/DM0027hFsgn4+Fa2N1vKTpCLXfz7eKlrAzmp8ZCxR7YSSh6MJ3G9l6Kxh49RtBysSzNohCpVE
HnLNc66qktUhXdeRkzY4BC+yrTfxyyyEQ5YonjFJMZXKiJ6QuBFsQV4zXd9A/MDeMDlZyuI6Yop0
v7D3fmwlLboVeWKu16DS9Hnt4TCwbmF6K2hcPPJbyboVRaQAqaOZ2OYcrQGCCW1dGnYbtIk2lVAp
N9ZJNewGsUc6rZAfWs6oudacCNzzzeqi70OicNkCOrBjSFuxjPYLfp1CLZZzIy+MDKOe748dUylp
LgP5yOwMD5ErV+4pFVUK4wVGAUJ1c4nNyIViJuGO1uOMtbSWm6shdrEFFkZp/jVm89lx6Mg4CvB/
m7e90rh344HE9LKE0GiAFbmjsBHFCeN3DHuGDSWcSDhloxffWRKiBzXUpmcPZbKGKi/GNahLFNQt
3/In1PHaBfLeSls65h3HzxemUMKCtOCXeTMgHjl+sQ6B1xCtk9W9BQML50mjFuj8ucMGf04gKJkC
/d38mS8k/gcr7cg48m2Fue1ho0la20dK8pTDA2PKvsMSOfuGsgb7R37ucEkDvrq22fLy42LEV+fT
UMD1gedjuJg3cWBTRcaPiqWsAuogA7SEiNgiTfJIqWoRrsZQWxv9JRACBe5C4k8t3LvVHtxJTIZH
2jiOk6HoXV7ldk6jWCeuZCqSy7oIaSWuT9xER94/05nE9SqlxN4G1i7riJ/J9i3q+CeCfAGw+T+O
Vq+q1r/YaneUIW3huLBXWH0ql1Utq5FI8cIiffpoyeBgzpyquq0whwQTalY3upskJ40pTmGx1xIZ
/Sv9OiwGj7+K9RJiZArtF9vdBYdoz0GheFAM32pSu65PyW58aCHUqJOAYzsQ7lMdqU4ZsMnHhbuh
OXuK9/ytRexqvCXQAxfKtcmIehlH+FAvwVTn8KEvO/s9YJPJoS4s4AZKJBQI1nPwrK+HJkvos3tv
YI4GT/ky40XuuzxGkKRFHSjSKekDLx40OrSU0E6pBeIsckFggDdzVcBJ7LdXEJpjb6oN1Jm6I81j
stPPteMUFev8CBaVOYzkfALZVRyXSpy0B7y0d332zV28Mn5QGmtFZPix0ZCqWrhR0vQozCpI7RLf
IYtQ6zy7zsQ1LOqIggrQ2iPvaT4C/qHGh4RQkuFq6vUj4ybzPVihPdq9IijU4iLJcuyepOT6mjkp
4vx0zojxD+ulMSdPvuN4Zu3K4oS+8WHqPHMivn9bglx9CDGeeVr/dmFFIr/Tu3nXOAzGXXyTLzqZ
ZMZE9Q0tER4PqouLDTNY/OXuea1y8KKX0LDcjtato4bQxUlA744XgVSpJrHmAnSHD7Haii1SZTzv
HqX1kbsldKHfcnmA5m05iFsICqvR7cbH+1MTIG9XkaPIOBZ+Bu4+SMiTQJ3foRQp0zP8IZ60ucKu
3fGa/r9ePc9T5mQ9jKH1BzHC2dxQTa3iw+1h9UwG7KVhBy0bv9DYX0tSEz3zD2uhvLCJ+UeW4xMl
+3pGo1SBGXV7eisWGUknfj8FehDlUt6EGZ7fDrUwO0Mypj47hJXewNIYO/XFZHF0tRuv5mEpUdML
O2Nbb4eGukGLnAaJzNX3yDZMsfJNBqwK6Ng0E8YAyWIDDd4XAiRME6u/8Z2ocqEjTN7lZn2mvmJH
TzHCP0DtUsoZHezrArhgLghmGrubqUwwE6clxyPbUhfiu4Bdz4zK1dBEoLl95fPYd5HnPUVGF3Sh
EQoAa7XfZM6xcSdPZ02yAhldFZpjERlKEoY7ZuCbZh5lWp7sclXNalfa3mYRyn63E2olFln65UGU
RLq8jnsIBZTPeuFpI6yDV11yqAryH3WkuFCVO++Ju8Bs00n2I0J2ik4UdJDpfjW1RTqawgYYyezx
6a0PVb7iISRXz16kTanKJ5/GEfKpDSeQ3IObuKjoXIxiusx8JZQWwXkUit4UPsCA8XKyHJMy5iBd
Zjt/hKhQNMsOg54WhJfQrx77y3MTe/Tm8SimftDhyKmnP/tylEoYbyidehNdVJu9NwyHaPvYBz7I
tRxBO0vTDrwa9qptoRN9/zIcZEQNX1lxz4RwY70SFXGDH4y3K1AA1rxGP6ypvz6HtuOISbwgMmlP
s+gxVU/80ZxcpugXGjl+OwGa0zZKXVo/8WCdDhjJY8Gt+TUYrcoHElvmQPHxfO1dVCj9pDLhWgCy
EBWpnvm4I1/GrzZcuoaln92rEAH9gl1Tbbq/kZ8ePq7SWdxnT/P1l5BQDXM4PRgilpm64uAl/StL
3Ysl9mEz0J79vMl7jcfgVeViPfxgs+Sx9BEb056ikPYWVQHA4bEg23HTBcj9oMJv9JuHSPyi6Fqg
eTcwzhL6MhHg7nuXGZpaJQFXULFzg9QHqrhMDTChVcYvlx4EI4LOewNXalwXy3vh5mN85D0VzC9Z
wzj6rXFzPVKiMLLEdEKXU1sbVbQwYK/pyelnXeWKFIKZHGIndTKUmR+19HaFEYqEEpqWK1dYOwHh
DqUb41yH5bRCO3mYwvY6Ea3rgIL2HaCALj7WXUhKzjLG83h9YLQ51GUmE61b0AZgneNCE5Ipcxfm
j/g+yHArJw+8RKO5i73V3Qbmw2DXGE6sNJQKu3OyNAAVZhMG1rA6MaZAlPcZGw5U/YwsooXIzjSf
6rmVKLbO/XVdPAm1NavAei10n4zCSfKpLt0Y4weUREzxDMaRXG189o2kEDkN+XYC/k42RuzZUZi6
o09eiR1P9JqDbOVumpt84n9ppjNvuK464A716wbZjfAxMAfJw959EK4N4pjxz7r710pw5lcbCAqO
2s5FWup4sP1TIWchhDxzmhL0zVVfTZGsiyP2SPbozgK29bvjn+jjEj1ukcPcJmApcAklgyhfv16P
8AerZA/3YjSU2q2IKscQid2Hr5BdZeNQwHVmh6W4bBWIXHZ2jCsFmD+y1JnEqXY0YZB9dmDeh/To
9Qjp6r4+IgIRfGGORz6yoTuvU5BNN1Om3Kb2ClvHeD07KtgrHVgnrVCtobMMB4ewUayevXswEIeu
AYKPpeVbpNpIGKeAVt5LBmWvDWJzzivV/syFk/PqSIlrJzYWRgciXyZ1qdFY9Savbb0Mt/CqlR5v
FCmn+J3xTYOh2g2Reig7vY8CrZuXVwn7EK383xD5gS9XX8mXFs7Ac78VYkdOykDn362wEYcXL3sL
7Qj5jzLszBVyPbLxde83Pv8jnyX4qMguiVCOm8SAsf9m9ac4Ra8HRSvfagQEe96phc5VHcq8Xh3j
rnC48FmqlVEGpnBwkDFhUkqzPW3yvExUnYPFKAr6L9ufuqoLXWWSeBUMQAZTX2cSnW4WuifyiOem
PKA3AS+jcDVPgamVk/dHxGfEzoFUr/bqsZ0ziNTk8JWJG2bke+HEw+9CkCkPcbNVp9aXGjuoj6VL
ZBKmOEd9v2LHn2wEg3vk7kglN7MSJ70hsrKBzZubnrrOuJHZT6FgYw3IwrSp83c/vFp5bOobJQ7C
ecCSp8utNCziV+d0RUcKIaPeL6dc+z2k102e9afWn7n1YktdJdx6QtEzMe1kQNSEqIC41pHHJrzV
bw9fHvsFeyrQu2URFbWuZpFVPzM6gyHTOpdBoFunQB8OrBq/+GjNpouGyjunZ+xuFMdpEcdcfz5O
8Vi74AKz9/IOUWnfnUUCu3EWJRQqz9IgcXJsqUuBx6hLX6araOWyCjH0LCCsEUt6InaiXnE5jO3w
EaOLwo/Z2KTl0OuZ2aK//+BxQZMCrXau4EWo41Mdt7vRJfu+Se7G6vzimAwhgzFr8sYw3kIfjp5/
ZQ7RHl5AIJvmWx3V+M//nmAmiTrMDMzQUF6lzyaUURMHWCVlLwqokzTqYc7MV7cSy+a2C8c1axph
zau8TkyYLq1X/p54lowzlLF8HGg5zHd15+SDvyB8N7n90l3sKnedS5GgwZonqGX4j04I5ZOjVkq2
VaELszDAbw6tftHH7M/dMsUhMJasvAVYydldxEvBApCD6zy8y0meNk7H5WvEb+oUcm7iopLPZZuS
3zPnFHyj4i3sKkYLTkXBbEpPBgzz2cwPTv8iy78mMZV4NCLNaAvOWaxU1G+jNn3Ai9YIlMhMaQHd
OvvbpQUQCrUto22t9lBePKK+YHqmX02IvOgmz5wW2ovK+yZKJvr3xrk9Zg1aW6N2M+344lS5JqUA
uYMQywXBpEZ3KhicJtSnFMVqcfjBL4lskvh40H7PdA4WBxUuUACosJ5XEPdaZuyzmvsGFmum8jX4
+b8w08YrEEr5PTyaWpbLF6a38+RXy4eqCO2FkM4gu5oZCstHNrSuwOMsP5lvD4rdS0Q3jtTqi969
39fjaJ8NmOmWqOLfenXskfMm53Ce+LCrIqWnPvvoyCIvkXNUPb0G1odglCDLmnDP/ti6PHjKL8sT
VBJ6sB4myPzTnJiISFjKHIwC1sYHvHPpQQRoWz2/QrLC1grb+WA+4tknYYYCLNuPn6TqRkPRcDwP
DO+M8yYYNWnzU+vmByLO8bP4sKNfv2x/Upkox7RgJoN2Mfvj8IFMmO4q5L9t0xjKgLq3PbKZ6dU5
DPJ9k2Fu9L7BNknxlj5BMsKsrbCeEjta75/ocI+QLVv286fzmio5vTcEE1FOFTfIDTXrAySIfQoZ
SZnubt/NVW7p3QA/1/astQV09kL3N/mmHNXDR4mqQeyVb62Y+cqR6GxztboOw4/z5l4wh95OBNvb
nFsn0nigVXP6bU839OYrGFjyXJ/T5umQnRhftt00GffmdN+myhUpcPTgMeG54mymPwLVBN9F9ZNF
3PA7OVS/kaSx1PYlgbTAHRPSZOKtjAvB1g9a1q8ewTM4dhGtYSmLm3v2l21+/4k4dbAPIGAAo8KH
FKDPkvim+7stk/6F+bnFfl5K0amf8MfgEnCyTLuTlSo+sgsGDdr/awv2S4I8WEX+q1vh3N5Vbdsu
iXBBuM9SjxaBUKNkb7D0E5xXcg+Qes8a7h/rxc2N4blFF1LG6apCdNike4ihfFJSNX8Tc3RK4BZ0
0FjFqEAie3eIL1BBnW+F8rvjCcoqzRt1x0y5yM5aEBGpmwMTxUqEyVhEWTzKxFzdJPVFAQoLHna9
7OQnFU0wdMh58vLa8Rl/fWQix8Nm4BNeBdYemPrx1Dm0xMDA5sv7gyy6C5LmS8PF+gMU/0CbCBCr
5+cFJAEmC7qrXivvB9PEIL7fXGYMgYqMdCeqnotrDFaneDeyZw5fcjhxTnT+KxdbozF1ameiALAl
WFiMqjGfBmoIH9bQ3/JNUhnx83PkvvLz0rFEc9XrfQdzO9g6fIf3IPKqOq6tPmlwCkPk5cjIUfRs
Kn4KoMqt7cmZ6zxGMSKK3+oJ1hTer+msEIPbSIs+o1vwzowVNmteVuEA7e5JLpEuUF3JDEmMc7tR
WztY1jQsHZRilyVZTdupbbf7ceqsH73yvyyf9mAJEmEpjZXvcqqcnulqAXQgVxLB3Og5iZ0+FB94
OkpAibquJe8nKjknHo2cbQOGwXaxVyTd5MBnux7FOJLbdfYKfcr/fhSFQpngNKNbZ7eMtSqG8GDw
2Kesaho/YRAdOy5A3YL9sV7D5II2jUlS7hwlBYkFWrHyH2gJyKql+gpcHg9Su+bRrRH9gBGpj4ZU
FsN+7okAsmxliNQX06fiWTUuKmYNy2w5gn5QRSblzJEjPugALlzCJiv9fgWt2I5rUZaIglaXr0Or
YRAXtWuA5l5dT9qHNMYC8OnQ7NxXPqjiKaztMDJFbu+opz5a1FENXnMiOzlGqzWi+o01f5ptAwE8
y7RfmIJCY/j6o4dw1ZfuHqtlxNz98JyeoR2VZU7waPnpP+lyn9UqiITU3PKZF6QwDHtDUmBMM45l
f+/sO/2GaRSE8bOKLpAXuWMXY+4G1R9sBnniwHbyK3Gd7vcSKycvi6vtcjeiY0vQ8qkM/204hY86
GkJFtgTLMVDLUe4caOUpYPEwuiuS+M1tYU4l5EGIzxqbiGs712SqkMjeui55D+KRqjB7nOtoWYWr
M8a97KpZjsEtLR1D5koNio5M3Aqmu4Rp6BFGdUXjfyq5GCkZ8msRlYxdm0mNfP8G49S2Y85TbKsI
vlG+2KxJOQp7ttl/4nemV061LX42Kce/Gkp//JNXMJ9eZGW/HCzisb3+Fwe3dNWzlcR26YFJB+Y7
w8QqdJ5QOVx2ukPA1oIOmbyr6ttiO5T9LzNS/6hVMUY+b9tcFcUZfrhZXHq6AveoKjHnq9XnWhc5
FipFxdGkgQbF89mmyJImJ9yDaVuxcByS5W1b2cmFZmQzRSa1lIoeV9t7wpsb3C2h8tqjE3rKibnr
4W07umEwOxavajN7eUh3PjFTPLUM0bK8mybup5zOG78WCFPtEQ7BC9VD/WfU14I/74uHJicdQj2O
lzna7GVOnIH1ILAADIWDSZOwYHSfsuZYq7pZvOv7RYbqnCoDpFjmNqq0qjZY/npixDHFwTDSaZqh
i8vGT9ekl3T+6SRDfKI4LRfPwJaVXmXDrskYa48lWDz5S8Jwts0MlZ8l/unl9BdDrZtVju5sJ2Gg
/PvyqsT7FEMOrLx5LHN5Otq56g/45zvtXqdexkIXbgX7FEGNqS9vQ+yOzgrfcCUOwXp3d2XHOKOQ
AkZsi8VKu+tVCjRG++KztLf/sgXe/ZqtnaIO3Qh8Y3PplRld6EUFKcArHWrv8WJELy6Aka7QCbX2
JGwz8QNyxlwAwMjXrvvBJgEEHNS0MVDTqy9iaQczl1FpYYG+K/TQExxQ5zE0ueOLtlaCPRXN/VeY
c5d1XkGMvWUyq4fpZdV9m5VQoQqRI0BzU4kO+9oR4U4blj83iNQr4wDcFqt+vkelmwfmabO/3twS
MNHr9dLIJFNHYwOjId7D1tUHEGgiNawcmonNLo5degZ4Pe408e382AMt0ue4iWqCZuHiFR4J21B7
r9lqPnwMi/MVtc7+6g9sanp9Pk+zpaRq+4vsObpWo5stcT58aUCCvwfWm4g/1aPR1+eNtXOfcPBz
36+mKuPpNtQiAXkGhbYUi5twW9Rg3ZWP7miYkF7DzpoPe0e+2Wo6rbbIZF7NP1YLns/W9bJN7fWK
LHdtAIBGejhydMFD7WlZ5jDKp2vC3hM8g+hVHFEigEVUX3BXIT7IelM4jyajl0CxwjLCuWdAoyUu
Ku/ynaEmA9WIOhNxTatQVnlHXwcuVcVyb5/EOfhrfeqN+s9J1ksGFL6z6MSDjpE8B1ke0mCjLq2X
huxhX1WTO3HFAtcLGZ6i0uGvtOt2NgPjgLk5T5LuE9fEdip8pMyieyoXheITc1dnOS/OALYfJtfM
12A31xLBCpgHzeEyW/oAEl3TWx9yIN/BS/NA5OQgs4mkByQROm4vXzCjp2O37LkN2mqrSz5R6sIb
CqxAVw7InNUA3Ng97iewE9n82jipeUGbbLBiMpsUy6ssmwXlQeuoPctxkmzdusklCDPL/1PLKaZB
EeuO6EGr/nrsp42M5dEIK+Sce1iNKrsn+D11Htkvm9wlf1i8IACXNKUBYzLp0p5I3EsePzM5rM+2
ybdlQNHAmgCE8xGr7kLtgghWWqoY5Sl6J11vg2EXWXmGbmOGGlHuUuUWL32n8NDcCHX0Na0Up9F8
PmtqnOYNDubW5x6z7Vb8ug9AsoGL1NgYoCR1Z53LB2hr/Vc2xMdAx+FXB1nD5ff5yJ93GgoDhDI0
n0K5fK3kTTuTED6yYaPQZ7S3VWGpGTjFB6QQmTm5JdAAlm7uZ31JQJLuYmuXyOduoqTKex3/l1g8
jIzVT2JIw0nj//QigitLt4ArGEt9Mn88uIxSbYJevQNG+4yzl++FNC0t5LkfL1mBoGaCD7ACOWTj
/DKtciz28GhDx/LP/HRiaVv8ig550VyIjMq586T1EwPc3kWTlmiiAXTSKCPZU85pps5LZbTwMFy7
HiGrmW8sJnvjFf571Sf7Qk0jIl+Zs/Fd4+03VzfFGwjoWEpMbgA8NqwsrpWTLWXP2dou7+z9VL9y
4yTM3KXoAx42LEsonGdDBTC0iFX5AutAansPjKp5QiNW1+yxVToRCwJHmsoovICwe1fw4zKwbS91
tvSlFyPmLVQYnwM4AdFlPm9e2NjN7jzODy4OMMriH/uwX9m3nfx23BL3VJEIdSyMCzG1tLveMi6J
znnUP1yJusQrFrlhwYfhhbUOcMt7U1G+8ubsia/gUMBJ8ubeOE0VHeMw38VOuE91HZJqk5ih9MhM
E4WJXKpI+fYR5sFmeJxAF0HvCT/Mx/P+WZ5Pl9LkVnQWvLNv0haottCzZ6RwvF9BdxexXcC7nUw9
qD1wgiNjgpBG1RZjpoVIl0ei3oiE4A34EGuOUaQJZuFfbP+YYq/P7QxT6w2F1/n8lKP1bbjCCRWO
7CnouUfROPEVz3PQjiWADs8dkido069KeehsvDm4PzKIX0NEWsPW6AZ2z144GSfojuCT5RuNERUV
W1zEcrQKoLKfkUGD+xFElLktmWecYKhOMilnn8TzMeJtFG7j8wthzFsATPVs/R/1Ta8qjD8DvpVB
n0Oadc1EwwypIImwUFQ9rOxDGWdc4g40Fw21c5cLqmhR9IGyEV5CMRZxJUawCprwwjg9YwICPTf9
B6LMMfeUAgcXQfGv7QkXewjyLc5axVmBWuFN/C4HW+oZ2kNjkRay0y90cwSywDe7jf31TlLXXZJo
nQkWpXZnM7oooQ9KM3h3VI+s8mxYbg8Q7EY5xCCNaT92mv/O6qKYOjA4Uhx10lS8T0t8FF54l1HJ
K21p5hWb6pXl1RlFuNRRDA5GBb9RTYMCo9f6Vi14fA+wZnRqIo0eD/w8xp1crUbirk41R8+ZSdB5
kXxfDQ2h/ub1RJfSkO7NUusQpdqTiN9kU+7FETFMZXiTZfeuHB5kNQGSGu64Zhof8jca4STITlgP
CkowJznvGjEMwr257chrPSCknhL9cVjZvB9c3KwaIOLcaOOhnY56psWrG2DCY2a7/GVnu1ZwKlcO
Iz5DwDZmWAPgfZUQ/8mOyAZxp2kWIoSdOfkw/2vvcqrnW1nFPYHsdxKVpcBeJgNa4TJwz3APUjdc
XzbJJEnhocH51Xrls5tZ2et13nrPNoAxG1zEUTzfQq+xmTrUmmOmam7YjRd7qqiq/7F0z46Hp4Vb
TN8dkAwdnT3kbKKLmiL7FcAn2RrZkOcPMqEOxyGAFcxkXk3SJbCtGOft33+RZsNDQJAzWWSm+JWU
2JlgSbeajHwafMYqbszmoQWgvyuWtr3eXonVtlcwVF2qNQ1a2+sHd022U6w2TNJiUkOPSOlw6V3s
h5PbqnwQanNguesyvDdDRMiZY8bzF0LbC726VIkltSXqmHzTEbJkI33oxEUwXVcmQFghJy3TTTx6
YLzNQw/ifivt5MC46yqRd9mQR6wcPQuC7LSkMaOXFG4BFjLM9FsLw+712T0rk+tr14FN8LfQ16IM
NyhAlIQVvO/IlEeWZ+DCRLUaoqPxhUnHv/0TnZDc91KwzfnkqAp2h1F/OVLs5nP51bLCD9PnWLKB
WE6daQLiXxDdWSVj8c8SUW9M3iIPoK6Paz1Co04o59hI2i8RJcB+91Tcvd8qcIcKvbKpaegF9aMF
fWc5Xi+NBRvnpkujQu+hyEJDZbu9IVF5CRi0q8zn6MDM+gLsMlKPCZ6lOTb3NgV24mJx18JRGkY/
5rrJYfyg0slILXYYN+VQek60mZmTEKYRHfTmXbnZElZrXOAEGzujcuJNmhN+xfCFiMJlihlOPohm
bO5FrQkyuqS5HpOQIEx9U6PejFpl0Ptv1gUGsU9EBsPj1G7XJeob3fkyA3IFvZ5pydC8nILBa63t
0uU47ZZBrJ4FLj5g9uYxQ/oD1c/iqAQmkFIsBB+w3U25Zfa7OQmAxWdxMDJ1RH6qjz1x4JjHHvXj
t+n37TTSc9FKrn1wIg3qUGI69s0lmVg66Ph7WvpRSWGfkAmiHi1nzhD85voTMOOqgzjXByB387UK
eqxd6cHBiu477nC0ioIvlcXNcgJOaUGVe6dBlFQkZI366qRGawEGsxyl9QGIWuRvJ88lsDByUsow
WyYY5pYA1dN2lQW6Jo7fcuOaIdLDf2r8LLzKm/tqy+XzzuHMizQDY2a0hdujMsidjfOrZDGj469F
kDzlOjO2TZiwENjr69SkyH2LtTYXI26DupsRd5UCmm7uBlCYDZwMXzfSlI1iBHsLtMRc0C1kDR8V
2pUCzDLUo6/nh5ETIvDxI4pnCfrzjsNJMW2WFWMJA+04jZKUokL3WHqym1G60bYX1Qyndcd13ulz
IEHEoYJJQ5i1Ks/6oORFSJDw0mxEV+s1WkX1KAsaFy7pb6abbTxgQ0iPwX3lL0W2VQmlx54ZLs6H
WVFtcrZ9FqVFxsyBlyGFM+JroYTGqpcrJsguSPCvPJPSoW8RyBeLxxHxU4gCnUkfkfQVWypLhDLi
Gn9WaLBQ/EMdWORT8gBNDtoYdB2QKGDSVaVyiixq+5PGYwGlBITeeLrQJciDWKEtFoxQm3PKTT/7
E/zPQAAOyntxibm9mbM49nITaRbkB293H3HzmtDfaXEI97ZoQXxkoB+wO01ZqCYmoHviLcJeGhUf
Fr1HZRxF+7kBhNmDbAJFFhma7uEMjgxAHsmIA4YL3P1fdGHp59i+urrVl0PUSwNUzSe7mwIWsrWO
nSh4vZUhPeeovf/X9ejImCF0iNjeBI5wvW+7cY/caQSuNA7jRePNXgtbEwKRKV/Pt5n8yC1csHps
3kUyBWU4am773ojjrL9nmSL9k0cALpnVo5nLW6CX5u5J8oOuh/nX2GNABE/GBWqSzukSwSSvO3oU
oly8eE1Y70dyQFHCIk/W0a/zN+69V9+VGuu5EwDaV20OkT8vwrVInmmyTGD/b4L0H50P2zcqmvP7
QKrHtH//CzKYHVV11kk7187gb1PFQd0YnYcwwCl/FTJ7XQFuLBmLQHekaupLZzv9iGqel5MjdaIF
HSYv8HX5/AlUAvrpAzQ1lPu7yHy5ysutfbbT68+4Fq9oKRT3nSNImMXJuyDarwJirSj+3Cn9NTc/
kwzeCBgHvc5HLQ0/QZmWJsHNiXjPnB+nylTNsYjgTKgC1Opxq3pdG4+F2azhCH5HPgUg0lBr08xK
BVeTQKGmVnd8JbSQ9yzjKhHGDR7kx7jKnkjAZx4RdwX9YfG6V4ACZOAJQT8HURjZeJP1OIagUaNX
CmUmrrziwfX9ceXCOG0J2G8XlfSfCvWnUQgCVOv1COP3Uxrw7VK6BbG5cvj6yapqQI6DPsErN/OQ
1SR5AtyBz593AltDIYLwR7P+R01mU2pcM0OtFulPEp5cKCGYWs27m4WGVHMNI8qIYSSjiYQE0k7Y
0rh1SZlUhsvIZfMay2KFh6IyS6OJ2KDE89GFu2UGDmSpuv9haqdChB0M1iqbgDqdnpaDk6/r+SCI
r6VYU54Y5i5fqS/JBLQhcP7gst3StzgRvf/vwrRv0lQ4NlW47dM87U9eeva5uptMl8+U4Kn95ISK
sLBstvZTmLgfKP0UjlHSLQcafdgmEcjW0l2tiSeX+OcG/XZUrwCF8hCiIX5TzTmkm+BM/+5334CC
3Bx3FjqEBNyEn+sXLBd4GdrhrnwefpUMDOdXRDo2Ekzu95hijwuPPpWDZ0eyIuw9ROj9ry0BsV+V
tKIfP+XrWjh/zMeDUs9TqFe2nLNa0d0X0qzIlnTNBJTqpK4hXbB1ikL/h2ol9mcN3I593bnAG2B0
7SDWyUrY+YPiGUgLugLfgwczt0EBphD9VDRi2KJmwjao3ZDd0tp5bxcXrKFDUPDytTeUnyXbwE8t
iy+M0N+8j5xmEZ1yWBCvRzKk1o9/ys7CKdNfJiUNOVRhYwWnCCuJpSORaRmDEhOVGWP1e0XQ6y6W
uV+SPnhDR6hOGPvQqEPoQ70ownEBjR9XgYHA68mfYwahETyxf57QWxnZjm234bBlfhFDvhDDT9r+
0X69DRI7yquEbWbaMqpbdTc/7R8z1SC/SDur9YV6rZ9Dz6umgI0IhUYhidenJb4YIENQNBP7REUH
aZ3ISMTL068bNbnVPsEdTabGGv4ZwUEa+GKTjmP/V/Um6lPIVEiPFIq+fD3Aa9jpW78nY+7uCuk+
RJLknwwWU/zLnWt63GxZ2gqV9bFA1FoSYhpcZemGYpj85X91jJZpt8C4jwlwnkxre/PN4tHamwfw
BcWluPXyVVG8WS6TIYqvdqlCa8Qjvz/PAR8ibKW7xMw9Hcnz3jJkypwA4xS9IDQiC+l3Grc46+fd
9hKBZH/+e9aPdZTJdtntV3iI9oD+tzovgD9L1x9Pb8eeT401CRKfwhz744rcN0REPHJA+ffBxQ4Q
VH9Rpx4ACr8EtDNXhQAWoJCydYFOaph3umbBerWPmsp7fZw5c3smii3RiQP1Y7/Royfmg0rBGQeq
BmQo+WtV439R0HsiJBtdByzovm3slsCIgvVEaVevAhCP8qWRJEq2JEP0N8n+kTydxu0HBZynoTXb
50nU117VVE81R3JImsYtn4vuXkcT7PE1KF30KVKtqU/S+8PIEJeACYxM5S7PwBkQaNdf5QRskOXl
7ChMK7de14yNNQnr8o1UD+BwVqmWWp3w4wSvxvsztK+cy+32kgDX5IW0DxQzrW1nOESfd1wMAp9z
FDEh88RuVChqNtnTgOTPqu6+tkgkjB4RySITypq0IzddnDoxVQrL2XsRN+T8XuH4l4V4BNzS7JIU
NIaMgO8DqOLfVyRaT0ikYeR+Vk5BtnGCWMdexUTJ5YoMa5/Di9xgG/HfP/GUIeZuJUph+VOkPSDJ
4nHIAvfeVrZE/TfnS7cEN8uRPIZklBGKR0h2KetuJcoTGlAU+bw3P3+oaJ7r8XO5ygsp+nTyIPJN
DkF1RlqRGpMNl2BR1vHAIB8PEXKDDFztj340PUiGrOeUXQZ7qIjZFXtnrRv37kt0cldhmW7EzE8N
mLyjGgfTx/P9jghKIf/CNq1hxIQ/mr5Z9LoTUX9kAhzZE8b0cP42bhQigmRF4ksJH7XnLgH31K/w
pDTiZijf/x8vxSiwi33d5isu7QwDxAA/+cYqhHW327G2mQtmNAow4qcEqgNYKBx1ssQdskxva2AH
3JK5hXhGlnm49jHHkJNmXyEaNl8grk31hiAWLU9F9+LtXvqUB/1FwKK99j1o4xPSuuK11KCaUFE9
7TGmmMZGj8yk1gQpZk0Byp/dyNzjdfIn01E2BIvTLIErYvgN4Gmtp+yAWXLh5EcAxRZ0Bew+0I75
g+oxOe5e1g/VuEn2YDcypM4d+AVZORtHAFTPZiScacGKIF8Fu/e86BQPxs4fqAsfv9hS1hmsDRlh
6Ztwt/U9T0Cu+GqD4evYiURyaAgRarE9OGOHOrkxauuwZb/Iotw9a76Re+3l5oHdWysqrKRTnieD
9MMhSufEl7r7xiO3rigoPgCts6wEJo0+vTmkABmVr/lWLMqS2gnz95TLBVB6m3wF/FGvQ46sWMCj
ZETyudz/6THd5Oli/VddNhs+3+X6iW28tk1n+8neWPr8peW+UJyFLszRUt4WwV3+uSUHFFWJoR7r
n4QRJb/5DaSHKRUyhIw9x1/3SXmc6lp77pkSZCp5k4rx0Lr7rMS4S2QxPeLVg07H4XCfw35MmA0x
uX3qXwxgatRa1sKNJ3WHy+nSQg8E096wOwWol4MmHmhhhmqUPSc5mxFJvJwNG4bD2jo3XtFTfH8j
Yo8KfdpYeUiSAyGZbdl7zipPN+K1kSpyeb61Ngg/fEXiO4Lf6ZOfdcGz45zB700Ea7biA805pQeR
PtPcV9UcD20a+XM58nrgqN4cVHrTNsmaFgcaRTUif/8AXp7PL1DFlM+WcTFGCttPByajkC+6Uxby
bSwn6CIRiHRuTY8Jkfu3XPMFQTKBcoQaAN/a92tD7+b0TDPeqa0jgVcc3VGyC9B2llcfw+CmAP2N
AJuobSwlWet/dxLM01ay4ppKaY1Q6Y+2Hdbt7jaOAyILZFItYgPzXdC5sOeq/issJGh+/n/ShKo4
53KZyFy4F8VRQdpUhY9lPHNC0wrEeO/X1tUEnReXNr7lnmLt++/XOXcnEVxvotLm1PUDNjaFOXup
/H99d0VQ77Ezt5wgFToDUVGKh/vpQH6mHZWYn7U5jx03SWCIlM9dbtxK6z/tHYIExo5T9Z8iWC0A
xSg42y3lKEUq4EIfKv5k0bjhlhZAZLrPQv+oHDNQzAb+2f7qkeCLSVBTo+AVyjx5ieWVBb3QJ+qI
6s0TkajskfMMCio2L3+UEdvD4ZYHKhJv5ddpsY7QRLpA5Vg9cVJsaa/ipzpSPvqunfkEyYHuyGcX
Dh6796zQbnqjyRGgj8k3RVWISK5/TVrkyHMUJXUXgunpSvO75CL82Nipb4h0BNaBeOnhR8nT032a
wYzRg7Nkipx3cAhIGUZqChY9m2gteEBuIjGK44tMSeGJKbDCTZ35cK8lfi+X7DKHIJlmCO1KQDya
WSQqy2ZE6OsgxbpYCjrjW8UJbsfl+12FSNCOWlLR02m8cfM7dIfJBjOjI7e+zggLkPKcG5C45kth
R+fFP+sdKNZj1DjvsOtjDCBSxM9arwb0QrvAzxfpRzuJ/RHN9SpwGvmGmIM8R6fcmI3ehrOAXWxc
c/h5r4/s7vmmRQU/h8ekiHG9nPMgO5/1x3KqY7rJnxypYl6A6lqoc/6pcpYM9u7o1SQaNm6YrxHB
/RF0Qp5OdPXaizR4EbtDEUm2YO65WYuanO0GOAGbylr71rvC6NP80WYj4DaFPTqxjQoGJ7j14v80
hk1dTeHSM8DyZdi5LBiThQHYTP6W/etb1NKkr+xG8ihv164CF5ZSBqwVBD7Limj3FpeE6tivzfJ4
KTKZNIe4k1xNEs8T0G8AexM6axaRI10CU/MNXuVyqTT0MW6UGmXDgM4v8cJmcx9SxyMC+uVPWDeJ
7UgKVDeVAHpgz3qQSyfuOYD4FchX3Ax/v2ihDsRKBxGdmOoQEejaMMxqVDvRMCWd4jIiT0LM00eb
5IUYWRHWRt0xPNZEAy1J/zh8CbxoHuPq/fRJE0wo2kzkGac+4OlJ0KqleJormVC+Q32oU52l/BtI
edslukfw+MnlyS13lQRvNXT32LjF2peQw3wuRaAIKB9BfNHAJMUoaG1aa9yGOkgPqsGRQdzJalXX
kArqTxuyJCFUqzepljb6DRt7N76XpCV01rju012hmHbBTr8hKqnMsLz2JoECARFuxwcJQDqdEm61
I8LZIoWy2LUUUlfieCacmT8qroZfmXbT01IWuIW5TKj7yH38rWG3IjB2r3dHdV9zP9DChM7ezC6x
TCUH/+15tyjY3JGZhTbU7c3AQk2we2j9i6ea1Tjff8XzPVfkiWGVLnHrBTqCN2O4ACxHkOzTxHgX
vkqv2hKOjMMFDQj7LekgasNZhAGbaR7g4tZqNjiXxF4qqXMw+okEuGxbxDH3JZ6EIImcBI4U80mz
oXxOUV9N5hSWPLHUCpIIXqDVadGhL+nL64VYQqc4xpLe5LoeBmgpscdZ35Meb/ZRTm6/gioYVLtb
Wibagb2SzRhZNKANfZqOuFBGOje99ujGI7yeCkm1ignSaLZsJD+GL4WzYJ53MpkrhJUr8c15hLNr
YeFL5UTjHk+8FM9vCH7E4Vc0g6DE6Ejm7LY4Dna9aWc7xKp4/aKkU+nQLiQbqeUa9i9lHLlf8mC3
kExINAn3j23ybVN+6OgyujZe1zv/ngS4eunfaWo7nAfMH+sBCU++2CT6IYzcAck4aNZGZSTTMi9M
lXgNPrOdUq5y3yhTMZ3s+BiWv17gUKaIeUfu0WZX0MxRSceP9yEGcU1vSRXgdpt9AICd8NxaXLt6
etBXZbQ5LWaIQBsPS7le6Bbvbd5SAsFDhFV+hRQxpsChlovoRMXpj/jXLXSDcBuOyYvbKsNGe0TD
cS+PRJfDqFRW+qZQrQwEind7FtlKwgx0Otq4HllJKXKv9ATSNHdO4RuJOZo/hJ/ndvnbGxZ6AiFV
PqdDrlfF0lv37kQRrDpbWCxo85y61k5FpwNGnxUXa8m91yXjvbGSTPqVl875fDu++I+FJLhmKGKG
w6+HM8TFfjCuGQVg91QLqnP0RVx8sRDMYKBVqU/tNOK3I+fnlSIzzwBNtg/8eFAmWrJoJFZin4pe
bikzO4Fi8pbVkfiy3VSQy4SUGA1o/re4muRcAdmm0mxkD94ZlfmL3Qpey2tXh3iTEPNnDkyhuEm1
vPwoaPsf4fxn9lhi/MpRPdWdzVTqkkQ7Rfim3NX/eRvarhQOGE34h/YsEvI5ALv6vRKtpmmEMPkX
fxB5H8OdhEElqUXWd+l9lV6f/KbAEEbpFLhmI2kDg5JxxUA/OIuqZ72zEFw2JvnyzaWEsdtVPNPF
ABSiXefIBoUmPn+dfNZs6KBK24k8lOchB9WLaydmuoFr6RTt34PwkqFOD5ldZDPT8hXb+Ix5YXd4
NzopLmory0mLDdgv/avZFJ4RI8NLDQP+owZMyGXBZLDhtUo4a21BAs230rkHsUgPigfFuZAoMZLI
kBOrsMh0NKLCArVLVfBg7h8rhT46bs5hR+5UdGFp6eoN5re3T95GJqrksBr5qaW6hLE5E9PY8IXg
WlLDb0IsmiA8aTKCb1SamPhga3hqWTGN6np/vo4JMTRFLMHlOm9HNUbmPuqfGjgI2w2EtsNP54k7
3DJ61kIPt+qo1E6nU73N2jnlcSRlf1pnfTtFwCPbB+MQhV7lNZTdk7imJXg+wFtvAf/lEpcx5R2H
XTjUtquE/t3tq9Bv7XRLIkFbGe8rBlsfcRv3Nhf3jw+a1oxla7vGljwfXGOq/sIiOLBqZo9LiVjI
PBKoDN+RPNLcqqmYIpC2m/lWnvA4y6kNxVGXXJQIpCQRREoQe8psEdXoP3cxGa0OEM1HzNScI2NB
ovL4DYX561zJHjB/5cjP93atR7okb07pu/RZyErCsWbsXLI6lZep7O+kYNcR6ropKQ28b7zmIvm4
cdLroRek5FlLrcK5RKrubPMt7uOdiZbQP5s9oge/Z1fBqA5lk+6alY/2fpDAHnv74XDbmmpIFgyz
wYdLX7B+vw7igkdtRgs2y94yVGyRclpC2zIzZHiAcpAh4UgZpx1zmptFYXFIxqNU2sXkQImEIQ4w
hMGnct7izbdBbaoEIfY/hx+gDGQhmDhrxNDrEfIzku4wnpJWSNAMvuKCNP/qprBgd0q4qIAiblHf
3tH+Yma0AEs1rwIDq2kfTwyq+W4zmXm+hvwhAvycR1sYI+1/Mul95K1RbBRhkGdD25COEN8zcr8X
015m7NXlk8g5f/NZgGgSms9n2wrYx4YQW3wKq2L6V6aYfsNWDe8cZySiriAmV5aUcOE+alkkugBV
OjDnUB4s9msqNFh0UEi3B8PpxsJFy8nv0RZSRAdZSUx+QVZVQa4+YHCeUeC3hTqeIJMR2Q73Y7/u
lYHB+ov1MfeS5Ly1cDzuo33Ganw5Lpzho6pccamqlULa7uvKUwSNglqRSXdB9kudzp4vbKR9Kymc
ZS6tkuQqV7rLhuzGzxl5rEUmY3S5YGIDSbb9l6InmtTdgYvQkhi6olYH56Ec+eCxDSXjivdlks9n
NDUUh2wi0YCyIhNml/xj9iNi8u6W6Qu9M84WKTPBCMukv6JpzSW7zyDPXAltBTiTBFNH6Uf5Xvne
AT7isI/0UJFQirkYSTDAOKgOR998vByiPK/TIelHQL9iIR7l75G0w78kFmKO5HlAofB4TZPwO7IM
bwbbeEIYoWLgMhzgB9kmnN0EBihE9WcnbvoSUK5PDcZGRWm2sNprGUvOA/RKsH53LWsWbiWiBMvp
YgXaTDZI70duP5baotR28ClIusoH3zPVjHm3a6HYRd3COlLHQueKhA6R8YkMUF+G5eX5ux7ZLn2u
kiqCCHU7Vo33e3efLtXm8Rw3mjZeTNHrSt3T0V+PJC1wLwmAaUYHM/lj/+yGLbBFbhC+bsX31cGs
gN5jUO5lFqr1vmgrZ9cygnp3HUJGicAnOnYFB94cUlf4mm1qXxjG/cfR4y2e9XF/Nt5O/+M9Qrqd
3QDSnSTZJ5748bzzZnMqRaBnOhkqnB6B4oiImrmnza9PKTdprodVMgJCkORqbt7I9hmMH5jlFvLQ
RGjyv9OAwESMkG3IEe1t7+WBKoHNc1E4SZoDDhFQbzKu+1ARAgsjwK01tY1K1yWHVyMVuesWhKdi
6SjO2WRHH+EVtDwskZX+9jEFlzeZYsDn6XxnLY5QPOmXvUPgJvopExhibG2XUJdMF7mNJvUaUPVK
WIKsNXR2tSGUMNOoG3W1Ow5UcBOuA9iszZgXRJXmmQqPODAIhoqxBsXweVHH+5bhsjqm5aaPnjAL
QCf51BcrrZ5kvUJU8n4QV5gojHTCspPvnFNU/7pUrtNJFKPeEvAx8V3FMA2jXmhHDF+S4egY7ztC
NM/A2/MJB7RqKrWdQmOWJe368CuyGUTJHADJrQWLLUgnJSEmrpgnYoJAmgm48hkz+3i3uOc/iJne
jgxKWWM2boE2Tq0ld5zoVG8aYxdD51JKIeP129jI5Jyfu/kAj8l4Wmt70oh4qy6+QbZFHPgKhu1I
ulFX2ub8ELSda1XiRrip075Pr5Jl3Z0bExi3oFL+x4x3QVSf4/81klLgEIVc1ai1ka+PU+4FkkCO
Cg9hKwC1rW5TvnSh3L+X/Fh8CWj/jy0Bp8WD1kCxgkVQABqkyJfbS8qPKgwiPwbDo+rKr8JJwop2
gxgmH1zSwF42o8s9omSScID6JunoNR2Qas5s1PcKadve1AnsX7DCw6V/9FbANM4+9gUbDPv5qvJz
gixvc0iB0h3TJpbkQ2gm+z0nbStUIyp+M5exLSMtx50Qb8x/6qa0r20T0RtZO86uqQPPFQfkSdxT
LBpBFBeSqb4nO74aR8o9PcivYrljNFoZrukcUMGYgwk46KPNhzTa7gznHzbPjejwk4frgAsJcUcz
TzvNysxSKSi5b1Z5q2tel66PJiQWgNYEXgHnL0qmkt3AW6dbMGb3lBQNKoUBHSyQeECEmnJbWF4P
JU3U3+TtyqGb9bPdvzJMgRL4Bi+D9N0UXQ26AX9FBX61hke2OCkpcmvIQKaSLLVL8H4cpYuPJfB4
w9QHm7BuWwuA4aWzRKrIA9mOsaQfmKXSpU2sf1w4D9QvFDIdzshGyi8lWi+2l2Y4rx3fQkN+ayFp
Xtvc7CLXxhMgSMZro8OPDKPf8ldw0uF/r9kJL4nTK1/4+COjmzVr6IPAqiSU4KOUh9Yx380omJnM
epM+2L2GDMtUoGFtS/L9sxDAVxxCaPtzFEBKf5mvCiJp0wz95+11Xl6zI0tJsC0Vs//COr8Zl13M
i8A7GHNO2JdV5DG4ddDz2Kt+4JY6nCtP2zXoSThex4HibUG6vznzIm5EOzzEFAgO/HMGx/MLPb8D
hxuDfqWggrFC9OabpBbhPROariuajeqQmGAILTgZNTOE/vMfCwHacGzN1b4YnrgnKnqZUh15D+fr
vZgbxnGVAvOseJpkOyc6hESBe5ZBCfeGZZMqFJlw+2nguA2alPSW1isbJ1R1QvFcpHDh1ZW1Rg/w
ai0qCbe9GsGs1+wfp+/uhpyX6J2XF8KTGEjDQG4jUNkXgBJCxfDqiyTO14GSd+W33RqtOLATKQpr
rhQTYs0LQXizC77iz137UAs7JfyF+UUWGNjUVvB6AjuzTEQIfAwhyUs/mXvbblq72PnxH03XN8JA
iZdD4VtzYb1K+50oDQc7U4nXNV0ToSqg3Q451+CQTveYAhctuh7efrMjsI8TSHCnppY3zh814WVF
HlUX5NCD3qCCD0led6HzWld1RrCjZPJ6Mcu7fc+59UlNsUK3a9KR8qqpT05RikjRwbsuO31g3PyS
z3t+V4L2K+mcHtCSzQmoMES2P3UCk/H6W93ZZZQpupX6vgYXQmi0qahBLdIbJLaraU4dAbIMkaxD
R2Rh5gocjwH9d4FtCrf9gfGQ4f5TwV1nOjvb3/bKRYBojij3QyQTvvprXg+kc89WCpeCR+I+AX1q
Wa0uA5HRPdh4/oy03Snk6okHjg+PtrzCQjYYhDMdlnt6+2SWmrJc8Fgzim4IvFFgrdFZ5ZLgOcnG
vVr0QfAbMC+tcZAX2a1sFyMAwYlKZH4FqADUFRNw11lgGyjwp1MMdUTXuUt21WwVDUh8w5reGoEM
nRysw2C2XyTTMn/luqB0UFrDqsDQhgqcrwIeA5+8CyN0kEmnA+YXeBu4XUWQ9bQuVpbXkGRtzFKO
ycDQpLHUrVBlJDGagePTvHp7dt5YzUyUh/ZZRlN4gQA5hlYclRl2LIngx7qzukHCN30cuTcDNfgA
jUXYD5S8GAVVUt6O0ekaJEILzJyK5z8XMdwgT0ASD9FiqJuTREGRIqXBhJa5Vil6KAkA9oqcz1T1
J8aqOMnB0KsWPlfzgonKtWnZXDAs/41TJyD8kK+UpQhOnfHARYWiUPWhGoqHQMte8Lwct9Z/Ss3e
rXbjdK2KwdiekQZN1OzTPfADaMYLo4k0BYhmcTLrHyDUaDKRg8rH2WWTa7h4iKxisqq+hZ123poQ
D09MHyJ7B+ALvpK0XP5iGCqtYA1FoGHkIj4dGfdzLWxr8OUkbaQzLzsgfEPYbw8efSrHcqbK+MTf
hYRBMfOWAiycFwpCvkhGNZbA+jFiPRgZPZSjNfL7BbNhkeDF26awlX6tT+IASihrOlpIvErzCnEN
JLCop9hpVWdAF8kaL7wRYgQN1J9qQNUg/RgEoIHyTPNP8avEOWG6/9psUakLr/a9E038RZweaCgy
LnRvGd9j7uavF3T+z2Una8oPXO3tPwd/gkti6WMUqtwLVy43mPkPS3axr8ZjTJY+OJ9St774K+ur
LHWy8fuIL7nw0rdZl/fmB5y0I+1t1ux/B9iGvWVn9jCyYR23zxm+0NIACTGj5AxYBUOUZUlJWq4+
TACE82IEvajMlGoeZ8zhieEbjZIePQ4ZaL/DCuwGVZujrICmNVRnQWuOPCrMpb3PBhHlBn/RWSL5
FtTDwz46gG7C5K0yeHqg1wuoTVmPmYclg77x4uQH8Q4vyAemdsoWL39eJdOUh0SVgFRhB296MMGn
LEn/oXE9itaSuPi08taJBf21Z0eIjVFe1hnm+FlmhAYmlvD0A5S2vNzPSTrCgcF64XX7gQ0UUHU5
Z8RqhmtHKf1cD25/kvM3C1BTtYHcJB0oonzRHjIPohv4LDUQ2WUAvXDu07XFXJqR4LqIK+TKPDUh
2fdkURS6K+9I5VuzyPCGxoZHNsXvd9REKmiCmdSwDaRLrPfCHWLvpyElFEFTF0L4jdpscmhueOFP
/nCXJLnbn1NiSgOqR6lgLb87YU4WyLXZFG1MiYLpiSI+ZNZTTCFU0edzGxVSE7fvIgFwnvVK1ndh
lUCh1cGsXzEA1X1jWIMrGZkKIWR8OwLhk7HWdAyvXxcwjhC2v1XwgHVGB3xhxFl7zzPj1TADfF7+
dpPBHitcCQqe4FwldeB6itKpAjf4Rew7HpxpiQFCOCQOaMPZig5IeSyu2RJNhsNX+mlqbNV3gK/B
NMqzj4JVL3WBgNvtrahoo2SHSIIxTLc+AnwYLlJUMXp0DYjTJlk+WKHzsd1VXHIKgNLR70RJ5myy
R8P+mEdFUkto6JA/k4EFASleapvt+RtqUNVvvj69kRMC5aDwcpvd6lxLmCGVCQSN2A8BuMFJU3Iq
51j4dnphSbH9qwcOOaohNFZvg5CAF8h/B5mWqZ1nqpkCGffWNRi9lCJAmG6FJtPUR/6Xi07C1YiP
q+/Ox5MnYnv6sKLi7Q1whJKfvHtjhfd6Xakk/8nZmx80W5JCip8d8du1ml4N77gMA7D+LuNzNesa
Efq5E8XPHJ1vZThYqiHD8SX34QN4iUn7CiDgR/pgyDOPhZBl89OjXlprepPLhbEwTEacQdSKf6QJ
H36f5bxsDXRizNIxUm5nXKFYRVhANzvYv9YaWzKGPD6J8Ah4lnEeAHqiprYba6fes/2T4xNmXaLh
HA1gZDhSxvP2s8Z1oWN3oqvfxRiLBuPXzCpSvl+25A1/fjbcoLxnCeuweo3P4ELemln2/cGIuLBq
OgP3XgxpdVHe/vGI81HENoZeEQKhNe3lksaVqOhDJLNP41JQzrLax92pbONi61xyEDZ2EzyUhprL
IWqcGsbx3lnU/1lH2FE61SK+COCLXf9QnPIs2mEeNt6rx0hy+leYvahnW+DfJKmEN/0Xw8XB5lqp
z8famy2tEscOs5MJH/7WhiuwJdj+C6uDFGHK570pH7OpoY2BnvWlqA8eg0Cgr+YNz1yWY91Z7VEB
kY83vpr0owbl3p5QFg3mX+EKqXI8a8/5ev7vvPsMfrbHOvTHLB8g4YcO/iReqQwXBAAlo5xKGXEg
lNajmn/nVzynvDd4VAyGTK2KaNTACOn5cHBt/GuexrPD3EUKm/VrSpucNZ7umvPib9j6jDi2ycmg
DOcUfkETUWlvm2vDHKd+5QsHiCUJGb1vqSKBaiTCdSaSHjpTIEiQbp8PMvIVfjKKeGWZh34HyVK5
xE46Aw/6T9RNG0GY7OPj9gmLy+HyBdOH3Ta/LFlKIHzixjxaprB4LNDEIxct6D+JsehBDQ5WJenK
8aABQvVWBCOuqChu9Znr4ic9S8TM5Ie90gGdRcBUvXzmBu7nuxlt9jkESfJ1KEARkjuQnX8VNAuU
SNeN2cnq36ZBw6njO4LEN9ZHLOx5QqNwe3UX7qrc7MDTj0pS3C8ZoDba973+s+ugc4zpggWeuBPR
12Ia6dZsgmTMuj1ManGf+FM067YlPMbfIPWjNnD8FpDKzyxtl8/F86DyLFFrDIcJnZkUMOrWBdpF
zFpwlsVTBHY+N7ccJaBreRpQxB17T1hpoiljStf7yaqNlr/D7DJ5h0+Pl8mnYGu3E7SrTHjxDPh4
7HXvqDLRF2DCwHQFEUt/GxvL2ZEK92SbkHcAIAtZmzIFORVZihqABESqOyPENUMctVfv7DIZF2Pa
fjCA048FObmJ7ix6JIx9cal7wnt+nt+M5NN21A4n2fcgyLE7P4byGf95ogHtb6Ri8v5rsEfqb3XG
S0YF5rJ1+xqT5+Ofpr0ZYODJqQQxZcO8puFVHrActxmMLVDHE0AKCtYD7J0H1gdjgk+v0ppCZYsk
XLzJPicNRrZWSjQYAc3+rI60m9tsUn1kb9onddVuz6eshOYoBjJDdQHlm0PlLwTBmyIFKgrbmun9
hyOQuB5zhMNSxjtiJichrdEf2y4zm8JIpPmGn7Fq1pTlwUBkoBVrpo2/HVUVfxeig1Hj1fp+S7ni
CK0QeLTLLHEvConataDWfD3Zcmqb2jZQFAc3G18BiTs3D67DRC3Xf+g261NoLyMTaX2/uaftP4iR
l0q4NyBgx4VbMhH1Xr/wLa6W/3SFrLo3gOC6qQQ9V3Gf3kDI1fPqFL4z4qfxyw5wqtHOwrIppSwr
XntBY9ry9JtdujBApuIQ6fTpWbU4z3o5XPpgLPZvWewnMYa8KZcVdvNy2Jt52PZDRwEIQfR8ggWX
ehiWHM9t/ekGGudO0u/fTZ/zN0+px2p9VfUSz+l/QTn2acnar5YZt3IZgD0iqEo9RiRGH6Vtcxr9
27Yn+junNPtDPH8Hz7/E3zuEUg6hONnxDPeTdLLcboCSDTFIYwxvoRwLf/344wUGaZWC3/mUbg+S
TH0aAdXjt2EfrxcrA0OmmEfWmz+PfvHg32QIQ4/DsZmpmSnZdC7qxacDh+bm87PAY45rTt+G/Hbc
ZCDeUVp7tHq3hN9rcqd3cDJejuDeAOpSnZHTFVPHy/nu3ya17eoR1TYzrR5r9dTZtB2u7SaN/wAZ
irHaEcgiqQoH1ITVfT2lZ+Ar8WJoEqHRW4CWzNTndCNISto/QauMT9oOGJay5bV9b1CO32/vc5eq
pVXUZatijAA04OQdoFQ8AL3LJrLf5LCsxfNrJJh+UPoJ4oRmJ2KYT6OVxd4/H2wFwSJaNTx42UE2
F0FImJqoJUENnMDz04HhNRqB4efapBT1Sh5nbhvF2W3at6pUGw9tGxAxzyfiujJHqYBzUr79uD4A
Pr0Li4R/+lI37o+USSk8jjAljcxZ3ybdBndQ9eNy3baLnfVKFCku9cjZMJMqw8w1QVWdaXE1+pI7
ord9N0wpWigseshVz72rwUWmmJDcg96QJtba8es+XRZ9w+kQLaMR9KGnezOfqTcB4cP/Qa+jBD1Z
X+nIxlEw9vBqXezLDSwoICLdmxGkAWY2a32X4hL6MIwbjOuPnC+MxF2E1pFz4orPdkkcyRldOO0X
5bkqbXzRqJJmqECeVFwvVfOlgRKaZ9p85U2OlieRIZxl/TJDlItpk8HtdxWD0bQDZmmuLLvVwW60
6UGIhYqZYq7NAQ9+c6p5hCT+hmgOcWRBFvV2g06mUUz5JzeuGZ7h0LEyJ2ux+nC9e8DigYKK6Y9K
i786YjynjS7yCrpPv0HnZYYy8nPD9Ur/OH6TEfSIOcdZ3KiSiVoe9cK5JGnJcZfWUADoAtbXfpp/
cs4nha2ZVanDF2hJFLwV9qs2hjYgcW0OEzurTng40a6RBlKsZ63VfjXGu8y8RfRv2Sd9KFk68b40
f8FOxn4Y1USKnSYQssjOnX7a31YAdzcaYzCOevvfZN/7NZAhzkso5hiUEOPz/VDOlKJNmfP8yxDf
eqJyw/nxIn2frYiP1+3MpgEkOygNkz3dpuMSGYrA35BVyVstoLRolVZ5tQ+8YAoW7pGkMkYnWnGg
fHlqOixyrrv7LJfnKHO7cs0xBU+htBpSjVPULDwlimGFGeJ1US0ABN3oU0FDRY6sZkcK7kE1UWw7
1u1keSfZE4U6BX75h5lgsDb/N45ms3yFO1oOmj+aGsw7YHj5ztESDIZhSgH/aMUgUXbRJjAuZDwm
IHOXP0i2UTxd54UXXW6iRYFZiST84YRXN9FRLUNevfJKQo86yY5hkLE3FXmB/EFhPjxJBdMjTBr/
stRRb238TpY4FVBu2Y5nP+czIUSSLIF1vr3hAwmMq6TwL2NKQwa4ur9a495j7dVrVbWNuQlhaq6+
DrhT9ctT50+RaTyY6Sn7UBuNG8vzjFNL+stgSk1PvbMr2a34JSfDOwrahYxTmucYHqXQYB4uUvab
yLanX+WKmTV1tc4UvI7UaA21JzpqmNtp63cBSeoSx+XCVWeusAIgLkShi/cnaZLnF1FQWIv74dtf
Nj3W56HckZXOJGxmu2QM4e+pdBGGJYRfqdH1fTf3YUnbuYOrV9dd7WDbmHp9O0erWPG/jbBDXB3S
xqvJy+yi3sPm4V0uCw5JzjiG/KZtJRSh8QQ30UsOkl24dK29sJx6uZjbuI4BKtEulJKdvIz+U5pj
UoK1q+zoBgjGARQwcOXE43TKpvDhKEIsS58pvo7Kg1ggfTLXiLAaAtNzyQ0KFo0MRW6CIEMrTDW7
lbke91D2bdUG0NREjwJ7bwIh3gQfhOeDydPMGTZ4Gszmwv6o223GSI3oRvlyVCu0b0MIX7ItJALb
JimRAVkw6POeUBsXB/u5ino08IxgXser+dz5eMxSxRVMMZy4+fDBa/OWNo/yyiTkQae8rclLbKhw
KnaATnmvSnDL3Qf2uB5sXsYXcgHLFcR56WdGiQsHt6nazNyc6Q4H1J/JhXsVNBTwfl9tREPLpOTv
6ERYQQWqcf3XSk80S18/3po06AZaxE35IHTlQseEccYRDHfuyMODglL0RPTd9znO7Qwmsise7Np/
/YYY+VNs3gPMU1A+4S/l8SdpFjeMT0UJmaWijlR08Z+4F7Toy7gmuYVcwd2ZJJwzuo0/rXu1e7cd
VGooC/JWyWzZoBJB9sAVypTlzDgC3JnlHoHzdjqVfEtJbvWrBK8cl0Mw4Szl0vdH0AxGMJr5RTr0
b2m+Qe6TYo3hRtinfDvuzuwP+WqG+BnKEQUB9KQEtWYMGTsHoBJTN0ylBIgg4QaBFgx+lT4Yiqfi
W/bCIUpIcwVlR2iGKU4Az3gaCsgCp3S8VqoVRRuO2lB1lMjqkRy29Lvz96z3MCPYVjQ6XlD4gt4H
Qa+8A4HeWaRsb0ZJK9Br90XA4bJZOwXnv9f2RToUrCwBjTz/gIanLjUlAGsx7q+TYkhJBMHtdCpX
UR0nfds/WRIcSiwJmf73WfHvLWv4DDMl1EtzrFDGGVIaPVkuXeUcNGD5wYMwHVMmuMG+ziAnr6G0
Ipu0Y/57y32xqAdnC2/g3AUWAoo0+pUGsedlgArJ4/+HebZjHDAXJMaVjcJTj90WgWsvLtzaUmI3
wtoIGDMDJZxg554YHv8tn/xc1JEXHy1m14jC+4AhrpZg+RfaPCJ2vHN8Pk1zekM5UDoR2VhkNw6n
3dnlknaMIwtkLcDbmnsWRLLX0p0gEJCjVYZLdpLbsOharjpYBZwm+5wUZeP6W4ZsA2AYra5+AZ5I
2Yy1kmqfCDeQsU1rNacv0g1AXE7sBQScbWSBOBCEBsJrkjJSZMTDxHe0lQGQqY9oBjrbFAQeKL1F
ohWVvdUc2Q1dSeytTy51w/pDqxUum5ExavHSZpV9EFsCdYz5RsZv1aM4c1KaPjec2qx74VvqnSVj
YnCdyK7kRtZtN0TttGafV1PK85EHS0IVhYA0McdCl9ZL/wA23fx6LaB1BtUKoEBUKOdyKre/dnvD
upA2HWtiQ2Qg5+9tALFcgaGepmC3xFJBwShkhEKbVcAFD17RmsRNhmbmisYELI766ehxYPyYBtZ+
FprJCqP1BsCwWOosLUgxHUTkPtqo1Gs91tGESxpMOck7qr3cBpHYVmRlyt/EgC7Eagl6KP0LjYDm
jLcQCCZAhqjvMLnZHybhJu9bfmSyK2kGqq+UGZrEl0QwxIA9tQyqfsbxG4ihEgFdEwRbmFe1ZSVR
Bf1JnBre6mFKwJPhQku+gYi3PUKEizgZrpF3koLXny9QCX1JcZSvB/UYyVRFKvcJJljQzjRuO3LC
A77xhJKFDkUrIrrp53YDK4NKOtAWGHR05Ms05kMW84PEAki/lMomMj4p/qfj6l7eepixRTfj//qU
qPkBCCYHtykSao+ZK1AYAHcjAWoQolpkZ+FRewKSlgbKzK/8KRCgnhsgjeud/KK+9yKg32h2eCYI
trBvB+0MBeacyRAJ7VmBwTXT7BB82L3E2QTRyOvTWwrd4x4jb9dNQPGH8EgvYli1QBwLAGNc+6pV
57vRL428S3RqROrFTGVpKgT9HGKWeVkl2eMtO6bvjsv4usFRwVo0HF9VhZcmQvzQuXZetF+hHXGA
VjcGdg9AeptZ+FYv8Epfl9GnVCgVMj1rJBY5XmLl89gB/PpKg7cugCdVfegrPlG9Kjio/F+nHbva
/YS7NEXW6r5WDElhniv/m0lnNr5GXmcJuRilzsbwND6i2hRaQF++LD00C4AnQ/5YubTUwVQg8On1
pgBPgptaBQFzJUiswqylSSP9ggCcFKpHHrDcA3sktS942osbFrIP7G/sOrf1QL5dVFE9hiFkqSSC
ThByuthJDRJc+K41zuy/KvArzTza6dBPxjQkKrINJ/6ruXQUKyasY02rAfEjfaHqrd6GH6LzlGVk
+2z/icP6eWNLJ0/ghG6UH4UvcXLBDwUZ5IX+jCEsN/wFGl8rN7ISOLaLdkQR+S8KsdZzyAjfttwO
klKZlygsHQI6hA41UsUK9KdwYvBq9QarsYn0McDFPCyJcCai7q29NP/stmNBdp6C+Gzzo36w9Zee
rAWoZdx7Jtzt+DArVB6cVJvCaK+OkhLjX92sDVYFgCE32NTC+1IKSjn4arhwmiMSb9lG8f6Ge2bo
0TvXLs4/VQ7+BwIDXLvc6YLrhZDIhcYuglAWb1HFt0JoMkmTXjA86S17MsI1aUCk0GjcrH9zWkzX
OLWEv/g5/mJW2NVPkZEJNV+6YwM+3hLI/X1JrkT1rmJ/aSw9FtnEf6SF4LyCk8tuslvmHP+lPZrb
vS0pcR6DwGfVRce2coAZiZLdXmb39XuZDDjrFw9yXJcqisoN5tEfBaVXt7D4EbBbGYvgGrLnwRjV
RGZ08kPgjVPNnIRTG+Hx0UrNFqAqTQlqBkFYEjj/GY+lWh2h/qaecfNrfodNtz3tHzzDuD8pqjEd
Xz2CtdLsYR53yMklKas+9ds4n8HAsxHaAmVgJlBXvw73f2rgh6eGQuHqG7hiPsQ451VWbwj45OXy
hhGdMZUVksKFnLlJd202gAWb/j5AoQ/EDcDqJr1VWL87pfAb7wK/bbrQ19x18B5o/C0yZ8BimxbV
kxwLuw2ZFiMmoNIzfLOwbknoducEoTO9Zywfkk9XqAG9gYj6W+56/ki85nH8HgnA6YknK96BC0CE
3TUlwrG9S58Z+wpdrCSwRtTVp6Mz852BdWyocszAPlRb+DTzKmhs8NB1X3d96DHj1SnSJDWahKEt
XbkNXkUSJJZE/5gVmOPj9hQAkFwSoFir7iz9hZz6RZvIwi3KAdOPCGl9r1NNzS++uOymgP3YDRbd
r/ltT8nYHZElEQ6UlbUTSIUOWa+Ktwg4ZFcNFxt60OSbvYueKZM148zRL0CSqB4ItOcHxhjIcYi0
sRLhSbei3Ewrx845/4PEmO8hnG6IAGLZKoJKyERaXQoy9eZfZDhbZx43L6IWalMYnXxq0xdWN73H
I1BVANWmcFu728JsXOdPeBW6rho0LM/KUnK7cbSkEmjCbafFTviszMbgvKoloiThYjvp8wh9WTY6
UgpzGuijhKQ92X6mb5inj+NMh2v2+owVPdXmOd9gE6Z9f7NXlRQ6q9n8yGbp4PuTBpG7vWq0nxpr
nhxO7dMYDHKNSOoI3Z0jzdsgDFA4Qt/sj1h3JTZ6IAHeobJhUDdFyf2Dz6EGkvzsjx1e6dAx9VpZ
KjT8nsxQDBT41rJPKqgVMPOU6IkiVf3eZRW6m94sZyQ4fY3wWM//KAWFJI4gWIhlLW/nBv2A+rzE
qoHHkPTc6VHfoHZKPySwS6f7iTIPxoNDpr7Xbgp2H4jAuF9JpsIzfdxWAfEh3zoaAEZ0FmWF+n59
4bD8i4rgPup4TlvVNO8fYiJboJfcj+vRIaOBPR1qEMU6Mj6gDof+Ydl07zywEIBPwIa1Nwftm0R3
Y3BI/dxcQ7w8GaIxPo7g8EwiH+v8GE7YXZW9QSZBvWZfyaDqyw3VWnYJY3sLbX6HrsGFNap/PBjs
Kl30eWcQP6amCg0NlnMNsxRLPhtMsLFC3ZvIIOICVIxnpviTyaXAITj4gJNkalS+gK+YTUGanobj
nJ7yCdQzoOSP4004HNswuxeP3jWbJH6OsKgXjWlnkyhkoJDwTyp5unVhPkwDrd+nLbDk3f2uvDW5
4p52bNr9Nggn423gP+hsn+XotoTb65tADwPEQKAT4kfAGb5fawVaT7UwNh5GqkH5A7kpmV8mNNwS
wPzIyCRjRqyk3ZL45kMwAwffdEa0N0mPtKN+twMQOeVErn9I8fmjHqv1Ra0JHGiGe32kTLgUw4mt
DR1TyNcS/9TUdBg6PX6aIPqT/Wb8JZjmaxsFs3KGKA8PpZSxQ3SBlYdZgwFpQ5vC6yhPl6nL9pqL
pqWREP2EHN7vjc1JE4cZoI4zv2G3r7Kox/lXxfQGKoF4A3LC2/Hb8S1STj/pqUZ0t168/JEyjeJ/
6aRfMLhwy9JpBAHPU8wQTYTCBbxEzbnsjNvlwhGxT8gFBKJNUdU4FNoW/oY0hAqpNFdi2cvBMKJ1
sUorEo118YyFlM3DDXk9Kfq6h44uUJiEWOqXlRBm7RpCj6q5VPawTi4rkhFWjAfi6qcFQhPOrwYh
sfupV5JsseoNJy2y8T8klkUxXqL30VnYrd66OSiznoZUsPN+YJeAlMXccvAnq2J/HkACA9wnDc6O
vtu6MpALNkIIqdd4gk2zUgyfYCaqhkeQjOAwRmLYqds551TqU60uf6HxK9T5YhbQwcNj7IvIsKi6
DLwdRuTHJvjbsEKoei81mYs9QOWDLU+GwtRBHN9fXXwEal0ejB+pLOYD/FVMeXQH/6GEoxYUo0zK
pgKgF1eMhirS1fKn3Ep126eG2EtAIE5NAnxuBjkXWTKa1Jp9Rz+P3r0Ww5DKC9j7HO7hDPOd5nRz
qfDFp3EhyZpNBEoWrLOrBEqxF6gbtFqOqJmc1r7CHX8aO+AowrqZ+W/Xw9BL9ENlKs6QGVKD/QG4
bpv2HZ0oZqzEUxLMFTBfS14e1tmQkeq7RKL5gSx9gXHu0p4Xa/8fJTiBl2VfAgtAd3K+DHWe2pNg
8IyuPx5eupQN3bUMgJpeKG5GgvbHCAP+g21qy5PxnJ4VLQh850+BtltQ0C1VZ87QQVJLf+I9mEXa
HYOyKCAJQ5n7G9+uNPzM3JJm+KNubesyZJQm6qtOBOGEIK8bV81edSm8iQVpbSHyptKcGUBf65et
1qyyEa3K5zA6NDYke6RRCeqcg1e4qH2DOA8QOy3Pv8yRyx147COHyIgm3Zki7vxNPYpYp048+zmm
wh2f3tz+tZ5d5K9/ygf1HS7SYZStl5nNww2ykJ8x8OJ3pS16kcodAMbuT8qXivSo6Io249DCx+y3
xYabGGh9FhbgRwVUn0ccsOIszbczWFHndyrOGAXMYgmlbuQx6Np/TvyEinpitZyv235/AuH/+u+q
BUdd6FU2CEBgxb71iVSvweBAgq/yTZxEId8C3grIeLyIaFtodt1AvAJi+JcVGYwALSee5acwcQvM
j2yETb+rfRSRz6APJh3iF54K6QP7BiXDoKrkOiF75MJfdYR6fsjBg0DpLBwZulvG6/qSDl85Ov+l
GhSjh9nUudde0m8ag04ivAf++ZUV/L+te/tNl8NEMk/RhF1XK34R12m02QJBmC6+t9qv6D6Nva6n
v1zjoFMo925bGiEwAUSIAZxmTmH7Qot5pZglkSRZgf4oe31redy9YR2MrKsJeRI17OEPZ1CbePi9
qrpbuDmBMVSgXeL2ffuV20ToIBeZxaRwoOwdpTjDtamkTLFHkzg7idhU+pOLGZFTNZ1p3RNasgzJ
YGYWJBc/zZQB/ErznLFPoedbqu9T3bBMBb/FicehOhjqf7Jb4ETwCwy0Oh4Yxy4kp/A7j2tGJ5ge
cQkV7e0bvihvcf645ZkIfSx7tU7GAbQcxJ/vOx42NzXDXs+R6vphiYTYcwRIUcd52LMaDmtBCMJC
iLeORDZSW0PUUyjSeH2Q464a/PIbR2kCj6R5hW9YNBKCVLjoepTqMrLgWDikyduvNrp/gH+PnwOA
aL+2gv6ra7svj+J9y7dZJAJpeRENAyyn05Ou1hEVHtS6cGawOPx2Zd1gx4BD/l2zZTE0eaVlRdBE
/SDFQ+HPOMJ/7gfWhHExnTLJriq0A2TRdgC1L1uCwl8T9ipV51jdD5VwGg0QSBhpUhhHohnK2yyE
T+72gwcUPPSlnZaKJu2aPOqB9ft7jxV+BBd3s6qLR/eTPyGIYEOCKs5h5IIK/n8fNRjPpadxDoQA
RoHdPk2JO/xX0y4f41NzfO2wM9qwETe7ZSiJ46GZgOf2rv0BXz+tyKMnejNFMg3mn6hXvVFINnm6
qEYo1+iSR6MJ2AfcP/heFhOqA7utvS0HR7KpCr2U4WV2IHzB7SbEubQ8DMdSJ5ue18b+PXEEde0p
LuQEWHdkrKs5rLTBazCuVAWNf0nC8mg5n3f5iUFhayD8MklrtBOcSev7EajztDNg+z+bmX+hUqqC
2dr9HTM4RA/JHzL4BDmh/znnYecUVan4DIQFGLB6Z4IUd5mv9zDg4DXmSx0qSaPtbeqOX4IwJiSe
+cbO0+iU7QN5rRrmlsqtyyeZiCXrYBQ8LrOoVgvpDthJMfNXYkMfyZLNmrrIGEPIAahvGhwI710Z
Y90FJiTHKEXyaeGkozWMJh0WTpNdfpZYK1MhWOtHb6LJ2e3P3tHBtRfm64Ok7aq4u1fj9WE18gez
psxS+Apr6YWYO+Rd/R6YLy6adOS/l2ouTOaGQPgF8R9t7oPfrlxZNsC+1gGT2rpX4h/3qU1M+/wb
+sDk+wOCbAp/JpDRU4BSngbSvK6TqBG01kq5NYcPVQ3ZfNBLzNlH7Q6jBvv3gpN4bNka90lHeqh7
KOaqytn9rGdSDowZL624L9MXI14Lm3yvCGM8KSuqOzU3oVPE/vbxbuUpU6kHo03qdk829RqdOhQD
IkZHTeWsJYf7nrymi3/m9F895drRKcmnubQXspm+L9OvSmrEJO55jsJpCBKYiurfo2Bn41V+SL9Z
fKlRNzBmrkgwR4XpHB8M/TmMBh4Iv8BMbw4dwW7ZCUC3FixpRSC5I9TRNHaKEmmbHdXjKYRLU1G+
AISQHlA00WGinO37p7UhNpXZSa2cy5M4Bg7WTjLJrdaR74XTmSys59Cr3UJB3XJ1v/Lc/VC6zzkm
hBOP4bGNpgApTdqkij4QUz+uCx+E64481cZmkwNmRv4KFU8YuVa6W38zOq8OpWdW8EF0FAjrcOoW
ioVP7Y50xgX7Q6CYqCemWzVq9EWN0QXPqzuFqpNgRgkIBck7CsNAhJ/VW5wmiTFUEI/fzxRxsclN
oNXwjG7qT6sfm8/43qn4C/JeGm3oCeTnk7Dzhjw6mIfnYtoxB0ILZbRr34xUFST7cZW1eYQcwTww
rQ4NQy3AiiG9mkI3wPI/QrWp8BytExZ5CTdt5Vkf/AzqIoANdJZlJS+P81/H+oAuDcw9fYPfkja6
lrtvecieUt7J6XAE2JsxK6q6DBZoGH8mQt9RvGvj8MFEU37uwKLQHXVfrqVgJTsEHLta7oP1hVkR
igPYRL1GTHsn6EX83ZZ7P8xTBWUjDnkni4ft96lI1TDzmlhKGPssPEJE2ZqlmnsLNydBg3phstEE
8PKofL3W3Gj6KbK2oygfqRBRtSvyfZllSgpJwbI/c9gG2HA6/zJSuVsgIZtNwYVA39pZr0OuHFvD
EyCwhnjGn5P6reCx9/99kH4SQw1oLSrVn+EVSEaOiYVbC9NYF5GcAQWTtv5wYIZp1uHRK/FkR3W3
6mjMrC+73KZySmm4ZisKzLLk2Ygq3DuFTy/kbYxF7r7bVG0wvSpc1D2fYSddQ5fpqdcL+UPNgBo0
hLTPW0Qp8Wcpo9H2LwGCiuqKkaNwGgaXw36xRgmRiniCHI9CJX6cacFbFtxgZqGEtgPuPUvK+2np
uzdwGMl9qn9ztDxBgISNjIxbOndr6ggFoYq0lTyTz/0MYmQcAnaiPk19Dl46wqs99SeXIRIpDm3X
mp/F/qxrzPFRxA0gkPPBm+KxazyPOme3U03vHm1XfbITu40d+sBcdFOHqJnxkZe7KIrst5tFv91S
0g/hnY2dhCADzbS82or8fkdzaxRCti2mY6Fyfo6uknnzFtGv/f08P4dFXtXGaqLzLXDqsI9MJZlT
5vsqn31I82zWHJKCK4lUyFJsdcURAtyo612F69fwyp7MtU4VI/LXMQFD2DZ9MUo9ZzfvXyh1y03X
/hsTNBXsu3Pxdli6W88KiNx/ZGyKUfw/JWzD4qNH8Tob7CntBgUHXQ5lEDB+WHZ3+dMmRTlJtFRM
Ki1rzsOx7qp+pNgdw0wNrp70v/Ngc+JvTrfOP0I/f4lrqq2P+M71IoNlHldDICC/4bxgsWsXG1xU
1ZTmiSINJHGHxLKz4z5iVm9xErOkV5cd8vTIXyFKbfzY2BGC5JUKNOqoz29X5fTUhzXoSwvTItBG
o0U1yusOeIhds4wW2xbtAA5+nFZMRlraieqz6QKFEMVz7qxWrIe2AaLT1Wd0Mh/XipKeWT6x5Nji
pq3YKhnneXS30g1bshG8yf1tKu6N8DO8XSQ8GT6oQHSz3hWgr8fuGd5xt4wV4rbEOi2WKChX7rb2
klqmsswLLQlv6xLZUIHX0eo8nQ+ILmcPpoFNVl6aAhMt4TQuGKQEElRF93MG10rqw8FJK/1b3Hb3
ffTeybMbk6qo5T4vWHuVLKtwfHLauYto7prWP3pJzOsAZkaPZSZNwzf4X5/EK8Yym3ObgUzeyw49
fZB0MYPoa3EyorCacOOJ5r1vwY/JFuaWRb11z7/6vQrBGXnWkZVp7z7LTABG+VDVYJ+K4XWWsQA/
CQsfeMVL/OBXiROvJjT6lhwYCOcZ8mKoE6ozzryRn8OdIvkAvrBueTnLvKvqs02Cwhu26Tj+etfI
UZC/Oge9+C6WtOgoESXW4qbF+t3ft9rTn6AvsYw0SMaTjNKJgoN8LmtMQSJXAG+aMFqaKdQ5qdvo
3lfwQw8IFwnUksSfMoOKVMlDpyCRSC9qahmujVznPZTNAAEU0JgsrNOB1AgZnHBnhFM+J8EqZIwj
vmSxEBDGZLmoP/SzuuTPpYq3J+Ui+nNdl/eHudVGAEeW+V373ugnygiLOVsSlrMS7NuT3YNEi6Uo
AnBUlrh59PY2QwTdHmGiM4mkpC3PkBOijdDsFNYsg0xpUbfik57P9vApbWcUet9LcggiTmUwOqgx
8fNb6UrAemehcewzqX80vCU9+ds8eM3FiC49IgDBNMfhOuGQjC39CbKRUQaBk6oRcP4Lph9Mx22W
9vvjjmPpDFc5ur+R3dLztW+N2SNCvoYCez8ff2gxj5ubHb7xqmZNeA+p1cXgymD1ucOBoZLKCifV
FSFhiW54HSOztSTn0U5hi8k8ZQkDUl11uafCiWVPJaHKrwJoQgKjJXKy8eG1y/ml4xm32t41KraK
RMIu0NQPe6Bu2x2ViwGRONgD4BFVbCmSKA0CK7Mafi0CE8LSYteIeTr8z2vPEYFeb4xSJwrRhHjY
q7gO3iZ123+eWm1r10jgrg562MDYNtylN9WCHPZ0Vrlt93gLY8KL7erpvCSPGEANdKHHUIaDA+oK
+AjW1lFnYQ+BKi/D7eaWWVhHqTQpKjNUXU6PKRRlaOnWv/9LWaa4QH6nQz0CtleVxUjH33SlhXTR
/YJIUBYBM9tB1Tw9Ea47ZcoKky1ZBes7E4GFJO8WQN0iRlMA9TK9vKpUXTfCGH9l4dkEQoVNazI+
uEx7+hTNZ2HtMBZBhstEFwNRbGPkzKLQhP+qgqZNJSMI2havcNvaMjGAQ7y/GkEF0yoXY1DB6Rf8
l4M6+GknpkAEszyzIiVmMPi0lH4MSXVr1YNfqC2p8ClHC+vdK/4R72OmlC1eCrBjcg+IfMbBLHBT
FYu3Qja2PfxFo2WOhfxUQojrvuXBURUUZWoe61n3Hq+FdGUBT2gBHxMlI2AlMlv9UuXrnAs3qEDH
5q/61Fl1zbLZDO4BJ/t8m3apgxnynRdEmZijPeOE1PwyZkohFuBQO+Be1004Ir5dOqNSC0PKVIY4
5p3Fr7pMTOjx5KIcH/53ldodNXJTaRYGxDys6v2M++PyixDe6+POsPFHDzKZfCYb6L0izB6oLgOI
G9FrXDNxWw2o16VrLVFZw1ewJAxK2A9cquSXAuS89pQuuYEp1dJA9jHEHUrTAFmhHxmC/kLEfStd
txrDph1aUb9LxwWyNtfvCNWaxvdhKY4whXkJ0BYTEw94y7T4U9Htc7/YhAIQ5d+Ho8T9TourXUmV
XPtj1ghi/Wvj4EWMsRTW76ItJ3+HSXA31+PisQJ4GUK9TQcBvcXn+Scs1BYPOFCqu1m9rlcypwkz
6hV5aP+ajaicQGAWLICs0RUoUxbfxf3q0+OUTc2T35NOUCwbigL1YVPX/APWSsjGKeOf6zmOAmz0
VFXs8PPwTWZXTit9deBaIzU7ZsBwvRoq4svpszshnBYqybEh+xEr3zCTUwaAOGTWXCH9pw5v4ena
keh/fQk03PcM6nO5xQjxAw4QdqyAJg0jnTFeKk5Wv04zFSP5rYRjLl3BJKIgzshhEb3xRG8ugbL+
T9kHhPG2qNQ9cVp9MqfaCDm54Q1aQQJvttsVv/Kr7nzAzcpm4P4ymhQlNMJPDx+9G90VF8FVvjZ2
fE50yBU9GL8lmhHovkN/zyAuW8nANaAe290DfbNogf5O+T/THEVZBokfK1RVG1zWUYxmDDmhTBXB
PfQ3qHDBxBF7Ew91AwXO8nPLh9+LYSaAPR+JEbTN39+V5hpx0AFVXQM1t1Mh4j+C4cVE79rNHgr6
qlCXLVh6sovHccwyko99vOGwlhgLKki219ByeS/4JBTbREM+Lf0uqWWNFqce0Wha76uZLfGbNguu
m/DebSpVkGzcjqn4xLvDRLImLLKNVpEra7BLOGTT4c/z7Ero21A/Fk3BRP/PuvqqUSgJA6jEpPYN
2Uf5aQzCwqxUbEHmP2SwgQxgc5naTWDX7c6jhlUX43XkeUUbjMVSCaOOrPgm4o2pshTJp7SdiSZM
ZKxBRAUpUiGrwJ5YdA9q9mKwxI9rAOKeObUzBqNADdVZVcvf9u6u1BvRakbL7TwGhbCtwVslHjJd
S3Rgvm3Arei/0uWekYDgNq5MFvyYyjt0dqAWbRHueXm3ZEh0WxxFwUVq4k5ok2mcIOcu4oYOmd45
shbJMkfrntdYzTafq0bJvaMVeF9msmwm637Bip7WffS3BxkQjuI2JN9r4Wl47H7N3H5XnSN4C1t+
tNvpV5j4lASEyEP7Jb/9qf06upKbT2/EtwXLYMj9B8lGa9FLQZrWbIO8KYqIGlGYY9ry3zLS0/Nm
z+yE8aNzT6UKEcMHLLiGT0fhAuwjbpRjI8IPjwQ2XuoL4PLMO/MwCcK99hFVjiTArD8sb1ck0Oad
i7V5iqj7iQ48cHSzZbEHsE8I1ossYd5Ps2p63V+UTweDuaHRE1dC0r2+s6qF6D8A4bojlo1A9TZ3
PzBXYC36qF0bD42TqJcic8bs1rMSKoXHustZRVPSs8vU32SrxW11eqAhsSjtCvw0GgiO+u9JvJNw
SwaO6Zt3FNa4/LMR/s2rz55ukH6Vy0JLnWrVIsyJXVyz0qg4mXm82i9kmjdQgG37bAvS8ocEEBjs
0xB3XIhQ70hG9YPbGULDFwzuKfgscuSlvBOI9HrtCX3slzmTt1RDcOhjK0FU9ioreHj3Z91x+sbx
fRAk4LML9h5nD/aNkQArfHmnwcB1KICdJ9bteyxVvUdaNhJN9YbRYwABPqM5t9WbZCoY90V3s/rQ
/JzujD7venFrWukO6BtiOsU4TwO71gFDxTCh1KuF24lFN9g0Wm00yqwCmvzDAzYnrftf5vBH5QHx
BnIgjQ+lxUkVi0niH4KdPPiN5zc8nLMYl9Anzz7w2x0ByG618XdNIbNtS19OWE8oUujPz5KnyXMJ
6vuZGzrgG9yMJ33GII1rYK7VB3AFv/7HgVcrDu4zBJxm3mMy/RJiQ3hCyz9SNvJ328QmjwD4OmwI
ji901g0o70dxl+ZvddEiK/4E1w5NvUJdsoasj537SSN9JHo/m1Jsj6Zeyf4XDr9wSxmtWPQtRJ1f
fHTkLwDGPng65uoIscBzRcStQOYDf6+aH61UI3w90ekvkNe1i1CiK124mCCx782/n9EK/3K3MV8X
7WOpw2W3AYciCfjdu4warCi2jcDwlxTDD/HO5QojZ6bsCOv0gNM1f9A6e5LfIX/5hHPKLNMWMBrM
WEgu9fiY9iegTOs+1GK8avoKM0vj76Nk88J7mLq4BV/Ct2W3jNdI0to8tbBWGo6cDfpZ0+Fr8W2h
vAGAJPRARLqnJ3pZIBa1wJpy8NtZxbJnRvz6YvplUevdHHnUEARyIqPgSGo6vnys/pYGWCgNMGHG
Vpsuj76nQQfBedwVaWFQnnPONZn9VpEsO+iRN7bsAAF98EPp/Je+nagQhpBi75FPhQI8uTJkllup
nbLYOMcaKUpBUdkWFQTl4aLvGOBFNmUP4Ck00wsrF/fANCdPS+hHtYUKeG9EhA5HvV6M4YNOC1YP
63v24ktFMDuzvKqYTavZkbbYbAKX09oCuPyTRjYs08bvxxRezjoV42Wy1wR54tP/JxpNNX/aBu8V
8WpZ5YzOoewKbe/Iie7R2OwEuTtjy/sCC79xRuNrkew+QNtzqPC7AXf3m6I4md7IljR6PWRRLT3G
ITfVGihicMV4xcHeWUVGw527hdrVsKfdPHe/fd4rY9oAUaOEl/WCqZA1w/Es7NbQGcXKt8j0UzsU
tShIsbOaNQtewDpgLKfaMuo62VmRthiNckJWmap1YP1OJwCNhze4ApAl0aptWlWNuU0QdW9wRZVw
WVGo01fkFmIiYoZNtY0dj4XmHBEh3dMvqChh33hOR+hYDg8g+/7Uv89h0oeN2M0E1lgHlE6sWAGT
Q9qkPlQvr2coxQGkgAS7zOCxaKuTUfdfKD9GKAWuNLotY6kdrxsYoJrai0bEZbxnUK7Kx5WHjtZf
9DQ7FRE9WBNGBh9oCPZA8MUwUopYpnZP/eIFyUJekC+1/75sUBpjdosCUA7yxnevqv7LHY2UJdbv
kBICX+LNqn6Dl4XkMIIQrDMfFsb8c7PHIzzYNRziunYneMLru6IxU7xBwOCaNSQEdToVY0Jyg05O
syTV8cU/HF/RmkRU9E/9zxSAbHbzS3Vpd7Xith8XbdSNlcs3UNZPiwIj6yMepw+hPAT9YQFHvmhg
SN4PBjRfkYXCe83dtANTKQER/XgUSb3JC0loZNF7GLHv9qi4XzsaD5jXxllryqnuhriOOie4tweF
M2gCyKE2YAhzO+7Hd7obcwpuCRNYePkF33/FFwcPzHLPlEp8UaQWXS5ZjW95fKM0RlTVSB7XHkrJ
1uqAR7KUBkLo6vR0rF9ZmIcppwrUMlxXQciqCHbZILAakGbCOxJw1aenJuHpzU4VXFCMZg8RAiYv
+cHCIJbnhSPLHgzGx+aLkPgr5FJbk8fyna4kv3PKrvWpI51V3fQvbkZpiZaUA7INC1fIWvwvJ1nU
MF92iszVln54TYdGcpAsyXwJzCkNRLA4LR7us4QzuOAuPIYDKouThhEONsht1hzA3SxsBAIjlJYi
1S64BP5BQvzG6WEKPMcQnni4c5Y3/p2T5i4TO0pH/OqJYQ2vp+ak0B1BoRbLmtQmtPhVifnmj0rm
lNAc+oueQ/ZBFm8901e6NleT3MWj/bGYndcTC09n4i+kzbQG5ltTWussSHZR6HzzUTFYhlnGI61y
HpjwZOLJvJroNSH+x+0k9ON42vCwzl6TXiSFPhXUyJc5DL4Gyac8GJbsnObkn5To9H9Bv1SzQjH0
71J+CuqkBT/i198CQsfgxOnaqkX/msQRPXk/G/0gjyrDV+JAmjLjowpCIqSBZgXsw15e+c4eul8k
U7Cp1e5nkfcU2ZghflijxkchJe8inmn9CNeKPV1tCLjMXS9XMk5DB4Sp14J4k5D1Nja6DiYpnfiC
ZXSqTI8kQGAlKNXIVAwCQ7XsbUxr5ptfjbobMVL2PfF84/2InS/7I9Py/JQ/uGWFqS72rmxFAJWZ
+sBf71pdIoe4nDUAPVMzAGvKF2aKxV4GWnZBaVivkD/aHED0SB13a9wjrzMjqDae1cEYrRfXuKxZ
6mSSeV8uhWiORa3ZOxchro8YzwhBfpOlLDoRRmmc79t3qbdfVJQ+/LqF5T+0c/oAv4rGxeY6eS7p
Oh2BtejGl5Wommpcuk9HpE8pCM45zqSkMd/SurK9vAyB5OToao6JkhaM+YA8xKgIAsKhdgzGRwF6
fTvWJzVKqGQGcjnw89oaB5u9X75uJVwEOm1QJie81GbhvbGvX53kW6hDjuEGtvQP4KuZDafqrAkq
Immh6T+fKr7j6lsSfhqFfSc3mbxCZ1EIn+tNtb1cyumKuA2cOsD/AJ8dFPNHelcmycZjLuce2J6s
DwOslf3nd/rRrlQ9BhjaRL9QSW8iEkRcb6YsjqClhlTfyyvdoxBOCGLz+JxKeyACE9mpJlXVOUyV
U9crf3QpQkIqznnWaQLzNY3Rk7XAAPG0oVQ8di2XGAYe/04+lB01Ke/5qrR4TRYZjJUrqP5m0Vrm
Q0AD0LIfPauBfjhGO1KcNsaA+G4A8R/BuiLdtiTTaDQPbQzSfZgwpEa0nDceSC/CUzT0GJjCqdxY
KssNtnuLfxISqpEMYUCgZSIedcO2XE7bxvwpyAh6r7UwF9oV31qYcCADnqkmvtFkMkBg7PWzB12k
mBUa4Yn9fBPD1wvCTguwcZ4G8Ocp1lHpM/l58Y9LSz6FntDY9OehgBc+7tGsfjw8N0BtMU8+J9HM
0/o4gH0/5luyVDQKTFixM7IMHjUcIDMFL4BgA/IPpgPFMJ8uRACg6mRwgKanEaYctVb8wnnItX0x
TatbBmguRUXavR7PkPaLTd4iLcMYwT5PC3+nBGRhFKPrjL2xSiG/Y+xWI+1rSzimA4U4d/TmvYYb
IqyszodT1hnmc+VyLUOVI76tEHs6Xm95r9vL6SnRCfPqmynmHNnsJQT8lPQNQeDYU+R9xRoZ2m1I
qKupCq1OZPje6MhPKEQs2QKjV37oyoPTBuI/jbJ6iJwh9vfGHkCk7Nud1QVZYkBEbcfp18wfXmLT
H+j+GSSZ6/+V22ZP+/DnLlcuhr8NqQryZt5iTVRNyPq7gAbtTFwGq5OfWLc0wVw6Xbgo0QaH6XRy
iNBWvERjOHMIxvQxBlyB06JLlazb8BMpcs6cqSFJvLcj7Yd9p4EMMcS9SVAdEIkYNXxezEXm0Fp8
e4jzfUGwIO/T3IoDcsGuKowHY90LbVVqXsqCiwH+DmeoXVS1C1Qe2KyssWU/iBT+PA4gTD/Mufch
4Uiu+znyeq3TQW2OrUq2r8Q0xPE/jPVNxoie5Wagm7Kjh9BI1RtCR41uplw7E1FaCvZM3noMTCdV
Yulbl4sK7ocnKA0+ANZs2hdEjmLnHS8LUqd67a48NNk8mOV41oKqzP2qPdEgd5795hdEYdPh0v2n
C/fiIerVaug4hDIM+KRXBDXdphhh6yj4QOpSVkXeYL5hyjX4xIMQeJC3yASJUs2rAbSY17NBEjWA
vZS+XNbVGcE4H2NNTD23Qi/IZjaJpnqqnhg1xWhoXN1zm5zwfxfvD0w1GciRWt7/4vdUAbM7u28L
Xqk57ede9QDnBj7gIJzv7kag456Mo2+DVCqkcoH05EGf3cK7wNFJlZaFF+XnW5tqDwntOiKlKBhe
k3XBaKPXMsUJUcZgyybCJn+v3sqxl5t5pmDjcczcZO5JEPphmOjw+SOiyK8VpjfPMo+drjfL3W8F
1ZI/xs873ImFlQnT2zM+as/vlx/LQksHZyk07R8wwc/PozpeYL/nNdNJfp0V0thvdP7oDX50cHmw
0FsBi7+EjlzSrrIrbl7VryBKF8UuuUPtTfnhFf/zPi4Uc1CUHPECrqIxpavzfOzNumnf4Ux7uFl+
414Q0KHuxXFHgEOw9etWWPcFhoSPQgpo1EV0OcF++Ho+o4WqtwDPKK51XpazG0j9z3km6ebhLSJZ
/HJYFKk+Qm7Ik1OCX866hUPUkQZRLoPjNRfd9+W2pDOYfAwbJRt2lgb44WQMVsRoIw4RkByfr0b0
kSrRLxto1E3Sot21nkiFhZZw5ugC5csrB5N5dj17Q/KY2jOSubsmtOjnkK5zcSSHRIFdCfJksGq+
muvLiYNZFlzsIMod64Yl/zzE9wH6OSu36zpj/LzVApx3/TkqQt3reAMy40ksfMUdh/0xcUVUhBLF
yPCIV+H54UTMF+k56TSc8TKEZqhwmKM1lf7DR/vzBszbgnfCsYyVF/WJGs+QE5nU5NeduY4SrB7z
F/swcdmzl7F0d4/MV4OOi9vOPUFLKACfCXkWptWaEukTCPOEVPYzLC5PirwWKTPm+UuM5dH0SUo8
fwO7vpFkOy9qsIS4ahrcYjp5jwk5on92Kv4bs3WdxjFuoFiINzOwNcz1DGL4owOfH4Gqnzv2Q4pn
OWuNOlRsCnYGMc69mqnlWciIwLF5dCY70yXBu4nwEgbU87e9LW/AfubPl5g/ajgJJz2k8E6X6w2v
xCNSIyOWdXOplwL/OVYZadEMCXQFz5+cmdtu8ifHc/JunSxfDJM2T+SPtXSDUArgRSJkwt5Al0P1
+m7UI5yzwaslyvtO6mxW02EUUApOs6aJ+YpM8JRmy+9r96I3B2vB+5tu86sZw1+WHKnY49ttz4Hz
dIQds+JhUlVdmq1Da8v8VYyrlpmFzSwe0nH3dEZAVjPp6yQ9/dACVackcl9gOpqeDKuwjPqTN/gQ
byFytV3cqQ49UTx3Jv+Jx/OPyajTT3fK2Mv+Nx9u3qPbTtDwbMl/y5BzILnk6oKvFgtU8v4O2SGe
R4k/Sv/+mJlpOXYAAAZX+6ibuUtBxbEBfxQxaOfGYq6HzGsivlbJY9ud6Vzyr2mnledqRtjU/6Sz
mq4JB4w/QPW241YAK6fj1PmTjPTN/dyixPQ2JBIAgYd5uXgbKgCdRJM4QdHGsAEOl/88Oo0ulsqM
OEikAM3rtsIICxKdy/XRcX1gd9tXZpnET5zNr/ShzjLC6huwssiSuwVlUHTm1J2l3a4ToUJS5zz5
/+3LuPExltvj1EFdTLcheVy4gPAq6pXWuiW4Gfa5ihPPxqsSpTFog/PxsCvoLDdZJPBrO8qw9T+6
K8zNsk8EWnd+bjWYoB26MCdUeDmmP82q0UjhtyN2ofm/nTmE6Df3vPNM5L7wZCV/lg9uCnBv+Ss+
zyg2sXcvO2tEPwPNbo9hHieZzr3NqbdOXW2YwNiUbNKnHUrIFgtrEFYex62Z4LcgmmRYk/SPBtDU
nStTJXRbDAqMToWjSGf6bbRkEbBApU7f96vmmmqZxRRMqt9q/KuYAmJ0cjuUAevVQR5+CH3wtk/e
leZocuRweEKFsGBQ8SsciK5ZfEsM9phJf55eAQzoC/Gm2P2eNQk4yZg6hQg7akK49srNki1+r6jt
qbFg/w3X3XuLCTJHtyo8InkPFMpEL49pYd0km62s4bKgriiNJhIY+iwmq1FtiVVDj1YizDXL6uFi
/gLHf8DSpeHU6WRRcxHkxyU1mGky9PaUXVR0RD7ilQV7oafe/zDhXDrE/+5DnQB3zGmcC9ydoDcU
LH2xApQbRftbkAmFCDihyXOvzlLpPOERtFzy6CdxK8z7JYO2V4oTJwW0+K1Iw0+LWjpM/jYPWcli
bSCdV09cpAek4YDUfBceS49babp93KDf772GBI9JzpWWdj1bBhXcic20VhERJq+uRwzsaUoLd2Jh
Y09dPSfnC0r9yt5wv2SkXQdk2dKf7bepIARZqHsuRe96Q6EBvl0PymY4liuQqJ4+JligVHzlYhCK
vCyyxWOVr04BRl7xpg/04ZXvOGNUvHYZP79TqlVFaF09MzeO2Psdl1/r2fGscMoL5z47xf1JCAdk
F8Y5CtsFQzkiYFO58EZ8kZdUGvLSlwHhj049g66UFAF+z5wGSxM1XCFuyjfUuFgA98s/I2XKCVZs
F/tbWu283bPWjIqmuql9K3W4y42FRoYhOJGa5aIBgfFEOjYvbIDJO7wZbfDdU8FJjjO1Cmwgu4VT
RlRb5yMQeDoydLtxgX7LgIw3oTBLgBpo/By68H5N1d0GxqkcQXM8gATSqvC0bN+O7P4zb/Qu3/N0
sPT3lJcvKczVODQWtCHg5lREpF35/rxy4YlVCZC6R/iPyhdIgOZam1qobLmPums5CTkvWaCcXu22
aunTK5ePWMejbnl0P2njGBYPj22+xl8ROfVKqFr1Zn3xWFpXP6iO6kBHRzQODvhkWe/pIK1Wq1hE
OW1e8ISrnxHZi3/wa63XiKDFUAd/jzKn2FM+mTIPKQFEilLsjLJqpB4YKy09/DBCWgJ3bMPllPdC
KsEpN98U+RRs1ABOsRJPRSQmkjwboTUzuj+WyAoJi6ial67g6dfIsU9g6tzyOi++O+qeaNWGrjbI
5dTTpuRJS/EmWdnBKPwKagEGBuSKjoClcPPjgN197448G3RX4IjOvk+Q1oVsw3lvPgzfGr2iu8gi
Nai7UKloPguO0sHkUFETyl/xYTugaV6L+DAcT11JX9bRjZ7Z8Zt0ERjn4qOZqd/mMvjgPjUVrD7o
CAyYju06cgeZhM3jiePN4tcip8A1x2BwdWTyLcqViIVIjhvbBOYR8TY20F2snOhkJMn4iKD5DvxG
XeC/8eNvPDuebDAANxLJUEGj5M3sy8Sd28opZ3MS1/X/tdeYFrB+f8gfDxXvC58YUpGE5jj1sHJ8
A58tvOC3W/rwDAzJshDdrHVxRGcHsexHq5cbnXOrt2ujrVw0iEA2l7m2wS/os04p3COhyNdbhdGR
FY/oMfHReIyNWMv6rgA0+nsrJHhSevqYI+SeBIhAz4l85rlu4/KzUEKLpaxQukT2V7j+XObh5meP
Gx6VUJfZVnVwcBGHCnpbpQcdIgqQlK0TCnOstATqsJaB78LgcmTUMnlzYFn5ZbIY3TvofK96sOtM
udSas76wOUaAYpMvBFuUtYAbpa0++5F7dGIS8EHn4CJmqrkVkfJyEv4ACh5/54n+jdPfex/J8SRU
51hmA47b5KmrRXloExR4GMrY8V/ojMHeXRMXn3MiOBb00Nngu7/+nRPL7dl5Byrw1jU7vNvLZGuh
xEmaCC1+radzkeQmy9MAumHpgtIVc/T+iBzQcXTkENscV+cBBuLiIGaSSVCKM+S0YDND0GUgGY3X
NE8c6l4tmUw68tDcAmRnPdbAtWKIfZVLWWAdgLd6qhBm9L70W/VwznaUom90Dhp6E74hn3cGP05D
RvR1mQb3rUq9W2exiHrsGaH4QcrqcnzFQSR8BFa4Dq06cypAGqPaJnVb9T+gAw+ZyFrbx8hg6qqW
46ame1ApH3JtrXfmNo/Ky+akGrRJ6dl0vjlu8lcZZrqz/f815GzyEhWiPVm5HVMYy5PxgcTOfvxS
80GlZ2sox9kyoOPaR/x3IDK0/QE06UwfNFEfV643tO7X5oGeGr8JgxLyRdEu3QtfXfVfM7JEX+6x
lK5IFjfBFWl2HP1FAhZxjsCWBNHhRRIo69klBo4dvtM3I+k8DolpVnkwOI5Wxs72PN6gwt+NMt6h
a1PfUDrWD1CtBojAPvIeKwWvVfVz1xqxFaFm56o6+2/npF5lQXcliQIb/HhEcHBvn53G7FSfhz1+
gx6LUmlr27z4vY3duDg48dM46O6xNNAvxDjVX6AanD2/PAmAWwGEXvgZE9F1EW1nAGpJJgHIMdA4
uzPs04IsP7CiXktjjKW3M8ogJY8bVoxV3PCpGT5QmSm4kO2Xy7CZyyhGrF3EPLJl3W20xPEifA5k
J8U9ICJZwYOG88hIlZi7861RRgK62QZSWzjO4+scpNiQuHMGK9DvcBNYVZEhtX+goDUz8AYVhfaY
3OqRyLKBssPn/ec8SUDap/Zv+J3R0YZp5HT6cfUlB6Gdr3NlQB4cUMiFvNTNnRcJRkHe32DXaiBU
zZLv4g1nEVdDWpiLCvpf3a0UCn/R9dtVQzFAC6WxsN/7emDgcX2uycl6E7TWiClpJ07xj7Bdg4qj
vDTtDP6tkfPdyVG+XpTIExjdFTyNX8w9u8Qr2uosMKqhrvC/GNwSK7tRcbWTlFn8ugeum/K5/Gz9
5BxiGDPCHpGWk59NxDF5SFfsNf04psOqdLVkkjyEB7zGqKvSbNQTFwPgZ16XE15O8gtebtN9k+11
aHfL2+TPBcZYLcJddddczRm/ZrPB5a/CWt/1JLrNm2b6jat/scwcyorffzuLstBDIxfM0B5xGhnZ
ZHgboA78uD3jmRh3cIZAX/pwSPSD4qTcm7Rk2N83sq1ziPlMFH62LLVJHZ7DwwoWNRjkrMJdrgR8
X4DHgg/8Uhiayb7C8RjvnvmUqlwh/u7dYuJYLBjY8j89lZ4sZrqc9+wc95BBQSAn2gSUnwIevtiA
8ZO78gzKkmimyhLKgDNd3iCtnOyZDTM/9aJiP8rx0mDXyYm9KLhP/AyMnFZNO7rZiUvgk53Qd5dN
xRUWioE9E0WDCaV+rJxrVeLsMWHhJaUTkbcQxDKcoWJspINQw1tpcv0IvBDR5NMow7wA91s+IM5Z
sMt+2FGgRH3m3xvnZZu8HuBNUq1P1E0osxr/+DyKlPBZ/qDF1bdexE0sWl1xWJlC35R3hqarCV86
qhz+ZOhk6MPd2+fv5nMAN+a6o5daKOC/Y/+gmxwMAdTCwkizE5iBN8XilUDj+kA3D2TrcCJb1kxK
10RfjLa/z4RO/5FAnbccQ6SLpZfmWzlrDufEnhR0yznFPpkztXi1Yu1Jxr5ajRinqs+2whfyoVXM
rASxFOXPIiBopGRIVswg3aBK1D9DLYtLiq0anP7dEmpgzxr2YBx3pcQb49k/ymHOCbrmqWpVFsDy
jM8bbbWSz8fx57yXRF+LjHp9c5zbsPoLBM+KpV1MljcLibxHqCXgXodNYbGVPzUpKqgbxlG+Fwsw
2PovWEUOnEXjiiJBJWO8QaiPH3UYwVWBbndAgYpTl1SFGqP47NQHe8iaRZp+HcAd1ClrrZAoidlm
Z0lcWusvnS5pzOh8Skx7dJSFeSuRR5+kscBH/WvdGDt/ziiYwZ+bpa4xMN6IxJY6VnFGJjRtNatg
9XkqYtVxK9x2aRN+bIZWQEmymORrywNpB6QD+KWVQKUs9JUmzyYj7ms5+VL+rL8JKjtI44XLQbMU
tg5k+pLBUPez4e4AiElk8FkoOmHp7e2Fh6ZvjE+xbl7gkOqnLQjRXjy0Zkp6aDEfatFqiS9/PCKq
f6a9TvFS/A76ukW7UM/XAJ4ShUfSfXNuDJqX5a1fIX/J4zu2NriEpeboanqqNqeoJpUPjjiBpxjK
QGDehqULRkkKas2qYWMPs0VDh5UvKx4UdOSlHNqN6YKTgyw/iFt47+M2S9SMS6Va/G0d53oorkG6
xBfmE4TplVRdLeIvo8r67YNH7w/zkUFK4J4Q2A1YlJCRPYKwUWog5IsYDfqXfDMj72z+yhEtvw6+
ZbeGzHJml4Ia+eUDel3KqBY8p+VnKK+pVnwLPzIhBibV29rKqy8gRWuvA4LWs8dB2jHVp9qEutV5
cjQlyRZla7QiGwJagO/WMYEGXPz9hpVycAHvJnvGtAeVoZokrIOgpanwjlDWxzqEjPUQf9xgYr/W
nxzewWwtYAJ++4czq4T2y9XI08kRu/u7fTHtgqA/INk2qjsjevVVUAp8L+zbgbD2X1X1qSdj61h6
PjHuCSnGbiq2UsaJaLPv5x/WfquE44Rg7PB7jEP3BZJ+5iWV9L4VaEAWUMZ3rV8EVN35YDDScb4p
jt14/rR4WgDtflhbw5Nuf9O6RtgtEFoAEHdgWLBEI7d4hZJCR9FtlSUtcvj36OndKiPW7eQJ46yl
wfD8/04aRxGL2OvMBDmhX2rlRLnv4noLIdYj7WdCFpD96ShkgdeBD4RVT45GTs3c1vzDnktmjj5I
RvMM6oKnhw6zlVKV9kNvuHUT47cO+HdzuWD5EkcrV2r/cU+4axW+gVyeGaMIJ10VqSymCpjrBULA
+fhvyozPHJ5MlfWKBN9ovI1nYdp3Ups3G1531YbnRLRnCJBfta6X/vLVrgoYangMTi3pbafbilTE
VvJ4CTx/dkIYn7cXL67NHgBSEhQ2wTcGx8sfA3Wv73zPnoWMEgAk9EtNfLFsmRB5sjTYU43jqkMU
smMCwAP6Fs8yvEkPnz66ddcX4mzsdKKFaTDcq5al4EidPz6bAOi/qR6gkOsWQDmMxB2DEEOhsry7
//kDCNKo656ySRuAh1GAX7+TGCcSQpCX5UX6CwaCULn0tEUk5wzJxxP9N5HsUsLYEHohBAWt2Nva
nSOAhWXklFavZNOSJvGwLvXXfIeQiGCwCyIy+YM7Jiusa0hADNFnzyu5zAbDCG8NsfDzaRHOqjQd
AorCn4v3gAuj5qr1+HZKcU5op21mXrCCvmS1AtxiLEJfZ7YT7SynYEfH765mmabHMuVz5ODrMNya
QPvDvOLN8C1vQIHY8YNUzxdSZVtJXpJY7Ybb8udEZqBAAEuH/sKVWTAv/yinqAVsKbkLtPC8bETZ
be1rYDgApuomHm0jAh2QQp01Qpe6cn90IqL68q6od4uIZa0lbqCwAUdxdsofdhQqqeAtsimeNBPg
L3J6cxRiWtQaiP7ZUKjDmJUAhKL/1byszK8TFFl8INDPkerxDNNY06X+Pb6BIQ2Lw6ghaqiJLsUX
mQ+V7dKpDsR6OHqs7Niwpbe/md1aPR29OXkaW032E4YXG5d6p8chHQtBS7nh5tlVkj/Pyf+aFUoU
HrHm6WLlN/kgQJjKqzBnagrlwSxJVzGBrNRY6v4CjAn9HtdzRtZxDwZnu7XCzmacsbIlxt45YeIz
6gadB3pMu2wjk0vLQFeHcWm8GFXkjgPcFOHB4ERFl2fSGYtYOqIenesRvMVTU+eD/N4FUTO1lHNf
/4mLkvrIHjuVLf1eotF+aL8dfpLc2IddvRvM4VMdR3Fi9Y5JI813KjO8z6rB6/0bMhUsSah/0wYL
wTcZMB03+ewDlkjdDmVnrMfw5Wt8j8hvnSfNydu3aTUF3nKTrm//xlMuZpT6o59G3xLyyaWeSXRP
41E+pNUMGIyh89Ycq32gG698mXuIM9w6yG/lF79OkgNwxsWeQWE43rI/UpwD/Ic4KenvVJQ8mvPY
dEpvL9cY5WTvoqK0jcTQc8VExyIwMcbRnatRs/cYibzrCaOgaryfXQpXxtKV2vnKM0Y6pHdjHkPc
W1YjrAijE/jgLoJ+/kGMGcWRfAzzRDgwOt5ESIcvMnlq1gwsnVXxWDXs9UYfBzzbbkdo9w9yx+Tr
Mx4xFX7+WFvsOzCZaMogikzYJjDgaasVVG/1oR3VIcYDkUQVdoefSmUNNgRVgKZnYak/kMJM6jCQ
VqbJaR10W+38sP3vhsszd3B+lvage3cu3jM1xa+EXfzoPWEeAqSzjXuy5Mmxx/Xub1U28H4/JvGq
IroMDSIrfhFRldKjdBCYdedTJAvJKzjSqyQtWMivPYSI5JIzLGOhfPNsmwuGk7zz0G4oAq3SBnyC
BoBfob6RB+XurhbS/7g3cjhGt6HZc3zDsvPHytFuOmZ7s3bF7oFQ/JzmHriJ/twmVTLcnZ8DwF2+
VefYxKZKT8uhwV7+kiLl8bkJDy3OTaj5eNmksLaTLZOzZKc4Zf+yVNchOLtkTl3tjUHC/Abmrs+W
PO7vB8AQhrbZwvVhXBST1H9N2dX77M5HyhRDZMIMRvIgFFcGpiJEuhP/t/g8n5XlfLLJ+mJRzeLA
oXmEAgU7PUEBSGPZq2AzVnLfxwnsWA3EPtsmAf0BclaigWOALKekWxT94bZyNTRxAxlXFjySyPfs
5MZjBMQQsjDoA67KhPvsYt4FD6HcaKyrPYy9iccPZpxeY0XWfq2FCSGCFKd3cFPEldLXah1Aczrg
OAxSXfHPvRBtJbOuxS+jJZ37bVkq452kvR+GiQeK6vsFZ0oVYz+fhypOqRvW2vFzifzF+t/W5/14
qQj41MuhvYm3x1aTNvAOvev9uT+X5tRlFQVwgwcwN1Szh61c9WDj0WRvmgxcwOviYlJoN5CAKfdJ
TfyVQhOZ9Q68Vf4xr/eM4EShjrSls48btEgJHaD4RHg6MiTGdalyzV1gXCD2jJZFcU9QRnJufbJT
DmHqDF5UI2NHklMIFNwtgVhr4oWAcK96oIArKkQM/PrKb+GRB56yeelIn4UeAhEDVA4P1E/R3vSs
e6NjvMMNrv48zZjvHal4d5rHFQ0QSSevAHEV/lInPx1enzRz6F/TsLup8uBfeS2XMxeYv/ZSkOMq
mZnZkZKets95+6Spxod9vg3kdmcy7kwsSTrGMd/1mlXdJ32gRbFnLWJzl69wzKjuA+zjtQdbQPrL
w7LfXi4w2JMsHq7o85Ccgu+iAAuapIHOcLbzUoH9WrNSvPcPctof1GxK+dvqtEy9sfcXJigzolIR
PjTNlNYcz2fu3Vf4ar8Jt+d8W8OwgqwPcFF6fA6eplykZD1+NWcwEsVgbu0RqADBSyvHFbcUtMZ/
BkG0DDJdbI583k7O/ayVBCJK3rimsIvM2xTqZkmRBhzKn0h0kjTBfrhXaCBqKa3csJZsPee1UubP
7XuCvXhlCj4FWphdTZtGs/gr+w1tHHpWj+xMnls2CCvp6ilUmdwcprzwyKpdfTqt+BZ+Qj7cImYK
kx+IBp0rQKA93GcLOGaHP88Y9bvDHG6iAGp5RIeewWlJrZAAhF+yR6gkRjvF9aogT496lRocRTzv
sxsHY5Wws7A37nllJ6qfJ/24o3P+Mg8IMWa8bCCrSvZ3NCfaHcbDKqA9Y/ZZBEBXLi4qiHRu6rdO
so0TtshtlMouAm5QSCv3qznOI7xhXQne4Ho/hXnTavBN1FORiaXxRf3GHKp9bNie8B7utvV6e9pJ
B+Dp9JYFDRgfbKt36xsjLTaaY9r+Rv2fGWrAvfDnQATOIFJANeB6W9oGqdEgBlc8NyG73iWSj+/s
Qgo+1jCkguHheqZ4CbSkUIp1sRq50E7ANF6uJmmSm5Ngc81XjqWryu7BObrSN5WMzBB/EJORbq2L
z5y1OyRAlkAg31nxJw4aKYbVDwWYVvXmJyJ5I6cypFDJ5Da/GjYO0vojhdL2GkO2f6BhdEYzKJs9
FLm5JZs211Oq+hePfEH7y/MRv7Wj7gSZ0DBpu0LXRiglFvw3bYCKT9MdwALhjwwDRvnfdQMKOCP3
426Ss8iNXeFNJDh7WFIAgaTK11GVLavqzz9SedDJY/xP/7gHW2T4qgwwh8yY6KAe0dGnrBRuAQQX
lGsxTHhABR/PfFS5sUW96z+6ZzJ7VX5PxLIK0X37bMrl77jSWv0VRvBP59bprr9Y+xQF1vN60R3p
Zk7gkM2X+TLH8KKDKGPPaBnThHqene27wyfjRtzqzWCIlTOHUJxIJ7MhaofO8Is2HTvfLQfMzr1d
F1PTQmoG7ZjMP9qf54q7snoi+51Rmciy139ICSKQJabl3MVpr//OegSG7FdaF1mSWzBb0ARUhX2S
K8VtUkm18OOPB2Tvk0IFFXLz+IknTOj0m+dlbFcnJVQNymSQSXYpLBl9GvzBnKHJvZNMTfJyxh+F
YUbCEU89clbRIxX99FpkblKjOcaEtDvJ2sVaYEdDdVMGWwpdhhh+6l8o3vzLgwLALgqDC8sK3i5N
NfN2NWlxbfhJgEtv6OjWLTwdyVVbtdSIMpNFSY3iR0mS0mAMjwAAKUdHzhVhP8iWJ6yHDo2nB6n4
62fhM5LSzjkL3aqUkrCsc0HeqQiWzoJ0B2m2VI2rHlxM1e+1Z3jfS1AaMYxpLwfkUYbr5qDr2Qxt
w5N5vTDW0iKMypRrf7gF8kaL9wtOsg7r1DmEMs3xpX1LVFjVrSu3vtoKaWMGZnKW/rc/yX4vwkao
jxkWkuy+Cjk5ywNTz+Dkj1VYcb0w1rw8+7/KkmVyMPxZnqcm6wHvAfSfVP0TY3Z3HBcANt5sjqrh
u4++6EM53EvvL0mkaxC0spGwWT4hXd/DcswWa0AxRYPwV9/3vsJcawmKOOT4r6MWKE/n94HKMGLp
03vQo53u0mLmZ4ijKk4CsS2/YaDGHqg128AYrWHSWjfRQ07DR8/vc2P4NW3/Sm69FSN+8lfHJDsK
f5OPr0FEByszuOIVpXyonzeb6wSMhBLYepuv71fEFppwY9ZhXMQHZqlUb05pCNMS2zpUzLxd7RcH
gCHrVK+Qcg6DendIHdgZ4psGcBpOcgOaZA3kzUzXBNBGZuIQxhhlzlQvReSmeAc44XZpeqJ4elve
oC73PgznXmACbC4IB+VydA241Fg63Xir3gGvKisJzeyPqZWnH0vBX0ZbUGhoLDZFZM0kcIf+SLtc
+eSuAegJ3MKPvMNpLhTfNrFI2F420ddCEr/40OoVZjAC4qTDLTZJ3FzLiEDl3sO+kRpmsi5JJvhU
By0WkmCKDFFs/CFPMrDwm46c2/2AZT2BL1P3xlRZvmoYNYrMAAUcxoW2nBrc7A+Bmukyg6GYN98+
Sz8uzwxY0tomcxBDaZrWvR9hCMmRz4AlfpuvaIz5xUUpe2F6aVnNsWM1WYWVJdrOF1EWAhIzWILm
u1aAyjh1uVTCTXYc224avvTz2wu4v0AaI/U+E+3WSvq+iIxHAERq7hrBDJL0x+UH02B/nCoQV1wB
Feue6M4992Eo2p6GxbhvENDhxr0Gu/PWuCeSLXoD6eKKxdm651JN4BGY+UZHqeSCfVkYguVjfeiM
U9JmKPfORdmuBObTpI0lmn4msyT5YjPuKscBuJNYs63Tax2MI7SMsn3v5Fvs7P2J/wQRuWRCjjUW
IuhqF3IihZuketZQZ/3zZ4e9y9DObcc+4bPCgXP5lFxNqft6dNQ65EUMDVuLqK4HYAWve6MK5nwx
xLApma7p6XsJatNj9ef5U0exMTF5GsA1QyD3iJ+Ugyw/Z6rk20B+hJBd84x8ci9qzRvweTsu9na7
pFp+nZ+xIwtCW7GNW8LuHI+vRS+EwioTs0Ans7nDSc9PmWhhn4WYvT4rx0+NiugAkzR2O/TZQuWI
IQKM/ATRDTpWwQL+Xv0W8dRKj4ca1g1IefUBBfn9av0W8iDTbHxIeLOTg7tORv20wbouU1WLWmh1
oBr+RxA+JNm8mEEOWJdC1iLrN01DrpbaVqups9e/Ub16lLRarkm/dWg0B+LICgrHIfPEJ4prSmf2
PHtr1t5+btVIxhjdnRSoqVdEavZorRtM5BvGyvHBIMC/8C9IAed7VXoND4eFA9aCZ6c2iV3pz7Zs
6db/BC1igsKwIMDcUqQ7k4cZ5t8Xuq24oVWZhdKKoj6WwquiXsogC1u9n9d6ADJaU0XqplnWzav9
vLXBX5J46E7keLeITh3GeAYuejoVX/7s7Tj2eC+EKBfJFX1EGQkAcjWLQHmf5TEs8Ix/BmoWRibm
GjA7nG+7b5ZWxOYKwTEuDyo2fhCOhih3RYAZS6Otl2VeZ0yIaUrUlr8i260JFUN9YVA2Et9On/Vz
AT2AAZSQZ+glCKJobYIOPA0J0kci5vUSv68BIDhr88nKQS/zmZIOU2rKFtRJKmzQph4my6UdktkB
vR45xbDLGS9Uk6SFUzcS6jtMyygaTv9jY3jKCRJOJn5tdWNJhe5a+1kPmMJ8lBqw9/CCJH41p5tR
gDwdA//8wgRnLHGgpfcv3yykRYmRNG9fY2K+N0ncxxKFaLCdzOWzJDVgoU91O0+tlp1s3hjYCod5
RBLg0uSV70F2+aztn9YskTgWpbW2cMTWHQ7cOkEWFu2IbkO2NEPAQNGATT92JNAIhfz0n9P0gIPb
FSdhDTHUA66P5bGwyRvoAw5fwGlGNgpKP9pYPFLHv7kTAHMlPVRZqiUkC9gs2XlzMvGa7l6oiXIE
QywYKkSCDNitRqLKdQLWENyeXqolEarj2LFj9k4JccnG1xfveXJdj4C7Wl2sifJ6aK+sYDz3a8GO
HwHFu0NyRyBKuQAoJp10VVAGyLKj5ucLQLyj0bafV8fz6zGuj6ctQThFhhYt6zrNzq0kGTnwZ/+1
d1t84kuxKVRP5X53Pc2QlVmaJ24Huju5EG9qROyKibUbhu4wTAx6SY9jRQCFDPLuRZrcw/yBOArj
uJkXXZdvv3hUzD1qhtiQbUOcsZN6hGktTl7bGIg7S9rv0JF6XitOWcHw7SC5YmjinOBe2in7IOP1
q9gOma27OVU+H6G1/ah8CMoyhCRbEBrEK5qhNNV2GplKLQmkSIASNRc9ZU6f+i/oy6Cf96T3ixi2
3ssjYTEbbwOsK/viOiMHyhRRAVr7Svx6D7wh8uUcOWvnYktEOjmMvzQWQVwiBvSnOxrY8eSpgvSN
gPhxClQ6xLXGuQCuTAmVlWT1ka1Ju8M4tEa52DOUwyKmgGinFNF1aYsSppssOJVmo4vfs5JNZOyd
H6mmohDMyxd736cuhtHmd5N/SjVD5t7QOPrLRmb5szfc7lgHm/yJ072eHZW/Kx276TWjWRuf7DcI
9JJ7xayIZin8DbEzmPGTJkFg+Ne88V+aYRIt3IjC3yK1tss1dFJ9jCpY/QDu8/6KoMK38+WmSxZQ
spsTQyYNK4Y3cgfBi1k/k6xasmS0cY4z/UeKOa4/N1isuyB7OWxRpt2KVlV2bAeWMuKVQe9PSeqz
FD0HvOza7P7P2AbByu7+kTqhNSSwUuJoFakVAboX4zx5bg4xfCHDv/qfTbTqFxkwd5omdclHBtke
QHT9SD2iy27SBkNXjFUNnCl8b+PqQwoH59ZETo2xPNIQL6i4mLwXNVkOj007dMbBFvesLxeJqOWQ
0lnFDLtG8TuCcmeoOy67NZqrIecGOvtLKI3clwOXLpVcZCcMcm3Uv25vPRYUCGly2CkjRr5c7Vaj
5ZCF6rm/U/JbmjYaI4bBiUejSAUIeQKO+H+Kq0O+MHp0eFP+F/pMr0tUbXrRdSIueN4SwFvcPqRm
UgtgWiAZva8Z1pCfiBGhkdRHxWw8z741h3xa2Q92dtY5ldFtCYQWjaQp45TKy6gWIHO3fEWfdIx4
b9qll7HKB7JY0BY+PUsr0MkY/Xa94th6HIk1WtPv0ALFueAO21qcQrj9153Mr2wSsZqoMHnkvJKl
5EEFNZZOKM+1Amde9IsHf9vmOKkjYFa9+Yw2cd2xvY4jFa4S+Zx8tkqTP5e4JztbSbGJL5wU7sPP
0TDbNx9xcZCJa/KGpoAnO56bLkX/t98GUQK70+A+2m8x/tyxuY9AuRFzmlhm+UCKLbNU8ibE+TUc
l3N8aheTixpobOg1wHyWKLxswx9p9GM58+PRDemika+tIV2UGRlbZc0GlBmjdmghBniu88ZXeJ0g
QquPUrsyvjbt/nSx12lEZgNVWl8bAvVksuxLc00N9NABgGyQeWMX2BPaGjBT0Pfsyr0KBT9QTvd8
jVhjvv2BkUlJ9AaIB47mnbSbfwpYwOYRy3jrXqNZ73q9JsfS71q6XhcvHW1VvgEzt9t3R7/o11R9
NnHMNBnr4KSa4C/DEqksdB7EVeLjQFzJ7xE4vHbXzleDiQ+P0E602Yf9IHaX8+PPJIhrNU63jyoT
sbliuqjPJBxKO01IObrr5Q6D2w4O5+0osr7CVPyjerNkf91JHrRh5hQTHkokTw5lAqsOU4uq9FXn
qVONCZ9Mv8mr4GwXXqt1vq8dpeoPn4LHqXpX2W9PdOUGaErKfC+KTqiWD/aBsZcVTvXWOZ6lQWqZ
SDLx3OJRfP1ibXoSllhOFueCp5AtreCk4MYjxuoSWwukA7ghBXahfEmc53nL95TjgONVhhXYt3fd
kPhM97iFKsEY2QJTuvxYfrXUJUzkaS2gp4oSOQXPdL349leWKpHSkZpD00yxXSHLvnnaafiSHkat
v7nWZK3n3bk3tntsBpiuWsKZLSPS+A/u5wILfV2I5ABgnkYrJy0ihQ9d5VKjmPSsFHRWPEIkXoMS
JQU8RYbFH+/Cpd0NMTvPjqXADXCSbxp73tDbl0uqwTzIXZcWkB9zFmVpCqW8wgZKyX/UuZ+VHBdX
HLtNh15ZfH7sRXKoPfwbsYNlYMF9Lh/UOjqpaqOFhsuongtHeUw1Y6Awog7WNLqQ5Fvudr+O9fYc
qFfJ6IKvyqhT8rKvItInvRFO0DhBGKTVCXnAQbgOzzGIL4TasooliOACQzHXWWPntF7CIouo4E4P
4RxQmUV3hWc9KukEjFxMikKBnl2rZSpMWD8LIhapYzJ7jWym4wgTdjHvN/tYzECNx9AaWBB9Spq8
9n2QVeFD1DAi0N7uwOic/gv4e52D+t6rsuQ9sWsNFy8/pCXU9b8lwANfDdhKW4AyBLTfrP/dcYKQ
ls10IvNZNoWcpaslVNNLbAH7WemSqLnLkckMmClqcVahVEeXNbQ9p7Aaaywmg+XiHon0b5YTR2+3
jRl3UIUWvr5VvDNzIKLBTKmmz1auxNUdI0OdGPHYVf8f4Y2hFbdeO7A429Vo/Z95RdRsV4Heh0TT
Knxv65JZGTJSB6O0CeR7crH2vCwDjQ5qE5CxvY3yofZcJka2ySTo6+GhZzy9dIuAZjRxN5fjs19u
Z5lE0VcqhtFhOxfQ+ZCeJ1qTsM6WPc+gE2l2PrkR681eYaVFpiP2NQBhOxe2AtkNYGES/ut+EeDR
6G4RvNlqS3baAimZ1blqU0wqzX/AQncaED/yE625xAJ92YIggDuj+MA5M84/afUqnZxiF5htJeUx
GDp5wKmqvTXozkOQBFJBlRZ6FDQibg3YZv0khvtWmVggBkWO2z4oGaCmJiCc2A5C3jJ889+EgAHZ
s5o3JEWJMsuf0r1CFeTFQfdWY8giB5LiKZA2nlCKLE0RePArK9X1k42Gbt5C3Dsv/Unc+9wQNNfH
TqGNT7SranPAOS4dxg1ZZ+nGVwXwKUIBpSNwXeCvaFE0I4rPXm8OrLebZrBcK1FKtQatjA4Ak3kH
ByIm4Ig34l4NX++I2YpNntTXyWSnewuqPnCWyEpXdWmFIW/yj3x+J1taRZLEvj8OoF3ecf4YYM6G
/bie0qR92gPO/dU348WNXXep0RRvT7KXWWrPkTDliH97gREfhtLddTXQOXhbkAvo0+l9XXCaPhuZ
p/j4OwIOvyxikcbpQcyPbBmSEhJAHqs9OrV7a7KRC98GrJIiJ88nXD1Ecq5t5d8imRw8fwEiruKp
VD74KI/xg+7ZpVK8gIXgrE+uloNJAYKKbmFe3Y4Gu97rPx04TNC4Vzjw7cLI66c+CPC14O52Slv/
tBiuGZbBVrqTkzWI2kB6x+q+diuYmsYQriA/6QimvsnA4zIjzbJ1rVsY2ADvVs4ok9yQ4XfD6OMg
B37Hq6tmf3i70k18+nAVed0/xmNpo6+PqOh9Xv5w9d/ZwnGiba7ChevlG1D5IqhElO4bl9TZ1BMW
ba70bSw9rKK/R5Mzl28l1vo2KQ/yd24k304yYRCi9kPWSiktOsSidZA5FBltjye3zRguIyk9onh1
BUizJziIonu9m/+gDbGnaeDgcXQR5JQZ61CkVCWJh9n67E1Iot3unO1TYeyAzrWi+HxdfnYWGAXK
YCrqsAyczuInAoWZ+yVa33r4gt/PrPoqJ/8bjYDKIZwXnx83C0tCtDmI4QTWvpVo/nsV6Se1SddP
RX9mXgNkiQhASHhZOB3yhoHKKaOge08rilCIIIxdZG1x7dX/jiu7q1RhXLLVRCmG45b34mC+8yOC
aACUUzlioVzMNaFnuxMaldfCrOUm1ZYMYMpX3dChQl12++rmryJe0eIhjeuX4SsnAyoUZPL8oRG1
Z3p4CJ6TTioB2o8oOKG5a0dryTb7Cu/6NlGnw+zL4l/KeW+ShhxOOzQJiNzw0TMAtpyf2B2EBTy3
of0LOb41POuEtlFy6CcrZDRR7bF9cXTJTojX8uXjIAgqhedfqZQYWkeCQDj0BWvbhzJNGT8CJp7v
rrkn6nBT1nCb0IfnJdoZETP4mec6o6I2NC7CFtsppZN8AwFEQa6WrrogzmtQRKXNymBNeZEOtq5g
f2/lGJmbYde69/tgzKwKO6Iu42vyLCHhKAG/VHMWDO/D+gDf96p7Q8LbcqGp5SBlS9CTbGk4hFwZ
tF8JNznt0/Z6VmdcDGhf081lyZn8w4yJR4VSjAxgdv7qkcFTSEN0MiqkMMyDPr06DOwGzDTKrDTR
llS9ZzlDjQk4ByFFYViRnQs8T/E7Wdl5VgzrXe/ZgzWS/nj9J4fq1JSSsvY7O0rp+H7kN2Dc59eA
D07sKpSuKWKa/Wuv6Eigmqmvfyfx/856zjuaC3w1mwLF2EMRNsyI4vuKRhUzNTf8o5MyFJVHCKxs
SoHAEvSH7qrhdi0sychhbLSDvce9C6Aqc0cqn1AfVXk9/W8uC6eGNZOviqFBNU3tAUpIoeQkYLcl
sgsAJbPUm5tuIJzu/R8MX3Xyh3IlvAmZtjgK4ZKTD+1LaylznvsaQqch3agpf891C2dvjvngjlpn
C/MZ/ZGjt2rmg1HmMwEHs0E27k6tmfOsr59wbAMGdzr07ByO7ThVz7Brj7tEL1bgwPfi1hyG0BID
7hmticmXAbmRKlrI1upj3Q1GXxQbpN8GVAP7LigbyvGdVnD1IIFQOeG0jSkbNuLNQOmOlHK47VqR
JSBze7uk1lIL/oNbGF213BYPizY2xOh+dklds4bmJGYhnSaj0EIXU79PYZt3WER36k2ihG6nRg2l
VGm3EClYx/FdEt0BFyI4EKYHWCsooVGs+9CJBeh52xPjdKIBrxRGfXpeHPQLfKyj8CGrXueAZJF5
XmkubvQvGRoxURIsQZ91HT0bbm5YrwySFVFzewRw9Gy3/BlV5uMpEkywAROAKy1YqdgDlyL/EgTI
KIyYO81DktEn5zAzJbh+IsI4HZpqHa9VYl06qC2gBdVaFALpxWJOnVOcqKtWeNt/AzQQxraYf9c0
Wu98CTtBlMrNfvezs9uBf/vCDxK5+Q4YgPcaV/7tTWEtL7qreDPTZpfVag7DdhQ7Vd007ObVb8GK
fwM+zvU05i+Tb+1yregYfqAt4xksXhcqFcaPcb5px2gdAhVISed2ZWs5XTOACcqwBAsAmi1E92vV
DEZd1l8HBNwq2J1XnVSu5tc/VUbJqyWUl007v+Q8ozvFB4rJcpdg+HcsXrccqd6X6xAMeSROFLsg
V+fdXOQIlhr42LxcjB6bYLH8M+a3wWpXq1wAr70sbOM4as9Y7a83vY5GvcEnrN5KM37qfmhn/6c2
DW5sTjqMmSgiha6Qi9XRKanOjmvrj0+aHFuM0n0IPCCF0iID3oA5GmJSfrPQKv4PGo76BtDg+UNv
24T9yTyXm+hi0VUxvcfeXKVY+yK6MfLJpjUYCtEeYXcKhuiYpSeQLFm5SWz0xZmHw0JsQmTBHyPk
WOhBMAiMWlKNPaZhv0tFdaB1HO1fHV348CCvWUhwiMO1sK6k0lEHiwVjT1e3LWtWd3cL5U8Jv+ZS
b9W4SDGZd+l2atjMZWKLTKI5qlHcvTyL8dsqdXvUKOr0b1h0d70lSZtsCPD3rIXzuGb28IyGKS2f
kY9Ogz+wiZrOrlUyvRa3YcQlSqSr6O9CPZui4k2nlcWWZW9qLLvN8fThgKb/nbWnaQ1M+1b5NTy6
iNOshjP5Ja2lBTJKj740uV2XJs0nrSLh+OABavXKPHUwZlBhM70P13wTqrW6o8IXYFwx9Z+wcV1+
RR5qA+KtwX7CAWfOjaLMtYV5ftCjf5D5S6Oeo4aVqbA8K45NgGEZNJgu5LaD18eNhuX0AVBKU/pp
Uzne35LiwK/HEzW+0hysMrJ03Unk9h0KXVmGA8uXwRGS9K+RkDLKdtMzUqgNp3YM1hEoNpWdWN5C
iQkA7RUO1Pnm/KMPcp+kq2VJ8mFPd+Y9De7ohtkOiFlUgwDc5w1upDYwXdHvLTGfY+v8UN1Gc+0L
LHl10IV4YR+FfC1oPw4iRthSlEytrMMJ4OMR/4RhdMIhB65BTRYL4WqoxxBz8em2kui2zbQnS5oe
TIOJ2jiipJOUY4v0ZifOPRD8OfUTmlWLk2yFJTJsQ7XWZ3OHCpk7rYWTSV0rkoBf+UuLalyzpOSF
WoKaASoVF/yIW7kBBKZv8XLsS1FV3VrCBzm79D7e7xFkVLAytZYc0pofuMB2lS9NcUFzRl0bWyZH
fYO8uJm03Pxnf0RZfaRjppNKhGg7jphmgxFk2u+8qQldheRyPOBOEgUw4g5GgYFk7OlDGlSYG61v
uHjBG/LR+Q7u10kbFdVQ78A/jfVyc7ZLhb5j92lG3A21sa8lFtg7QsDTtaS2Ensp3yiv+N2gpAZ4
+w4VOjnG8v8KBgzlzjL1Jcd0Z9DXRTFx8Y5G1TxQ/tmElct965OSDE971D1YhZo8TNPLCC86r9e+
BB6AeSxeAvP0L47+dh2P8dNmqBz6wvhZOO8Jq0gpzjs4BsDnkBZ/wGeb4i+Rwx33rLLwwh2NugAW
/ZDNe3kdgeRLp5d4ZmDpHg7ozMLGZpUeTlUfeIp6Ba8nrog2Qihu4Nx+QEWIw8TT8rzx9xC/OyKL
PUIV6iwEmWvQRqRMrY5vCzwHbNx8B78A1wlsImr9UBgPICWKAGqXgezfTCeth32gposQQqlemc/N
yMmYRLmbbaqsYfc9MQgDsVzcNMOxUK8BI3fOrLhYnjnDXntMp/9sQ03y1uNIGSdRi5nc5sSEsxuV
W2/wO61Uhv1bGO3nlUMxSm+EXhKYx06yfEUG7CchAeTzoYDMaoydoMd4kPOdxDAaPn1eWACKOIA2
4/6gxk3BY2yA97lW/VlHbanjka4lhuG323fT+Z9XbBb+386AtXfgzxP9OTLaAEeHojBbatXQNBeP
Z3Y2cYoIsuleiyKdMGhzckP03N6B12JSpOKkL0C6by/poB/nfyqIHH6tw6GIwJXrymgxUX0zTwc0
Y+eaEyKiuZutd1IRUs+sfeY8Wiu0pfXTjHi8Zrf4AJwLtcwi0kkh6ukc6gLFTg64im5zpKCTyqSp
H+mT2+z8zZhuiaHn3j6g7ZgHxrv4okAoUcvwKxjrXXSwOxMEEqFw5VshO4SyKqeMjvzjahZIRnoj
3yl/GY3cznzwqbKovoWJDR985lq4mMN4aIVHkDxStik8r3mo0r7RXbjasvCK53Y9pVvgWEHnSFku
ZKiqWOgQyZ3epAxA9Iz+2TKMuh6Xw8onfKXjHdAOqgQVEGyeumm7g1p1iMRtR4RC2baSoC/Rcily
yywScEBfq4bGwos5L2chAxTwoqekPBfHGdtGahj5x0Z1zm6HUq8HaSyzLK/6BO/jQLJyzOl1rbw3
dzyqBVcvQ+IBB0pC4nt7BKi4+7FqbuZVyXpfok0Yg+vI4QmseZYfehy1LLgO36tHSJ0Y2Nd0bpug
bZKgB7KytCFWdxOVOtGPAjQFCMaJNIDDcFHZd6N/aaMQYRjs9EMDIMDx0GYv+z/PX0uF6tqbSqkc
jld3yHnxVkARnwrqRBVcndWor4swzmiAmTdTgJ49Gg5xak0jUYB7u50wv4fJC5/rzLmeszn07SW8
TnzNZshekBV7YV+5Q8ysVp+Zkjjy0jnkOl6mVIpJNgd8dTQjY8+fVYxG0MENXxiY4KpGLUysgEuy
xTw4ovTHiLnfi6x4Q/MuvYlEV8ns59TWM28oG/5g05jhePxAP1bJdXb6bTRc/hISVaixVuRgDfbB
M6aOydvIPEWG41G9hVjF+DYoIgbefmm8vs88xjmNftqlRbDXrVvv9xtckmWRWz8VbXmSpkmvoIdw
QlfeR5SLCbISWTFel0p0uBhQ9w1N1o8V1Opw9cLSa4brDw8K6Ubsbc7ebZZCrfApXbwiGRmopo97
6r/RB+3SSolSGancAn8VH8zGZeBWdrVvBT5ueiJ+EJv//myuITl7noMPTiXY+pBiwL6kmAdnGtyD
BD2+zzMi49bTH0j+ZdQeRZljp6KGL+rnoyyqXKdKGSIRrhMCyZHwIWZORpASf4NmfxI8WzAPsr2k
E+xqZtdyY35zlafDb/G3W3RghwdAO3IXgoC93QahEcAJ4DLgEQ+23itNfqUNR6PGZIWqNPKUG+uh
ANpNVyGJ30wT61z4a9oAwaSn0qHBGw9cXCH8pALFKnLo6s+lxexdmu5n+DjTI1JMf5oX40iw3Z54
0V97/C7iqG9+I7Lg7z/kNCTvoL1126MrHpaRJYgFSdzbG/XkcTlPT3MeSIaiZ9DpFxxK9obMVBWQ
gau/I2Pb7SayAqLNlGOJfHbfhCzK73KTqpWgIh8Ilhgk2NX7kopYcJrrjKKLBqxs51tndASkO+ei
2szlpno91W+VwbwL0VP59kbVffynLU+IFBBoDq0hXIHbpsyO1ZxkaCMLtSZfVOqdRZswaa5KmDHC
YF/cTKOKu0/rKdxu+EZkJ/zubkD4aF5PydB7FdEe1aoC5PIl8cNmp9JqEHgoPobDa3fKcV1m8jqz
UU7SGssU/ZXcWJGSg3VzhuDxC4B9ZiDeUR8ZqiZXmgrg8Rs3Sr2ez3S2J4L5wv3a08SRypSSwVH9
QFe3LNd1Q3IXXnkB6N3vqFf0AixNT2xMlLW4l1h26cSerJigIwQe/Uw2TwBqkryrQT/pyGgLChNE
x1YhGMqd1ROo772bVBZ7vCHDz6f7/J0kFuyMyS8rA46UE++7ZWyz8L4ZEjR5p8SMWRcbcno86Eym
8dSvsVvQqGEc070vCEx5Bby3i1RRHCBmvb9lJTTgiT0xGZILNyHmj83mGwbHAuFqTOqzFdJIuDp7
HF9nagtTyjKZaHJ0xsRghMMxI8NzHBlGr+ucZwKt2gcGytWGMW3OJvtHzRunz0icqqpcY1ePwIN1
QeSOFdnWupXVU6iD9RiRheWVDr6kktqWl8tmuxqHn71tY/tCGnx2ergvFK2OCMYF024TV4SOYJ9a
wPjaiY4wQCssqsRM4qehu8NNsg3Bq/MVCsvSqSOSQDrh+Kd8J7cHfMgV+hiRn8vhHnxr1AEB/znh
V8QKClHaH8sBgNj7uy1r5NPOdTdBwXTKn8dPnsMA4O0qWZftUj/iDFONy6Wl3DcyAAdeYdj3+br7
448ubWvSTaviGaEkxYpBJgHx99kFZviaG9ms1iZMfPyyapQTPRFmEyOjTey+E2/mICP/nEzvp70e
noLEz+bpFtXPxficVrxqaMlwsJdb1yOACp2OXi4g0TdoH48xvTte78oOcpFlDj5oAraGhcaSYxwG
n7V4PaTUzdxhJeVptqxosFVBlwztR74AsH0P53vTvCknsteGLXP4CbFXRZKvxY00I/esK6pXEnId
ElkeuQm2zmH4FdClLcFr42LXOWaiAZZEJ4Wa9LIPJVNV45IsRqc6NQn2b0z2nCRQ7p09IJLb02xE
9k+hPILGCGVf5QMaFlWB4jx2yn/v5Lb9Unnz41XMwuIWgx2Hko0P/AKukMtEYvoQPz9JaRHOwYyz
nvfILUsviA0HjC0X8CqQ2AFpOFrLSxG+5owzBtg+JrfD3lrRHIcjLaeB7Eqox89Q4ZRYwolzIBJC
uNFQ9EP5mZ6g2feGVBzJnT8sW+3IX6TQEEm5ayiJ2oZ1lHKvMMmM8HM+DkyRN2vtPJo+/yxK3TG5
dSUNua8BR+oFZiOuf3qC0rrypNXiaEtw3lpirYgJ037FGtmFcHJD+bcKSBeMy7zG9+SGUWF36nx+
u0xh3d6b+1L5vsWdftZh+31L53LK7PJYHw6ykD8btea9zn7XunDywrNUyRuYqZ+ENGs8v3zI9BZ0
4g+zY0ZEOjK6mVC+Xm2nVPyfrUCmr08El9XkG01vdGL48x5oKUWB86Ly8Bvji8d7ORF4EYAdQPDf
1MuafS3HUHZV6R2WnykKyXsHbSTJQmJC+kOglUjZvOlQgOqI+uCABn/S9GTddCr8o/9EJKtNfPaU
x1fHJlDLFdrb479AgQ7ue2w1rPiIIuSZMTTaGGPypHsQ1QKbyhnmo1opvwlM0v72/eX7FKtMFhYa
QJZE/Xu9CES0wG9s23IR80yMHVPB1o6k2q0CdMwtKN6ViEr4h+RZ1qfY31vD0zKCcXhfIUeG4NiO
1sa7VRpWmWgEbYUuoeys5VlQum1/jYsL+gADY9/F5AqAntdD4jo4l985qwmmksTKzgnyd62RgwpP
fz1yZhJKINWSCF9uJCobQLLw46Dkv8QIZWpv/Q1aSn9VWn57RdIy/omt5amTa802c0YI4a29L8Gu
Q/b+1LEHxhSX/jM3qocXWFQpC1oY5CZf3OnsFLuj+jnnUd9Ra7YTEJzBjD6t6bE1Q6THLtliIK5L
JWGYU/0lwYCxNnAffNtvADnCUg9fXi6LunMjHGbfCTfKw4xZXj0O8NUeLYl8fbYHNAY1yVR4w4o2
PpmstGIoWpMemrUGjHUPXyrReZy/cX1WdJYTKrDg10e7ACYRz8SFSHJPOEEVJfjZsz8sS7hwJpR+
nIoe0GZzHgXRVpKblgF+VvOYaAB1jJnMFY7/QJdkhK9DrNGpQ+x7FtwdVKfEX7AHyO8K/2KQMyUG
E5D2MiamZklP6CzLWvY4zxZCwRP5PsDWDo+9pbyeDcD6APpy802B1Nbr2MQ0nCCQNKY95KqtCKXu
x6lJgqjF494fM5weqJBL/T2rjPWPfZYAXCBvo2UcHXPN0sAgKajSfoWkUMMvJnyif2qdr7kCRuMv
RwPpzjgShsE7QgTWbmDIlRRVkEZO/r33afh6DL8w/szTnT64DCM7vtajUkM3Ekj7nPsIkLV6917u
JqnFktb7WgVKx0Fru6NQ2KZaLPV/FawS3LkPXtk+flt/rqfV3XsFV3A8+Gyr9prOZrsdd3vZKNIb
XAEhDogJk6jIr4/ndLCXvO67bcd5if/Gm5HEDtlXVu4Se3xCvjEEv7TmtXpSmt+gD3qkT9zOIrZZ
ae8K8I6ZHh/YoqA0LvP3NtrRDQb6noC+Xp0HJTApOC0yRnccgWISrocExDGqRuJmlyY3Q4WVv0ez
5fVgK1iU6mlJbRPaS9Z3lNF6oGcJlRjozYiRQkuxA4jTIDSCtz1FP104JNUGhyfqKNAS9v8H4L5M
SFwffYtshB6htINGLulcP8MU9j+De7U+jl6AePeO2DbGV3UNZoGi/bj4PPmyqEG3U3HR+bfX56Qs
vdjjQWWD3appXrRjojYBhScR448rQV6SHWrUZndViT2kYQTbq7Qln7wwVvhDzUSu2ApFGo7pXGH1
9xy5NLiODwnRyQQCFYIHcs/1tUiosF0zTLA8ROKnHjSNB+2VYL14c16XIO2p3Jh4cadHoLtJ59yr
paanK2B+HN5cmTfa6hbuj5drHHVw7wFiTi/W7kuSxYGrEXBvuQUlOsFcSZdztm2UaZLuh9nevoAE
5yEQrRGhdqPSqpu/SGVr9Y5luD2e230Ml0tIN/CgRD21tJqChcuPLfzqeUdgIPk61sGx/1CRKij8
oLUWmqhBhl1E4vCa68mpz6g4iMHEXj8xA2abGYszpyBaGiO3St7ZYc9sXTziW2NmXeITrEBAcRdb
D+Boq0JXCdzg5vQsMdEmr1AuYkfdDYbO++aPwK8PlhddLMlNz4sPgVJAZVZ2h0SOMuZUUD5/3bhg
VhZPNQErkPC8njSJ8ljN5MC6Fw/mlKo7nnegBujCgclk0YJX4uvypBvMOE6uxIygpr8+43Z1ZRH0
5AdBQEZeCwhWo8iZqfs9NPyQocfGVHXAf91zsQkw3TklMm3rTxw7JCr6WDxNsPxOCfAm8fPEgPNi
MzynfTDR7LuqarYM9clZfP2ZBIBQIj+HX8HV4nvWtGzJBe4CmBH3sRgvGE1sORsiU8D0uLpVcP5V
Kz1IHBo8TmGZmI7UH9C/7ihPdNH5IM7TXNiV1coPnm0DpxWEtzpw8U4tO2eWu69DwKyZiV8yOCbI
9JiuVseznuGFqtCW8uJfAWLvgedfakqLg8Xs2EC+HvE4jNAB5IRQ65ITTcPJ8e5ZiHw7bhy0DPwv
TsNXfN22R1HEkofpsvb2nAU6a/En9ZNBA5SJLUnVY2wFg5EN+9u15ilDVCCsHhAG4GUYhQKzvYdv
MngD3gXuP4Bh+GS+tDksSrGxFAmPM2IuIoEb/zPiAhX8KG8WsoTnr+5fslSm1OO42dVIniG3RR9+
dDKYr7lvlYKHuvbJWXheKdwDwmnlUXS/T9OZRmLWHBm3jPFETiFIGzEi1ELfUW6Ke//TkzOgtfg4
FYuiUDN2d5Qp0hLwxjg6Ns/ngkvsnAIjlo8Cppex+gkBp55t0wQHrUxrnKq4YBOyZUt5e2F7sVKi
CBcuDtvm0XXm+aafS8jVjedep7gDZuX3kjmsmFNAMERvZaSxAaPgLErhPpJZMx8EsQV9zEZfcT3s
Xa4oEUV2wdJY7TbS25zSQcuy0DLT37CFaLgi0JroMoA1G4xFsX4KBL+/N4fxHqFfyDUe20BdWe1a
YCYX4Hvd8ToiT/wCQI++6sy6BwpUVjJ2Pd8S4+LeNwY3ZtYpaxhfAmbK5yUNcsdolqXYv7jMaORc
1F4NPybRNbHdIZvadNBvcB5TIOFYOypgSvXbM6pBFLXZFOEKgGZ+CFwDPFmGAFbuiK1Ydg19D0sg
5SRloPNM9xcZf6OpmWmXBFox9sIy72O2jqAq6DzLqmlb631fCD/OhR0crPMZasuZmZO3+Z7QF11H
XGOYWkbLzTMBQEpBO5Dg97D2iq9vNziQ/Zu66EWTMo3HtLzwua6X9KEcUVXW33gFazsGdH1tm7SO
wr1BMSrPm6JdMM8v14PvDsUddVYePBXQUmV1u2LMlxfbwL9xVtbD29GqzR5SKymQMzSLf+vLRev+
iWIhdwcV8glZsGgI6Lf9N1FUvNxoUtdnxOJTDvRNU/SqUZewPlBIfkey2bbreJL99onEXZQE6iAY
KlR7+XG//F0lq0J9YE8//5lA0uZ8uaCTjyiaH5QG+zVNk8WVE/C06skg+D7M1w0oA1AujFF6Crd5
25lIZiCQUN1X3DnIltG0MVF1+LdvS7a7VlysAkPZKNT2Tuu7eYWI2s42f87l58FaRa5E9YSt+DcF
ZKNkuRC8DQbr0vvxDo4Mp1L+eqUA8RNfcCcqL0pfSeU7S6Hddp30Us4+MANK2PhlsWq2Xt3I4XBz
dVA70k8Wm04lvc2HKs8pqWABG48aEXv5k+4JhFc3o+1nRsEGL28bdzN3FKwOh5HQ7TDtnMrTNMaC
WR6MbQ0WK5ur8g1VWNXTo7iwy/0zjPCvAD3uHmd2pKLSfup1BiqDgZq1IsCEJu65syxBIJbF1wE9
1KqB2bRwy+vN9mebgudYyZuR31l19dfwwz4lqrY1sH2LWikaPIv/m6u8zDjAjXbu2XEsjM+IUthp
Kc3SAHGykPzeVhJtIo61dot1VunMb1tQW9W4UDOzQ5+MHpw2sZ7I4gEFMDuaE1RRleJbKlwvUECY
fnWombh0SjGUD01wKRbt78mDlmnrU/25hscpIXmsKRWdeOdTLdTl/2VlUJRbMViV/PzSjUthmEcC
9Cm5u4+ka541VbDGtFMs4k9JARSsdKG0mrBhj2tW44h7htdsgjf6PgDVOixUoXtEQizOGhtTW0wn
SEtePRv38fKe9mrhgIG6YCc7z2NxQNT3KAjnSOiJAMxILIDWqlQVNf2cjfTbkMEwzPRxRV5pUxaG
ZtqYyrFWqpJp2NICoIFcYl+Qlcer9w2wWjCOWBz3Nue6Q/71dIWG/wifzMhLtIYbF+GMYtwQGsRp
p4y2Cd2EGlYRKeZUTGAN3rIgzTbL8hvmZLOkEqAeO/89quU7zji8NKr3pBLEMHrDo9neCcrR5rW5
+vK2ccC0/VI9HppzydZQdtfsvN+//tCbreJemblS42ixIHDxYmVK1OK5SktixO8JMZrj3KZQq8VO
M+3ECeGgb6rqAhCqM7wn9gDkPr4VqINjLE/00Q+0LHygFRgp+6WJ/wiARRWqwszwFp86f1Wy++UM
T/V0vEdwMSIT1J8MIw+YAHGxx9/vsZ1vyFHcQRmxv1+2Vwqo0TOhusytagxmNp8S7I8sjHIrEfpk
zP8e3B5cViXv1lVjxmHtrfEIMnr3Nj1RVUgY5Wkf40SEe2gr53I6hwj+Sc+vA6ILT3sOZAbnqCD2
eUe2AzLbUX3/u/FWywOQdi1wvlgN0oiBDb6iSjq6SYksl4tVMyxjSzQQXac3ITlTTEJRPAwVvJ+Y
CjS78lkgxrBzoRyZa9F4XmsET92eXm3JZgoIdHd/Mm9f6sS7mxdF++B8kjvcnxRdlVoiGebTHruL
bVk9gYbD538FaMXAnFS5Fn9oywSX4LtybAXouOUdoQ7M2bLkYlK0NEzRGICT841vyJQ+vpRT+an4
nshFGrw1LiVbYT9iEfARpLAeg+E3Oh+Io6IeRp12NirD7AAErIflF2mZ7SFt8GrUDM9g5xjrrwVx
9QjwAi2kLARSP1TgM+UTF8LePUeEhvnb+gtcmwYkGEwn886wwFVl/NsJZefMbtr2erRwgp9p1LxJ
jJPUEdLMNS3+T8jswQNulTLf9Yzyh6xraL65uaRA6dJDBfEt9b7IQj9ZZvF6g8yCe282uPAJvsgZ
hd/Oul3LxYt9u18jN3EwOsCw6oUaHnxU6Q2VloPF1rpFALlXcI1UmKN9RP8TZ9Osbq/AodgokSV7
TNIGKdPMVPE/Pj5qTjQUEq7b/DJyJITpKo6UbEQvZCcUINcPb6yBhAXL+jHxj+G9I4awrrIMRbvT
5zdn6pGJXZni/4+pXBXqXRZiXvMFcpx+e350vuD92HmxJZneke6DPAo2kzIeXF/9DwSsdUeo0glU
lrIPPnpSIGOAY4WHH05lSPYfs+jxnGB94+BdKsJJFmQd53li4ObQbD8AHoxtDgVlZ9FWsSxxf8qu
gKm9nb6NDXXw1azZMU70s8scB3TnowIwbkBKUDxBZKiGdLfws1iPXSetNFU7r9ydKcSJFi/RoAbT
49wrPSSP6jrsrSoivBQs3ShWI1jmT9GoTismsYc5SMnIVsODeVd7raGkT4fmNiGFqnR1poAossg+
IGhXjb1HTcuAx4MBziFCaGz6BKFnkKsSSN6VYBSc5TXA80uTyge1yTZIjpBZhRJLvjELrO3qj9UC
TVH+Kp05UwYh4VXpWxZui13NYec5J8Z7/BEJ1pZGrna1r8v4fHoZOJa7zVZuR8dbD7cRuBPgcwEF
EMwnyy/TeN8i0XjZOINyTNjbeO7NzM6++IAQhWeqIIG+8zXRJ7wgEm4GlUH5Jxo0foaXx4poat91
J7R5VmP7kxrKYHvyAny4FVk36NOqv7A7ID25ehOT3iXZ6MFPK2TYt0mmL4+atoilLqeqITs5ujK5
yL2SGaIUDuK6Ny47Y0bbVD0U3TdmNtaZycEWb3OjvmUzt9z01KF7cNHygW3ReBDy1PnT9hFTTuwT
gGZO7Kmvjuc0aKCj382bWote6Y3GFr5SUeXXk5ZnMSXWsaR+wCAX6y/i4uR+HwH0ELAdecCoBFAm
26A/VrtB/IUQN3jJC54htROMb/ghLkwEvW75LE/sBvyDUA80HmofDq0EOarHErwsgY7NNM+NSmFZ
ilw1k5DeaOMGDYEmlDtebpiZKakc9gz84ywEANwRP5bKB6Be9Kpi6VrmeeOa0KKbMJ443pcKd7TM
aI9mFM2ySh0RECJkZYVyP+pwxUQ+jRHm5HI+VJ+veKQcuHE3+6u6WvgbLgEYUsgwqvBp+4VMAdr4
8D79v5jk/oZ5iMdD35k2v6982zOUvf3oArnXl0LzdgohSM2aH9n4RasscEUj5fTh7yT6FYjPHyvn
LYRbGhxY/07gDVlTKUaO4gWWgg38mxaTjpqmC3pmLguH9ZgHPfkZ5HfBaHR6KTXaB2BfW+LqU4nz
UqJ/OcCEte4Ynggba8LkSj7kRU8fD4PIuFoo9crAXXETQLuGKhA/32U8w/frcSRKjgGawT4k/W96
hPiwUzCv7mnBrFiiIgUkKip4jDE94fkHJPCf6IoHEhQE0Hjq+KdJimuegInkdBi8ZaxAHov4hxQ3
VwsbWw6zhNqzMM3VO1cr/sznZuPOF29pz0qnqqZlvjyAetz373qkLF+tpuRbSkmX51lOncy0BHuE
dlHg4qiJq6kT7Uabq94TWj2XkHSo1SVa3jeSXnv9YE2ov8NyoFMUMhaHJVg/i3yS2PsRn9rJqKSE
3KFPLzZ8bIHBxxVi52irUVxpvLCCQxGAu8/adE5NTK9wO4X5ejZpflloD8aALIGhtkUAvsqi6Ql4
Ss0Tgos7L3CcruHc/q1FSnMOIxFNqJOFK+atVRpxrJ/qn84AxPM5lT6jHdmdLxL+3d7AJFB/dg/G
OY37i1VGrLErO6XUnMG/H7VlK6g7GU7AUyHPTXyVrldx0ftnvCBsGW2HdJ1MxxgdWG6DhNvT3P5r
gXjsnt6L27umUjkKDAZR4eB1gpEWEv4DOm/kw3Hkah8ED3+/oMt5OR3lDL5EEk5CbjKjszC4B8CJ
QC+4ShD279SpVXQKFktWyqL9LbfHDI4ogNE/7hzh6dSAMsBb/lQkEkGLH02Sa5cHPhq25E5Zrqty
Fv+x/DkiJTAs7zBtJC5kimmOn8GwBVNBtRwwH3SQpRdbORhdoUXJl92rdvNzCJ3sOQQ5MkOmElZQ
dL/MEytLfq13BNlOm/0+quT3Bhlk/GZdEGHg1D7JQMl5lWcugjWnoShoeePtHYX+lMV/4stwq8jg
3C61RmgYNtNYaPo9OqRjiwnYMUQt/qelpKdroyP58AuIU3IHyfZW/wLBUmNVBhU8zkoYotXyLTsk
DNTrClJHpxFaTBi8Oq+oNdnkG2i9s0OvYg7jfyK99PZ4s2MXeMIK4u/KlqRKowECKEiA0to4eeo0
eVzTOEDAfzpD5mT7v+8ULRBJn8jRn+o8aG/LFnnJyglV+xv9zjEbbwfsKqC9HZSt38CnhMx9WCTp
FukrezhII8e+FeyME5919Vw52bjzNULQLD02UzfZXD7k2JeW1VBkDdmL/vVM78eMBt7mtokYjvxn
OlTkQfXJsaXpwdRhecY9nyjNcKVo+G39sJx/yDN3D5xr+kqZAIXgXQ3f4PVTWq2P+2o4QZ8YOLBx
/6DSvWqJp8AzC94SvcBBX+O0R0062KVkJmCLakQtode37pGltpTJmAmUD7UxC4BKvHAYlpaYxmDP
EIicQzc699T+ZPaBykodICqtC/38V+gwQQjkBb5eP6BNUziDaStaWumjungAXPKiX7tAOm3u56rb
NP3gOpC3OjI/b6IDhIYPKoYzGNz2n7vcAgH61QAyTGoWi6dTF1F8GX2wQqWh/ZIRQFqe0wW6nASj
LGP4R8uzS2Ib+fzCO338gp1CqVyPQWH8lEFHLV68C0enx2laXiwUS6T5nK2fLmkzu1yMmcqSn5TA
r1/kOybR+qZOvURbHKNuKsGqmYGtClvJ048fSI4XILX/dg5+w78KH2xgQGaSaEOHtEVH8tgtZHSV
kdJgaEAX3i1vawdv+eOEZrL9RcIcx73BFbNTOSlHiAoQ1zoD3C/p0La0tIB27dUZAtlUkQL9SKNX
rD/z5ndYC0q3hr+tlx49N3bXTfVz8MlCg+NEpgR9Sr7N6OwB8oJ79z4q49aVbqN6esNo2dJV+5G6
zDYyQBjDL7QV0+C1WgBNuKgFReRZG5NlgSBShy3TZ683r95kelBonWkUOLCjL1FF6/Mo4z3D2Bzx
XCoeL7AdSUm3Gnkh8kL/E5rSyVnnSE86Wjxv93k/jmpuHXpkxpklNxv+YogHoVQlWttqUic11JWM
J76AhnTL+JE2OLSVA283gw5GCNll+6k9IS5PDdBIMcH/ZDOV7cxhk3X4RGEEYza0KgYprdiCuhlF
zzEov7NTUnPmydT9LlM8m6B9LgF5iZ8W3vHWME5ncEpCpAn87GmqTBfQaxehCsKSLo5T+dNyf9ue
0cj6zWOtZ7L/sT0vx4ofVq9DArI0SZbFecIQE+uz+dFXsbelwxIWwLI5b61yX4g0ysfTiQeD151Z
309Dz3i5XIOhYfRLKsQb6NSIxjEF0plmt1bFG5jnl8rf+4xwAWVgTtHa2XKy8OmmC7l9lOogh6Cj
QND5bvyJtp4hLP0MFZOPY3CwuaRBPn0uiHXg2T+WunAjf+NZQoe2RC2/K139vUN2ok17yVgcGxxY
61ud4I7So4BXqI+yeMQIFbmnUC3kFpTzjErhQxeiJUu2KZpWKM2p+LJS6Z+CPm18KPZCTqNIveTE
g14Et193407qjEByusQCx6wsitaPPLyC3Dhex3hfxE409dguve0YfAP6Mfv4oOnbQFq8bBxWYHq8
cAb0itClbdA6/KptDzJ1R+/Q7fdv3IBanTrwLb4/5unu0wa7DY56cl+ubwptQgDsabHyNG/1C+Jz
W8t1Vx9Xmu4mtEGvYzWtwCjFr4C4mdpW1/ybwVm+Cjklwef4LT6egeiQK6GZy+m+z3mdTB6bxU4c
po0Crw8S9R+gm/zIucK13ordBnvbO3kXpxkCELJG6VNSjiFSxMMxshJgCyn44/p+vj3EMhB8wz0C
u7tu2pgIWQVW9JT1OKwqkr8KirxQB6zxWdRNrWWe8KQaY1rzMMKSuP0dp0j0PPxKZlNMk8Zg4ik4
MmQBUzaWr28ZDmh9fkpl/YK+P48TfdBAlqa71h72bRPoCxJgj+tmIzjnx0ZLLEVNeb2pNOMUY26C
87tmxyqSaCEDILNjB9zp3Npsy3SkpignudXYiFLAiofPYy0jEwkfYGKUmQD2YSLjvNVF3OFYrFmL
9/GBsGeNhGPmqt95oOXXjzooAtrTwsdoIgMnfzq93A8M8Slka8rX9VuT+mufyRtHg7ye+b0F0yI+
uA76dhHDuUgEPTNVAgVvlecuevneil9qao47oHtPZtntmuDlSx4wbkeaTA1oHiWZ8cVLfi8gN24V
PQE39kS9oYHofS0yFeG8sHC9CtXnbjzCU37JZNiiuPod6T0Ya5zvgRDGcysURhxxIHcWQj5xGPJP
+XCAS8l7K/Cyt2JE3k5iXEc+5A5gYg9pWNL/KrDrKsF15/aE0LcVonZnZHQusQvAbA3j2ZBEk9U7
sSdagv1lCk8rhMOM+kAIIRtciClLoUP5kUtaG+bJO5JKNXYR+35EGhEuJAPN2VtC0Y35giM7mwDs
JZhWgZwwEp6v03sEGX7SbCqDVEx2PAuYlSzfTqTtvz4b75YO+lFogkIHtVIeB/3/eenxLkyaLdOl
eN5y3U5/wo8X5mVATMUSjaBRP9x+Btj1sMNTbWaXeJGgAUMbvPSRKwtolE0nFTKqDKFXvMNiCock
4IMy6K5D6GR5BXT8oOvi0oCecu2OEKZYzOKLZbrnt3aa9WPnCQPvnA4TKiMtbCDIb/HFwgJ3n5Nu
f87AiLPoehc96l+tnOE7HVaZKxfPFpErI3OHobvlSBkVRwibEutnB3bmw6IY0TbRMypjwYLTwUL/
iybEbKz8CLZCl66v8eBQ49cduxYXykwAUdlxKHSnTOFFf+7nXAgGNpmvjETONuSwpPJqQuPyIbZG
MeG7ZF9YwGMUBRWEM5OIZqZyUR5DmmfwHav7jlR/DFDPJfvUiFsK5QTiYo7+LNqPALzE0H5tdXoj
BHPd1++b/GvvNUFO7b/GJKz34p49mNI791BZHTqEHZdj/R62YI1cbNPMfrHMbOAgzwUkzNjc8IXm
Vn0DLb04+DUYzhmXxhkWf0OGNdX+AwWI/btr4X3YF8Ee6uNHqBPlS5JWIiR0LjA8uV1p2iQrMUL+
8ismmxhDMDLgoLxnmYMgYQs5Ozl8pQvxj2T9o+cQBb+tY58V31TfDU/1VPGHOPihTRlBlP85xlG2
OYpBjrhm1NeIueoFm3huRxYKCk3XmlO1lf7SXJ3hI3zsDDc3/+G901sKc50lzYaYxraitraNvIJw
JmknZcbF0GcC8qQu4mmF8c3S6DMbZLyNYpi84jwf8O5hVS0eKfzJvSqugt7M1Di40xlh/C/ck3g3
5NCR3xNJWzBRhGpXuhrr6HOVodcJcGOxurkWpyk48JM2vNbQgR6GBl9V0NUzFp8lT4SjMAyc7jrL
h53cjtUfFL5AMLZT39DZsqdjBHtht1Tp1J+gdXkOUOnhiMNKhMsVZQS+eM/ulXx/pxi7d1P3b3ET
S5XdGw6hto3jpNrKghYDN0FlTIdjs7kYORdPlRSx7Ao51GYH6l+AnUS7M5SgHkqgFX9Im63zy6ey
IrGiNktvcVUlvnerw30B/u24rfrZqBgwwVOzdv6X2R0GlvjgS5ihXIr1j2agP6UPBIo4VQeOca3E
RJa5j0P66O4cIwl8cHTr8jbf0rgn5aL6GxUrdpdQ4jD7xRrQtjed3l0rSn3H4rnsMsugxgZDLcI2
JZOKXxp9ciVB3mNRH9rG1QsjQqoTxICScU7v3a2K83gxKsnukW3MSffY4Hi7oe/jr8DzaMYt+nGi
PP+lonXWWZBv3iQ0e6b7+Hj4VJNZu2AXFH0OqygTkKjq5t7PVU7lHmqhwwUFXNaD+on2+0z5ZmwI
F5Rmnw0hNGELQ3YRYPdtI4BRjpUe5k8ZbudOMH1SuJyUxz2B4xlZxRxGDt7hqnB6WeW7U3st3k/W
l5Moz/FhzJ7ZkLqzH3AChp3ojntTVAg64jhUFFPnlKZf+hq6xBoRVXeKcnc67H6A/DhFGT5lkZyk
SN5sQ0jE8fqok2i5Y6jHz4WHvEQjaaV1HewL2SSi9Of1tzf4/tIRz/qcP4YfCwNcF6oUYb+YwNbB
iBHvJGQUsxbKnftbyQuKSCWeea9vqPN0BHHCGRGkKlSy9u+rLaZGwUuJORBfinJLq0qXeNjosqwh
0DnACl58P39TtF9UuIiIeSo5/la5soW/usCbutisxwBLWMf/Dh/SQVvaWxAPbB6OCOpXnMDqKGHB
G7ikuEiw7R2EI0mYjkH1EfV8HGGXBIo57I1glG6lBHynw67eucON5Ywe414IgstK9cxkSeMudM+u
p7dbjNAV+Rx/x8LP6dKtugM5vip8Xxsh7eddrYQh7I/kLog1DUn4P1mbkZnaRkLZRaJ4Sv/1sZiV
Sfmte30yDIa2kYfaoF2yp5lZ3OI8SIJGafHQAtZeVAhX6cg6bOR3FKJlaDl9YLp4Ehau26yXiBH3
I9hzirNrph4aQga+LgxjS00vij2zwJWGOQ2We4QwJWa4bVLoUf/nEpHyDhnSDeTDPKqEGQlJB94N
0+94Y+REl/HB71CpA8iv0pOrkxKHUeyer2rrTNniaIwhDnE/HyGPqJz/38UQoojnwb2RmFo9vIK3
t5chsKyFIoGLmtXLL0gS6e7pBZ0GnoKOCuAHIs372WoisGzWbQRRV+uhITnccbbfIUlFkHv6s0IN
Pe1BhwW0yEoSwiA8VCcN3o8nstyQMvggfVEDtS8XVtTfxXwJUkGermYg2/QBTa+3nJuBp/Jz69ER
mauv1np4hDNCODf5CPvI5AZzF+kxVyzoOUiBcScXTekuOA9mVjh2uZB35k4FBSW46hLHNrM+Rcfx
i/wO9SrUuhFAFnVn8gv5s04v4Lqh1fufJqHU9Vw1IitLZ51JJj67nYgBkDwzOSNBSYxPWAZInEHt
tcYtkpK+qdbnDpZrwyUZiBHzsQb+T7lyyr3wmJdwlboJ5GiiC74gy+ZyzX9ir8ci6ty7wd+FBuNl
rKV9d+8LWXlIamdR32+tFFFrpWFe39sHkA3x86oO2zD9agfpfhUPJ4GasSJQ1FeWG5/iVqXn2Ddi
elzDY6desjW5yHVJEBJThMCJL4i9Otn/yGYfiCpa7azDygAf1FXFaWnJ8mkiekUzhu9b66G48NRf
QCAGmOaNVGzHJI2ThQhDOdn+M8pY625eLIjZS+x5Qxhw7/FXyAVSbQToVqr/iw9UkMEjRigUhAR5
iMZg0NqfXKrpR9XDXHWygECDxLY0lrFsSnWoV6lPpmaFOCv1vMjnBupKQvazFHIaei1dSb80hHnG
wOhS/p5+lyvChMQYeNWz91rr2Id9TB9GB/Hml9ugBGEgaSXcDQqsyXSOq7uUE8j3zyyJfUEeXUi8
jwcl3Hc2ZDFPWcTQ/xCA9dRXFAYiAxar9LDNeaspTS6FO8AhuaSib9gGRNDQgABqGYxofnOezuk6
DCJuy/vZCsuf3CdhV84zAMY90dHxC9NzR6ft0AImTpPbIMs/rH1IckuLSpKSwg/Etw4DhMectdz9
wSy/bYgVnFSGSSlgiUf8N0oxd45ghCxXkcOjiVPTqS4jpe/Qedo4SukJvUM3Y1e7Qk1LT6j2wVbu
CsfxIR6Xp2ZFK0SzSx9xiqIprz6/4sdYsVTaKVC0odRL6kpHZCDiWF9RYVlt3f7NDrqGNCBHZD/z
fwQVqmum5PkL5QDYPPrrJiPQBDY5fWHP9X69y680UxI5ygGPAX55oHN5u5IWOybAxLkpkScZQV6U
ggEz8zddIgywCoxo/SCgZggh/8/vVyHnsjRZeJV6iT5ml5xWCW3JAbonosTGpL0b7bldPAa1kUnc
vklLh6kUVKTJORCK/vgsaVZMX/QY/+ZVkOkUOp9Vwv7FkCnILLdbXcpOLhIuJZ5ZLBAb90UTsWzF
2vgPq592JC81Jq/7PmvpUbxmugYeBk5X0Rbjp+dsXXRf+J6GFPtOm9OkDHEU4Z0XhoRcalWsTJb8
QkNN21iDvrXm8B5T4peYn4Jw7b8PpCFKGEfC6i3PWshF4KC6XS+uZ2DK4hWzw+5S+HsAuSs5M/fx
klbKU4Zm50DaSiEPOnTrzleqECKYl04PDwa8/rOK5FlieJePORQx8clevoW2F2nKeSb6QVMfz1YF
Xuecqe6flH0mdptGOBdPhoskYDpDfAZZmoXv2iyK5CINc4LCrvXu8FhWKFdFb34Khzxw0tk9QQ9i
ni78a2CASOerOah0GZjVNh5jb+9eGxxScNXS9u+vI9uWpPMXz1UI3o4j5ZvpVXkjRpmLPU1hAe1C
d4jkcNVyQGx4+CWn66O5BzlG+Fxgztpq4gTMOmB4/GLfGIInAmFD5kqIn8WhWchV0k2xX7AdYXJn
XZ3aI9qCjPV90U/WvpXnU2OG8UNSD9/f/PJ0O+ZcBymA5Q7VpcAbs9dPzPtUYuBtpeLm/mqtAgD3
BLFmaT0wfrDVWnZ/dtzMhSlBU46QsMxmStcu5/QeYuQBMyCDarFIzI7V9O/CqduFQ+bO8RR+8rco
kWcAObaED1UY8geJx3UG6Lj6aSSaxZv9V2ox3QbsyfGNWB6g3OSgzgnG1Q3FLCM36jgJ8W6uiDKv
7OHUOLvFcOFb+tzh74sYxbRziWZ8ZSYPEAFRKYkskfFy7APB/jh9o0O1PQuYJhLrek/OcsTcot1C
rS1Bu6Mkcl3DJhBd53hNBnsXdSKm1M3NmYvbwMsKE+O46qyJ+BTrFutAJeYoBvHDUwEoh/TaK9cp
6vsIIdPPhdJyIryver/+P0KqWpJTRClHrv4EgBlPCoO5vX1WGJm7xkroGNEvqrZxL2Am9HxiNX6Z
Jg84nY6SYfHmt8xvRIF+TN2gAkkA66gIKeY484YiOh4Vvwrjwf4wldlgkXCzKXXdcEv8kIqPdJ9Q
yQJ/Bjh7ujySOLyHYd5Ho0RUzi99Tx41+MHx/R+lJLKWv9h9uDJeqGQb0o9lEmw3AgeCaWKbzXis
X5423+7NIFJX+xdFMkoByvJTK1QlU3MNuoyvEP2LTdhpjFR+rWbALZOh8OF3UjZbhrbggcsaudoW
VEOfy9vHjRc5EFNe69ol8Q6oCRD8+WhujiFXBAIs8b/nmv7cDR7ogXfB05f5cwtjNOh8udoUJH9H
wunP7J0Me/E/dgKwvqsJ3BG1ewd306dwfWR8Yupw6gDQuY1DP9/V+pxnz4vbDVgxeRIiGKJS6IuR
3sGhxqu7pUW5m2SQFGGhrX6ZrRrn7QZrifWmLZOVqhyR5vsvUZjHzijsn1LlSExmLwR1Rs5RB/K4
Oz+tQg9ezTKSDTmTpOYEjG/RpV9IQqV08Hv+vMK9IkTBGKTdCqG5OgXsDlfyt9ztalBtE/lw5jjT
or/kABmfM4eM1fy7Sjk72DnuJTTK8P2T4v6mSwK0W/1g9X7jBNhquqLDSYOqJ8mHAgQvmxr7uOyL
BJNFkFmekNbmq24zt4D22G6JTFfhS2gBCbycDifm92shGNvaVeZ0rT4/xpkBN79SaP5vKML+bc0h
XJ8FjnwIHeJ6ia8USLU5BUNKG3OHekDOO7wVlcydmzFGVbmvXVqvEZwj+aqSHRVgCb7So2MsQLtR
rlfrVW1zHjOv3kWF+2BVEk10wl4ccxxwAgJwt4pEinndnuMVFux67aUiHwxnkgmu+Eln5f3KnnHO
6NiESa6/l9jK1V7NLWt3534Ecd8n3qhFgHRk4iN/NHm9/ophBPgnEBtq3gncePsSCRHHFLcyfRDa
0LkTKW1Hn3WYVlaW6Qj7vV87eRM1Gzkq3DfN4eROP6x134iizMt3QfkpKSlGluY4Ph7vnc9AoR3X
1rwAbq+q2aJjH/usiNKv7X+uMdEN9pBvBW466bDzdeMv/iU3dvfWt864z3yZhulzvetqhXTQ1f8f
MPoF5YcOw+4HX5Od9dXrNv3PrSQYWi24vaRK11FKhDr9xvVppfYJvwKgdk2GPjEoaoL7cbeFTYkx
YpHsUmNgVh3dY9E2B/KTpD23g860iqVBjy6rcT2ILtJhCLa75jRKozjfhe4KMvVqxDl3eaSoGxJp
qwB9Ew4JfkBsB8WSoCMakQaPec/2PFS7JnLY7n3z5n3Uhecqn8prEAOTlo9QMVBPl3m8hp7OtwgM
6bHqOxEs0aDmpYeBGqwNrd2QUx6HQ/XUr5Ofpp5tQAz7w80zMslljvdojJ2sEByUgdh/YVKXyMkn
X/6tL/t5IvyMFmrsZPSAvd25HJTrsuc6S0hLei3auZ4/T6LIyEnCIzWXEX6fvXbnrJCMqWA2eEZ+
fQGPBQGSHXKM1H8unrSyUa8HmCYv0ftmJd2w0a6gUY3z4pvHrM4BS9IYc5ftIDvK0xCsg+tMholc
Oz+5e+Rydv/uY308J8xzOU1ir6UkemzkqMCAjishbRm/B5kWELmAwub/DxLw/211p7Dj2zO9vdm4
9xKjBpmYzXkzhQGkEDBu5HEcbIpo7Xjo42MJ2K/ch79z9msxYt5P3C2WolKfwivUd5b3qAMqxWif
FCUZHfVHQzyroTkz6hXPPfAbXy3hNGC7Pjuzl8MPEXiqel1Twl36Gp0lF9dEIqOL2SUWtN0+QYTm
X2mGR1c4kuvdvBL08Fl+mXwOAa18PVx8HOB7lrb2XD1ZzBqlNIb7/xemwLnItoTnDrzmkjfRNRsv
xj4CMdnYacmITwYJrZUVRxBlWAcbxeSeGU2/psKWb2A6bl0VBboPjcVvZtw13jtdpax8peo7vuW0
eKOIY2DeXVYPRnClDlIR934xQty0383QcznQPE8wsL8Hk7d6KGsVwFn6j83e0YTKMCNp0rBBAMTe
33FjpTn20Y8w9X6kKEY0gh0TxZmDaCOglkWigZhvG+AbCM12ryUAuN1bQs3n9WwqGot6kwLirB3X
ClOCF8CZKRHAkX8SfVhwrOFVt5DxLvER27ooPza+xsDNZS3er1uiMLTxFxqrvL25l5ON7s7jkxKb
Q8Yv6ypOoQtzTeJ1ut6p4zBEB97ZQBdZeFEch9IU3Qxlr/7rap5B7VopuqRVEf7Q4l0bkN2Rrk0b
B+Nwa5hj2h7lc3vYLu9WwnQ67SIf6THSMg2nuOir65Ue9u/oBFwsYKAcYgo+4Aq7l9jLADI+7N6R
X6uaHi3hHNXaTGOg11m8+6F6UiPGSxnT7d3atkYrNKAHfXUgz0bxOMNQoPGSiUjWoLsu+et0K/K/
qCnOmkqPmocWdr0/zm8TJS1CLLd/UU/hv5ZXzW9toeX5BuLDO8cP3uVYp3RR0CHDXB9AD8x0BEMJ
2+3hxS1fa4UOv55AXuAUCU7eRKDQc82QeE7hPY/LwjmAonvg1bMbfkFqdwFZlP/pPXASGO8t2AqO
YKQNY199MAuylWyiXvKs5KSJAGXv/fWM4yukY3XBTg0KL+hEYWqayybrqReJyk+lD+GeEeGuHKsB
qr0RGl8e8KefWXAlVwQgDpCkAxJ0O2MWgfPyXO1FxmFQepJhn8RV+r8a2QodW96plpGu5/iadRmz
j4V32eehFm2861RldccywrJv7Ei5g8PUCx8+0pwWsqYeBYB6KYj8i4EAfpCvDQEZteaCZ/wdTQ9F
oyDuAq1biUCGAPQHZG4z2JqhunIlR+bTg0wMOu44U9XsWuMloK8/uXKqYTJ3QTpZpEovm2WiiIRF
3VsiiXD+E99WF1CD1O/5l57TYOsASCVp8skSHnKXe3VL9tfwgOwNuoIjTzIAD0sB4bXpbp9tLEGE
VQkENQM7IQC19eoaXJ+Ug52sallwIYReyPVANwozsNan/RmgZMPLzcXVOl0rdP+9o4ufmMN4eZVH
QMzL3D6GjOOBpywhQdS9fU9NFHqU5fU9BszZDaCtv6eKm8UvJf6D5fLNOy0nO5E6ahJP4W6HopTP
QvAy/smGpu5pgFbZVtZj+UN2ThMnZxIX7TnsORtXD0nnm31PBwjGDg/Miqkx8ROFlpW1OIid7z8x
ppFPCC4VQaMaKqucHEhN6qinBvF6SYJLWyXiyIsmUwjns/V22IVLXWdaAs5PE2iDBUZQbnSxFpsK
Map3bKRYlTkZwfN/fR5fZ+nDo3rhIoRBsgl2d53C7uiSp4ecx6Y4VJ5Qq5yRtQfl4veUg4bQfdvc
H0jhC1opNmA9hni6CvWx8M02CbCgwbYZvefuw9KXrZ5kkPOFKLSPpLBeI6MPxJyk2BA2JdPKm4AM
ZkIN2iRSyGQ/6n1EJTQk+2Iyf2bDHxva/n9gReOaYCNOMXnIhsbYV2xMhFAsNc0SM3k6Hf3hh+QI
D0ZBglU4lYxNpiTyv8fPnpthRvAItn+dU4luUluDpdnkM7fsFQlwlOhkseQqNfY3bfbFVIDtuk+L
2+y6tFOUkKT3JdosSGwVH/52J5boO9rEEhYklKLW7R0P6WhrFlGrRyKYMxCx6KgIZCvPJA8pR5wo
Hlazn3IVwCmPVQNGjKi+1xfWEUp1Sxy7DcCwl/u4qxvljf0fFibSkKTt3I3JuEpu1XlDTaApXBLR
+nMhCc8gkm3Sdin+E96tOSl1hAwroWbwgr27lqYxBM67nNexge6sx0t419JNxncyuXa5v1VguiVC
L1s2kNId3yoGWnWA4YlmCcgZB/vh94OdYdP7Z/MIeZR9RnJYYWbJOP8x391eGjGY77BHSQUFa4dJ
OW0z+ZN67Lnpb4qTwlLNCoXK/CAP2tUJmRrPUC6cLEAyvtuJd4B33DwPH8GHVBeswGLnSN1D3Wpx
p1jIa9KW6KpJND2noZEKEUyHFXCzLD9gDz/bQ9knlPEEWFQYa+qCThp+zLq2Vsq8ubDZAWs7jdeL
Ll8lSqVFA7WMWuvJbZ/vvuHlAK4udmeu0+mcZYvR/Skreu/GHnhexpBjxhpG9ZH0nv8AiZ4a5Ran
1A7MwgiRnd5Ntvcx5pghrTE8gXkfiGA5hhbGtT2D1Q6VdOcsnC9qctp/xXS3z23cMGqaQcCkfDpN
M/kocLzD/nAmNfdO91UwOBxK06C9qpKHCxaSln3ewlCDrGYfXGG3aZIxO+dmnf3vqHi/dWsj+dPU
NQoWtCqXJvF3SGeLF61ClwLU8l8gjP94bC6GVObg+9aXSNAeGoBqe3qvY3abaxLMURuSrnLrdsiA
AxJzF/zrPupNPvcC1qcyehpaqN/2wI57Z1NEwT3iPEOR7no0BR2QdSokWn19naEhvaQqq0Y26+jt
fva+pvv4s3PUqi4QytMtVtnn97k7RjNu/TvB8kecX9trNWCQGPO4KSkhFPBKBpw5CrIDa7ud+bcS
3eXTuJPhfeSVuRv2I4QFCPYPuk1cNQh4ldAfYf5gEZfNIImD+lazdxrh1fD22P92NrwYw9yfG8Bf
95iEtBhtfPyVQMDXT0ie0oreqDQRciEvwWykmVegpjclWntXCllvHyw2/s9iFApJKlmUot+Yuw9M
F4WjBnY2wBAc/TGx+BAipXXdVo0z4+PJQHOBFaH3gaEnIRbD2+oga82Pl5ptc1L50JFZcmL2ZYBQ
kVIamB5NFd08Gdp9wm2sJrvLyCWxcHY3DJ9OtnIbsaiqCJjGJT3vfBsIlTAD9W3nBu10YS94PpuE
EesP8JE9Gdhk8YE5lMZlU7hqf+OKTGe4wiTVmmm4KWhxQroYHK7LHWRGGj8z4S5wEOl2ey3w/7GX
mqwIdNjANaxxEjXZ3H+t5JkysKY9ju9dDsWst2U5Na/yLInffzFE2ZTe8lAHjL/cgEqTO4G8IBGg
9j35Ji2oPnC08Q6icidxjB6WLsPqIKCGRoEbphF2DQC9VXXPxqKkdLgloDxQ3TzCS+IsO00axyYU
pLJY33bow//4FEP3+TNNA1DZ9kQDLp3qJkrGu2dZCQodRiC5VhPyHxs0qfuiPw0DDPK0AjAScIZh
wCZV8S7ucSe4Dx+89dMXlU2gHizeWwYGThzY4dl8Y8e1Cef1GZO8o0vEg7KfvG0jQUUVUWFe6jEJ
ezuwixsT0OQh1MRkDmnPaWkfLlWPoGDcIS2OXwoNuGXzJUd4OodasHvA3383LuRdd+kGUnR6yF0y
tGHRKJaQPOJo9XDmD2BIM+UBcVnPVyd91PBEXbXomYdOEsAd1gG/V2FSCwiFVf4UdwQdTlBN7Mrc
7ey5M72oU70/X5Z9w1Sk4lBPs9nQ2Le08ZETiJ0niim+TeEaxFsT8qnSjoDO2jSa1vTSClr66WnD
K1oOYUMD758vZyT+xdwDHCIWn1GRlN+S44ZsUjw0Fff1hzm2TpION+Xxx8+BSFMaL68Gu+MUxRrz
TK/kNVo0TkeBBdGpVYU2dJLtriuk65q4QMcW7Qz2xynraabgkIyR/7adD1bPwR1ZcCB/7HYKelri
IHXVlpeP9Eh4bbJ9n0gqZuvojkKVQE2ti93416e+ujQ+ym+kZftjX6nTyHE1C79jE3rK3KMqjnS4
nWenpMqL9CEKZGgW0rhYsvfGAmCNRoDNZyv3CrU1/e32ey8p79OvlmqPNPb7rIQHFbRGfOofzBhi
BbR9U6RnL0Fm7qecNT6eF/qz+Vzo9FDYbSgNYSId0zI05sU/NkQYvj01wK84q9pYLkjPwcAfJ3Sb
3udlDY2P/7S/qzhUoLKcO2wDS3/yV+658IPyumEbp/yh4CwqYgabmC+fyeqAiBk8PbJAwVgRKrLw
2QctyGmAKelSLcpZLw+UuhfEA9YpOw0cVt2mz7GuLzygrgBaFlIuvk785NinQAyyNeEG7171iYEI
ek/RIZTxR0yS1WnNne2z2Df6IyGXisrm1MI9wNFVf+8dxHkw6k4Ap88nAGF8Mw5CBtn7ceFelUcc
gL8CYG6+vacbLp6a1U8gFE2h9ZMfIS/+Hd32aeVBk/ELpr9v0IGb0/Be30BoUd6XgrCof1jztuVl
8gaQQcmBwmfXZLO1BieCjfsbUzuW2D/ycooplc1i0XSYFJoRg3IDu6ugVikIpU6CEXujZzddvOnv
TlKbLPgMD/i2wkwrfagalQ7oCAtMXzEEMtXflSy+LGyEEnl31IRcznhOuRgYUSxfFyzs2/M6HtrU
NaJ0GSvQg6xn/RVXPQSlIO2LpaAmccu6SZVDnCu5YCCApTQnXSWfKbMHBQxvIZWpZxk9scDvliil
+HeJH8L8GSWDZt7rrC9z8bgGhGjURZH9RClLSNHi5uPJXJNapCHuc9E9BHm05CsC9OG6s03b/KCt
eHSQd0ZexixZTsfveNIH9zdgGmo81YhGBEHafyOHtF4ELozr4IEiRPoucCKSF5XfmjSz4JDuPGBY
PR0/K1xkhzpbK2j44uLsUqXysfjW/2+qTMqzS/wWpqItOI7eD9OeVpCdQ3mv6ncHZ+8lej2T/mVu
a8hRqbaFCEk0NFz6/dIdabBsIaQzz67IwuIWcJOtVfsYQ+BjUZE1fEd48hJ9D6FELCWzZuCJwTRG
TTVauG3adxymXayKAOtTB+t3F42kzLjAKkhEWIZPFdU/M1aoufNyB5ObGSId5nc1lwKKHCkLZyog
Zzo7MZqx3ZRxut/UIK/dAlu7TfK4zgzh6NrgzfEabFx2tzEJ3TpmT8mGnn0agQtLbpRHVnumSUBe
0daApTlkSsv2DQ4DAN/Z1q6HxS4clnUwsWhMxC8fPqQCUHtYKyRYlFldOMo0TfmmEz7Mg1+gPmC5
smuNRAsJsgd/XotbFtb2VLtcO+MhgR4RiFrQbWuwg9KwV3XxFeQbTMiFOMKbT/YRG22qDP5zEYJV
tOx9CeVAaXnyeUs39IXTjamqqENqRAxQtmjkJ/e+DSu5HOYn9reLzk0x4ujHLxTN7+UjjWEaqxlT
bLKNdKDpZeEmQPd+xmz1/Qimc7jy1Rpds2hFTJi8nAmctjkd7pZFl4Pzpgl8E5cYtUtHlkCzA6zv
YASimAnUa94nXkcVFjts6NXlS3NpJZH/aZmW7Zf6blAVNMoVRRf5BpFtaChrucZVmr3N1Ny3YcgW
wOC1sNwsGB07B6+Iq/qGMpvJ9QffAKbSSX3kTWVds631KXAFyLDDtupp/XCCiB2jSwRYkmMO86Dk
dF74Y/DhZxe5J0+U4HvwdJraxGYg8EVrI7jq9Jhii2CeXXTHyCzs9k7RLkF49E/N6SzcYSX2QEUc
M6b6cgKbVRVhBAeu+eM5ZOwMPFF8yz+AE8epk73rzsiunnkZS5l6e0We8Mi/ULYHTM1/jmBjjPJS
79XDDpsmYtHClGp9Egl0dKIvcb36xHwSKOuMLNesZDPgpnl/681L/3dQsagdnY0T8VJ4BqxMP9Cl
ppaGuyy25L2gPq5Cbd077NW/nV7YHNQKeJPmqIWdjqDH5FUWitx9SolsPmY/cs4vzNYY1vSzZel+
fkxGYcjSGiflyKlYps/ZmjSOZj2s4+0yfPTj0G9mSmFYojP99z9hi7nAMbWPdTF4TKvFDVm8ZobY
cSS52PSFWvxxQJ8oYYOZhPflMn3OxnhkvsMgEZaffcYupfRtPhQNBwCrIY9DCdW/4wslo9HoHWzP
ikG/bJ2/M+/xYGvvJpktMOh3O3kzPxXg5sN1+POxXjr/WTjpqLUJflzjtjBMBCxkSWErPeg3hAMu
YoPmknXowWRHcHWaxZ6/agpmTMrJ1r0oWqs4fLTpNzUDtxHtZynd5GyG4RJoYnSNO9yYaukAMxVj
XpSv23zriiiG3/8a1uxxGcx+cydVA48IAD9c02OnFPbCOFO9Kuci/HgunFneFatSsj8Da9NuFdrE
wEn9wEOQtMEVVPK/OWJABJIBsGoPJuNzWSocYvYaJiPznr8/u5mrYIWLz4Fvb+4MXElfKILbpYux
Dtbx5VLOLbwxUCHuqUgArVpN820KznbQZcDLvRNpBA9L6wxmZbE4SRDl7R2msvXsuOkqU0dvWcAt
XM840KcZi1adyLVxvZVYW4ZVmAuADMOJNlx4XrsJym6aAl9XNXofIbzyIh38xikuy6MR3MJf8dsq
NQYFq+GfTYAe/ScE+qIH2UB+Y6ZVdAsgzVQbW9SE/6R0f0fOUZLKehdNpwhR/sFLMqn3KaCC26r3
e66XLKVRoU/V60AIsLXRAhqvxDzT5kK2DbIop8AfU9DtmY1ndU2I+gu3ysYFEuj4SfPg/g70ZxrM
rsYVcm5nm5pi7A/6jAaITMmAbCsXgJV23O/bdjPQ0P9PBYvkRqnEybn+/57bSyp0uPoLsM7IWPS6
eBryO/vgILZCEfX72K5pTz+Nnyh5A0f5TtH2RGDyJIVf0TnPl02/XQuNF1U/VpPPu6ew0oV/Jve1
4yRJ2gHNjcy9rtwr0cg4H8dG96W2MmSXbZ5JCMUPDHOHS1Ij7ZXUwSD58LBzIzTpEpGkM303NAyr
fCz6vrYgR54hV1/FFbvwoPCAN/72dqRMl4cRycRI/WJO7aoy2ayVNLuPOQOsn87PMgwVMpN1ugze
b792FkoHvRo2h08SItEIsdivsDsi5k+wOaYMeh2eCj2NKLBD/ltPSsKTjawhlOkUkka+aW4ZKtns
yYxTGr+xAE4+jcBW8AEaxE9227v4TNDAHir4P+5Lo/6+zav4UVhZOH4oVq9bDVRI2hQliMfkJ5eC
SduSwIxuIhtagQNfobd23KGrz6SVG3clMHdt6QSRnAMn6n5Mwa4NDirgWtIlz/cH+1/Lz+OuYI2P
6U3yVp8tfKXTTcuIaVipwJzNGQ9P+o2KduwQsLBppWLR7xYn75qjD2KSmblwpcD0wgcghxqZ3zlJ
XnrokqfkTiKrG6feVLlvncEsbmmXy0ivKX58Gv9nME1/XqOq10rr7yMd3R89irRLXZRYH4N6myRI
mwFmS+W3xpjWEcX78nuY+6A0v+y4anZMN+83/gcJ6wwxHEHnt5ZXTZiLZijyzMxNvCUWPv/UwVzK
zM81IkV/Z4XULuw6D78cznwSxC2uhkxoTcEG25LtH37FSAnTlJ5Prn8EKGM9dIwjGZINA+zH8ikk
EmUBB1OEjMGUm6Tdkm4+/2ifcySl9cYnFQdNSwuKE/+KFuBNbJhPTquKRblXuFV5NcjV3UMMNlVE
r+UFfTlM0t71+SQFn4o4Z1ccp1WxcNwJsrp21fGNsQV6KFA3PwtDRIGns2/Ylc/QnOdpr2VJtINb
GzQz3AhogZsHhaOIRVJFzf4dj4rMGqDrtpIcewxMC0hKeR5SypuxULv1cGKUJA5+8mYopOmtMom3
mwCguoTare+YHJMxGSRFMXk8fRFKn3wf5c+cxhHvWZq7ySOR+lm4sNcMtWV7udS39FqH/BIQsK2T
nStgo+mzrfrADOWPzCkEgHNIZdYa4Wsk9Pg8yJnlJKUmgFICvL+y9Jl64XcPQhvPBq53reS50FaT
wUsMGjQx8w3jOEPYj5BRtGwpCTZ3mXXbGp1Z2xtvPNr3qLBifBkOD9FtXWka1VbndliVgKZwD9Sf
SNRg7eFl/8YFRdv0zPw3g5x5zG0Au/VDAiW6veAVdj3qIS5NWcy/ilIb/rj2aCM1fDfyjZg2c/Fz
jbzl0FwqN+Pb/vwWeT0xBffNRxRmFRY+gfPM/h3cYKwIZCZJ2vZv6++OigU1FcFXV3O0wEUA8KDr
5GmWj4hwGBotTYaw8VCLxWudqBCHuRwME1xG1Smv/DcswDHBMfrCqd8lnPijZsVT6t05BYZXlOF6
HpmKJmKWm+la4Dd3MGr58PL6acK531qY4BVbSPvfygb/s52Fyx2ba04cp4Gsmg7E1sLl+6l0bmkg
E1k8ZhAUbJ4UqlW97PrDAjmvGyVtBrTCrK886U7j6b8ylbXErRNn0y1N9vwquVf8COXlL4ZrIISO
Cxi89OFDH8cykhuoVYvnTmS93ulOeSh4nf92MPRGVRmSqEjpwVZ6BASR25qzAGDPI3y5OKVw7cR8
qNZi1MZ5lpnUonwwUrADUnzOOuWbf+0GkXAYjZ6DrD38+dHQ/2Lmm1D9AsawDtTpzyYrhw4+a/Gz
aYuPhTOZwR/Hzjj09gQ0Ordvhn+/9L0qGn/rydz7J90v5Z6GR1oT1S3UYKsvx5HL+arf6WBjPZCV
EFvVE0oZJACM9Mi7OF1SAQqLVQHI7K4JIBfH6y0mKwGlst1aPjgXJ3PK/eF7DoiAvqq+NscvyXlh
V7MZjn5sUW/dQPKGfTSMijxWlvkK8Ezft/4OgyR8cwMXocjhTUGVcWHPuWKiWN7zkvMJYeVuYeel
IvH3DRiN/wsPtmDQtKlXMXvmaGa3QGe4+jq8HaCMGD7+W0zVcCuEA369aK0Zw6Hv4AHKitgCLnRS
Fao3MuEhiiQV2XKagPG8K7ujuGeXPoRuAT7sBuJu44V79RL9L8vysdE/FsE6HsQAWCwimhUgA1+g
dr09QYPou9o/VXya9VwfOcjKwT1cUm54bp59oZUISVDoxQsZYAs+dzLmgbd4VFpP5G6kV/f9+htW
mlzYEaWDD6dYfu4upyTAuyP17xMhu5ObcTQS7d/qmiiXSYTCyfUVfCc6Js7bYZfrDg/awVTjN/vV
+tjrLt308zFNQ2lkgDu+FPJp/dFlXkSXw7F3RdBtt1h5lkkkt1cAnjaD1apdYXsfIOi4VTo7PX5o
eublMEKe/TFAomd1WjYCH9g/794sYl3KTvHmymCbpotzPzJl8Uv1Yu/co0lWcuqkghTxvsEOcFg3
nX6zEs86O5MEMrLw//XAUWQ0bfWbUozU1qtgudp275Ef1J4jEpHFe7hjCvG1rliDYAD7oymt7P6n
BFVz2HOaBVsjXjp3JB5eC5VKmol0QYnmKwelJAeMOAGAxV3oes91a2qo9/jvqpAWup4HBFjMirZm
5EW3I2dDeu15dn1YAuUsnvkc16ngRhSCmOrdVth2w3yE0TaxfMQGPl9OMGRLT4fLEhdytRXLYoaX
uULkLIb3WlBiVxR7jpLlP64C1g1HUQKLU8I0fbEH6Qh7T69gm5wG1YX+VK0KkMMt9zkknr2PEQwi
l4He2paf3fwaqxvuKB74OOTDlKNt2MtzA41zXtXT5cQqybBax7CruAJ2VFcU5K98cHNSoDD1HMjY
da7tAqLcxdrZTuZ5DNVSUM6hAECZ5ugbgfQeRLG7rq/SllM8uSPJYiBb5N25nh/76BJ7rO2HuwMX
SbQcL0p+TuN/YFSma5PBogpTDoA7wEm8E/Chzemf0S4VhYGbDlXhBcc4w8Mou4ayPCGXXo0kP835
CeWNNdkFiY8TbibFhlprZjhD/4j0gt1ojGiOoLID6lTz/rOGcMtPSvRcuPCHN0ux9/CMvjbajepm
MUQ0o0diOtRm5IfrKCBqHu92uHfMj6vG+Thug/gjupJJcoQQYWJipEk2ZeOCvHAhlPXXpQCWcSJh
Yhm4q9DMZ9OdO/cA4hEtcX378yeQa/Sz5H0pakq1bwfunUw2OzemJ7lCiSaNFNrj9j4KgYPWENuV
CX1c6UjTh4Kwk67r0HSpr6xAAyJU7WlwSazjVyirwRDeMfDJkWf6H9Y/lo6P2onQPxAzL+AKR0++
fwVLOIiCYUcg6T5nu/6oXQafhtMRKa0ffm4nKhVXmJ82i9B3gWHd+XmlRjrL5f25GSZSGbMrWBem
3z38ABb0kYE/pb+eOb4wgvIAy2T3g85RheMCW6CnWXWzQyPMHc5kvBjycpt45sk+CEasMkfQZgfN
O6iCDpQBEBVBHW9XRjGyjjaG4iGXyGJje1J3FsM7+lvSVUJIK2m5+bBnj0BXNlN5aM+OdsbzshUv
tgyLpx7eQTidhicN3fz+y1SMMRVycC8Oze5v8dN1pw8j6dvIYoUrUmMk3EdwaScssNtuLVDY6SIH
h3efQz5GsRIvhF3eb1vHcdHNfcrsNfx5e+2g+3psTVD/FYeNJyOM1kS714Bu6KKdBQAnmEDJjgR3
AGeCT3hTWVX710W/iygFoLi2uadrwkdn/5zT6tvCmtD5cGr0U8Fy9VL0i9sgNQ6SP+M3yIiqCjMh
oN/wTK7+AOMQP6D5YEs+J4m5EIsRGXXfdbxkXAiz3jtrxeUUl/5yvgnRvnwYy6ilQhb1Sfo7Yn5j
2aVaiOXhREuhoVx2q1Jl3hjvVjQP3k3ihwTiLrt2oG2lcmOlWGFuHKl8rjpNBy82+eXaToMlgScb
7vPG9IJzRHHSyn7f0duuwdpEdwfeCZNP/YdYzUPuqXeVrDBcNVRq82CPprLcBhofzFKNmEPxrOzh
RAAsQecrCxZ0A8Yr4TzO76r3vZ7vPno5EBRzUIPH0Rd1/Bkr/egl4UuBB9IId4m6Pp8IEo6tl1zB
UC5zHjfEwlN/vAlXty6GoyCNZiSZe0K8S2no03p73WT6musFi8Lr+Uyj/CoSJ0Gnq8UdH2jed3Eq
JkUut8KBwnAKb4wrKHdQnRg9/dyHG9clZyzViKfUGIpGeUhr6ZP9AQnimI4vxtyEAvFGKzxfhSfD
hVBLyNLLFrzR3Z1X7MHypojUnEbxObW0h75d4HK3gpZj0czVXllyysqXasCu3/5XtTXqDXgvIpEK
RODDI+3RTc1faVzZeYVrInbpKakcHmsvi0QttVW1iL+njU4EGuHaV73ifXpoDLQ12pWKiM4oZ7Pv
EDt4jgN/ZPbdEKMT9N7mNOz963hyxPzkEQRA9/OBQ/l8T48j08zNbNR73NmON9FweiW+3rV2AlZt
SSE9zOZRWR8/7fVeWrfFPtuCxPgQE51uxWLzyOxlcTeFlDodw4x5/EgJATlv73Q0aGK6u2oFJ7ma
rzBCjBeBvASLFfVHyGabPc/aNZ3RVBlFYAhfxUSkuyH4R2YcxrOx4/5OSSzbd++0PURRnaPsrEzM
6Si9ZxV7R2bzRWzR/CYxuiO4+vwuo3VHrlC3VIFCHKv4Vv3q4aQtpCkzlGFtHwU4jf/MLEBnuO2W
l82lJscSEsq4/anttHUh9zHiCDhO/RFIJ04Rtd+EDFVshXLPxG5B3cvw0pBryz4ALYToIP1S191B
nBZLs/fUV8QYftN3/7S4rTASFC+wBrfluMK2Bl3zrSKFTbm47Vw8RcG22Dlf1pTE5eWZuP69cK9f
tXkpLPqmGWKA0kXj4aPV6UwXtyXFxT/xhZzgW/vrljr2/MMT6T+P4nX40Nc7D9vpN92W3w2r17JM
ZktkpI5uB1ZFLwQKG64WiE9mvsOCqTIKPiyYbkS0ursx01b/g4m9AQ1iMam2VFkyeiadS8IGpfS2
+yOSsXrYgduWV0HOTCn8PonfbFf+E5r+616n9fL01c8c3lZ7rqP2ayulDsNB9sCYEp3YAulftnEH
r0xW0IkWpq0KTzoyaVYU01d7z8oAPXP55/fAkl0wK47pbjrh5ePcO1umhQtS9JgXpJIQqoBJnm18
yaVPc7T/8Wye5LebQafnsE/qZSXoXoN2y6wTacHwkLH7dL+hz/xQ4Sy71/Qg+Ag5dojYkiK0xHvS
OE4hDHVkPrZ0aNu3zbyFxzpi9QOpA40K1ZeGYt8fkaji2O4OmOZ0eKoFFWQqgWjt3Qqg/65Ugoq6
F5vOwR+MFWDvRr339kHgyfO4ybQfE8YNABmPSrC7fkXJFLIGrsBzkK4OoqCwqvkStXVVOZ1vpJC5
yz8VSFPg6OsUT3FMoOlprg90yuZk87GgqzKGr2VBmNBSkvxlbCbF69XPEO5OWT8exZ9Tt7L8NBug
leGsN0ojdKn3VlvGHgW5E7keeuju+JPGvs8ARqnXgr1ViUDKPObAF0NEGtQqH5Hn3qQF1//Vxe0M
FjNClXe5p3Dp5HIhUo5jpVCWZpIF1++I75Z90qEqfhhzwzBLc+wgndMqFw00JeT8kAUk4u3iZ0Dj
YxURCQBYYLB9jmtdvE/ioblFm2407K8t7mV0H+OGqw2b0R4rNElMTJbtrpre7AFX3KpOFLBPWl88
UA0VP7aRmSS90Wtqvr1MZdmV1enLns9/eXppmR5g2xukr4+mp8YlmjEepi48/h1rXRqG1keWtR6G
8s+vdE7FHrhRxBMrKCkebi1x6zY+zyMpwvAMmJJQKjXD41Wa6aAvwRPPPCSmBzRHDEf+A/OgxZR1
uTRQFMhhzBWdhs1T0lk7d7zov4aHNlqiJa4RIYOhxT/7nqgAj2Qj6gdOwtLmdxQvB9ZSCMMPeGI6
PBoc1KexKnqoQGbQ4L+g5506sarCwfsDYz1MaUypM4Rko7305wPuAkD1PH7Jx931FH9uphxOSMDe
OE+Qwf0QoNQAJxVMO4yKNSpdUZwtegV5lf4cMl2Qrcgoxv29Zxd3MjK1/FgKYwLpFt2sx+QqEegF
m78bcnTNlVIA6ChVh52yMyGC7Y83SU4NRzr7ymsEKRr20NDPukRyFMxKqguJxJDD8bCR90COEb+J
aSOpqhsRzUCF5Siu7PI96XXcZ05YXGcVkSCX/l3N7cS3auqDxo0ZLE7P3ZTiUuAzBAH0CZAXk/L5
yJQV61I+YYK4uYqm6MXe0QpncbJ4LdKMexNVyE+U2sC5R/3BmQWZmniCP6NGTawzY1lt/vHddA7v
dQ4QuW7cVhgV2yxASE64MRx8a+LBpAqdtem+KMn9KdjgVIsSGvQr3W9Doo2WYF8MonXb0gHdQ0s2
FiVPvd3BNX+3SonSI6UhB5fk/+Fq2ZDWYgBRH7RfCqe4rRB++JrSA6O4isNMLU63O3FCxMKz0yqu
YZJG/xbksMx93iV2Jnv8VK0f2GnMVlUauudqWMUjo0xFhxGRzOQDRnyrqMVSQLyELEPTnw7Mb7Uq
TXY4TshOJuWruIS1xcQxRQ4Pcb0l3uVJlJ0jD5I04vzzYDOYw/ABECT4ypURHgMQtzQCxppAIvr/
Tr6OYB8X+KuoUGFC0cQIHRttuiJGGR4Ji3w8sRFjfPctROnTcZZroyOtCqDwOWbeFfo5WWknYEGQ
lesAhvXWN5Y5IAwQhundVvcgppKKeav5zrh3QisLGSwaBbtTWmGIW+CA/eA8OwFg+1VB97mWUBQl
SaU35p2cYzzWA9AQsqM4xn4fTGNijIAIe/s3vkS+1DzNbsdB8B4lRIIY/X+7GnIhc8vnjCfWt5tv
nn0ujMfzjOTsl7tMaOVTUY8jo5wfqHeLXe44VIGRqL4+xO1DFhlRWcwGO/DS+sgxTsS5w1oNGyqK
WfIrM7z0mmSK0ILu89XKf5D2O6yHIiUS2cT2g/GwQpEQmRDhA9Bk8bLMUhkFAxGRO/7V/MfdAmX/
hsABr5/W//MRS+G8PELQB/1RIB5RwENQ2mG8PTggZ7c2VhuMsspmmiUFMSgS2vnBOGX/kg3iQeef
dn8qr02n2bYSHNMAPe7Y6oh3IF15al3YnMfkHH0sb5UsLJS4iqEdJQx8Hfkl/YjFFkkYvSoQAaNy
vKOwwmSj8Fq4Zl9SPy3aSg2q2HY+j8wwblabk/aByBAhiEfjX76bUIZ568CCETzZzaFu05lBRGII
JBd25rGizUMVZzMVthb+uNX7CgaYGoRbwnyXDphr9xEyzmoedTXAMWXAjWWNkr+YaEl4KcBVZX9Q
VybEW206tqLYdrtC8rBpWwjyCNtxtLCFNuZdBDm5l9Za/H7pytJhYJC7ifT43gAihMaJbMUP21fs
S03jXbpaHb2ANN0knFdiCu5XHg5K40tAqln5p1AJaMca70j9+vCITRuSh7JSfOfPaeCnq7M9DFiz
qCmhzm2lyZJk67IhG4QI9k1yVa2RxBQmXAAyl15y6loENGmKyttP575hZ//l23Cl4M5vy52uzPer
aeDrcTD/7I70aKFGFaqn3slMtONW6CicVcX7laryshd2lBCq4VKN7k5iMt22KdD6tjVf3KJHoT0X
FDhQLn2+8SmTvUJYrlHWt3iXTxqS4Rj56BrIxbALDbkxtI58HyVvo2IpaztkEo8n+GUZ0bUcBkKv
AAesSQk2dTlyYSf0QAJoLJo30awkaMuDBFpQf2pPqi6Dwnq3e8gNY688aLiW4zhlpJ470wlzGM6q
mmCLecHvdo+CLCK3NwBG71cXDCMz3EWeM3Bv3+F/QVKT7ajDz3ajNm61SbZCYu2Y5ITe0Uad9lly
6x+Nk7X0yZS59pRbOZfRi+zeU1dUQxPMDrz8UONWQatjpDh7ik5XVoTUuwH1QbeutVlc2ob5J7GG
0K0t5U/SE49zssUIXz9vsuKs5iOrKJPPXQkO7JDBa03VKDgbIln0WoSSjhjT8quDOkMDKpSZi/PB
dztVH/JckfJwtfXNdpMMtdMWG7230g8vHjzC2TUNIAeuT3Fk46Ktya6sBHJmp2Jc2P2GWsppbtrr
aPrkqckYPfoS+jn5T9C9wZKW2QVaaZENYP/R6pZJtfi/2krPCzhJeF+ZeBmP9A64ezFyB4nBjy5m
mypv81gIxo7t3CaVlOcuK6G0RJ2sHtvKm1JQqpgDeRlcj+Dmd0vGCQnJvf8IBJj0OSwY+/7WoRWa
shDitrxofhfri5NbBvtIMORME5nxOuQoorEfRocNF1BdWq15GNXV8u+OEPPFU+Ktpb56SduXLEBj
f3p6cqBFRfHrZzNo4NSiFJRy8hSxbgx0AR0SxQN7PKAPOjs5lc3+l1m+BJ2BpdI3sh+q4aOWnOOO
epHBrjKHYvoM9udoX0VhHaqRgEPRo1y1t838Gizx/4ATi9RJknavj06cFiRsJuYJdJo0BLbMiPKP
8+VKfbd1A9wjxt/34DZ3Fmjs2XNqayY60eS8BWe3oGe7SevS8uRKZbKhwgarhNzIG/rybPHWop7u
LGuajBvtx/7f9VFPKA5NiDPGbrlphFzpFkpjALEk03k5aC6mLzPTn3ApwxaEZjQx9Tce8DZutgtJ
Korj3WjTMHQ1FEX720q0Z6+aOlc+IvoqUUKnGaNZKsMfAZx0fcP1uSWxuBy68mkENXtg8U7B2TS9
WagA2Y9Weyw2wLV85efL72h/JEUoUtA53qOQYHt7t0+PSkfQ84rGhiToekLIFpkkkMQLqob796Xv
uOVZO8o30mHHOfRFQ7VId/8EsKt/ejN1aIvWouwFeab/GCWMa/GTZBXLtnTKALAIboZ+HcqMhUiJ
NI8KJtF9UrHxvJPHOFAnkCFSaB62bPm4VL7ClVsDZay42b0NJTKN6pVCqogAVfxUAtUG/o7yeEec
8IWToF2iw2hVLu2+rDUMigrRD57jICuk8rlsYhz2HLwsbrY2DV6boH47AcdU1eNKSQ+nf5jVTU1N
LANMY9Gxlux5oLjAbeU/+DF2PUfK4vq9Sw9lXwq+pEr0cyVDR4s+XC/+c2LigLgrCTOlKfI/zaOY
c9t+jua61sQZnYbUUM4d0Qs+yzivdj02lHS1lnBjLUuExijwHa6S5CEnwW9C5WSrYdINbZKhOXEp
JWfqrAfBRk00BCAVKOuxjLAkTdC0BKRUqwi3zy7jf1U5fsoAW52GeVawQEJk+3YDayWhOOb2X4nU
P9L6weykbonGqWJzSsZduSKbrM3EF19yS0TsrNnGYZp02vC49SYpdMrra2twpNpaPU19b6G3m+RQ
cZIV6wMLJiiLLSrpJmY54+3X8EeE5eThHs2d6BTYTzE0m+V1w1Aoy2tkIsTWY4LAOwnHH0q14MPN
RiuNwxobGXDRHXwwwzmg7LeSvgeZTsubnJ6kTlnDLICY8GARIQhQI7w63ZUvCGoF5s2EQDUA9abb
NVf0/uE4Tre7LZUMBLieMLmY11o8kbxTL6d1d0QxU/OY58Qr+06d9oM3QMDT26gs6rmCpq23EZDD
yftSmQMN5Pw0vP413tO1CO95d0pNpFlRGgHBA8yGkg+4mqFMsayxEK4HBC0lCw9gme91pPpn2mYU
T06CQrX3NDaox+WYRPyTWj6UpHI+mTTbGVOq/3KyI7T+Y+jfM8T23M4A37l8D/ph0L/5tlSUEzjn
LQClz0He4gt9l9NxZGd5+pI14Z69rP88U9UD1UzAZkwW30mhExixiIrcyzHIdSMP4EOy1VLZY7Et
MGd1iBgToenwAWvkEwkcX1x4ShP70o1/uc8NkkmDZWQe8VkE7+rqeaJOWjBqIbPGmluJRvO/E4FJ
mMD8nDbXE8+Qj+oGidV5wtdAAfC12jf5rw19EcMHTZmT6Dylos++lLkJY8Mc1K4SD2P3lFyM9RmA
N1URyExRyL2UEZw+9kdj43HFhkq/FAjEaah2p3iJmfjn5qpOsoYxzqbFujz6KpqD3LTq9Z/drM/t
rDmKKJAhZ5iN1ZnfLvTl95QvYHOuOgOfj2o7jgcu2sBPopCmn0wisNR6PZx784IZdrN6wCknpy8j
vseWu0siYw7gvZ9yorYh4wrA1tzA6X41aL7ss+87GECYPRVU/bIBGnQ6V7qctPEkzACu6nJBk6ll
L4G0B4IwG0Kd2JkHajctcmq1SNKvifbczklOOla6fqwTcDPa9KfmBrhEVt22yHcNf39zaDBwqn3V
WPmBUNfj40XZFXQ5oMYkBQrehW3mMo2fsgF+YoqvVbAQNZIOfuECNWmtSF8We/Hl136Vu9FzB73g
VIZQS8rdSu4vKtCt5ySkTRLFNjKeWdCcBCFDKh00ltn226JN7AnRUjOY+lcTR9HmsKYYGYhW8njq
QzFJxZZ+nrHsQ31LKzk4LFJBYMQe1pmFijG2Kpdql5xYUin7Dz/4/lx4K1wXx9n3viGMDCkheeCo
iTOj34GhurmimLdlOcelq7vn2w84ytEBIZLtlzofJZTkWqchCAqHtecxRpNdu8L6oC3eUAQUZJDg
/TfZN096gCCJKH65PAHS3C6q2UhilH/QTi0OiuZDteVxuRsEgA+iTpLg9TA5CEYlIG+bOjG3Y2xz
UAKF0vSi6mYAQv4jE1XnMv9FbHallMq9002N3AxDzhMbkOc5rgwGrysQDBNNN6Plywybm/MLynZE
Qma5YprqdusEta1ik0LknIQ56j+Li/F//U8Dz6iyAmYqNvt2WplTJjPEE4DbUR6EvwjntnBECG9R
rBlCA6KKL/y6SuYhmksJhCR7XOA/7OEbUfgyflApxx1NWiEvL8ePdgPwm4hz/oqgVoYWp5dYghMc
orrcHHdBIl8YorlFrSAxhTbdWSuK+O1lOJxBB3uKXsDMqd6485y7E81KFAlb0ozpGAfKO/bIBrBy
GOH3/p3P2vf6M7PMorS7yFbbqZw+1N3wEx/FimrQkS40Dv2f+hr0mLQZQvyWq/ocO6+bvhSm5C37
YQYUt9v/8Uuv5rlMqZgOBVBBL8mWkzPhKr9yULBCFBqsWQutkhbsI2AlPfEpcZO8IDkLB56dyTcF
yCx1EGj11i7MYwfhQGUXA4HBiEnAn+KZVf0W6FUiabVUM6THxpojTo1o/qpl1TtaA5J82Z0hkMKG
NMp6Rl4I/b+A98elWyp7M0+y8T5EAYRQWNQnBJUrWxQcNNRUbCt+ir1eeoL3P7qxGDtaN5P0xE1y
nIBz5uyBCN3mEjnwqw8KjQ53MWcq10bJUY4YROGYL4/3jyLJ3V5IfBE77M3GhN3zyHqzNzJHZUur
hnFsIeRYwsHbOTR+qI+B+eaejY1u2dZy6zTA0+mYMOVWnO5fE2wNQ1ixrTvgMPAgICeS/d9z4kSH
JTPmt/IOJrQpil+x1mY0BXAaHrmy+h62CIUBe1n8PFzUxqGsctWb7IaKL4V7AkXTmhU//rR1zrkL
7kIHVEQd0Ahlc3+qaLbMDqet72thyQKCshItDti1YhRcNsnbRYeCN0XQYhXNduWawYlKNBF8sMVQ
HiXh3ffK4BRyoXZtjAiWad4Z2S6OGxbdnYG4gM/SEUYkvels8Ji20GjDn8xGySWzfCHAA6L5LI06
obW4WxjqhwRWcqFHyFWoKH3PlH0yYDIONBzTL4Y6DfI88QJt0FSc6sCluKWeWf58OvXK5d/f5ums
MpjiC6/QEstJsNm6woDtuRZkY+ewX6Y7BoO3wj5UNCgrOHPmk7nw6kt8bBii5TylTyoS7hn9LY97
flgQA6WMabplzH7yC5IiJ0AMI9MmTpwVaveep87oFZ4ZjNtlLsQmYieEYd4A86UdPf435R8shL3n
vazyjlS7qlVU8ALZcmN1lVLKK+JaFmMZOXVQVP210B2/6zJIpZgjsYBrw9XGS656cF2azu95Bw2x
XxVJYVFC6RFXZPJf601gz3gtox5Clmx9PClY34YglBTa5JGW2jMotOxgPgjKM7TcGr9CzmAHsOYP
pqR+VCKh+H9ZV/3LtQmWDCI50rh/dUAI9UArc/BWWSHaWGQ7wgm0UETy+QIp0LX98PBJpoZlJb7B
sXvhXzVFwbYn5u2SJrqcVzJGT1cB/DseyIeinCsKxoBD6P0aouZHTkxohFpYQXpiqV2VWa/AWiTO
K/wRQDOxDjZraQj8nxX0vHE7oSkDTG7bbz41ZCCZsA1ock3knpuxwWIbIr9Aou7mGRpjoYmHeTy/
s96NPxvXxBa2yzHQQSNq/jgHAzN7bGZjCziSnvmOOP8Na5MGdrzbbMDVyR44yWbBGZu0zfMzjh9D
mkcfCAf7dIb3ICYVVGrk7UUOI3CU1VfCPh4E2bxjcRAY4cYLq980fwseGEHtvbsjKSvHxW/6MMQK
ZiOssoxiPh8HGFqzvA3yiM5FngueXF8gRNQZE8dtTGG0BqRqaGvSP444gxc3oQt1E98/HnCu7+lZ
HC21mSAqhsTaIhrSdKRfzjaIAcfllIkq1r86ohTdkVi6t2ill09+zbpepkwLi9qz5ccDr2r4uTCR
jz29LoIR3F2so6r3GWQ6/K9N+xcRhr3728ZCZLcAFP9fioX06YhiKM2M5xU/+8TzvC37ggWctPMS
GuHfqNcdUlwWGI4VskWiL3P+Iov5X6ldf2rdTtU6qmZbvamhiGVyFKrwgpzbcUyhj18JNQm3yho2
ZLQEwDa3ge2SBQGUKGAsujT3PXR63+gRNqLeBMfT03dt416kskOqrShWbjutflDKOWvGHpcRYnLI
rN7mLhGfn66H/a/k97UOx07evAsS6dt9NB6RadQMbr7tbL1n/i2RXV6+EA0CpyHVHuorYiXNIxHJ
Jwjl6qdOMvIQg3NRSXYFZMfQAhI1Q2Tva3bEb8F7TcV9c6NUVsxozgYTqTDjIU2f0yie73v768q7
bQOVj0dZCQQbTgvmb5u7cmxRcSCLL9XpdW7dotjQajMcLbVTdRGzuTgE9x59gb8oeklB2T3osxMK
HsvXAek2vB/AgbxlTSW02t1QV6YLfaLGR2zG5mhoWH8ubg18SgmH+JFMED6tmt+jZHLbdGXN2dnQ
+IcMSJf/xsP7jt//COMJOj+JL4leUXLSdbzYygqL5RE5/M7/oa+XDrEV4SOeOJLwjhS4rjUNhX0A
VEclJX+WLTWohKKtJpxPB60BRcgI5Sej/QUc2F1DAGCWjr3y2ClKziaMvfOHMobwPghxnu3MbE4b
1QD82y8rYEkhV4Lg4o189YDMsf4ExbPbn8diBEspf0C2uT/Z+Y5rygMOMozJFBgAxtPH0DVoAI+H
+XKduLrcecK63ol8xXg1kDiStW0J6mcs/uL1Md6JjTl81vhRu/gyL3ziYPnpHeOXYPD8GMbzYxFr
SB+FYIxwC6I0yR8Z/Opqlc4zV4zqBX7o3ZOulMM0wNkNwkLXS0pWKqfWillKzIdSA3Ljxg/rKYtF
Cy5Oi/tbWst84uQlobtasX/jy2RsEPq7cuf90hwktfgnRZkdwCLRR/5gvbKOOzL1iQhKbpRTiiZZ
im+7D0nfEBsBTNODKhYL7zPDQlqrzmgrjYtjSoAhE2J7W/wspTEf0pYmhd3O7VqBljjZjAY1OYUQ
G5bZT8lpOi43oNVPzaZHl7SVMizUPUC117sgpHPnvi1DdOK/T2a3SrLULImDmOm9kYxtO4DXiRUX
GpDAAaayvtIHHpxdeenNeGQVoQVrUh5jUYr8Lrte7hueFwSE+M0QQhVQVUnbcV9HCvDnNHxQXnfF
H+IKqfmLMJ42tO9oACsbSHQyXPzjZ72W6g9nSWh+3TEJi0xJ0pzWi8S+/wnYE8/ffaSRy2jKpQhF
LrfBXiXyjRnH9dXrnImiwdyrq7NHj8vJSAB34WNZM8eiTcQwNFDldGRhjldzpTcsHGZ1qx4EUyGz
QrhZG8BMBTakaam/P9WiuFOFMlPeLa1E1+vYjJajLTU28VrVRpHylcalphiTkYJNtcyTcSGuZ9hM
yL7aJiJy8wNckY2GXoxs/n6h1Wc/1nGyZ0V57WnyRg7HSYwbe7BW0Cv7ET3HcHmqqj3YgBDdD+me
0ZzLyKBippvpt15Hagk/mVVrA4ntPOgDiPK2olb6OP7cCHJd1wOwMHl/UEuVeIi6U0hsUW+PD6xg
W/I/s83TDJIpnG/7RtHfoMmygbOunvaeCpaG8Mhyw4VKswDB7B3KN89AzyeHVWkFph3bUKc9Q/xv
EPQwIHKUAqixXnAiO0fD3F5kK84YtWkAgXj+Vd56E3PYT0fwni8vF3f2g9147VNSMQ5FsxO4JDVf
WHjntymcya20ex6+pqrHrJySp1flICtp3gI+M/CQPnxk+UlRronZWpFr82EtcA4sW4qRTEZeO9wY
60j4r1yR8m1v+54n3cM359rOEFjsZ3pD0KpTvXTTDPb1cOGIm5p61nn4GtFlQdWWzIyMF44xogDu
5zzJcWI7Og84uPitWzlPgC2b0nRZmL2K5Shd8cZqXfTSew1hSMHUsl0VawIKKuiP7jeppJRSv1/I
c5yPDS5z6CbkSpej26dxm7AZyXBnwgBXsBIj84A/PaJDmC7Zdbrt2zkGHSQew3jo8hTRGuDkxi9a
SnRHytWX3e9He+HD7xw8r358SXcj8293M4urMcmLsZw0Fo4e7CiUkQsywI3nNd7zYjColKPjXPbA
TlMYByP1omiwvEghidPr+JJ7K49nnGGN3AELtphN3sc2OeJ5X1PFhrpmXqpjMtraAJbMzILMNSyE
RDcmdt1RKPlv5sok9uvPYSXQPyjm4wqiXhD8poQnjohqL1CrIjCxi+u3KRuPW13/knOVn+H0MDEI
b8UtKnscRKBw/A9mwAfstrJvdWzrCtxrjhZ16ahFoxBPYqKPT+vvVRvHhQhcyrJHA1Wwqk4XkB9l
Nt1fxh9+oX05N1EmrUn98J3DZaKmD3HWgZR0ZfPHiSHR8A6ndyLDZI+5VpJZ4Ckt2cWelTTBCDsd
z7Lk0eiCeT/iYvaWkNoug7sBmUJUJxuwKWIAfnsbxpT17w/kkX8krI6r/GydY+i9569+3ts/Kot5
l3nns/5woz74KbDDV99wv7cx86KcE9AOVzqLjmTWGnKtBMANHPlEeiepyCpvgj+lsF/Sb7VN0G+x
823HPQfWUXR+B2FSeMDCaeU2dJp5mhbjXTNIdnfeGsKt6LaGWH3Xknu/Z23v2O81u728aTt8x6iU
bbsHMzOUxmKboUIO7535sjiYxXzmGVps04UPu8iErZ78ZNjkW3qamkxsf4tmz0ziRAIXDcqb9aQn
VOYUSX4ybFPrlahVgxekapE3RfBzo7QO6xEUWK3kkrz+nIBwaM6xZutPNPvPK6q+gaL/Guuomo9F
oh5WDnL0meD8s6NlzyEzJnOQ1Q9ZXXS+6w/OmFj5dAGB+CXSrztTyvGIOHM1y01Jz/NZCD0th68/
8QUobue9tGdnxVEsJboL/mjqye3TIA+JPFKjwhwfgfR+wMBC8LDf2Ja9rEazCgvchlJpccgKmJOZ
Ty4JOoZCNrPV7UetIvmU+hqi3Z2Z1Zyi6RjO8rpHhBADBmRql0zdREdTiCNB6/vK6u9cqGEmSk8w
vKF7u1i7fCcYZZp+M0WasqEy4ZBSnwxevNAKNWXDalBwa0ExBtY+vAXNSkehqxpr6Za6XDrnLspy
0vCs/tegbcyJDWf/83OPiOh5BmzioemOmViMNp30pqoaueZNrL3Pcy8/uIYJz4sOlrN+M9gEPZUq
cGb3NYO1h1Sdt9lcUg6kxS0jc+twccO3cxGou7OGua9XCWeCVmD4+fA8nsG+u4ULq82yYyUOpKnY
3MOjYZ0ZqSHsLjJ2knkV7MM5YQNShmm22oR8V1qiaG7i69o0An7rLCm7K1uX9cIFrYDtvyEVPRD/
Py1mrLkuOhFveyXoTefXRriY/HxklgaIyHm4se60Pblz7dUa9Mywj4SR2gYvsjU/7Ksq4B1L/otk
NI63zJ66ZlCW5pPjy5snJLqXDuPLarPTqvnztHx9eDAePDNbgUqKajn34CQ5C6WUc2ktG8yfezV+
vscLL7vHd401hvUtvYUKUHtDja/uWvPUJa0U/TYNE+NW4yprn3/T1QHEFP/XxhtF5RC+mA8GNEeU
iyExwDOwgYxcvFKKwKUiM5MJH0b1O/Ba/pXoWiAshUPYgf+DorTs7Jgiz4vQ2sP3tawj1/D1/qLj
Ok4Nq5GvdMO15J0cfaO2owOI9/DsI6D7J5iO+8WLFQZYXjXVqp6yGThKgrc7Ca+zu67RZkn6wG9x
deLv8GbEN76hDZyV1UB6E34wf7RWtyPh6E6c8GDlwumu73n8JOwl8iy2u/WqPkwiucCGmUOh55K8
kDFE7Lah0CsawXP1CCS1cGRsyl71jctxppODcuRV+5kG7gPUelhV7bNOr7Rq/0Q9WKmii8mzjVBA
UpQUqgBj7h47cXlhQM5qjDuSXUDZAIT+QhQ30ONogC2gsYobXqxhECIKMYKwZUXlCYmuUOUt4kiR
+Vj+tN4bajpgp8iCthu7pUSvbK5kqb3G9zuTKqa3Zigodcf1y9frCT6s55uEv2FjmyG6JT9ayxi2
9eIr/Sdd61ru1ThAtG4VmLdsoI8UdLEZVP7fQ7edSySP4+gGJEkADrw9d2GpE1hetZEoVjLK8Y5X
wo1GokbUwAsO8ZwAbcMhWOC88qxPOEi7MrhQ0eDNQnzLzlSz1vuCtGqpjSQQT7xl53vn/mQ5u32m
OTjfBqClGGIYOgeBcX1Jiq71CO7mc+Chn0jvtaYGx3LhdVSjnsEi3RhJVEeoqhzrR+AuFRRexBBe
AHdyNoukfTboELo85HeIVTxMZPY4YAfpMEvLaNOB2P1y94vDYCu/rxwlkBNsn5bNjQaj0N0UhkEN
a2oFZOy7Vfs7oyCFTlxOvhUBZtfpybWFVKDrMDbJKXSe9gEU55OXnYUGtyDnph7WmQJwY8vQkOk7
DylD5PYdqkRWnOa+N0H/sL3AsX2aZ6yXe8Lu7NkhmWhQ22KDJEozp9dih4gVTPTg32+FgBI3lf2u
/rvxhInLc8L0fx9onaqFbgAD74nMchRe6X5cYUW2eT83Ua8kKU1Nlu1wTCPX3y/PJDuDWchS4sbK
FIUr/+yTjrH4+AQCFuT7UmV13MyKzj+GSejjlYMli2Ee477n5nTbD8UV14MrQcQK+A1VDkPqzrkW
i/p/jssUBnJeCgdZT/FovSMhFW1egThX0Y8BW9hQ73JmkK7pnqgeQ9Oq1mlVCAwtIyP7VNwRTi71
FPWrbsJXhrze9/GjYdI3lJqyKuTp18Q7HVNF1XzsROq7y+jv6Dm9T0nfOV86vUAYDL2jvi2Ne5dr
F9tGQpFp3o4HdXIazRvfOs2R686VethjlBaEypnIBN6gfHlPcqaUffEBWRwXQYWv9kk9CXiEW0vi
pUYEf1ySeX4+Mc07sOTiOOUrVWJI3D55Jy/oB24mO8Kmt0PFX0ryEt+O1aqgKw+a3SkYRNDeqTDc
mWlOsL2f1qJzYXE8mIuHoysEh6A7AA80Z4VJozHyIMiZonMoHBf2Vr+goqN7h8wwPDmZ8iBHMijv
Bflw1+7AUmLG3MPz9F2og5yo9OQ8O85hqy/00/e8zNlpsWI9Qyuv6/Yp7dMp0UELDcza3VeR1f2T
uw7VBcY8D4eQPU3FNT40JJBZ8ljjlhGDV1cFQplxn9HkQEygvIKU4wD8Vubt0rAVIGmTaHB3yS4Y
lSRWZfKBeYsh4r3qusr6vnZ7FMXobOvgUy2j86UjSLx3Odx/aQv+aN1MZWAofAzriyhpv/2jGx/6
6U4zZ03WOdCJUHAHJug5PJJCNCri/1/kKWSQEbsp4B4U00tj69T3qtkfhGB29UmOYuXWEMi1NepT
Ujts9xoSrjFKGsu5dEclWnSAlg41dcIwYVbf8B2sa/E3HdQHJmugaQ+4WFv+azRvPZdeJYT5gTS+
30ZlBwHzkqtt2GUVvUqLos9QCgDeFunXBEdxmqAq+Z0pni9bBMgpHEAXagXSKXbuyr0BuS6oRLhn
QrwGBmSdhrWr/QS+4cLZxd/fPM99/ciQ90IYd6SR1Js2SGYPdw1t/9yY/DVWWu5CzPV4zEpGSOvf
HE+JLt4iPdasB2XcPFR0xiJyRTpJbGheXjlmov5OyL9uLa2Qfnd2Wden49kGmj5+v2v6IVxRHNPp
Nzjua6bX6kvh3oRvx+y8L0ANcAR+SvDIXVWsVZ85QdXQcL+rKRzvM06bW+Mi4hXsOX86f4OYMuCb
+mjWP0iH8ywfcyxgHx0iDb93EmKWts+uLRZmcurvtNR/9j78J5Dl4hRwXA2gJ1e6vB1fWyXax3Le
7JT4LTN48V+0cM9teld5qXrpYDYJ6OfBytRuC/3K2UG+VpBrbnBjnQDpdCf8WDkG9FQcL8Ug9lpH
a0jpESBgGFcZRIc9GJb6mVdvaTK3RSVcvkPmuVM/r/aGS5Ny1a5IUWodFfw2z7691hzNYsrcRdJB
Bw4xtVQHgs4uws/HJuBCly3CINVppC1oxKczHEhO9vNS/3sDXTNR2TX9iRPW2M+qWLq8B2iLAqLw
889aFx0Y8qRBuhEY2bAfTb5u5ygDucOXUL8tD+bTHDrLLDVg7SpBXUSGWJgtMnOf6cn61bunTkP6
SsRTavRaI521hoZRX1+erII1mhwx5M9GAoTxJnlPa4pCstfXefqwMSAulkJ1CbU/wIxsQ2iEAjPK
yb/luOJruHeX0sBMmD9lYZVTPjkDZw0lmFp0E3SLpVw5B+33sRYntBqQQDcZ7QMN15ecwOGeoal0
nlNulEnVTo8i+LebNH8Pk+UFOWR4Qn6vg+KqZQymAeoARkgwVj9oIucWS/MA4yH/KBGmqhi1oES6
mlCKzERgmmygfLgzisdv7WHS7dgh8uJeL0PFWfm2bV3OP3EQNlPSAi3D2jpC8dL0UTmjoIjKk19f
3VinQHxim0Re8noVvDRAwB/xO3x7h0swkOlxmlH08VQd1rOwCMFJrOyK1d88GG5UTO7ChW0FgcX3
ngQ+bNWUgvxWvfWguV8RSgAeqas6R7GVPGmgkvBcs+wPQaM9cYNbClu5esxDJRIW5FVOxmjJ9YN+
SqWjwopHLd/p008Yn0E4ntUmOJJs+J9VAoGrjiL0zEzAZKohupjNosQ6+heCer/d3YAHP8R1P9DE
TUMFmxjHmQi87seW/nq04X+xfUqhfKyn5D4RvEjN2oPEyLA0NIq6NPKV60o2sKiMvdfQai4+0xJJ
YOfy+lgPBiOu5N4wz6X60xdnQgGGuOBEunbU/jN6TG3S25NfvYy1hh+Pf/SLAssirHhDpHEdeKXU
tWvCRbT6sWWlkPACKSDtTBkJiNH4y7B1FGzXdvR2GjMfG3NVZPgHTnb1eGoT8ou83hu7uFCx7qNO
s3unUbB8znpFcPmNybPcTTURbyIWdpsB4OG3Cm26zjhhAQBZphpSyfmZeZC7BOAYyTXiOSkh4nK0
qNs39s/htwKBRT0F8/S9DKCechici20NQm1FFmXxtB/kwOFuUsSG6//3Qj/9TQ8T2QwYnzi+sA5O
WdFn9gtWO4X94vdZ0wA0KUqPxH5PRsL7IzvCfMp3Sg06hDJzjgWngveWN0mkZPSp1h/9PWSN3NFu
loHd+kdI27zv/Gwma+XxmaNcUgpOtmIFRxXj3PTYJFUDMHEED37VsnKsgBz+cUxzy1xuWL708cvl
H5XEWexl1zNrOF9aP1cmWuTs5lTYq5V5yrtQkiDKp8edsUdvaVnmpwi5W0S2vxlTNcMJF05HQqxC
W8tOqwqy0FTAxSAmHO0avzuOLW7Vn8DD9cVtYr4TK97YwbzXZgFcmW6KpGNRHIKLkcHAkbmy1zN8
rKaCsxGevqulswMNZLajxbZXRQ8r63EkolvZPMFrLvhBudnjgPpcpIlEpKUiR65tTTqLUZXD8ZYU
UT1QedwdpNkuh/YFqqe+I9B+ZkYXCJ8n/GZiPKSCdaO0sDz3aCxqHSJE5bvHrxwh+91IZLMCi2AS
IAbyOYuTOXYT572serRw6EVToP2YlW9SzQ84nKjWZhJe+Ficdg0VXFcr6F6J7mZs2uKpIJ0ybAV2
WMS8ayEOdsK9UpubEKGSBxazSCeYRuUwtEhLNc4IdvvFdlNm+FANvQDnq1XYhzSfZUc8FzAmeU4h
EwGtzht4+JCEzP7ZkxwMsuIqyYoDPHyekfM06nw0u6TXfabHTpF7pceHXh0RxjUfb3Phwp6c5aLC
tmqIogAYiD0WnC7PgkdiJIjBGBgDbFgEJUzJ1izyCwnXarTJ0qWNujGwoDSD/USkxMAOkJaEqbNE
Bajqp1g6HWlZU5GRUMBocFBce5UeBKfxOEA3co0NptVXPljV311OsLvpqIfI3QPmenb5YfYTOTde
2UUF9EVLFetGo9Nri8N8auncRv10tW7ToDTyN921YmKTvY1rBA95dVqQPLFDb+IzXb5RvsDcGEQX
8xFE3cLU9IJExX/jzVmV6o/mHfRgKXQoJ1mfbl/cVRKCXBMHkb871jpIzt7QD8acjN3jwazs0Pel
gxnHD8bFLBoEvTuMkUXBxWkd3h7PtH7ABhz1WOBXcu6vVJrjjUnJTjsKZCP/e1/2p4g/XK7KQglH
xMlhdu91MTQp0h9OFCmt+u2/Hiev4Jt4UzWYE9mi7/LP3Digep6QoIabYN66tCLKKFt2MfDSir/O
FVY60pKRikMZum3onk82TKBHDDblGCw8BMpYULaA/PsvLMaq4qfIbZEWYSMolvoTZB2+/d2j1qoO
E2QDXB+txvYUhO5cn2muMuhPj+Z3rbqCoY0rR5+rnh/EYyKoTTm8rdH4dQAWb4VlhTra5GCPM+eJ
fzMTGy77W4CQcsdYX2Pwtrg4LwjvRNoqyOFzHd2EEnTDoP6Fr6fFH0soijiFKMvuTAzq4XzGEyn0
Bp3QnqLheTMkmxlHuTthF0E9/e4T7lV1vukwqS7A/UhyT3CXhaaJx3RUdZhnAyIRTObnyUM65WJn
vyzqojahYryrI+o2tSXXAN3pUSvWOhp60Xm+cQNndH014xxgeGbBgUcBAdnHmkxlvGVhFNL4m1Fh
UZRKWNzAhTlJIxofsyoi0+vyeSaWc0biZa0GomEG23LP3DgGwch6dYZtFYbVZOa0aBhqNpTF9yLW
/Qn6zDfgi/zJQPflqTxauPI09aSFDBvx8NDf0LSjsLhngPpOIwY4COUUZ0WXPdB8tjyCYkYSH1VR
I2EiiBj6nEL4UzXaS2ajXGVHlnOnm63NkgfjiE558WO/2PY/yUXfN7LcUrzbMKExiX/wzxcWytCq
fYQ4O+vO5V98Vdz0t22p5OL7iEFI/k2W43XUqhm8tjHwIibyzLQk2PH5SCbhhH+2d2mXtgvML7aD
YdJIF6+ZoQfHgmBwb2udAWWoSDY1dOMLUfLW9VrpbvwC4oIMXEihm3uesli6WxcUCr2j1U2xhBdB
/rscTVVXUNkHYfijil7/WHQhNN/PlN+XcY5ZSAh/cg7J5HuzhrEQg6LdK7mNUfK/X4YTFin50nbT
ZRmHyhxMKD4/hx1R54cg21wG1c59i2aqI1BsVkTPoGgXLNu8DzRYkkfFzJlC6wSYkp2nDdZ1d3Ok
rMV4G/agRLmY2pCcLKzEy7RZEONmotOCt8z8pEFxMB1f6VnVwkiXhtbrOD0VVqQz5Q9UgyrRdmIJ
WAqdDtm4HR9CU9CDUGRL6I+5KxlSVsZ2t4kR7pG7oBqdO2C8zs1/Wp2822L3cocJbvvLfHwXYQZn
RT6VcfRvGwReSL8vpHqykGgKmiIx4s9vEUTMbseOM6hbOKXYn5xIr84LLwT6XtSpCgMBBaofnhIM
ZyeeA5vsO2PoxhaB7bjVPIRBXGI712Z5OzgrqJ5g0YXe8YXmrzW6jY/lzBTG0TH5gtNQGkeXYqdM
pz2BF6SRf3nUy9RNzpM9XQ8Ej/4AbstqCozSN+2pGdyOdUpgZ+pQ/GmJ+GXkm8zrA4J6N2l2z46K
lRzfDaAbVWbux855DNb8GIs0IvyM1/rih6qUWrsb4Lu1Kbp1kKzJJ89CXsSrdi5gbBrjG/hD9NHC
UU574sP6FZoOOSZE3iDfLTPazCIaopLzYW9JxQJ3DPw0zQ2aDM0fnngFHnRM2BCybPWQ4C/9ihke
KH/U6FrHLycIGEqPZ32rAK8/TxEzEy+Au/gEBsQ2lXXOEowOZMsFvvNSgsGEvfd31+BelrrR2k+8
rUffC5GUzcGlF5/WuELTFUWiDwAK1Hh7SF2UWg3afo8Xr4coHHUGYG8ARUF4nMBYMn/eYSXh7Lza
G8Bt9JMxViKOBC/NPI4hYHHBUNrl5xKcvp5hVfFcoU5hE1uQpcUzsx+JCpJxb/TjR1HCnSO4HG5+
od5KABZdw53+nSB/2p8fPf+/3W8LlE+E+iDtxXxhZFwap0ApERPHlYT1z6AQt5KcZuKP+2mPvirU
lZLYXUSY7jd1ECG/ElOpatOD27xK1HESnDv3+XyNrNqvIZCHileY4hbdkaOHXeTFqzcS84m/D6nA
xRsLumy8KcUAXt0CEl/uRzgHIfof5x5zK+euwR9uGnOZqEPz/ZdHIIsHaq/pCBIOiyARzonD67p6
UGt+rrtClL8faFD6WQ1b5O9smqLGcq+/m2S4yOTMXLvE0Ed8fv/mOebO5uw9cNcTw3+jiPnQDo4b
EWXQHT88uxF0d3qy07UqXZeiNmeiunhsI+yBMBHn6NN13qxJuga21U2tIPlzoFvHcLMRzCyApjHj
IvEpMEYDN9EnAvhI1WjPmXI2L69ONrE5KksNQvmyXLnU3GEQoU7phiWEiWzLhyS8daXHay1+V0ak
PQbQAmvAv2uQIx61i4J05oPoYsC53lBueO6DTHL55jMeyHbzWl4ysDLyF8WK35kMuSjSMkhAS68s
MmgFotc4fNecAGr090xMK9/EwixywiAtjdWZY6aNKT4c3LWJ+pockjJJbiS8GkYZM4Uj64zli7Oi
VVsNdThBBzBDAY45mDKQZ4ZErMPw4NfQBwvkk7FF9YtbeGQ59DHYvmWgjRqzccL9D4AurkkSRSTs
e2Rt0xv1CdFjWJ5Gy/QBhRsttEAtRN048fZgFUaG6vwkT3ysX1HwRoT+/54gMzIugOYqB1BjxJTP
/w5rCxAnXBk1KEViArsOlljHPhvL0ym8woa5RAk/p9xDAwyPRpTtKp3tfcIm3ZgtWELbWHSHdth4
WVo/9DJDILHHZk9kFBbljJRinU1GIRUoVS9xDCTdgVIrg1W0Jyn67r81z3VqBFGepePR1GBn+Uoj
liJ6B/Z3ZDmZ9P2YYd/dDmy7HCBAqR2LlU8hVwaVZ4EUaKs3Hn2SrmBKuaDdMNhrGu3gW43+UQjF
Jg8uDqz1cbW4VaYw51ENH7F+g2gHlKzK76L+F0CO9RBHFgRTVSWszPTzRuTJawkqQ36W5RM4SmbG
mPdJLGdKoxrfECcp2RMyeI7gltueHoFAYAep0cI1L335HblNO6lwkHZADiN9vyPuc6pSFkEmZiEe
O5dg5DgrrAdEVRfLJysB7kJPJssfVyiDNrQgxd/7m0hQWXoipiB2oYrnsufE6JW8tyZjE+YNTCBj
Tns8wzdRfy1QePIAkx9xJP2LW/SHRcvjqhQerAjrSnhZPtrgQSTfcyOsx4FhQalHB7Tuv946gkS4
NSyqhxbBo4kkQ/EDdrrMFp5ysQX9eq9z9PFwRwSZRLpNEa/a+cb/6nZ0ZnQwb60CFvWCNpyz1mjL
AYqRZlfDJSOkXuHo6LsSwHK5CzMf2Od+XCK+2Z5W4rffhU5Z99eTgdyIL3N8Vlno7BWthlqOjiKk
4AtB/GmSNJEDytre7XdVgQ0bMZ9R0Ku+d4GKzDvDX6GyfDgLJj6+syn/Fthe8ChUr/BmJzG0s0GQ
pkEK69k8L2c00h9diuNMlmiikXNJswQ5Mn2recyCRaP0pL+3/c15Ks3+MTKh1abQnlQzxJdafCcY
SJxsy3+Tei7xravyzoKXmHeVcc2MzJvgDMKW/152bEfxBfLZzmnC5jlVs6SmxBxJdUmB3CmOju2H
IDQpidRIKnosBXA3E4+5U0EJe6chi6AvlIubIgPF9q0CVYi3uE5x7e1trcZHqhbht4n3TJZD0Nn8
B2sq9FoeZHRjXi1ux3h5OVk90wVKQOogQhdgwoquXm9VaTqQhUYbPsjy2JUDUH7g+tjnrNMZzyaj
DQGTFZxKba2daodYixWhepRjpY2OKxh9qvQQU+6Fnrc9wiX9Fp1IUiptgOcxQa/BRjR1WjoLUxZm
MXQib346tGN6vFP5yehdQOpnIZbzQijoolUCTn/840ccGVRZl0L25o80bWVbc9hVbhSgEhQwOWAK
zr26yCrVYfYR7lVmNeQOtIcgTyKgmGvf3SZnsq4ac+Xz/MJuNVauKy9rTEiy3kCq9IhOL4lgmfPx
IqGORqcmSxLPtki6pHCOE8FO5cQ1T1OyuG0q5VplMRXQce6ri6AEb6LHm08mfleOg9Scs2kBE0I/
p/LRn3BparLePvVrY5Wdx7hsA3gB8zyXpTK7YUc/0ZX0ZVH+pHJowstd2cHIZg6p4L+RBa8ShwEf
SNp5MepWjm7936IFLgfEm6WTjSmuAzy8KlKXtTe3t/iFnXJzQ7aswMHkP5zUgKOVgooGN5veCvvA
bb1R0mGUusNo0pxwRp/xTpJFg5sDzJuzhVVhWux7EBSWTZ/87K9qufVRpNY1Cp5mq8FNlc66ZNxm
w7KlzWsOFFynPPSiMf2Fb+AkaY/7p9bJerQDTWaVQsmehsVOgoPeBOCAIpv/8eJwMJd7p2pPsk+m
uwqBxEucG4l7kebLwJiUZAPUyBOF1Qjd4N1p5J+L6nECBX349+PSgru5n13GWdnSRRq0mZwEwMGy
xJ/V+xNASqOnr9vYGiyZXMIGSt+n32pFddYg7jazqQ9sStHou+GfPtGDpiMPNno9Nj/zMnGNfITs
CL0EOYrU+ufpkjaYJQEsXba47LKt5HRXHUqg76YmaNIadCufnx4LbO9A53hZM9doufKE2TE5VChj
9PqDB+Kl9dWT9dDbfOY7Myv/g4O7AD02NUV3wJZV/V+smSY253Vet/UG4dSfJpsokQE06XFaLq59
5gGgKaosRCelW1zkHaZMCLbFnX9fEdMnDv802QL/3xTWjfGilGY1N72sLdl36HSagHwYBg1IxhSA
GtObQddUIhioCrqcKkOEic3AnZremSCeFYg7Oya7hi6exw3vinDEgFSjraUdaIDJ2VkSRAwjXIMK
xG1Ix8X9HKGSPvu1/N9dtv42NP3aTcdjsoFWjPMLPNIuJnmloG7XJHt27mFPqsBXIMhjpUsy1u9K
Lifz6ZigVEMJp20dmSMTaC9zUffJvjeYq9+QLAYPlSr6CrcrqPLoW29eEsYHfOFtcPV7GTQe1saD
SaT0VxI7OI/0Jq1Np5e5/e+wxv9MqcIJiEqw9o9bQPxvzHKBO/kNRc0hrkxrJsQYKxO+29nxITTj
VvwJeMjtrZttNvponHDPxM+Ms/RaU0rYmUN2uSo4Xojfw7WQ0ozIMfyGRI/7AEJY9BsdNHAt4oti
WPofhJZQgnP8IL8L8lbJuN+NzYAVKS+2qcxUTSVbvcRIMbeKxM1iKtwDhhfPlgzgg7nrKkQezO4I
bCdBJ8zuLKPAc1JUu9O3PBPM61bKIIuYOmAscLloT6dW9y/j8CQc1KuMXusyfixQ+tp+xvEpOX84
AFBLf3OU5gsInBIbnvnJUgNVJ5c8/5JY0KXrjOVFWwlxi7DyK5h2xWdpjEKyeZDNwA9DxgnRtLuf
F4zrQwovZKPmEhhq3JCaZHfdv07vg/5Bb8JHBvBAENMejSYVjSy+C83AaUMe/jDz2eYRAVTG/vRx
0gpDcD/NL8G60DXRUhXTOS5kMwX0IneKa5JOCwRNnf8vr6BK4pd4lG1kolGuZ7zZr5nulr7FFWAq
Pcmf6gYSc1sqzpvXC6EMcbzRF7hrfkC92EjV77lTbT2akRKrwAONaO2SPtUVXWF4PpzRmXy58xmj
XBpovADVhrd1SvmuJmuZbQZ1fd1NHa7TLTgbloSyyHadfJjTyRpAUrY8U+okYISU6Iwi80XQ17qy
mVXO6iDfQh9X0RLu/M0kTPLAJtVSgbIgy9U2rYEdsoJsERocho7ieCZFEqYZKK3LbHck0pCSOL0e
hEcLNt14mhUqJK4+sb6QqnN31PtaCZByX+vwl7koWD46t+ZGMoLGUZTibzFXTiABKhqyah8Cc5wc
28OLkvts0dZ6wUwNXguACOLLthmLf3AmTDKBcpx5fxO6Ge888aIyTGoniGqxu6vyEibpcNl7Rkue
w7z2EtfMcar/00Va4NPSxEvbiGQRM0vqlO1Q1X0KX8mTdNgm+vsCm3L6OVNR8EIgO1U/dwMBi7H8
OdUuUzuoptvYerOJdJpkfSO0PiRHjjbOh1lY6/5W7IzE438b9cTBMHCYidy9wQ/PP5qn8q3vT7ts
dZbKFp2ubrSGP65HF6D65xDXEPkY7GsCLTpUFBSuIytDZHpV513bl5RlmWhGSDWYbJZkub+Szihr
xERTp6EgZzJH+HA0I5PXptBei7YxJWtwe7Uv3kunb0ApZyWYrxWRQ8BrB1mtKreadPAo5Ma5k5fc
fRt1sm7/Vg7aa5IxQYiepsLFpjBgt4WhiMphioXTAuiyxIPEpgQswCWLnYKtNGNAypkn/cHzv1zz
hGREwLLF6Nwo58EIqsvVT/n3pgyvjkeKLFD/BoAJbn9YPpzRAoLVExo2co4pwcX+/nvuCVGaTEPM
DF7ZH3/VWmZ01K7zzV3a//Q+ZoiwQ93zieie7hW4K2qjg0t0Rke5LHLl4vElPSLK7b3hWkvIoWbH
Qo9NqDK6LZydGxySScVz+R+8W+/PIy2OXFQVRD5SE3rm0HpXojI6dlpeoRFE1V+ZOjXB1OlJTtd/
8U6F0yAe+kAKIesPm2FS2Jivm2Ioqaxg66n82jGnekl9FYlBi5ORmDZKQzrXNONoNxiidoi95i4J
VX4Nh74UwNbJY/6xo7Pl13obqzuSeqZfrX5uaxUZnX2ttRUpUe4DZUghMx4wK4iCafsYniyCP48K
D/0kkeTUuFKAvlrZBORcdUM2NvhXVQ71r8BLpUFiXtbLpRDj4vZMZJBNKkbX2lQ06NsAxhYYBy79
x1a80kuZtv6Wwmt+lOqBadTUqhN5w4m8xB9tw+NFn42AIJUC7WBHvWsWHoiARutfo8KakVjYxc30
D8sR7Sbr0eAD48LRgAgkxX/qmzLExq0KKST4ZDTLPVUy8eDVei5Q5vhN2KbxpWf3EDo8a+bHogTX
kuhXZx1v3blsgZOsjyRjAZKaJxulhEbcWSZ5vnCkLfH0T1hXcAolxxVhECSfDdTHFp4GDTpbq6E9
mf+qm1SCgpctGXRvlyQRpCr2VlpPPCdvwYFGACyVIKLMBcmE7DbZX4zH0uulJHPVHf4sK7ogS5lw
XH+vAKpCtL+QynwhdGIfbRSjl/6cR58H3blOTQG2kobP4u/Xu3lJlH/uKB3OD9RU9DwHuZljOgG/
Wd3tGVA4in0Iwy5bD+Pp/OozMP2KQLhAJBmkO7EVaGU6Hr3gOm1a8jFqRjzW8ZAfGV0touMZTIQ3
06gekAL2WxicSBYeI3nIh9/PfXgs4G2eZXXE5OYsCKIqLeDMUzotGEi4P/IaUmPA0KKYhdZz+TUS
bdDTyGhWJNGf6ug/EwqgJJUafo+5pPvXw6wgZTx/AJRWTOzqAKSIwmyqf/HFnZq+8Pj+ewFSa3kT
bam9/WxGeulOcPGScikJitHDUts66wT6qXluwGJ2PGftPpCa+0zAq6sOLJROD1LVfOaOYqOJ6cGr
ASexJw8Qn5sgK5z+HsjQ9HgSfOyYDx+zyVr5qcDfeT3Ki39GQ+/VldyiuSVDlK1+VEx5xYo2Zyk0
fKTSKHfzsRPX44Dv4ty5hE7NDkNpOncx5aI6cEi3Z+Z7hdWZGHD3LNb1Iz3F+eGpJS3iPirxNQ9+
0vgSwu1DH9kRLRUyQKBq8juQfwfFEyUv1q+bsZaE0V8lbmifl7Ik6cKzPcHCGbhqMBSGXhvE42fd
BC59ldGzL0jlf9dUX2DPbynmrocfS0FT1oGzJ1U/BK7e/0IrqilKx3ukYu1KikWCY3G/aX8sPDrS
Fc8/o2TViMWbKOftB9SUu6sHg0nIzn1Pivpt5IaJh3jtEEXXoYqkxFPjXGcmXaAHLiyDT27QPk/7
kZsKVtx7Yl6qjTlnEWOAZDbmHLzIMBgi5PeDxtJXDN6JxVtFA1dYFjpO0KXAsJtfNln6tIPTUaQ6
RuTOZpsm3trLISd/6/m6AsXKcUdbIRLGtIgZO53HRECAMQcXc+17mIwUoVcUYL1neo2sKDfuPdv1
xtLGN4aa7x2G52NkIcZIiK1y+vUCVWD5XwBTKOgSsSeNU1rEwzOsN+4TaOi5iyTmds5aJ67deSKq
O8dstv++lXG4p9HWs2UpscIyA3xV9rqwGrXDuZcDZd9eGJ2p9uInyCSzb61c4ZIgXxoi3fPNa5D9
OvvRy9Ylf/ZTmcTvQxVGKQ7R6jwcxrzPa99bwSjZx87dxsKZfpmnGoGB2zf1fDzxp9RwdQRTZ/6/
LVAXee6khuMAOj+FSLSraKOWBo4ZqyVp4aRB/Od+xqC16Y8TObNCK928qYLrDnpOTiSRgeoNCl7f
x0/uig3Zi6iLV3zbzEnCpMQ0plVjWKVlvmMvpxa3kKtdsObW6WYzUhYgmuAG6QnakwXF8J5MpOrb
fjtnwTWlbPkfg3yoYNvNWTdkIrQgF17xUb27BwpfSMj1EzhPu3/IP/kAwyvcs+2Vm/el4RgIfgXU
d7uZMcLV0b+A6l6pwTF6TratPajZZBtbu10Oy86ubzF6PwqtUfCWvN4JyZixUsCGQI2NW6qREkiO
JyyWx4hSB3nOsTAtl/6FlBdKS56PXNcwnw89FcUiirg7cMAAFOgR80UN0VnTzwrBvRxpr/Ix+b+Q
6atdAeyfdQkUFeIvnAtMOEgLxqpZTD7SHJUiUTGSv4IXb4i7rKy0pdxy6aG1+ppGIVA5D3/6attc
9RgmMamItO04LB3BXe5vYz5eDp98CF1HTyDj/mse6o91gtSOn7y5etJJNA6xVZqtYFnzdMSH/SAH
U3Y1TaZ8vEaNXxdFQnrczWcun7tBUnV61BeDOiOKlv2ZvmhTZhLtaxs/Pj04M7r/cf/Rm0+b3FiD
z12sh36ycFarOKIsF7WKnjgPNotoEwQ/uKZPqCj78rdfKstzrbbXtJRnbQKDVAjrVdUWhX2lh6TB
a7tZw/dDxpgiLp7UxUzbQuivGU7zts8qcuhKiVauxyYaf/D2copfZR2Ha2fJ3ZoAUeaVDPGrsUkG
alvzm6Gq0BbHYHaM9m3JQQoz2FM4bZRDZcrtnjUZBx1MkSI+OB7r5+3lOh75W3u4uQOkSK0gGFal
jElfKSgjH1ZrNoHcNlXCT/BrG7PZvF/uiokW8Du+snb97cR3G/64FT4V9F1p3GeNUOi1QmU7gAsX
RR3a3mur6NqrJnrrBHKkKSdSL2X1ifzyTPl2ri486rY0d9Mu8YJ4XGMWYxwUuQCrK2oFkYq95ptt
pOXNOHrhe1Y5BtexbI2FtUMB3AdBvEnNFWiK8Um1s3QsghAs1p/oLgHQFkzxIHdpjZEdyG1qNOOe
0Ov91bhwmtBprZ6iWG2Y1H1OyMoc2SugyyWCrl0BIl1tXIptUjX31sHmpZi9AZHRWwwHQQyJA0qT
ZbM4QI3kwbe9N0MB3yqgw4e6xOGrga/he3IIpx2RV1IWqz5JAdPNmq8HOuR6Zk1eEg2NMmiN36qb
vl+kwmvs/2jesHl+clcZ6Y/SZoXFioWcjXyqDAzT+DXevhClaYlByR77ED5rjN7/nJb2abod7z5p
xBL7Dis/kojgew8TSuZAv8bfoMOxhMrEKy/yXgPaX9gzp/6NPEvFO8odD3RwsWwmjcocMbGTZGQn
O9HJAY6nt1DXEFzKsrFHhhrfIFi7WNgA7lFDWd5d9Gjt+V3tHDb+Cd2LyOAWRRkvRlRxoqH8RWij
45qUGR6u4h0vjyThVHxiW/N4RH4RPHqwOawPdKoZMJQ1oJtPV2I2NmYPkpg2B55RdIUcB7owmVcf
f/Rld4NjI4pQuBXotSwC7brTAdQycArSzeMN+aYS26Cv073IF06dvz/m56To1ajIBrM6zbxAzwnr
LLNUex42Mk5aqqTxHU2pcDN+kRVBORQ9midNnpUF7ImExsSI+puBiECs2cvxnVRJ36mp0X6H+7Oa
nvEvnTI+DtWfhpW9aQa1AKOm3uZ1dWdNknPC4mSWA1XbFh4yI9EWEzv/KfLibZmxTTf1kDkBODQQ
tyzzxFLc+M+e29RpqpCtVB84FQuyEGiY1NTGo682u7NFxDl0sXBIPLNT0K6fC5UdJ32BYCMI6+WL
r8wId7+WF6SiwV7N1lqDyZ4bH2A3lkGOOUMIT3IPmYsq2LNd6c7nihC2rcjvK9gjjUWpWjgVTcWb
1Is3NKdYhHfpr6z3MIqCDq/zoSZSkY4pbCvZJ0XYJjgKyWVlFpCzhghIaUld9fq6gWlmNZ+N4PTC
4ELa/Wq0Kdts4HKMExQBN7MrD06gOXel1YeERZtcCsD24UXDJR4uMZzH9KQ0MSD5id11vqMu4VzD
lt9XTfJUmLrM6moNAINL4i80TGAP3hH1CqX/cprvd2G0nmPls2lVy0ekMqqvIma7z1UGwei9CIDy
hbpo14aeubzdD/8EwdQzjk2rGjJ8r99YQbqW1MRv3TJjarXs9hoUewCySfFLQn0f6d+9jhZUcW+9
EO53a3PKvV9XLUgb6Nfi10PIQ4CyDzr5mKWsElVkvw13HQGTV4QPPH+4M8P4/fC3LrTnT15ewyju
dZyvSf7lhv8uzFynOxXiH1wg11oVJi5/5700o/dr8eF1VQVihnn2zkU1FjM8TgTv7oMrsaPYEAyB
VgAR3QaK4+HRfzJpO9ePvaTslcaz0KSdRh9osm18RFBnz77WjZc4iOAEr8ND0E/w3Ps99Du8N13Z
l5XUImlvjRQJQyLj88Vati6Goe5/9VKdL0Ug+yKs86rOCtX0nCmCr60gWi/gIywRK5Gt7YgqE+mh
XUNoNER8R+OefNEkfvB13++Yvb5UaVnvgkkz8hXRSFHuYSM9D26/WdNoHWnMxa1DQqyJv9nYWdFY
+xWjcVNs5va3y3o23Ga1eydCbajdeJ0VFtmEI7N/hz9sIxc0dRdf77j915Jy9US4Z5m9WVOsSaM8
fcXTAItHyYYxU14UAjvudF2shaDPfgaKoxsVm1bEkJhEKqw5z2nSPm8/wpRighLkfDKP9rXP7zvn
jzVZd/rSMdW6x1LBSPrb1TDiGiigJmFaQBRQHn8L93e+f29MZ8BzSct18dpM8JEpZ/XZp7VYdfKh
gxGeblv1FaYogefJBouXC4nOwfOjeDUT9YNLVlyBXibNf3Gx3ewcezS8ByvpzD7YdfMEWVoAsQSA
R1ABYS5d6ZbE9FKgILzYBwBaummcbWYbA0J3NcbWq5jz10k/L91U6HVi0PMHXBVQrfT/1Mv9oXLh
/NOLDDQgsrdjB0v64SAwjbttD52LpX1ei7FMbwTkPUfZZuoCSZp7Md4cfCdRCX/Xr4mMT/+czglb
pBzatYOY0LC8LG5LfHgBsmu2lPxQIPCqkFjpKBOnRe04W2swT6oM3oGd2Y80vwZ92h67eb0wgKVM
YNcFDMLO7iy2eBGPT2BncdaXBgYJYXMPf35TTPRNXOo8qDzJ50GJ6LfYpIbe9TmD+tSIkw8u+2o2
3AbyXsQ+qwjbPGF3Bve3M2SjiFfdp+DfgxhX0pZ+nvffRF8Fqg7JAu6n103i3BTciZ3NsbSuGmcj
PsPQQGI9Oeg8cWTRPoancAVJju0BSQVZYC0sr66kSRnReZx2ypTn8B4J4HpjwiJiHK+54ybJv/hA
ieKS/XC8is2dSp/Cpb8e3zjRiDOexhGSuMMqrFoXfkaoror1NZsgajbbI4UyxAwaPm8y1WzOGCIt
QZWfCZtdZide9lF4u+a09ojJ6FX0b7qIRYPyg0paAx6TPnoX6lgA1GKVPWx5n4ZPKOcos7b22ngj
JwEtLIM1aXHJ8sp6zxdoFWIRcI+uAaBNiRvrtJwzP23CypuNy2G9rueFuHVdK+u/ja6Dpua1wZkU
tDs7IePGpM5xAWz0GIOD0RXjH0vOUtlgZxk3aLXHxQYy2HZ3BvGvDVtlTb703ZYtd1Vux/vhSIzR
jmO+St1lCCddHWstoDQ5eKC5M9Ezk9DLIRmNs8p/YYLAJchqL3dHTjNRAjpICRq6XgeaknUpmAzW
3JjeEB13wLKri8SB/86uzdwz6bDkU5U6jCebWeOyMp87GpKSzW0BeRZk31zN52AzeT6wMxclykMS
vDP+3r0yR4OnMdHy1ct/wRl+0guQVUATlv9UcoeA5Pxod8N8w6dqVrUkVhKeEDR8ee12/1BoTptz
KsYqbhl+lOrz7Pm/XPrjx9J5Cz+qRNOBC/wg3HzyaINGkfjH9ITavuWFsREKOXOs8NHbDWLrAXQe
KMr+/1ZAcVmdd7kdgAeiSi8s5thG6VLTGIpnGGuEdaQHuKmeOYd5/o/UgNOJBBjyteV793ZAXY4C
p454uaVJFPh08cfmKjN+E1BPZuFison2N2cS46fon++Z1FTZKZYy9Ig3OcOYcYoqE0A9RaDT5urT
ZSlY7Li4W3qF64mpRaQv/R7zShimjtTdCz46F5c/I4vwRVAU4YFGTgA6ZBOOkMMUhxUfRuhmMSsk
5O5nC6tLVcwQe7o3wlUZPgqapKJ+qYJIXWnnfdZILFY8Bkz71mRFXz3Uth5v8UFD+NrWQZZe+P+W
p430ojy4naGDrvcfQPXV1+F4rflMV8blcjQU8omhysQ7ku6lVC67Gf2FRwe+feo9nTqv9+uePuCd
LoSuPbNwa337BrTQipo6T9F23XtNGtA2cn1Zeif7y9Boqi2fC1hRX0BlmI4nwZ1MWv4+s5UKpdx4
puDxDPTao989G8+WVEcWmc9NXEQxod/T+cHmFbh0xzrkHnnGA9zNYVRH/2am2153/m0zuZV72u4t
/BDMIWKvjr+XcAidfNyqASxsBF5CaItCkRFwBhF022uUTMX5ZKEiAp2y6VHACYt69kFyXAHD6BnZ
pLz1Mg+3rWHsRmD9UVzB5jtb1uPFTfItpyg5O9FOR5JOI4p3b6J2A9q8vOnFffaB5Hm7GYUjr7pq
REDMJulwVBt+pdMgx/0jxgFqoNGUEoRRVKpdPfJRGSFKmkGED9hmUscQwdZISz+RJLqfck98dC4Y
1UDJt29D68YHPl2Ocb2z2tlU3aGxZbjX4auL4f6XXqQl7//LrcPteBb10N6gdNcnUmdAKi6Tys1z
OhM84E3V8nSGQsZnioCTpATR/M8q1dfhOFIKIvZWvXEfbHVn+ziNXpK38HhaPzqad5X3loPX2fev
ZfoYz7WZvAsIxmkXwjgnQ/Jf5Wn+NsX5WfpINOpebPoD5KDu9wn10cJLTJl0ElykxIjERdEMQdFd
LhtyKfq0tluCHjVpHLl/wQ4CaxNNn/Xltk/j6JVOiXLPTK14+uZ6Zfe0hmApgB4uJp8V2yErmN37
MBp8MppKn8nv7GG16I6zQFaL7FXkZzgIpcUyCLxFsXsIQM0sW+54pK7jnFtqaxXBBCosN1tWAmm0
sNE5IivTgwRONLz2BLANsyB0W8XE/11KxH/RgdQ7sVdeehWQyx/LMGXKmBti3FCcJXnslqFrpRvs
LPTKqrwmlbfM3oOH6wBj0LxM5xYq9Nc4pSAORgtluLbEAX0nHItpr6tO55pXjx5XA7FCxJBM5nOS
NOl0YYj+/KqaTX7nhpCYcGeLKk22U7dDVQASKYmrwS7fDO9HBKXia3zSV9bZ34rZ8e0clNbKO/wE
za5/MnFO/Ke2eRmqrCRLCwxplYYS67hmZQokQe8c0NxvUK9ZR8wVIshe3o8RvIHEWCRbRmF6GH1J
RfXGPmJF+GUV1LwcY3aOi5R3zSCvf9SflZTUaxc0WJooqx33mR3JOHQCFlStlqiPogknDvUJhIEn
K9SnaAaXSjco/vOCLM+wQTa2ODmjiiEhD2N4axiEFqzCjqzWCt6rNYLTgTCHWlvn9Ojk7r0AaDNP
p7pOVLWMvZOOZOOkM1RJ9G3uLxJu7e6jKwPFxgziofh+5OEPwp9SP4sseccm8wUiaVqWKX+q9w0Y
jjQH6a90/djqU/AB6TRaDNNMFldsnjD6rCakEoay7QZloIVz/Art3z6GULvtCB3vwzoD6O+NswIW
f4ivm4YswQRJlWg4cdvtv3hXADlPm7VT+v/2c0Tc5CJEQJmzfaZKsY11iRucBLhTLjf1KVuR5jbr
5bjKrMmWy4NocOpBGHinQavXnRwNbsxPec9yF5R9i6Kpf5/5HR8qGtXAnsXD6nBiqL5dNaZcodUt
Prn7/Da3SsuZY+QfWtaaAbOBkdCXXFN+VWb/bNt3wW+g07f3MwOUe/UHQuff8k1hMoZVDF31wU0A
ua7xG6eyeiBKrxWWRxFwumRIbcUM3u9PzlNBAXkKZOOVYPKsBBrHQcORS/wltu06dtvHBH9s+YIV
bgnSIObVvEBkgjtvnJLeZaeuv7MymBswzLaZRenw9pOlVN1V9b09w2vbEpDlQMIMwfgYmh+AVnKU
lBpR8iaERikKSKu027wxswp/iKDkkArgfZIhLn2UIclyKiA2KrqsSu1yzHxUjWovMhEk/tqPbYOy
LGcSIlPLSfImlDHEp5KvvxtZeLDi4f0GhWz1JNHn4HDG80jFHTg+CTHFo9FMUCwedkvCpjomzOk1
Hn+Phy/EZ5qQk5zLC9aqw1PDPmaLuKx+qQQEtXsTejmC8/DWGz9ka4WmfAJjrJRwcrAg1wqp5RlZ
FsqFlg3KDDuliHFXj86Y+FB7bRm2BePxgiOSuxmIMQ8BmEeroqKK46Nu/ZKHXo+QWzB2nA2sNKMs
7KfjxZ3b3VsPSSkeQz/9mBYgHLi+GZbI0Zm7/OOgxFI4Hp4uWCLFkLnLP9sHXAePxEQcCRQL78aX
sHPKgJNnGpoVms+PlwoMFOmDcJ2ib95q5EAZ42TzHDaFHRAOWg33I3SRUDfrGxUpCrF1jKcrPBXs
l3Gp6eriq8N4dpHz9qLOqDCrkXm8t0HFQK0DfN3sjXu9MhNXGR0ddEjFPJog5OPWatBvL64iQ4fM
sd1etWfHJwfDDsYdZ7Bdu1S5+CSPvj9SjLdeZ8LZgL9OsRo6rdmfHkO/e+MixuwY8yiPWOuXXzEd
LUCOFS2Fsf86Fsl5r9zM0GU9VtJA3eqEvZdTBtSd4XbXh/nUxbURHnJWCy92kNd14SMcvE+IaMEZ
esb+jEBLqg00uhDepmUSWJZ4Oirq3TKixV2/NR0ZyOuifERSxXTy5IpU4I/Mw9iqdUVm8Ao5IyZb
YPEPWU+SutIM0BFoFDIfXquJBhm3AEI1gjU5E8eiU/XWl30vsS4ibHcUqd/6MY9Qj0aGBVK0L/zy
I7Sg8aAe9CPJKv+yTUL8ql2eM7x3/4n2hyRSEgw/tV+4GXbXWZMvKRuGpSyK6yPzdzpJZg2zECCY
CVPiqEY7DleLvl+UEFCtUxURwlc7rk6pBgFCYaGIzPY5ZNkExVz8b7vshRrm8oV1vcfvz4dnNPzH
5hj8RUijY4bu+sZbOcWL4wVptERYz3nDmpuNqOLt8izDpwDilq6NfdGb3GHJgDB8bcPpeU/3xvX4
3w1zFchtSHQw9mcICDgck5Ln1SFjpyYCxIanpkOpZttthxUKXuX/30Emy90oncGhJNLXblNdsGgY
aosobAXAg1HN0aDNUlLetFt5fGptzvfmxvSXuiFXqTYz4tluNnYiFkymObU/V07NMZiusgajDQcK
YA6ehE5aqSTMTOk7KuslNfdJVlNrILUak+YxIzJO0V4pLKzzKt3e9wYAkiMNmmq97+26bfqo+1IN
wLyTNI9KmjNXKspeVDLIOS1dB7pxIdn/fbKaJ3MBf8dL0A3U1SuxVc5ZQQcc6F6lAHzDRwHUx76p
vw2qWqm4faJdoiFFv6lXcPNH+ntzhwY7i7XYPBOhY8BvsUPPlWMNyR+eFm3IqpshIlqIwb40IVI1
myvvX90ULg+390jBFH8Jm7aA2pWeR6tgZWlMMJGevxjX9u+WPwIF5MhzgJ6ANQ5IgleDvuXSqtm1
bRAi7YwPZU3NRkmOkVirsBHOEWHAQh+CXV7la0gZaHpNtWdE503JTXprG2BwU6XscijQwnVp1VTi
npLMvWFYibgy7acEXsy4tP5ZWHMPerS7jhD4npduQFDAAw+5WrC5TiuJ4N+rBVV0SFSIB+k1pVWZ
5/XXj9PNBUGIY64dgVETDzXPfKO86CPvweRA2pwIJtQ69nQpzhWCw+OROBUcpwIN7C+Gd9aJ5ElY
yz5T+8xM76E6ZMHK8PPwI7wCzy+mgpHquMV7++9aZeuGoZm2eAwhPZxcI23ZGkFyfXCUV1vglrzC
3FfwNdUHE/nSDawP5Gm4VzB2TGpNFjJ+oBSKWNUoeqWHpaghSVjrEsVSggOIZ/ZdjcdoeStAu7G3
kDht4uN+zGqWJNdPOx9M7/pf8Ed+mo8G0+JcS04DqoBvX9gtjvWLFXXG45Fnf6aKqB/NSTfZkFf1
ghx6iHXiOdMYNikv9pnxukTB7Nuj0gkqpux28Jzh4Z9xt/vwfSj96A1yQSR5bjTQY6mLVmMNvdD6
LKd/ixEvNuXCKqfWBEtQUd1F/l4aniyLxGSYJkeC2/aMcXOXfatKRdSQewwAyqk+bZetJDOeuvlP
n72IgVL0OTXxI5W2NlTcAQycWoelbkaJj7/lBJxmT9J+JFkl2FBNWrdoQCc/uNkS5nMIX2EpDEn5
WB4dbNtjnpHQr6K5iK4nxrIHuyCpeXALAdOY25TaHtfyXWvIKehN4gsXz7X+acia/8SkCf57DeJj
bzHb+heo68beAR1P3AGSePvlkrLRQmoxfpRCkbGc/DTRHiT2UsmRcQ+js0ARUj7HC1O+8qXtuJ7H
0dCtgGuMXGN94TO2m6qAdfBOIndZFgT5Njsj0ZtyTcww5gPDLKDxGrZFi8fw7vqYB1Rlh4eVl6Eh
FlPJRUpHX3Z1LHSJzbKweTvft3MQ7WAZA+17NZN8bNpRoMsWtVD6Xo4N7DWJAn8qxxf0k/ifMgIf
W+kIaW2h62MKg+n172SHgl/60vAREqxvz5t3nURXCLJbrIBfOjwiwIHOangKFN7QgsgTK03hN9df
QDuwdDHOo5q7ryDPvk8VFGiyltqjagHMNSOoGNrhYnpUepjUYVDGvxLYj91P6NY40DBG/TGlbxT5
hPOVydclt7+JNZnHSRdTnHgpPmwfXu1ZTx7USD2ON4gt1jA1YQMsAz26033mYkS+KJVaT/fmF5MS
iJ3m2EgJoWNOy/q4K8PcMs0zgGKMElCjpz4xYD6c9TzEJxB8DolvuDRjyx+R0Mh2aaThEdS9impb
LMX7MnOC8YGYgyCVwGF9DIRyZsrGDnqbPcE/ecWRfElvXJhhfysLFggKU6ZV5GJJV+cVjAUufone
YByU7JGv903KznCIf6eNpEFPxXfCXd3P/1R00MtVR0EzoetQqBxRteIdOudwB+rtFY2bDstHqgVC
J0qXJBte4gYG3OdblxwEMSHeijyTLfwuXGZ/sHEEI2YcQgxweT5Gs8LWqlurCuCmYAyKTOUEvJrd
akJBxl2jrs4tRXs21VttZi0bxaVCIdfciLELxempX9qB+tl6KGvYIZG9ErDAkTaVztg96D5sYZfO
qtz4xOsL0mgnF3AnBRxH7w/neH8j8bzpSMq/gDvcPDT63/FhywWsYs8zlamozvkuIkriLVRv/YrX
1a0HgO+oyryxrvgBCKPeRaSHE/yxMUS8JOLprDvEh6ELgrLngJQ191VhsRvvqpv1/y/cQx8b+fes
46MDfb+NSyxxJ9ugS47bQgCX7HKsqlpAaNszo6nGcmcLyCnJMTC72Slm9iup3665pMiErW+6n6vT
7f6U7Bw6iMeO1eMKnAfzu7A/9Oyi0nl3M1VQrhzRb7MALtYGFHmX5yUhKiVhEnUOI//rrQ27srlM
wJYsLEaXZzzPAfZCd4aIZkf8kq8IQabw5Fxo3eLObaYxLdtpTAs7AjPa3AZv8B/tBKy6EpIDLsNY
mnEJsxOypn2v3Mt6XiymCLuxO5bLOwQckxKNG4rksVgOV2M6gSYucxGupcqB5b3glIVYPvEsMv3x
zpnBx3IOZozVhWJWjvKxOs02AWr8sbK5cMrIx6fKksFweaZvxEakpEUpyrfNPgQrrzZQAGxcGIrX
9Q1tN+mRGH8fCtOJT41HknXdhxSzFMdm0DTKKN+PlxbU16hS2STqoHmVuJXrdtleoeELE63MCTs1
2BrCLQc4f+y5TtRL/xQy5rXorAae5GXN1Q0wiSk9hM3Mq0jEyv9fbtMjIyQfxel0XfB1McrbxcXO
zSLCyf8253PZ6tzp/PFykbN3ZXvx17rT9jfaHiNVQbNulIwNXlGLdyTBPCtW0GGx5RLwjp1uLuFd
D2UGR25BrkMV+v31Ih7MLgb0XHF+4KWN05A9VDV+bj9elhqsFCbFwS1AUSMNrzqw1Uiu2ECKYRfN
H5npMlBnC1tpiWw1xuBmvhN9ONoB/BH13aAQSDYm/DwXTEmG24cxHjlSb/Vvm/mqnJ28VsSkJHjA
U2d/oR1TLWkknfdBdPbbMPg/aT0Or4WunZ+bO7+bUKbpd4hzer7AGXPjVqSL/xnJYPRwbyBdqFSN
82jbczENcpY1SufWWGFFsZ+eeZEH62UlELilmdAW25vRztoBw/K/R1F2/KZg1J3UrsS5gIckUHjp
HV4QZmpq8QoS2nHXWI4YMO5OcKcq4FJL/mRvIG59thBT5wLFIDpPef9BcCjKfIN/UomoRr1CVcb6
aOGhT8Pld1wa6BouEbcbAYXNtsoRseNOlAl+IxxkaTyG03SWqXYFd3/uLCKh2AkmAsmH8Bt2y4IJ
TI9NKktTse0tyReDDmOWtL48m1AZsZX8QxNHPMRLg9bhb3hBLUX9Y83vMwZPTlAOsI2xdd5N9+7g
N7AOQpkmn/fxf/l5tGoVEPE5DZ+LgjhwxXVZ6YPYiO7OmjzbqVaN6QMaAPMv1p5flBR9YgSXp05W
zcrIFCJ54Ff+ibFzGhhdJ+oCVLX24ooz8s74JGNh/GGDIIKe6EVD20XfLCC8okhHc2knf2+Hthjh
jYGXnMImm9XSeYSqSE8vaNaKBGbKQNObJA2NAcCFygEF9N/bpsMPtl3NxDt2s/ae4zQ7hQpTDLA6
xDBtF6aAHH4Ozz2piJIbvT0mnUtMBMfX+b9MUmFTTWVxfs/K7fIXFLDuJmCfEqWbFCTDrNQLY8q5
6lAwlrlkp7R7UmxhZ/4VOF094QSfbAB/zTsi6hFeofHSNhZjnBjd0WylU+1srfpj6sZLSA2JdsBk
zhz+1I8TQyR23qwNHkZM6NOsNEdyKnBo6v7HDdnL6wmuNLHlJbFPF757SDhxguaGtKvGeYTyqkit
6C5KWv71n3BCUm+DNSLsSPYB/OuDjVc1SOlcMobtxx8GnAb6S9B2NALhe2agM9fnYTXt9tbxpBfz
ryCopsd5SNOSC56ALrERhPsVvTC4c3t0UXAnZNLHvtnHuKd+1JGX71kDnP2DTduUWNpwoy7MtTth
sbIzh2Pe/GoJiTxAOUL9BqSFskQpnI1iyrZPlcvX2/Rw/BMReJYAv+yE5NtVG5U98iLoIhoSfiRn
tsQtwNx6pQDs0ct+v87Kxaqq57NGs5mRC+6tOchXKiEnDmuEYMxxnJ4W8jWtjrjXqBmJwO39u5x/
kQMAy0Hqjy961eRjiYtonG+yLN+JVt6yjpbqEB8XV8iuoX60JVLN2JEi6hKQlLgyhsnwodotH7X2
Q3MM4XiAbI7tryRw7iaunensvFSL3LIOLiT/pzCSWdqi8023NmVVxu5uxueGuiuLA7a/0FtLoh93
CgsiEYq6AssG/G2xPzlNrnlHZewUmtkCy/fG0VtgK5UHEd6rjMtYqDlL6+7bzZLWQYd+oR/lNOLY
ukKjg+izA7G55EoEdZoEtXpnxXRWWNxIAF7+Nid0NQE8lcfQEiek2csS9Q6NqeMnBKV6vxr8pWeT
zTrUelTqGjjMm44Jm7s0kUR1Dv3qSVdn0WWgARlevanFrTbxtBlyMa46/CKGUIBnpXcRHWNI3VjK
YZ/LIBw1Y2Q3uwXF/LzmfMvhwOP5o5CdKAGdGBBLIVFqVSC35xfl7bPpxKu51WWsTgvWWpo/eEsM
0pE37AGp0/7ZuDZJQFQuSBnelQ7zgpAd7iHWg72ZdQSnL8sSqW4+rw8yCr+Kj8bZy0IYWapc10lD
9UqWtyiOzGkeGsySKLuA3Y/PI8r7Ai/x0t+wN0T8MYH+gN6ypy8Hcn6GW+XNHEkS5NFtLpFCYDD3
6hAmvqT32wgk04z2Dau0ETnTi9Nhqd+O/0dm1RadrptkKZ/Nn0gHzJYFfqt+M1lIqD53rRMsDNOK
W+RCQA265DPGnof5mY2Wy0Fc2QOTOi/lhe63p7fkqhDVtWeMDKuEr/HwZ1geyFvb2VA6lvgd410N
wpfbTx0Y7lkQqZgPktwVEQWsZVHmeptSFiIRCJMSLrlkwsH9bP8iX05sVGwkP5ECA2IeD4owtsx1
SFeq+oDVi0Ua6xKo45VIG3fXSx6Om/q0lw2LyK4a1bLAHgKxHjLcRTRuDTYn5NqwTyY2UcMeDK5M
PK7rxrCNR45HtD2mDguY9dIAj1V6wq9XQsHnjQnDOPrCou/NXk8ZffMwJKMZ2KrzDp0sNvvHjLAa
scnG+DYp8zkFbAhTkhunfE3EAphEvB+79RL1/BggW4uwyCYsQO4NYYBITgNse14H5KQkbJj5Os+y
N+zpst4lnGCETNaWa/hC7TBBXCQ4sbixZ5SSA1K1V6gTnVvalIIF09mfA29OcBcArkq93Jky8QCt
f2RfTooVpF8vO2wEA0ayhqV6dve2gy3KbzE3JKPuCevxsGmkbkysG+4CL8ozl6dvBhGa2mkWVeaP
nDf7tChTo+4E/Sps5JYUyn+RHNQis+d1yesQ+gAae5oxAbthT3/i3+qom0L2ciAjqTJrD7LjlIVH
jQHHiVJJfxqNpLJkk4fihgqWUYnwzOvUfrYHHkdmJvta6NysUrAhafwQAcEAQfcklcfCSUEClx8+
sIgWyxlnm+EOxnwzcpXkNchKoRjvWEOqM0tsVq4PQSkvtd67PDh3FT8NRTXJEsw66BtwGuTek6QZ
/3pEYnvNI0KwGzToflj499PnDzXr7ZjLwIH8pPXJrCGytpnN/blgR1F6H2surwpKFSS98r3D1URO
UxrKvdXomTn3SGmn2WS8DdD1bbq0pknc+0+lv6uQFOhiGf3dz3TpH9HQfo7T4HqwunncZCYnxDyi
DnSBlWNG7gBWpIjXN8ZAGs1GeU87j4Ru3T0zJpi/q1i9PJFVmcqLHSzcnJhJb1EI+G6nuM+aZWvS
Xa1/TLXESMInsgdd179OPpugP6qGqRUDH74Mh5F9xMTRw3ccXOO0bNA8rvG7AOmtwmIcvm+bmREw
Gx0hE/OlvnibHmtQm0fJfoFUX25XcjyT7z9XAt0YjPAjNu5Ok10I/8kdXnxjQ606esgTayravMV/
BJQTnw8YYY2izHgK1xsK3H9rX1bg3vDT2iMwEgsQ4EWSo/2oVq77rNf7PxCd+bjL6zUZ9u6SIuBv
fNh5Hv7VZzh+a36iYnt8Q7Kft1Lm6/7S9moqgDAMXMk3emy2Qj9gH4jWyJPlL6lEMMcDDmXHeG9V
myqKV6nk07oTTW1E3YBXSZApUla+T7Gd4x0qfLXKxsYPoGLf72k00zAjcWCO47zQ4EhDG9qu9OEr
p1+n1xPVMehNkqpifLxhXBID1S2oZyPCXNQmui87rHGumZu9hke19jueINGm7AbcO4JT5rUMld94
xjxzWzBBOd+bfZqgCs2uB0ctoGsiBEgyOLUrcolsmRoNODcAokkMkm751HDw7hRGEbd1nhQvtR2+
NKGBWZg+nJDqJtYB0nhF+Kde9GPg6YNeg5WBVvJfXjjRy/Hgs8gIzGxL8Il3EZJjKZm3ObGHJr3V
Iol5CYaJmGaRxUjcGhfYSwQ3XRiSInMTO+VxOU5WybVjMx+ecFv2N8zuzt007WCxSDI+fPPA/IN3
n795nIBI8YYevlMXkU3wQy80bTLRkGc/sMzXYyF+nehLh2BJ7HaqfsZti40v0b+2/Zn/GJybMlSm
XiPoZauAzHFCaa2DuhEms/LzV/Q+I1bZkBfWyF3tkFdYpHz3o/3hCnyFNgeM6SNMwtiJvsijp/4x
9giP976jaGVeY/HpgVwJJeS6UwxSWHMYcZPmfhGmhKuxGi+prPT4ldR4069reIBrNlKjYFa8oW3S
dc6nAqt9LU7OZFfXn7stsyRswyl1n9vn+JLaIbqbOXFhI3djhDiYQ0laqvNbbcrVoKvXDUx2GhBB
zmRLRiWxUUgo0u8qSSHeac1idF9H2C3nXY8k8S5lEVc7y7bMWesTDQ8mg1phb1V1zzH31dFhNRUE
6lqXhN80MfvIRmh7P2DYWLAZ90FQx1ilt+mL7fTqfZWjP17tHZTzO9DPcywvkSF+1eDfXY07M04l
lHgVCX+k8IWyOF6jxuN9acJOjU8CZAwpeXhbGVDMbfua943oYnhuIbpl7XQm34G3rKD2JrmkFATL
masM8+Kjn5u597xjKfVEF2m3B5YBZyQQjyp6O+9reCh3Cv8zkj6tDiJV3bQcUhdCMY5RE3ArFiKc
8Gw6V+e5WoZnfmk9VADg3iOOiSAoRJs0tL9/exxt7iM7h1UpGmAygoSIw42fMvFE4+M9rRAURElu
w3369cbD9egUsEkVkjedqUCr7968oFeurqqhOA33Jw2AFs/sgduL8vIwW92lS5rNJmbqk+fmuOCo
TkDkSxpO17eCRZ4QESuvrkxe7rzYFapigEa7At9vdG9kljqHeKoQoACSzGBWw6Nxr/OS3iBbLnzT
QibsWZ1tW3UuiBQ7fl/Bvfnk1qeDrAHfRGCaPe86DUeOKRax+eEdQtGqCUeTxS64xbmETGHoYTwr
SDoopw3bjUgPA27HjxmIxDz2FHWwLUcf+RgYoRE5MYsYUnSH7YA9PnB5LNP3rqyYj+vck+hfpVAZ
oRYjzqs9xSP5M5QcdOPY3C7L7Hym5Ovbj5JTVOxp74+clVzcDpuOWLoGmsZeMModwrw09nF1+Zu/
uCaOwdAwRPvrMjnVDjo2SkiK1l4LNOVEmpiMmQeDNsWiyoUyqPbfpEQXtiLRXrWw74oaqTIAjKNJ
E9ahU59gI40yoNjeGn+ZOgppOuylRB+i9dtYXBxHWoMOIc5B4lnamBAM+3YNuJQ+I/97LiBTioe3
+mP5hatAIEmB+FmS4Sy4RKpz9yrtlaZ+CoV9W+wNOhCW2NDYA4DECrshTnvABZ4OlYzCJC37/boF
DxO6kiIzEUvbaHd9Nb+5or3vhrwTnfmKgKrHuVZhHXK29ORZNpZIB9OdypiLKIR7NRLPeadtsHfP
Nm5rH1HBiMknOgRFnhj+ghRPiHem7gvijlTLlrqeYmNsx+TQY+p+uMzGxotMjM3/NPjs2QyOFASG
y0X1JY7su81p0s+NkgNBeYMR+mlSI9wY34KxErtoTyAfJSajQzaXbpPQ4qET3TwYhAqhtuY6ov23
j/oaK3v9oBakWvDarTxlLMBRkbypyUiEZ4/EPGHmOh0/khupf5NiJernD31Ma3snUT+bzZRp252w
vVm52qk3sl+sOCQbq74hPOePjrE55NOChN/RQPrKIPFXWnZ27z7xq+0j5fzaVOg6wsZYQ96Dopmp
83q/RirxkyIG4vy9wxQWaDYXIqKngc7fASYl8G+7gBpia3h+DvgoWZkAYHaMtRBjxuaJXdIpa4yG
daqTgNu0/mvVHSJRvYdjWNgsrWM97ePbtKGmrKIHxaF3zSdkECX6LTao8qxWsnMWxPudrcVlXKeQ
WCFb96SFSEU0wAJfkIeBojzgCrncQSUE4XCqJbf6K8hnvUOmpDHwQqmkVAttevuuEpC403hONkla
Rid3ZLz5bVnPsPsijTq/mfwHqrW8TNQJDYYhOVd+v9/0FNQ05BcWovY0gcEzBFcfo952SIaaJ6es
nFpViLdUGT7Z6+F3kwwJ2Kc4HukfskOp4VijMjtYOVLoPjU4b5NIsWXFDbXniwRdnbMeH7hp7LvA
eZmB78AVRRAvMl+XjsJrlRrdJ/KDaB8uRI8Tfg2PDKLR7ruzZw2g5O4wIDOPiOGPr7WPdj5LTTbj
gKaUcJzzSjGY8QJ2jDg072enq/NNgp64BtIoX6462uUe/TfJP5HtIXmKW0jaW6laV8WC29tnPAq8
1PMB8AZDvDdP+3gZyaVFKDtUAimeOeoV1MTr4usIrQ2rfNOVtmZP8SHPPKL8gfkq3VvUw8ClIpiD
x9mlOtOOLYRC67/A5+OHiPYNldCFXguQGjmYs2CGCr3Ow9oA6W9EgbMV0qAUqguSou+zlJ6jQ55W
N0JwlPkPJGhFXVRejAfi1BDCwUvyfqR/rSHt8IZ1/Ct3GVhH15Us6UvvZqXWnwvivWfpSBoTGXCl
7oqWpRoDQ9u/aLrv+qtn0nw+OO9kNz5SMiJXOocqvqJSG58Hlmfky+OSNd/W9jfGLRPKUsvufMOH
DklUkt6+F14+e3vQSzkSqoGqVdTFY8KrdmP78w5755HO6F909+ZPuLQK5fG8NxvkuLwkBKvHrFZY
Q9UDJ/gPcKJW2ue0H40tITbrd4W5YrdZhRnZ9AYvVaNExcGWv1b8qv6uo1uM3sJHpxU3Laekxlf5
N0eA7gy1a1lbNy1EZOv5gK5k3picr4UHEdnAnUw519UUoNDxLZzEcKVFrujBvRJo0hDX64TKUPdJ
X5CB8B8h3T9fusfq0A2WxuRrdZOClbb3fXCK8obdnQ4la72/XTeRaGee/8USWn1+O+y3Nz+PlZi+
/pJWyHz/z1jTgLiqYWPJ2oDrNpP+sxfE2Yak0pmavpZm+Ybf6iqBpI70g1N0XUVh28vMo58qtLCT
/fTn6DckIYrQ1aqn/kIIxWWAe3K4F2UGoQ1AEMx/Ed0Oagh5arDhOIvI/4s9/vKRFOvPUDxfqJMR
rr5m0lBhoHqA932wZQAsuC2E/A3sQDAn9H/YKpMQiAPdLsTov/UNxTeB22woXyNcOGKcqpqzjxNm
9AINm9vXhbEfixHfVHrvn9ByR0PC0g61epLb0sPrtVAlaW1/7qFCgT/qRE/djs7UzdrjeEyhQL80
ClslSm78YlQJRM/4ot+c8X3KOlZYWWMn5QNr+BWt0JdZTklyb3p2oQejdsZZBKHSKNaln+DJILyY
A4I3PUcZGEczmI34AHoE0AW3vI6bqMLu/5sOlnQQTYvy4Ahhat6x7AcJVssAV6G4ypcZcRNNme8L
jAv7j9Brmtsa2xolkVvcZIHto1Nv4ur+BY93r7j3BND0mJbc+NtsmTP2k5m0nGnQkmh4b0WYTEmi
QQwzcSBWXT1fVshqE/SEy/tUaHb5RRHJQeX5JL+UR+N0WL/asxKbgP+bjQPaZFmu9IcUIGJN69Ok
yJA3KKK0wq0JXgNUQRX2xJVdeLbC0Z0Kb+wP2sxw4TOImMzqbtJVnOmv3jaSWQvZyY+bVJ7Cnn5v
kBtQUXpXHbB48VWmTfefPWTLSJ3XUSm4OcIkxRh17/e2aX36gJAB/QBA2Lg+nCwmhkeyhZdHss13
8BZDt7RoOIRcc/LlFt0WKvj7zHP3Ym0gMJEUZla17la5ZGR4PqnFBnxq/xXL1RDHuUiq3wCEnesu
9SSg+cori9tE9AsOIXUBddn+upapPih5ZejLlVnFxTVPHY/NIZQPluH036NU0tfcMo5PEZJ0qvtI
BwxHNInZPmL7WxogCxfHaA3mMUcgWWMwn5wvAQJE1TJ4Jc06aD7RwbfRRioT+1AWGonj0acq4G4V
56v4GwWkrmMUCP0BnwadoGcsikAPeQl5scWHfF3IptOn4Hk99xIcK4aIMs68/T+uLkf5hK+hTpsQ
JVqbrYGX/lZ9HE8MQ5aDkrGfbInFau2WXyx1E1YxRnDgICsLjgpF5FnhYgCqVo0kSYpeI09GYl6F
gGahGUJ85bPZRQkTIPUfbgImZp7CCgytNCMdYNSnKiX/ahvN+V6Qa2bvtuQeJE33Um/9XEAaxwJu
8Tt4qXEWx0QjPLOoFxAK7dXWJlIfq2g1NW6gNQXoU3N4UZvzaPmpmgN7EB2K7REVDqc6LSCfm2ev
IjxyKQUStO6r9Y8Eo0zanlKFE7qKTd0Nh9r+nuXPg7MH5qBiTInIE5d/caS6PB1IXfE10d/l+lEd
gkMRjNdO5/4oTI6pgC9DqZcI0wtAm2POf6dL1qUenfLrd2KugIXHK7VpYplZ+QFDKcw9i99Pf4gC
1BYQ/PbtVzZJWaIjpmNyyQ+c6m7q+5VP7rN7bRTFddTULEmPDv7RcAmkHsrcifk7d+J/SyCMW5yg
nW+43hlLA9C1pDFs+5/E7vb/INRvYXcKqYJKX67iURwaKeaPqBEHxjNblH35A+laj4CpucjZMViH
dQu+4OY3nUj2uTw/9WP57l11EsPcWkPq5eE1DdWQZrXVXwULfTRy4J/qXmRTrwWFjCVk0hjan3pk
uAWhfIrA17VyC0ulnO04QN+OrpAWNDlx7x/hzz8ohmldS4MrdsIDH5Iv6WzISdquDRLdk3GmKP3N
xw+58Z8yv27YoyVRRArWu/sun6Kpa6KjW3oXhcVBrvH5NSUtSMde5aIy1U4vzWq/g7JV7C7ks2QP
IwLpuSJ3P90YzHiwWQl0p6xBguk7K4ODSvPu+2eeiQ6pLYOW8M7ZtpfnRHtif9F5fvZFWV5OtSHt
Mevda9jphWo8pp/QDlb7MvhQNp3pG/HXSWbe8mnwVayvfx/IUsA5txITr+ZFPdCu+PY9Sam7JVtf
UUqeaXnqqESWMlAnGwc/9qRKQoGJegRAT8VWhqBy/u88NRwBF6yyR68cZb+cQfnY8CfbwvxLQbfM
c50oEUiGUJYCptJeHCpJ0c9Y5rCxspA8BSR4K1F1LjsjArtRV5kVg48qMK2XSbybBxHlV/hP8nhW
4zsFM1Q3du0ob9RNSZQo5I5CJfhuxMfe6KM2farE7iXqMzR9eULhQr32m3aCcSsVkYqmbx6XiKMU
+je0ZlXg1krKHcCLLNLXk4w/pO8sgNm7apbhHj/XWzZ8hItsNstEhMzbbMpJII4ISudYaTBaiWnh
a1UNYEwMI52P7et5YJQEkG7rJ65FUjU+l33s0bkwEd8XXMDEzwoKgdBOWEh1ByLdh/S+XFmJxfNu
C1itJXecU+33fFRhUnTBYJZn6Mfg+g5hxo1JGw+l+GHszbTBidw5naEwtzjEg4uerfub15uARGRV
ViKeqrwfVl70J9REo7pqHMZY+pORwIvrfTBdJI8NxAWAq+W/3dVWYEWxneN5iZMSaGW7d8MA5XQb
koHKXaXmdb96YdwCmitFPue5QeXVBgtYGItYrngDdbxGmXOkuhZeWJwR/ND0LHyynN4cGgHuTomW
Xnw1MV4Gu6X+17L9pXO6UCbfOfZjsmtGLkU6+SwaItbbPoSE2TndxeuQvA2sDK4+2t0Y30S+W37/
mj743Tn9TESCAiT2J+NBH8E2S7Dx4WvBN14rTNHZZaGiRM++ScjcLCRI1A+E9hrw3z00oYi01iox
YqffcosPINb//U/9bul3UKlhfoU42ABQqLA0ISHO9Ym/qwhbLKh6qCXuIILQDpuIf66F2pdUHZ6V
lUBaz0tvNtP4UHij2oYK6A9PNVYf4oaX5gn5Xp3NxSVTPwaLGrdX7Y8P006VNSrnc8lMkTcZOb1U
IFcBSOdlysXvISmJ+iB5JDdE9S9MRwmlggZo0vW1eYytspU2D9GE22zxm5IDxkOvWe8hN2y31aUz
KQr+7R7TBUbP9kiVEPMD53iyqSNuwWYdRKJ5HINxA91pzOzyvAMuHWY6rmGlXxHO5+Elaw+LV00n
JqjX4NTGFotk7Lx+s0BE7bPruNBEc1Mmionnpak1/HOEsPCju9g+/e1TCyUD98mH0PYgiyubJv3Z
qWrABRIwFXQZk2Bc04DEXP3Z7H8BgRNsr8DbXaQIDpMKA+wxn0Tk1yZm7dX87uhn5xR/BFqwKwwX
BuUmXt6/lI0eWtjr6EK3+UvfnvavULbVuHMoTFD01gFKEmGndbkaHma/60Bc1UI6WvQvJuCOT+he
pJfpzJWkoaif//AS8PFvGgVTA2rQfZ0OgsXvDjrgN0P4edScZIwTm1+MLf68I0j/G1LmPNcSvJXJ
m24EwTwoYw7yrEBwhEBWLRFc5/OOwi4lmVpZh+7SQKX6XkjQj4vAaqsAGWwwJHvfVRETI2QdhAPS
1Qhyn+kvxQW4h5Yak93Wf75i5k0GTd/0N1Or8qTaUgvGR5gr2lMjpaqbdKSTnpLxNNus8mmhTkYd
LizpILA1TLYkuqidev+hMdK4rxJ8HRVA+8E9oALyPiv/Euk2b7dyOU/+NTeDjQNu1mvBzHqUwgAX
S0s0ASW+NnpepFuF9VpIWhWw0MN8QHL+KY5mj76hodpFnMFsxfxwIPHwaGpXeWOWH2msHBho7fSv
Ryw3iwfJ+xFATvYxgJYo7skxNEaeHhAPNaP9vWa22IYWeHfidpBfW+tXwzp8+f6otUF6+fsCNtLa
0COOK+NIrl/vM4fKs7W6C8k+kMHTa8+nKupAOz69dNl5hUqolMhBAVZUdzK3Y/OnHKfE80ZrgdY7
n49Z375bCwN39a2Ck2NIX+TRTWN0Ah8C9yQpP6ckJW7wOraHi2cipjAI7AvW6CXWEY0ANQsEjXS1
5qO/d7G/DdlK5SuXXAUaUJ1NsaOtJcE74X8Qly8C2M9N2S3QUNZryNarABVW4UkJzid7r/rEVG5Y
4ePQb4qL5TGcrYNoNjtBJUyhherkciv/DYX/SRKLlEuFEWJKN1LKAbbG88+5Sn6Miqptsk8aWpl4
1DCLDD48RguF6blDeWu+TA6bzGmm9cF41g54UMlBMGAvsQ8hprkZomwTJx8IqBYtMp+3mILlGJZ6
/dxE30ilBwEk9tM7EP7c262Kbxdg62zhKmpIrSacdhsxOwZ0XFHdPwd2N+LBZdySFsxf5NuJ9KVE
lI6+3yGK8hju8AJ3A5fyt/wWKFZxX57KcD2YvVw9FVrSUHdVZqkus0UAuH8v100Xldc/LhnP43gB
DfEDt/5+EOHa4wVPhSnZjWpOGY2UBwI/Qbcmu1flbY8iJDDCd9ano6Med5cw9ivwu2oMOQlzwwG+
XRP7Um/k62Zv3nIrs+Y3uIU09oTqjiQtfzUS6a/Gjb40ROSp0xpUDLOpKPxFED1BOv++EPEHp40M
RBv6MHPjUzwLWx/M6oL6POhAYPIsAqjmXMSb+nAa6Q/a5iDo/1H2QWanClB4HtSj+v8tpVXYym/s
DvXE4NPCWK+XpiUPiT/4X9ti9nNWrd6zvobFyKzwtU2rw3MSJVo411CwGQkoCJ0nMGD88YMYg4H2
C/jaV4vHQHxphhtm5sMqB9RT0/1q1XLK68L7XfBC5+ONTmytXtMgX4BWTWleEuyKtT404W3OAqxM
BVtTm1pNYnBnQtdYzyezlPsfBl1iRAiq94vFGvHmTlWhhvDUwQH2zSdPlOr1rb35soDZJKhtH3/6
KIce4gKWSu/vEF2/cyprDZch3otigWyovkviBR9/zfILao5JxYYEC1kmN1d8lhIkZW2MhamgvuLQ
gKIsLuCYLpHIu6LcM5g7JJ+gfglBUBid+14T7C30jg+7TeTQ8VCMvQpUlqSbRoZ4AmlUvZB+hXL6
nOaFotH/kVvNXw+soo+wSn1njNyMIKZ9lPK2RFcF+hn+u891b5NW9BtTw1njNko4I/HsEoHErSvt
hXtS8ri8zxVlkMj2e4+HtlJ8CAk39xpLGE2E9wTkH8Tpwm7oyp0iowPOSnLMkf38HuIyFrHcOGjc
dn8WHSR6HYBlwjr6uXtgOzuHdj62PwLD4jZpWdfKszoB60ZwxK5KlfF7Xbs+mfE8t9vqN+EtQ7Hn
dlpRlPcBS9G/mI920CHQM0mcTSj0+9sg4rowe72sOm1rMLyaQh0sphmHL1H7iBHTC3oifFMM+1SH
TOYUz2G3E7PVzielBaUGE5F+kv3kPPftq7BlOLBBWGWtcG0gSzA65AS6dSO8RqV2TI1Zex0IcfIv
ExMjWGhKE3UDHsqwdpjbSA/L5yWse8r4IXWBvMLy779caO+hbPIvc4rQcM6aagQsziPHiNAgm9L3
ZyL/VG7tl1Z7zjpS1YPKoFcSKxtsWYNHIiflLPKKMCnjctbD1yfbowQ9NxHXUsKcdgngVdOhYWMu
u+ThVlGC3qlAaSZP+F+ZuXxYcE5YoTXdFiu49Ei6F2O2pVkdj5t3EbeoOfFAmScdoFXNJ0DabnFv
522zNHIlCE2PDPGsCoNN3oSSElzb1uSN4vRpvXzfn4r0EDxeEacUqGLBHA95bjTfFm05nS6mEVh9
mYTAx4DzZb0Y/zVPzw5Uh7u5IR41G5kEOwWKHBJwOK2ngS2ZFgTecFIDx3GeY08gVyytsS4lRAAH
rjPxLAMzxr2e89qziUU8jVORD+ss/hv+8eUJKbWDYg7d9ECzXazbcEvz0/ZhpZpxlyOstxVh9eDJ
n32SpvhWRVK1I1H2F2LRxU9xa14uWqror42W+uAM70kU1E0RUgV6Yc4RSlziiwpQWflJoZu4Ttnd
XpNaPgK2zMPt/EC/KYGtzkGz9L6zxM31D4IRilVNxJko3KSdET8oBl+zaSCsrGUW1rXljN2afW3r
PLDDUSlkV+N3PcrObXhIIMAbQnnfa3RtMpwgjvJhhxKAeXQJYWlciKmIInn5acHs/P1wI1hZDDBb
R95jTOhfBBKJGWq2aGeegS1Q/avuifpkl2nKyDTur+FTjNitkSagkQweVrNzxR4C+CZecL0IaEbP
jqm4QY5JCBbtvq7EHmDzuHT6r+Qa+OPZ6DfLO8o6jY3vwXV6WINnxFNAQwmq4s+1BXVhhxIDAnJI
1moPwS48CdFwcYdb8YwQr45fZmhLpN9h5d0lFYZfryL52cE1UDEp2piFZIMziyCu+yF0k28hbnXT
Z5+INO1K4gnvhqzixjaIS9xGW6HZfjR9ubzIn1F9P0S4OCxK2RuuxHRtxQGY/o6BgHJEGf9wkVwv
tefXkBDoHR/pie8yArGIB1efgID9CCgCC2VSnQLdL968nSBzkHVrSYbuiYAxjMi/ZQSi3PwOYdwX
QF/BrAnNlkAnrbxjYcrv7UJVvr0vWIdcY35TV5I1M5fRE0mcCVX5rEA5/Y+n9Ewu06r7Cq3ylJED
0FUl8WSENFUVB23h9EyEQViaNeMG1CJ0R6Hff2Ny7c/l36vPPW0DR2nHJei3uPGR3MZ/eKJuvv3X
wPfkALG0bo3fpL5zx183fjWjusDmXZjri9GJLaOtcmK8NZxsRerjGQ/cae8SGhrMUA19vvjKpzG3
kZqfsH4SvJb9ta0jyf6I5t8YeyNfFDclPHGzzQzq3OIR5j3v/wVLcZKa0jod9KxHaReWv62o+2pE
VvjULKp9GOSpxWRv/sjoQ7r1KtSQFypjPALThH3g9DY0IiN3z3MPlX9FfXGJqizO0Qsmmwkg8KI4
RzH3gMyDQnm4XA/nf0e0IUcRCby7uvlaOQMqsNgTfGE63Y3mrPK3oAIaNnKruS7BREN4l3rtEIuy
WZVwNN19xp4mKAjJTgUAEGaPgqBvztqrFSPLFLBOdEqSbEPDSmjNjoYTD4Sa4nRPwbOvivrdEOEV
U0Xi/JlMrOXzR906ZZU2gqNtljYpo6VlmNMyCmphXfE/tZPvjIgjDOzZG23OkNLP7+3zUEoYpknD
jmZhXdwh2h0KxDyC3sqnBWpl2Jc6cDVIwdKa5JXYdO2OSbWtBJurYcg8LKgtU4q6GAt6mVw5pTrX
J58PM4Z+NyHhLc78JcBkjfk8ozOEWAlZ7tqj7K3BF3ZaHimgB1R9sL+kCvK9TT5Nyh2id2Tnkzn5
rgYlH0XWjp0Gz4rmiSAFZU3lwBCvIEK8Q8jQb7fogNmfbtfbtNJussKK9r6YUoCmblHqOD2A+z0k
ZHh0v6s224fz9HK4hsz0WQiB1dow1bTs4sG/RgeesvUaasIxw8dq24mloLU/A4uZQjTHZpCynAkB
VwqTAX3YzX1zS4hC3m318pNWguP2RdPjc6oZdM82h4+PcQt7KCvnslg4KV9jdu+bS0iWyGRpt5CL
0Oiptj/CvwuiAE7qCJNZey7rBDekGrDYRIvh9fjs7bmOzqXRemiRiXqjFD0UM6rtS6gn0J/fnWnN
ZGo7nfuz5hndY/8ggKTzth0NgPBkJwbo/XUm7Lw9++14p9rUirUQ/oLO7YhucDlf4kAfVG/2YMix
iQQ5WJzYoUqI0VjDdJOgZqUYVhuE+11lplj+v1gW3xiyQIw1Q7YPHgyIat+MvZdIWjP1sD8hHjPf
Eeuhx+Cy0D2DoohczHHEQwM6NTjtTWtNrOIFKGyn/ZwlAcRc/kwNQGRmmXcKHLGewnXyoLAthmjH
IBSkJyyPgZG/uLbJOERHo1S5IkyOm3vVvfcX56+yADukdtzYSvuYLcUESc1bm8VCrDE2Wlol7iuV
VLxMbbAbXXaCpfMPvA2BDwiFbL4rW8nLhudcZX8YJmnSxnG8hMqv94OpzQ2mokOsa2IDK+dKMczn
M4VOpk+PggRxUYSBpwcegK2BiJ+szE+GTl6+viWZbNFVY+CQwd4MuXQotgE8O6u0pFDN4mpCnd+3
uWVQi49vU7fj7drT/qpoKkEXAOTjvAIWe7kImiR64mwcSwHxL8SRP2oCB1KNfXgFDtebanepWPqO
GcktPlV3jAt8usjpn2jZR30E7dCrVhDK35K0y6MCJhi/rHjJZr0KB4WUPwWRwsmnEhXyTBLiI2o9
h3AM+T1G4FjjHnIuXX0LmvlBifDGE1LYrTkiSQ1GcRReqH9Q5lHYsqvMPntDL7GNCGtnwQDkQ1L/
bP0LNom8lvGqeg77JzZhM7rgU/AFsnb3xRjj8IxerjzDW2DTCazeSk7BHhOdRYV7rvZeP5wtr/xp
kWTFOJR9UkauZWC4rOchwgs7EicH9d1esbtjGlocoRkoJD7RzQR41wAqKSZLOjr3tTPRNXwLhhMX
/GeK5oPN5EIPZ0v+3UYAOCiGFsAATfaTQrZCLaE+kHE70e3unH+Edcy9psW6sqHWgpxlaVejnaAc
hlUMcd2buqj78qLSy7VlfdfdMKvsovScABZmyjndpudVGDTkUCdwtP/0PYNHg3qnkW/7kJpXv3d/
+WNPX1qCPEBJ+DD7aE4EHHM+YrM7TiJQ9t0XoaKsmDbtuP0S5naF0IHgU6PQiyQEV3SX6BpRJpTK
FQpooQr2fx3+U0rM0iyFdzUKpBBeZ7r8E9++Q7Rohb0V6+HPLsEQH1Nz6CyWpxNF/JwRukf74VnO
s9jm0PIvEcy8OkkFIiNjmblu3pkh+D74NUvbQZex32NMybBLUmNQao23UvZimdg3jHuvjfKbQ6/4
MdSUPXsg8kH88MjAlSwm9Ya7CmLAfMoKaZ+KFNegicopn5x1RO8yuXaMX1YLNp0cuuUDKCZXiGw6
azZzPnXZnVJxv3jhnr/8HkOipM0ieBCWXiYRFYQx4fR7QFwSrqptKUYv6psNJ/jYcEzrU1yLdFUL
ob65q9h262otjmdPShL3c5xPWH0Jk7OAmgQOnXo7b/2Me+VfDy6y6606SnsDc99CHIbkht/4L9dp
AcJlZhgzbU/0mxYcxbSeCdp3uFgQ4wUgqrRRrliulDuwbb6q3NIjV2uAT1Ti33C9DwHLPHqqBand
tl+0U1ajhsgcd4YEK/EL/4TSvio8Zl0mP5Rq/9U9D1H7ehJksuTXGjOqqV004cs4vcG03TqmVhac
9MzoCfykP98KEh1BljK0kE+rKoLlz4cBJLjcn6gZc78fTNYiTSlzlAcOZUpbPrUro4y9ji0q3Pv/
eti/KZmiyEF8PetU6ktoYOONeApmdPxu2oM1JQETSeDNvAUHCgMTh6N/HocNTU2iB+WOcAIlZMoK
PoyGYkzlSOdlFkfUhYWtc+ogCKn9M07u9+sHkvP+QLrrzFepCIPB/Jwjl71fAjzYpBnI1FpP8/0A
3hktdApTdxrJyKzQ/uRm7MII23Vm07pI6qKbamKXJ2ktvQAbL4bfRYvfIGncd/ngseDq7QYSy/CR
WWGeMSyhcNok+T92iBonVvlIh+bR4QvcwhUuX3kIvL94LnvmUsLFh/CbysvKgt8YWLqqP89ADHsm
PSgCTaISTFspha/IVfy8KGzSMt7k425U9SHhbLN24F2duPADEMaEXC/orykOMckzjWKjS3scbvgd
BSlvLJqIJIC0hmfb4ALNPmp4xhecm6tB0gCUbNlfN6/glqVSO0IIefzk/xncFKLPYFZ9eMw83V9C
x0XV6KbJfV6uDn7UYuYI35vT0Cv6Az7yhrZIM9b47E43ZgdDtf1ifbpKtIjm2F6ap9QkgRhqq1iB
A1d625gC1lsDmHdAWnKcTi2GJQV6Upnp6ux8/mM7qmDUePZBURd6oieJ5boHpRHOcanPP653nZ2P
/2ooEk+YRdDd1F1OFVuRvEw7oMH+MOPQaDAtI5rEqCoyndw09/w+EDm10WxrieBh5x1nq2K05WVH
ErtcT+XlNozHxNt1Fja+F6VPE9mBTqQFXIB/TEq+TTk5D0KNmTEjt3daowMONrZRvLfQq2Zk2XYp
+itTdS8PgPXOZdTfstRXzVNTDtIuKGs86rZE6gFLeqb+8Jyt7fvFOclK30UAB7Dgh/MSWzQvbh1q
njzxxUmieW+M5EPfH3RZfBxI68A6IeRODAIAdj2eQK7Lqq8TL8Zjt/PYw0xqL3UnS4t7MPD/wDDL
2OW0kTThUQq0Du0UJw77LenO/WPzx85ZXTg2mvZgKyYu9IBqf0VTnArDk91psAV2QxQU2FOfEOzx
sJYth9Mts8YBFKL8CoE+FebZMfAz34+jSMDDdJF3ebH6kaLM5Hu69/NvxfSlCoa5kKKQNIL/Cez/
k7Y37Ymq7fRYwTbvIldyhwkg2fS6HhR155qGhunxtaanctGegU2KijEFF5xkLluWYStII7wNMZo7
o184KY7wxIH7hHYOO3jRMXnbfefJdE4PTxCL4fTQt8sV2dWaw5mKO3d2LH8aDCgaQN/DHk9XnBQm
ZLk/FzoSDDo1NrWbk7+cszn4Fk+CwVx5BOZ6ytM5FFmxl6dHQtPq3Pv6JEhsu8QKaXndIVzvAHdZ
4dDLYNmcHcXjTaIriYSL+T6ZDgfz2FogDT5Opm2IOX56+48gC3b/7+CQnAjidLjMiHpmMu2WQe8d
J8EOSN6Xuy5E37HVsYWJdZ2+WZgOMSong0l7gWsqfx8J8LE2n6IjZ1xcJogm/jQhfLo+Lecr4wYh
km9OfSrjZzZ5Um3wyr+TDGZTU41E5xelkfvUbBNQnV2sd58QNUuIjdHx3bzDnH+am0gkRH0Rcbdf
4ItCOeqkU0BzxX+Kp2jH7lBe7vy1vbkwY9xv/dkfXj66urL/5OY9HgSqz6b14kK6o7fXdraWfXgI
fIVF35S9g10qF/JkiM3gqi9W5vXOs7htQfRx3JgfH9kQ7f8SjVSsYp/Qqct6n1tmKJ8fWzhvfhd5
3qFjkOHHfXHKGZjoJGQvcUQhIth2wA2YOIkHVAU+DUqfvgT8Cn2LLhY9KU/4CP2A3JQO/tqPfTZq
qlIbvO5e+nFttqSMx9OAj2q3cRQKnvCs3Q++FVYg2hC2liCoiwuL99KWYAv60GOaea3JK8+Af2LI
78TzxO3EnBqWLz3D+o6/hbAFLO61cLfQA5cGabX0fUKdJMelYFCFK74lpxb794ks0FLv/rjvkRxy
SsBjKOEUHTcVzftiY6p5vhdLjecML9KCSluY7fmrGnSygLQnXmZOC4XsY5RiB2B1yCG9RwRAp0BC
ZkRvo/WrcPhJg3rtRwrPJOeYgslxVruljx+C+qMvEa6HBZHoltAPBUOyZc8O8ACS7Jmj+AbNY2iP
YYwaUNPtSdoW/qiHx7silPFvo2S2/q2soOD/HmmYGRxwnh+mrD5AyEy7H4QWkrUfzOCulCUFf9mO
716kE5NRAU+7R6v4p6TeHLBCqXab5UNba4I/1JWOdAnMKJIrm0z6uFv5qGYsT4Rs6txfjr4Y0iUx
tWF3tU+jfw6KD5DTBDXVpDe6fbkJ8NdQNsLfrhvvSBWo2Aoi3/pI6TPHJ8cF1XAkDu7RMIwMWOCm
qv3+6weRLhm6766MHjCvlGAPCkxqvxjTNr4ST4aDb0N5Sxf6Mdj+DR3zWThcI/LbRumjfBuzzIIq
EPHtFSQJST60XLubs9GebvUqUeXo4PIrK7UXSCUDMR3mxm2XCLYEI86PH/AeMHrQcVZen/IwrlE9
thTYblTzoseT4uZOLGLDRw5YazGgy5CZ0xyVePLHswdCXyWKLi1rldGP8fUXAkBeGSTVgj74TfQq
oL6z12J9zCLEvq064hU6Mj3Q6q5+RcFE55F8KPkclYKjef8BFV4nex2/uztBUzEXg9UAa4LJefdH
PaNo6iybgVOTAaTpGwtrSr2ZX9cgs7exS95WI0397V3MB4yrQXb867DxbO/IaI6eE37yVOdSAPSZ
/aDawo79q4k3nwxrQZIdICKWrGuPd3C5UFeV+bMBiO844cSmMGNV2iQ/49ynAwx856iVFEQ/xx86
KU7+ukYQIa24eoCzj4Gxpz0DCrac0gQ9VJejF5bsOc40y9NgF+t6Cp1z4mqtDGpalhRaOKGvmfk3
i/XnKIq+9yePSTh9kEml1Cn9Bh3kAdmgJo95bcBihKp5jTrSPzlB2J88RxGSgO3pOOjS+Uba5XTC
NMQuubA9U8I5dKauKvAQdxAen//2D+0s/RPXQ5k/WnVsf/h0ZK4jFMU4sS0Fu9x1bfYoFay8t6PL
3QHC5J1JhFfC7LgKJOUGNOXW9glLiO4U2n/aKoVUVZUXB/vxEs36pvcxWpbKd6rmvvhrlwzi2ovW
x3ueu/PSqq+6uuunSahAJhacjT0uDZebAi38DsF7jEMXGg2mdUtGs2+lDGZeY+5bfeBcR1UFkSV7
+IBU0SZuMYu7CIGLnPQaSumb6gvmJmwJwYZVW9W3nlZ7SiVCWrXr4X51q5oagl8t46+ss0cfa3ec
7APdFh7tgckQNSt+94sXaQv9saFIDGkhe/EW2VnqhkowJjwbp3szc5ThaVArP6YQoJitf1oQ1mv8
aNzY3bv4su1GZuBciTezBD64vxDnIECJbuSlXBFoGfjzizkjez6ZwhjoX+YQEVj8/7pqvgpBSUZQ
rlCAN5F08wtn91N1oYGRtORFyDKPUgi6wD1q4iIwPYV7xAGQLq49FDO4SVKvROW5aQX4PWs8pGzn
8JBEzZmsuomyo/vpnyRkz9jHdOE/ii3gtQETv7nR1Lp4gnz6wUPMAwYkblOQOp2UOcPwTdH7JO3M
SUJSNZgv2uiPaAs/gdisHHne4ASe4ixaG8+74RkXD6/lizP7FRNQNajOxtEAtzyYrjDn8wQJdKYJ
7G4aH2yHq5do7gdll1djtN8W50y+WFS2RF0QTDQ/JLmPy7skIFnnTVQnDQe0X/FDiN+RQEqRH+8X
bPvL8fLRtZfBVKcpSnLoWRFriQ+Xtxmzq2kX2yIKSrzXfrMuFJS7Ze8f3Xnybsnhi+AhTfvK3VgN
Gdwar/nVOF04JmzauExKHj1RzS2Oy32uKALlsiP2FueEVB/wbc/JOS5ltBVm0hGWc1wrYDkLLUha
cfzNX82AhjbRAdZqjiJVb7V++omZ0jYpgJH+uXq3XwSt53qkzTOgJXNVVLHESX9nro/M/VEYLlnZ
vCch7VAougQA9vTG4E/YkMCGotrhZh+8lMolNXJ9kd+R5DsHMlcJsVTReASupnR3KchZF7CvNe6A
RKHuSuRw+sYeYj0vxtGFYpu+iILPJX5Mr0DsFBWU6Ul76W8zQUngpHrRJlN+9KZOZX9fOgBjNxPf
ORYxJqQYJINGb2H13AWPBt+C7tJZMgx4eSo5qo0eRB8L6+U2WOYze6U5aaVCKCjBrR5KKzkwx8ys
Vdtkll8weDuZTb54HPHo9UHDbKcCsib/9YOkh1cAu28nvVtfIDFPMdOaJ3du0ocW6ZvnuB1VLacZ
36EVwLAeYOqQN7lwFs4wN3gbx09JSVyogbHwDq2gbsv1unteeNdCseZtgT4roUq9Q2fDMatGo+Fe
BLSco6ziYghTKg+n0Kl7T95xZm+chxo06cDvRsDCQ4b087/BH5uE1vMYrTPYSG63pQJ+LOqy+2Tg
1nVJz02hcYh9QPVm+1c5k42s3+UEm2+U9EgShWJC2pKarDipik2KZLXv4PCu7pverEMBrzYROlFg
SLpFJY/RotE5vQN1WjmkWtKeGcGJEFUZirOj7bH1YBi3w6hkfh8ix0w2iFA+HrIHBHjSj43MCkHr
2oEGZQUbYXtAZ77ZKN+bEyzyQFojtqJE7C6SzubHTvdGOrFfuXtVT7z5D7V3UehIyktaLMrVndfi
fJc3MdNwdwfGERQg5WZXS/z+nRlD74cca8ncUnxL40FUJu9DHZVOKZXuySO9qhaZrGqmDwAD0eM1
9Pzmn9MFcptxzgiQsWEgT981cjJyJPYl7cIQMPAVSLF9BvwampZ8yWwvJ2Yn7/0UU8okZMxX87Ri
jzDKjMnZxmLLCWmuhyYiqjG5/w2kKBP+0E1xxfQBRR62dxBUD0UbcQkfSISiF/Pcp9WDUJEIajM4
944SLWHM8mAFirxtKwIH+HCtg3nVAusO+qdXNEjRCBIHYdCwLSBB5UZhgOaNpEIhp/MujgRscQOZ
iHMsL8guSBCK6gs6zKwfeRiu+C8tU5wFhXhqwYBO1E2BxwHHc8vlAtXZg1C/CB1AumcbRQuIvdoJ
ZiNdg0RrRm52rVY7OYnVWXcW1Ey7Wp/nrkOEJOAjBj6nssymotMm6HEE/kHx44bxZzbSYJy40ZKX
mjc6xlLzGbpkkPGyLRSvv+DgiyjGeyH+fpNIFlrGuFnGYuxiIsVkY/R6NtjcECZBNSZ2J/qZLeCF
wnFYSbv0hF9qbQebRGTMErI6znSWnaOz+nqkTBsHxhY78PMrhCqssFJfdzRmT9r20GewPzpmO5Rb
zGGD008t9yWeQvHkjMB883Sjs4HRzjDLrqj8PN8LXdlHggB+TFglbo2mEveBAcDjWDJJBeTZZbVg
3+bc9ZySd6fPLYrW0GORN5o9jYJgWphi4Dh3X05ipt2qSaAiqAVeEkODEmxPwrAbqBHfYgTwU+Ml
ugRhUX3QCPkE4jeNu/9UqVh4f00g+e6DHAvi3dJTuEzYzia+T/hn1rgUFYdxhnEKen5PJ6e/D/6D
ynn+KJxyLIhI5Qdw87iUfF1BhzBf2FDvOtm1pqr9fR+V48CrQvKdkIAxrv7UXVFhTYe/cyUnzwr0
Epziuon4vVXT86QX6Yo8pPtvVzleajGPgQTZtzHcIjc8pFLz7pmkbu2bmzn4Ib6vc/gFVC+eZNrZ
3CwX9r5/vGAaguxbIB4Qci3yd7yjP8waGf2kCepWgIn3vAcR1fg//IAIfB2kjd8fAWfLGJBY6U7A
LxiS552jVlcdGdNf3KV/A/rUZFJpPajYq/FSAbOoyAuoKCvWBB0Rws5OVNDwsDqW/r+w/5ipD3C3
6/9kR32cVl73UojD7Msx4OXeMwVlGCKc68J7KwmeO+Ou2JBXu1xVdjJQpb6HLropYdlitWOttDxB
A50+vMLd8PUIul6bYCzxHeYQza5OPAfGlIzgWxlGBj3qPU6V3LSbqRpw+lJVBeJ42UOZOuKEfHts
zkdzSMyfkWK13sTZhwtYY6+wBRq6xRLZnL4QgzaVR82IAd9xX9MR5Owrbr8kYoHEQCDAfU3ZHIHL
j0KqDvbZokGe+G9z3IJhlK9ncfdABWEneDL7QE49y3iHDeedUgAPKLjr2Z0B3IotlJAWXbw20gsw
3cZv/jBWt6XVonydVi2kWCM2+5zb+MfghCRk3La+7PZgIUS4LkEqZAquNz1RSzrzMYskHTQXpP1v
ETJsMv0VMK0DPfC9svTJb6QOHIaJWw+e9KqviqXCK9omIFHRv0508fQpizGFPSYLDdFd5DYciDsw
irlV9+Xk1rsCuZ6orAj/9J9COdHKFmzFZz+AUJzT3rtWAec3he40Urg765FS+PcnFGMe4OCZGDgv
aFPWkR0yz1AIkwqAwKBIq7i5h+Gw5tDvnpu7zrDCoBfHKpRq2woO0WOozry9U4Exe9pzZYYbhQdt
NPiUtdakWsFf3V5eHI9KgKEtVG4hp+SlDNXdZs87ycXh6Y+67IX3PHkiTlqXJj0sUeoh25GJdvqN
KbQL/tgYCv7O0hIPTQf2VHoyB6gzotroT8bPVKn0hYVoEaBqiSFZFCmifJAtJ3VsGxngCOo+66bq
L9p5UI5QFUztFiDEU4RxfKyqxw6TrFDj1DAexlsyLGN9RgqLhintAV+L3j8YV1pok9cbRKttU1QA
JIHKFzNhCzHcaJqbJHSGbXPJ7xfM3P0vDQyY4/SY4bjzPTCP7yMxlbBB7Yagbthw+S6O4EOUCEAq
TmUpMIMWC6F7eH0Lq1yXTNtauSBF8Z7t6WJ49gH5eFUtXd8cTgywbnAJDVOfGBpZkvLMYcyx+r1b
qlHk4MInHIeW3FBThApojeTm67FuAd9rU7CEm8R7yxwwHN9TlSYMexOo6dUnTFvk9yn2RfnSoEy4
wJhXRrLxhl0zGF6TzAUV1HvHTlgWYcUm9q2vHtWcAzjOsicCllBxetNVPGFw1Sp4+oXEPzujSVQn
6de9ckvCTH//2wzU8lXTT0q5xdSWYL+pSyZkYVWFQ4dHmxt6WxpmaIYRtUFC5GoM0Az5xAkwIIYC
DjHW2vpQr7oflU/57Mw5PjpGpIxxJf61KrEzDp6dEH1d1/anz/GU7MZjYa5Fr10g+gAo/0zl6y6H
SCxMptiGmTIlw6ELWrooo6NaOHN8IjxhQwsD4Q/+xEPdEq4ORyD/SjU5yoNaaIdj4OJPdZyxNqsw
qxp87RpFL+X8wE67gkGllgx3w5WruRGiTbCwFzdJrtRc2uCTd2kceEe6Pma9g267Nfc0ApjRRvgI
/OLiRsZnDLnRKDCE51Ia2z0zYLVCI1VdbFG+QXMVdoWFlDWVi6sePXrYLKBXlXv1W56l4LMwzQkj
11rVNVopuQ2LQjaHxbenYz074PA7uqkmtDlCYm0ltDJAXpPqysQDnHysoUFRIzxJ086hneUw5cgO
wz/1sH++Say+VDpq1ee+Y5zT9zTZl8GtHcIB+C+rsBTBCbYNe4aV/RK5/jdvlKmuW84SqEmnuONS
AEbIVVsuaLMfq09IDAW8x+lv1Iv6+rZEzQTr+bRtKjbQhcB4ONSucLy4eNWdGyxTzEJY246dyIuo
cdIHWFgRVd6A3Udups0b06ln8PItpemb2E0kHE3pHmg3NPACSuzxY3O0sMwOfYuySJnIImw4C41V
Zxb38cfV1kcxYFu2D/lJiJJqnpg+88BMZpcc+sIyXlshkv+FrddSoqQxCP8VlpYh2prFkP4me9wy
SFjvUVJTb2eS4eg3AMK316iMf9vQfW3EEVhjFSB+WWm489U8MniTrGzgfX7l79yxbxzEvrnZsgfB
kwmU/HEzejW8bSBbtgHelXgKJtIM5M8UaFq3CFezFIJ5WhrqHdAlV+2wPQCYsq9TEsLauoFr0xEl
jVtFJfyOWUVeiEz00jhVYTQ0ctFcKQTRMGcLJvIbxayGXK4gzhen3x4bx7rarwAiKFnKQAVK7PRp
OHZfhXyxVNzJqnVLklL4atgbrT/s9BC67bjIcEmNJfzSJpCJmwNTfGE1q8B2s8zn16GDRR2eu0Nh
j6D+zk3kkL0O2Y6Ig9zx9Nrf9dgILe3gRkc2SQGdMfPx3Jwd80Kd0T22lCrB5+Z8py1RjzILbLK2
BF+AMfN4lgEJKA/9yK4R8i9UtHHvfqDYZR7V91LPbRQtZvNuAjGwxLurKf6JPwPQSNrbb/iBuY8L
4OZ2j8Syz/Rm4456sQ5iCVhS4UElWWIV9waT9aQFwB2Y5JVgPYxZ633pzRx+08TGy9xcxPySBev5
1AqvICCTv75z9qpTLIW4kUoyYMECuVJib4F3akkk2GDGZYl7GkywpY1tKOjAhsss5D6FsPXmcjGS
T7QoudIOK4O+Acb6RjDcScCy57sm+yOw3tMlFFUhiP7WUzDHi4TK+ndy+y6jvLTO0USSrrMBDtEW
AKIBZnLy7pEnJ6okWZQAkXXqWiix7TWHk37YWAToPWtQ+lhd1472NKxHwnlTXxbDETWs3YPjl1gM
i0smWAokxKfLkD6Tv/unzJzIB5gqo+Plm0wVztD4rQSg7NbHRYo7nxXppFDcXgXFltBhHcPnJBGi
HotKIpO4RJtDYMILAN4E5mgdlyUOAInK4RrqDdB4Mdi4mJTnnckzFqa3BDtq6BTsPaiBr5z7zoyw
jYibn9axtL5DvkIK4BJkk9LmZwgsT5Tbclr+s7Om89r36RpWWrE2oByV6PaumagGCn4nbmBm36X6
YIjbXetpllNJBjsTHhXEVtwDLrcvsIkM/U5pY8hU1PJbxrE8h3aDXrbGu52D0CiiY+91o28+lwh4
VgRfjyeWuygrwDBLSmXkYvKRsriQOBrz/z7kjQRlM8C6CsPJ4vvKaZj/kjfggrbRYCy5evRmymab
wJBeqTwzTmtWw3Krf/4II9p0FzDq99eXXJ8dWXRyF10PcBOtG3xjN4OQ3KplCIlwoRDr4nrYLq78
Es2WoZNPWGORSr+1uSV+oBbzC/w4DmP6hBdBB0eCHk/ncoxlQTRXEzqtvrhAVU3iBPFG6WYYluBW
UIN5gnqaUGEaTm8kKy2EAq2X+X/PHBkfLZ4F3m03AR8JWeArxXfo5HTR7xuD1gOXOspmglCfQ2Vm
6s/6ACW3qn4vNr6Ba6qmA7P5zGOAQC3QyZaA8mpcMA6porPdYot9EejSL7P642yhIYx323oE2Vl1
RZx/LwFGuyuKNRGWqIHYpox/gBkXr3P3Svf+izNV4zpf5+saZVxfeXIbi5stuPScJCpTGGKSHhji
iYiyAI5I0l0+ii6R2ARfiWN8ZNypcXNOzkie8QT3/Uw1G81Fu9inmI+rb5YYoJTjzHL6AzYOtQKT
XfTC71gd3c+aX0M2N/4IjL9I1vpW63vzQS0c3YuqrbCzFa7fZBgDEiIhw9lS59lOwNyYRnzDJMsu
BSIP4Z2S1y3deN4jc5lnNbwUOEs7/K5szVqAlsK9D5HGok3BVhQdHmHxZRD1J45oCFNtb1/pR+Fm
ViSm+kYHgm3WXYz296KxAz59weYMec8fs4spGjP0TLtzpV+XE3bz+GSVp0BHZR5KXfi5vIw7YDdW
55copNEyewOfNm3mCc9K1Ku8pOefTArVX3ZU/zCiK03k9psmduRz23nIa/bvBJWay5oBdclHJEoF
1qSHePc220Ho+tKEGmS21Y05V15f50RjqZZK6gaAiaxMLHd9AhCpbKDrwkhxlpYChCqUvvBosKn1
d+njYQvzP5qUx1vltflzgz6dBpQIUvc5kdVfPVmYR1mwn8KjcYbnn6AXMhNQxCeBlfhO+lMDT3fZ
fwXegD8HQ67tTx2W+sm7dfY0IsbdHfRSIeAhWKeiB3Spk+XbJIGadIi3/XVhMiWNTWBxsSUSDwxG
89YIkJlzWCUEiIcVf/GLQDr+FfNP3fESeKdPc8fzasUZderBzG+bCwL853vNGTVtT0vjBA2Z/lkf
Z8rnQpIpbzuCPrEXu1P+JTmgXKCvFZ0dEzim7QS4RCLaytjesINkH6sAmfwaTlckx9et/UenaJ6m
74yYt7oauFSp29MlsjVKaFmXg0D6d/jwdSAO/g2fWr+S4RYshKSqN0hRF8Kqh5ouptMVQbBFvm/e
faYpKpNtzeTtLsA6YsRq2g+1IjSRRXQNjIm9YgLg3Deyuf4zdffqnuq49XQKkkRl1xblkCIoWTds
JhOhiwxo22Ad1APyug7Vemcb3Vrf5TCSt9GQVXQ96DyqCcuxQa/Yn69tE8THgqPfas3rbc2w7NcR
knRMKvohXhCew1MnU8dtw2OFvqTZzCmxBfbxDzGQLnV8hT6cKEJnPh+6Z7FngT2yGG0rl+fnIpTU
wN6CAwKHG8VatQlf0rxFyD706C5cay151iZ560RYb1CDauJjDPPzUH/aTLxuJaLWuiZKN25Tti5y
KxY6ZpNw39YJbr6jq1bJbKFr10jVT+wwnlmhKOPCmJxcWSSaE73rs9Dr4SuKCgHHLXUc6I60x05Y
vvXYi5PQDem3A9J+dj0o/QGovXwc2p7oR4Ei293Y3CI60DnUB75JBMMfpvOom3w+vQgLoBAsxxYe
XNsaX0GdKiVLAfx0wg26FPyHdgyM65fOhu+pZkAOtLDjGOJktFoF6PB5GTjaP/7rQvF4NvNyGpvy
aVJjO//wyRxLxBdqoCbBPpx5pK9Xf65rskhk7EMU1kC9ssfLYY3LL/Zw4u/2+aUdsojZFgcxkv2L
cqiIaKD61s+LIiY6M0/HsqE2vLZmi6HCgzQeTSIJBUpjrkGSbSxCRm5/d1CLwzH19WIlOKsPhZPa
zzZreQYuzLmT6lHgk02C4R9RO59cbR+FwFCL1cjBz4H3zn/w34V6ZzA0cTT5R97d0wnBfZloJIuz
DTRlW3roG9pH2VvDeQwTKKIxx5TbJEmM/XpVe4HNXy0WxzdPsOVfkYGDMpohFtNPXYOcNtfGDRRM
1pPcuynO8ZZDgr/RqXo1WPL7oIQsUhKIgTg5olK9VHSpAgSZeuLek5pSgC7kN8vTm26pANcHLkUh
XeZR4WIEqEICYk/lBLfSFk0KdwT6Ph2F0PHGufxHYgzdb1xYNT1fYrQXNVdb6ExsB5CVH6sG8/fI
7hhCG1fANmTSPZ0ptVS5nr0FI1aKfgGEnKw5i/Dgk+jlUKNRjeCjGPZuMrLnRuRlu5pO9Xl0uZ4G
Y4okqeD+IFtcHgs/yevyh70gtBSpubtNwAnT90PeHKpFYF5HlfWjCR/BqAmF7O36lD0pUmYkT5LS
AbedFUqPrRvDPUnkgEypR30ZOX13F6NuFaasW8vIYGgHpwDpt0ol+dVZRhZsy185rNepxo714jg0
DE0goYTE2lRifQzPCDbYTsvMdedm/Zl3Bj9hoFqCNnRIbIC/k7GnpLYxzJCn6Dau0LpzTmHhRucj
WCCk8ooYbB2Xw58hDsQaawAKiMfc9dkZwSeHtFsmim2uyGPFL79uDedWzAq+S5CW7JD3lJV+kuQZ
SqdOd51JXNi8W+jb0qDgDpwjRBcLtcpgQ4Y48ElL6IkSRdGDmHa4RhkfxZkAL6kD/zF3mY5+/nBE
tw4RyqGp6PkSorCMvFBcYdGXu13uFHHb0w4yKUldi/6LJrOSV5QQzmGZ8+B5MpKYJjkK5Ofp37jg
c3FbGfuy155dQhEiccTdiNeFMPI/vrTyG1KyWj2Ut5SbHfP+zf63IHHjMJPRrVQuY+xBcM2YEaKR
FwPTSC/Gfhikg/aXZmBQ6P5m1PMTwxvLyN2sr71wrZs7x58QEUC5hUMSjpzR4t/oKV4z3hu7EUiU
jM666Y8IRyWW89e6QhKcTctsXeKUVnPn7iCZwwjtrdFwsTGAoU3KglCL+Jd2ZWc1sGx1X8iQc7cp
O8r5UOQX+BkLjua5zEiVRSMblRgpMAptB28Oa9tDY2NQaRlAS4UQ4yqJve7V94f2OWDp2ZyyLX6g
wDs4VCVoc5oScrZiuUBPTUs2paw29ZlovOqvzuGp73unRFIxogYwAMdzLMyeTLGna3h2Vk963T1+
x8F4DkdlY5MvNsJq7pP/cft/RVYOskPkn9SvjaTHlloLh1bDVxzHQ6+4fUDrkIVgzLMuh8Jvvg/r
ay4oqozrVb6VEJpKhr5PQByKenq7B+nf/qr53iM9UFdbLj7Lk+tUlFm1QXzOQJMKdB276f8HkgIK
fjEQKGp/H8pPlQDYUG8cY+bo4W/3kUns3wO70DxQUkQDeOe5eIYuCK9i3LbnP5U5ezz83fquNIup
YTp9/AlupoSNhjfjf1Dyfvz91y/IGu+9H/YEHmUy/s2scLGNu+1ZwZvGz7qp05g9CsaNFR/He6fv
dYq7PWdVlqWidR/ocmJ+JAj/PECK+l58M1oITxNXI676Z2XQZ/pkxzG6Es6mp6t5E0W0yMu0+vts
LOrHqTjPlsGijGqxARqYLt3LmXy+YYpZcCbtfOGjtjG6xLt84XgtEpQGTZk1XrBJayYyQy5cF4ql
wytRBvZGwd9/BiP+t1ZsacMlt5xWVjmYfamxB+RcvsLozuhRJdjsxPdoA7Zqsthks3AFMV/BFbhG
E+3yX/h4kXc+yD7TT61UB9jDp+RsK8ol8W5Je1dXEGNZz8P5BtdrFt1qQn6KwTQOmgsyd7cbeWiz
ZfLfJnxPzW7n3spDjYXsBciwa1q7gWhjFC8ybiKgdRmo/6S1ue1JPihXzG84JShjyR9MWmJH8OKS
JDUG5b4Q4EPxhFsSfJ1Xt6w/YHRsL8as0UO3zIEq/R77KPtoXWrGSbuKWXIvcR4lDrbZ6aRZweCu
NxIFsEihbYF+7ai7147f2Ts8riDoRFTDXBOOPRXNLH9SQn0HXCvphesVa9FOade64lMyCewSzEhF
Sw1zxrMGqorCiDakIzi1nLIUidpfpHhjADEwc/7Em6NNVuoduq9/+r3PDzxrLDnOkkcCIhrQPDer
LHj/BIctUeUlHPzRjv2PpM3r4CPucIWrSxaeWY+OE25ahah5XEios//LxJFizcx6TScVOkugUaJO
KFbIed1hL+u2oR3mCd8zWpp5luF1xE3wWivsbHt0eZy3+xkubwBk/4SrF+L3SIw6EWUsb5Jhpok/
3XFzgwciPLHROFSZuyk3Yy4AvpNsQgv1mnLeJg5DI4bHv2FUhu84pdU36rqNUGA4dRhftC8Af/9I
djaZRV+BixksqKe+/qgBOZ6rBmBH9im6sNaYcSqVr5aQOLdQuhzRn+FDWBDGTD8rDhUMDYa87lvp
lpedSwMgF4559I8L3+muqR/gHOobWSLWn3l4+Wv7NgvoL7cbrk+xPVZEjoMGEbg46tGh85c22fZs
QwGWYF04d706BJ4hvHedwZL4K072EULI5PVTAH3qpU9kbQhdaPKjc3ASFcujeYUH5dr4DEOmd+Lf
J+VMB/j3RfN+RaKUFdXnEHlnbISkLFgwinElb/ocoGNXtz9GmZCW9/ppl3gPmXx/pF8Zlr1roIzT
yveWcwdNg3bSjuRXOoFzk0Y30Tdcsd0+ZauHzicpnrBErx6LvaE9IZ91Pw5tXRtGseMwzKZgSBT4
ic90XTx7SfUhJpEuqrB0ZKVebDA7+Dw+3IgmH4pe5nzjYU0dCo9hGYapgL0iPMgxNlXvpq4IX5lt
BtSuAichI0w2BzU5YV+2hGYSTHBdZGQ0+Dplh4myAQhC11CvV5l6nHKIxxY4C8eHp7Ac1a8uonUV
A4DXJYe1zFbIabzfxYNTE5j03JeYtGR93iLtMRuFzYYjLFyTGipLqSRrGnTT9ouMqLf8CR8tcb3U
wMgdpwmtusR9uzrzobi2ReF8JAe7fHiwWNfw/ObcZFerp3vWZRYRlFZb9iajubldthjZInlC97rk
g2QGQnXABK8/In9/4WVWtmgtr4Dsx8yWsrDGsDFF3139xJpnTu+PCjDTf8T3iWqtFoswW5ngpkh2
WaLCJgGGgWVc+dVsu7FT+eJMlsTb+Wqz8XVjYBanUlJVxZmWGZ1WdvwYKxixXh2llkO4ij4DesLW
AlDXbKz5wevsxxKlZU6uRGyzlV1DHGcdcrxFDkpGSIz47JQ1500aYAz5b8UrQ5yfkQiLhNHfDeCj
p4IJHFQEa36RQwpIssJocMBrOGHyhIdf2ra7NegNuceH1ULc4hHZe+4+H0wxrYcuAtMr0dyxzV2i
GjNDiI6iCFASaz0UCMxbPQKYDEsWLUbsjhJ3/GKWRVos6fjQHJ5jC9RY3vBqYkwknj/ZG3GDpEgC
nS4JNAYrevvumYAWkBGYiC9ROeez/BLuJ7VDndd349xcf1J3ZLnsU4zpgFvQ+UVhTR+FDf7ZPdZo
kXLPa93Du+mMZl6SUhPJqUGsQWQEi/f9lIx5M76douk65tT9WonZiJf/6fVyJiaqBujsCp45xPae
E/lCPOoaESRWRsXjTRAHifzuPn4UjhxQTmsubJ3Kvd6bPCeKokyoPDOtrkfLkQyf/c0qPaT6U5Rx
Gatpy0Rvco3r4cyXef6ZMapEQC0PnICEzSlRINtc9sCfH/KI0FUo5DZHNe5duLRHYejnVI4NNuDj
5REcmOc+Y7xnxUJdzKtkHfYZqNSFnQYPHdPAwjLBRQdMulV9ia3Jq0lMnepgwlr5QGeQm0z7F8TZ
cg1yZ9D1IWmhAhBBhxtk+rJeCcyBTa5Vh4DU8h/6gz62vwwM9EvU04xUikP+P+cUdulgprXJFwes
Cqta59nTTkh5x+uzCCypT8yUjEAs1uiuilG6A0uDmfHAL7iySfL47lr/O31aZBNIe4W7cj7vRMry
SiXAo7R0ONp9iNhtLCSasqT9WOAuai/GYc0+U93kGBrySF/40U6Xa2ydamnIkMPgXyIB7dqoWcW/
0YkdvVpP/WvfbWv+WdlUItHLh7lQbmAv+XQAOtAX22/d0JNG24Sub1ODexmPzRXeo76EjJQ0iVap
mGrJuwaq3sLkPRS70KGSMcXmyXmncjVsuTje3NKRrzXSXfoJPkghpgVZJGYCuRXMsUUFlOOAIGz2
r1/29a8sBBhvH7kINuh91W90EA7OrCuXKHlIAl/hwLmjgTvc300ZykSYABszXIn+bi8JT+Qv7dGW
4IYs97b8qhD9tWEdiHQ6mRlHvcXe7ukl1u6dHd4XB3p6glpgU0Bx2gHk4OdeOjduMnDI1w+HtR0C
PU8IkAVqrxw8J8utwAVMAKvMJUah2LERJ1WT9okpDEb8Lz9HekvQRXme+R3j5eM8iRptsCumQXtj
4kN4YW6+bTvA/P/IEfKEWFAVlq2ajyR3IuYr9NXBwHgXlwqlyScPFOh0wKgXiODgvM2Xr24Pi6nk
svaotF5nJGhnByqYr+nGAZoElYWAGLkyc+DLdJnx4XN46gG72PEhMaUxmkhFrxJ4W1+Hb/TwJ2Jr
9ZNGy/qHQfkwfqeQFdLVWmspecknfcF5n4GhaKgwPD1F01udO9kp6nqVgfcIDt8j2pzWbsy27EfS
c/5jFSMKdYAPutVg1ksisaJoY4XmXhfMkKdurU9rHV/sniKo6TrqXgzw67jk/CLxfX+qXOFpy2Qu
Iayf2AK27Wj7ak+n99ErSr914wDy++lPUTGwGPM8155KCoWexkxfklBfzhgZqlgtxKxLfJI0Pl/m
Ly1z29onbBjIpWXrCRrLLgEzN3/9yarajedxDdNjGyFyv+fk6cok+enzn/zL16Dh1vmRHTQbzwqk
NG80nMVSbM6Ig5mrA9xjGVY80krODXyYZonYXGeOQoZo7/Ths32UY58SwdX/cyCsYJvgKb+wk3Bd
aCKwupJPPljnLQj+cXJ0/4/e0Ke9IivD6E+L5dONR7sLKg+7SKgyZCwk6i3EMXJ352cgnmNOeG6T
NAbiVoidq1qhSr3KMtqe83hRdoVub7hMxXcfv2toiYc59pNxl4YXvqmUx9FdKxxJts2Avnm4KefL
46yEpmXbKQr+3nGEv4Wbbt+fK6BUTeOEqtDS4TI2crkJNSwohWGVVNMk+nnYzWdRtgJBmNTZARYm
3AsTdNAeXp48iTSlU4D+cGEWQyXLnk4gGsTyj7eiajOrbm1w46BQc/gE5rViiaXo7kuneYDj/afS
b4GnIN4lHyxuSMz9kTXOPSl2SVUP6jnCzBTvPliCHXvdgI5R2y0dX7SUR21OEZJJs2mgFTGTFynO
Mt4oGjdDTj3nLCSawNmhW8rfX6mPkUsbjl0IRe1M+AIONuUIxM6bIAyS4AC1zGiOdv3UtHjwrIqZ
oWHVX8CtPbiEYcPHoFZDwspcCn/GipyS10Y8egfIsFmxqHtHOg0I634/LYyScaH6Ho7h5YV6l2Yy
WOLsXdl8F+82/FC81RDIrrOiPH/R7m7yBz4KAZlTfZpokYVHGlfSUbwHVYxQs8JlNRBr4hT3J4dq
d3wbUAzFIL5rCyCFaXDt5BwM3UhVAwJBTfAP8s0HNvw81shU7gUdQWXDGqu3cHNYK319/WgItVtD
AKhuZnA6RNC6aQt9Up6SkkcvOxN6XI99uK22A8L8Yt0M2K4NxGqyesWcgTYom7LXMYoJBKXQFU36
RshVNQU4O2DwFs4mieV1E3Vz997ZH5Qu8xaWfQcOmxZjKxhfxTsVk1CCo4GkumrumqfgLN5JPWSm
nk2h45KdTSVY8IgO1cdGuAo31knn4pjATeNFNkCIg0wshforAEqe4iRZh1AAv2edqZIgBo+WwC8s
9sXjS3/FdSm04a8ug90pShC3N+HOyosFqwDHcBrMuwVxpS1crGY2ZZPMFx/G8Ze5k6E9ZtjfJj27
YTcOU0jHBGhgj2wr+viF4L5fBXOCFEKnDbY5enkMA9ukpkZ18w0u5h3R6EgU1hgNgHH0r+lIdS6y
gF65lUX4mUSVVXO+bJV0aodo3zZNLUfHqzv6iQBSSvSFwBt3J982oDYTJa6r0KNNKtcrk2jPda4K
kzK4dv7rZoza5xAWvQxc6rqj66OuLn3GB1c63aXguje91lidT7Psx9M6XLAevdybM1qgfIaUzbJg
+B6U2Q5alPkfAIk5EP1mlHVm5AYg/cyUesFMWF8ZXOIIagY18yhikVeCoc1EUkVQuNVHavWx+lis
FNGD9LXhyzPGypcFVc1cE0mNHnrO2AZqLqcPGsJ1O08m2NbUvs6CBReIAcr4GgsI4VdjAYKfCRCx
eKGOKD+zfompjGfukq0sz8egeMud3DzR6BDVhfoAQ4/8pqEJTt0Eh3zkMECxlnAH+gKI5Tonz/r4
GGByLx4+00jBYAN3WwDlf+F9WyCW8laTuPLPBC2dYh4Rlaqhc/wNFI1XcWh3RAPG6uC9g5YXkqHO
MDfMmQCC9TII5ju5icelptMiwXXgCBbsTxC1oFExcZT7nRIz/HmmvQpMlYjs0ZbrUeAQ6UGMbZRK
2WkmBX0cSoeorEFLn06PuLk1eqSTtmIZnph6RlgRP3qsVrqIgqZ/9PxiHAm+3ok609Vg1EkELgCP
t4PBH4+OnyfNJ3Tt6gCD+CnD4nkZCXl9wP3nW/rq0Dc1VQ3jB8BFypIcj6XwN8Avmy6AgUPtuNGM
0Yuw0IPJP3d6mjpu0ypCJ3mveZMce9Xj8RlVX2GMLCu27cF3/6m8e1b8FbLnbECWi0uDY2YHTd6z
DbQpKxWb6r4Tg+sogQ/R5LT3o78g2Ielr+csUcxbflQ8fKPFweRdN+cKjEKuMHszFgro3LfGizIV
5wf02UcqQlKFeIrN4blOV4fGRPJpFUTYwCsHm9NMKHzJ8NRX87R0MhRM7ycBvb0DE5K0WoV7RUFr
H14BOYYmpPOpT4pX6M/Rk0Dw9jprBQEiaisQKpAXXdb4u6Mi9gl8M9DpkPER+9+syLwEJH+JjNSO
4Ee3s5yljYp0oxsgjhf3LShpuuj/Z9dGaiva2jLz30xUED2fPCjyjAbK6VfLL/ji17VTmM8qhbNf
5hEwK3M+LDEDiIiepbUm7afdpJi0N84U4qwLfcj9hQIqbNxYZBE0FVUHo4Bg89+RDm31bOGtTLRN
bjpjUoUMixDMOHzc+3fqYU2W9HXQqibULS+32UyD3koNFDORIphYYtJEecFurF0zyEgTKuF6wF1b
RAYrorQQlxx0/nnMC0mbNeECR5PTRyrbheZUVZaYdwwvVG/Rs3oo3oLU3s9uqYv1TEodA1K2Y784
IGWsKFqDOBmz959M50I2ua43q3oUwRIh98f9qmw60OA3SuzldfVyofEMS1n2/dCNBEJg9NQFAV2t
PhK1r8XbyiaaVwTkAQsFY26qZ/KRY5VbXvA/SN27M8nT5XoRREznFdXWWvjz3YhlQH8DIuIL5jEW
4XBWb6nCn9EcdKUaGjbB3jFeJLlB82TSrHT6MOwkYDXIy92FDMZwgnXt2oG06M0OyB7P39Mpe3JV
U7uISK4/rFMup+l9RVy9L5aS7i0EgjBHTcx6YI7efCnhUmjMlSUE9j0Ux9vElEjtAptsko4du5RL
J+JKd19ujyCD/9v55kEFiwPe4RlFzzMRE03aYtI9sA53pLK6Oc+KhUdVUsO3pw5MShBNpYrT43Xf
2Iz4S8I5ZxcVeqEQbyroKEMmlmF5s3S8nkif8wXmXlYrzh68eTVNcFjuKJJmmnQ2wSTcejmxVyvd
/dVCguenLkOxWtbXZXH2mOVINC6MMhz/DMSbUQrs4lzu5Kxk2ZL1wKSnPJvmb5Fm/nZtDhK0T2N9
GCQsxVia7H3M+fHLcwiYLPlN290eG4vbSxi1ODfYOzhnqPENfClv+6jWrMZECSiylyhNSht72Rso
RBGSo09jKZNZpu5S/kadukB0QXXRSEc4a2W3F9zhlv0bijmNurc0EMw//VCsxaHQEFCSq8cOCNDe
VrbM2AaQMFnfKDHkjrvfp4xZ1jrsFEoFOtp1AZppbkT+ZWrTsZiTu4oES9BqS6jc7fW2L32pm2gg
wZIdtGB31iQavepdLF254jiOZM04kOmX/2iumh77C1iQIFNxG9F9Dq21e9EbeJVuKsccAtVBUf71
VlrYqwZYjXFGzli3gbTUMYJfYED6dYf7kNNZsWU1BHkWzHyZ/Gn7KZ+9iU2HIHbSD//E93GGb30M
LGLTafG9dFxZVpC1cokfIpxOUmeZjxRU0AMAGfyjYOvRmsIiAH4Pn5wpmz0mDdweizynLaEw9gq4
sZ1PoKS0VSpnz6lcGpLlnxnYmS+lTvakdCRKqkRSFmVE4gQcbFG6dyikqlZSRLH52ZK/2hqUgYt+
p/m1OmpDXbQ3STS5b/O09rwTbqaP0meTEPGFkKPRrMAw1Rl6kWOMti5LK7ku3hrFveGBAuFdRiT8
TXI9P36ktFQdbNM3Y196JnJrLoJGOQr54sTepn6rUlRboGcnGZMfrlfBd/WmeLkCmWcDKsRFbEHO
8iS0YPTZbWPwrnvJsORBUouKx6iXmKpu6IJG3OZ6yccfKOLRnCAcqs7RgQu7eZ4dikukq2g7h1yx
FpbgrecynWZMWLTOSPV2XOaFOQ/GE/XsLEX8r9wLZah1Ubvt0mcotY/UyIML9Ii6LeH8OKX91tt+
FdmlTs9vsLO838YBcL/PICXLZiIFREfnh75HdAurYQVcmp0BQrX31lWrNnhiiOEmBboYXot7rTF2
joJN97UXWLhmylwelvX4S3TvucAgISwH4uihHPuT6CK3sUpHPU8OuW7VEMPHH2xiKzUk6DjJgdm3
UVYNAwnF4ScBpkZe76JDjblnAhTITg6lEYv0okXEvsrJiV8pyFS/Pw1p2d39K4MNRiXN/tX6b651
l9aGrprXjyzjqYoHAqY6lOZWvOyeMpx0a0dlv1TXCiNiyJ72hOCEXcTxf9Kkc2dN1bYnGwwy2AoK
NAhFVC8b9s5+AtU3/cF1joJYeCekG9Xg8lCfbO2Bx+yWVJdpJ4IyXz6svU2lTVBXgbELeG2Z5j0a
VGXNv9vVjVJF+xL8Vye/dyIJlkGLeqaXWnY9pL2ExpsFe4YPKIplC8mihdYq70hcFPu0EldmW04f
HbztBTYG33As1sJBvsWZGfQXVCTREaEy+j/+shVeBPstZvK/Je/i4XZ49DHjYMZu3ZIxgvSfsRQC
Sj3lAfTzyxdx9llHbHEWfgfSdW3ASTafiYwFMA0qKbAC2KCbdXQTpQUw8hmcPA7HLoir93oRyK+p
CENeN2RvjfV1/7OnRd/JtF15k8h4Z2tMRy17ltHdYJvORH3vqz9AlxLrpMMifCywkIZhhXrWHpIw
L25dsSTQjjBQr4d98+btq8ainHydFEnkqW8eG7FnbYE5d9w7gZFGXqfNr7gc+WTqcdebUfdZSVsf
hCDBJHVHaEjsy2DwN8deshxpNXrX2V6JKjqu29TQJdzmIalGiRyWXYtkAUZgp4W0sD5Si4d6DcFQ
pRX+/268MKLbAmKQBI5V+8307LPEJKOr9onaSKvtLxajD/C+Stzmv/snwUVHhRHRVTRiK9nb5bPe
vRsNw6L42MeGBnCPk4dDsScypQoukLUUT1LX1cJR1KMAs7GJeJkgreg00z051DbKZcKtevGpkrot
tuyJ2Xo9J47yncdB81iO9BSDKD5S+CwDCklehGGcq3sULIyLSsRT+o4RUlUPqV4stHvzF1rcu0BL
y+d604E52J7Ieg3W0E5PrJKei7bgv+LajB9YCdaYB8CwAnDnrcF6bebJQDzgTFpro/6QwpWoCC49
aiHYoo8ZwX+q36zf9dJXq7o4zokjyLi2NKdDZdBA3wFrHSCCOl6Gd7nV3GY1tzVNfn/OXg3dbG4A
8qHtuQNd9yd3+3Nor877jklSd4HJxhWoig49FOHscsABO1vl9Ai7sMHAk/e6M8Rqwe50qvyGlSnJ
+MEyaNv1O05nJ+7lj4hmze6OEQgsrwKzwU6OLaIo2ANLA9HW3mPw0qNc0DMYuR6drT6kG0GjXUfz
FP+KVI+2D+upPLx+C1bWWiwe2ISgkuL/fPMdjWudZtkbuPc69cSOp8xxXOw4qARl6NxwRVlurp5b
cqev/5P4KbBSz8jIDAxmoBDFxtHZrmmT8XUJHP5udugZs9i/sHc6UZ51DYOWIuEYN9MbrbK+So/H
uhNnPvtAR+LoHI0OnkvtCb3v/jG1m6VWTVP21RL92W34GWcaKJlDHtkFHQ7reLT1iG3ynCUPBG59
pgoA9LxnBHb3ANxogwJL4DxSAu18fEyE0o+xxbEG6Df710Vz1EofLhlD/rbhfbO1kKO4jVB1KKv7
cyIg02YjTcrmXyAcA4eS7B71dUazE2wOMeCFN2D6WVHwp+FwUXgJqouDJvFGDZVU+cnrVM1G9QSM
Z8CtCb2LEx9oPTDnIojGUm6NT7grpG14Y2Vd1xegNF0UHi0j1YsLpT/B9ri40BfLVpn8gH1vVBKn
jV3bN65Wgo5UYo28DU0NRJ+LV4KMvqf3cWFBXM7/Y9wkvic15fJUXa1dWIX0xaDA2+wHVl99u2dN
BPSZvbh+1YyjlGgbSJVP+G6DNRpXZJyqXYpIyiQlOB+mg06leJYvKRJ+DKVHZBBO0Uc5R1E/zHCy
bBGuk0jEJQZ27ydXXH+QhMC4geIoJE/xHU55l7EdccTck26uenfGl9UTf+doXv5pMl3I/DXmRFcA
IPBPCPqDkdxhK02kmrUSJr6SdCDGPmO8DDQaocEkKm2IVhV5SOZs1Lo+LT4LXdkDdAcxXyelGyzK
lIOEqpca4qi8v3j6mghD/sYRwj8sZ178+3tufsDYcjx1wpCZnvOMWLvKF+hM3eSn18uONeF/6V2O
4DXZwK2sWn8IQ0mMNf/toNBL17XjL1Qbnir3HZPC5g78uZ52vzcrBWyrPx0oZQk7BAtnHYEGv3Jf
a1RPrnEytBBDiz1YrnihlhCKUH7Z37shg15d/H1NHpdMDarw9NNpg2+h2ldG3EMQnEwy9FN7apkR
e8CbdyAcqSx2nJXYA6QQW37mB/YMgAK/RYMeND4MvVGCkWGCopJOtWqnuebiijd3XLvtoKOIzPN/
yCMqqqKGi18/WPc8175wCMolRE3RObNW5+4cv71YK7oTMCSDxssMu8v1VL2VhtRgsvtOh7FWG00v
QWBRPLOyrvZUPZeUqj8S0Ohi9G4JOttoz25XMhZaTe2CVdQW9QVepcSH2rLIfAQhblaXoAfkLNOg
EOltfBFe4Vl4u/sI2xlXtzD77Huwx7HUMluhO5J15FsFS4A5DQL2XJsbLhgsQauh8nJ1P57keesK
7CA4gldMCfBcAAD27Q6oy2cHhlHIQBf8Px+PWM4irj99RfdyPmdgxzH7NHS8CPkTixysXmDisxHG
3bpcmGJH4l8o4KxQGjrKwkCvzpgtk7hwikxXUtAqQE5cEjf5Vk3Yji5l7lDzieliuc0vu3nj1dh9
h2oFlXlMVv+OcXjm+aVh754HCvneA2h0YRbubBRgKyv2nKdU2r2F0SE0K76T3lpNmIYcLX+Xytis
cfmksQSUvJecNNVRWVmrzBSSAj8dplD1O0cYjwkJ9bvrYtcER6O8ZRww99THAEFwH7zPYTgIs2SS
0veDfdBZshhoS2tEFGnG1ykC2FbOGtRfjfjc6BPZJNCUD7k/FFHhdcs4+hCOiU1s0Z5fFXtqx0nA
8+iPf75vxqoBbwFFUWJMxSZPpom8P/uBeaHyv/rRHQicWJ2QvVeMKS01H+Ohme2D+wqKVasX54ro
dQ57e/edwMVCBvNBjqwsJr/Gx9C90uiST4NHmDfwHJo05K1feeo1GrxrXcuvSKoRVks3Nm7qcusw
lltOlOlpZqnrMbFNfbahmmbmlQcqFHC78fOHotolTxLWsZy84RtUyY6lUIF5ClCPqw0341WrFZSV
sH9QM3eYeupCp8JQFPc9fayfp1LT0ksLpoMw/q93/qq4bzak2QpSLqFSmvNYkCoD+zIyVqIk1HG4
0HoX7xrkEcb30+FHQwgz6ghdSLje4T0cHsuhPrpdJixzWVUR22JOI2sZBg/ZHmhAqgf6W8048tYA
HqmGon06QVBIoQfJtZTCswn6GpRHGefm5BN6/8qd+Q+RtXLao9SXyAyGRnJVdIWQbnNmcTgkNaRh
lRC9FFWrSpu110+LzKBOLdu708BJ47SDEI/NL73p2PlSvmjA31Ww1g+kDsylsKAmkbJtO1ION3VY
zxEds63In1IQObu3K5yScAME3XgMmgwVKDO+ENwGODg7mCEPhRLNwmhBJkV598dElhBGO1RHlRNA
opznT29q0ZpUydhq5/tM9bCIZSa9T8mw5BTBC7Z0hqrZiGB4EyEfv8K11duGrqzDIXfwFc1rsjmv
XxZkXbAPyeGrp20cyg6YktQHyHZKIJ1fJ+BRTUu1A6bAwGYQ8NoC8zdMAJ+BOGAiY7ovbzDhEJLW
JrFBhFIrcmm2W8hmJgDBKdpsZCwa0Cr7ROr4QLglf7PKHgSvQZJnO92O+a/yPva5NmzL474KRsGy
vUm+OD9tD/mj9uAdYddblgbTiR3ZXm+/BI06Tdo9bnBHtSkeUsfvOXkoiGG44VzixhFcQk00cpfG
xU9cardpHu1SJTIyvFHSrBlUa4m1ZvFmt9icanlbpU+S3lsUDm/itwAXT4A3WlRVvwBCxq2YUuuA
QG3zCFZa9EHP+7uecyRs+VO1+60jdVn66nZfpAkdJ8dqv39QV2m9W1JFu303FoyPz8Krq8U22rSq
4queucF20m7oZVnkkmHCV375Oglq3Kw/3dY/XvW+RX1U9eeEGrlLc2vMmX0iDwjd1liGOX1F16yN
Ye5vq0GTbjSP8HyNRF+Hrva6EuzEEA8Y4wD4vDL8d9zerPbjSj5KsDOYSj5L7Bkd5DUDHygkJ2lv
cuGYMA7HdP5T7UrYN8FqDwYdzxNWEG+imFtjcluCjj49LN0jyUVCLOWdlFUwt2+CkdqFzssdu7JA
JvH4hYqOfJYq7IeW3d9wUWpe4sKEUv0GOKhULtIgGukZHVjX6X8Jw1cSfpX+7jdXPr+a3i0hmTaM
iRe0FyG8mPM2uR2GKedXFBG6NagRHRIevNPlaSWGv2xBp1LgoFIpfL3IKLM5BejXhks2NaUYp/FC
N/fB+zQHjRZfDn5sHCHaVKP+IaPG6RbU+l0IsEbUEoUn5M8KfCq61LD8Ep9DWDRTcJklAZr7BCAh
7VqmfaTIPNgvAOxUJwYyuzCRD4IOsYKtI5oeKJqFWtFZ1OfB6sz2pqIxi7AI0pXFA8D98eeoRYep
3sPvNMnJbXzy4ZbL4eAU0zFV8dob6TY3a9TkZPLGbR16YjQeJmC8gqKds25Kc4VI7NTtH+7atnMP
iKyigMSNcrPhkcO2vEQUZrjopTIGD/ABAejysLS+fo/WD2NdKMb6qurtHenxJSwblgLjKyBJ179r
xuG8T1ybsRhksGBYAR5Eygu1FrfvdkI5f0TUJ1usObsrc98l4wm0xLKgeqm9zt/QaTBIxcb0r6ey
EPiRvSekvQakhuz15dWFv/HdDiji+gKwXC/vYe267KMT5YLKXFsB7dOmqALrJ/dbyIVZ3rFfo79R
QoKWyA4iNhktJLRVTdeBdDWoCCecjs9j52ogBG6wqns00JSqj7IedcgHTeVupyEROMGgwHjNoVqv
sTWVW0s0+xiCuTJqN36W9CNQyevqRlVarJ3cVOy0+DBEvc9Cej6wp0urguW0t4L7Q8FlGkR9019A
2DqbX2LoBPDzorgKmwe3KeWzwrErpKwDznwsEtlHKyv0wVGSfrfC1vCoqOA8pKNMo5E9Vlaog95d
E+KyFXswaYZjLLEWQH8JOhKRFpBwN5IKd3n6F+gWlKAJO8jHYF6ear1joUeIdvON2IPZ7GjwCoTT
knPYNTUybszVeZrK2ktooijJiTX8zX7bXJN8tqntz7TCsaVorrt+Jsj7c8kw/Pkq5C0uKYurbGVj
hWPqgm/ggwGyMEjiZqa49h24ruNmCnV1O1YIA4LPIejtGr21GCWeH9u7zxGU4TyiQ6+ebW+/SngF
0s3140Ey9TKAqxuWXeoXwHMeBfUyLdhu7K6y+p3Y7zN78clTBLH9PX3cym9pdYVbVTWB43skiL/4
ZnaznByZzQGQb96QFbpb/o6vFICqLUCHK366N54L5h7Zupy1A3yo63BT4bSlmzfHp7w+Fd4VEvRV
IzfVem7cp1apv7ZiLIa+p1EWeabOS4qS5uSnEywPDOxumABvf1UbTnxiFnZ/x8PlFcSNnN/kzrc2
pSg4eaEv2raFg5WldKCVvjtA2fe/9yQCkgJ76aspJ3/NnqHBi6/qWi424qunrzucjfQTHo4yB1SN
M8vLKEVdmgNiMzXCEdNQhxlSsOaT63OceKGU28SN084khGkVY0PtAfnYGcoU3/dNreYuSxzHk389
y4MXruJ+r3FR8lvCAdAHU5XbKBItXPIUiliU0i1zbM8aD4LkQYTgYY3oVpOpMe7poTPjWxbeCe+4
cDYDD7B43l6Ll8BnIEXbCgtGq4CHCi2gRZeRApp/L/RvLDDRA8YxSWgYwh1amZiv4umHsIYHuvSi
MAR/MlZTWQsb0AKKxWEj2etcQ3WFuoqKRfI0t8+2MI3pHq/LA3mGa0Sss0GcIuwfg6z17Y+7U1bY
NyQb2moLXZoIuVIeHurese9EVLPlRcHroTopoBKJPVvAm2pXYAVFCBLUnnokp0/xRPeP9GkLhkJT
cEcWGdgcbftu+7vyUWMLDgK7wZonHlSlsPufaGIxhb68011FrVVfMTI62ZCrQxSPHXdd7CYJh5y7
0caUZiOI7/d2aM/csSgyebtIwhH+etkQz1VkDmbSTJ83dBeAX04Bel4VOue8xARG2BI+XppymUaX
cykXXvzb2TwakemfIchzHFAN2q8vy4qNOoGbY6XM8BPt3j/dpbId2uWrGTL0bgKOiAcW3Z+W9o8F
XeQtUbk1RWI9RSiKvn7aTTMUbDwi46y9rT8o6QZawsPsvFS5oJctZ9YuWfTi04T8GiGmbBh771el
x1AtTGGU+zqxKKEB7oSyXsuEM+lPTWAiyMidjeNSL1D7br4Nwj5mcvgS0j50z822l2dgogQN/Lsx
+76V0jdDkhZS7enRYaEvspkhrJW7Oyq4qJ56Piv/VMbORziEHKwDFzeSKMjiRhC1r0CJHWzi0DLi
QInb5kTNKpNKzqk00ivnBCtRvKN94j0ymLKYAjVD5nKSwXwzVCGroTd0ujepJwox6D05Yip2RK9r
XwTpH2zi2SldBHWw8g3M7AZKbRPOyges8ziN4Q7sD5brr8WtAeSwDTqY8f32MRdJ1cjrQqAEBMVB
VVe0oYOPwth9BD/Jybk9iwWQ9wf9YfUr4aZ5UC0aPV617wBrrL9X2p6Vpj4QnWYVJlaOb3b7W6qt
Skik2NAg9AzouUvgx/SiC2VdYDdaIwpxQw4gW4D4EJ9oQVA0koIG+2RbnyKIhN1gLLrdw8ORha0M
pRRD/Zgo9tFRVTo6ThVQSfimwbqnDcguRMJXCzPdhY6T7YJ13mL+DLJ9LVC9X4m3b2+c3ARipAdq
cVjMd9CNK4UbhwmzEqeWNcaLuYafYxsEnep7QGBYCEWTMmkUjl/xZu1qw0qYUp5l/t9GtCHkOkAy
nJIQd5fHvcEVnEx3YLj4lrpdh3YZB8CjED8/JqajCC7r8nn+UlSf67YI3Cf2tdbopVuY2Z95onKM
Yn5sjtYgzyR6zZhcKuY9bT+z3U9mZD444MNqeefBXHgic5nfAV27v7BSQE48iupEUVUQtWdvgkS8
HGiNmvc1vIfmKA7xqVdKxlyfW1YKupX4WFc5qYtMFg1pB8WwyUA1ND1l/Mg6XThsXVrk07u/P01y
S3V8XQULd7wyaInfzmQ81lR9lmO8MW2020LIX0DjRiAIABirncgEjdmJkr1aAnYl2a7om14W9CQg
7GLdpCk24mT0ju5ROW0W9Lda7UwMfm76C99hK1EJcG6G5zK0eIor4GLV+ncvdE/l6eFbKo+FOg6z
HX5gxRCX0o6BqGGndL1LeQuoxPQ9Fe13xbG+TsEu1ALsjOWSq5doB7pVZcavvW2JNjG0eVNIqxX9
MO4oVMfSgk5b+QTVhSFE0wdcrfs+vbvFUae6taGg7iVjDrX3cCw0AuwEgrFbElo/wX2THX1T+tpK
1s7accLkk16YvLiKJbOSHRhWgnTdnKxH3tpWrbOa9mm9+yd/EwFSzneuIMogpYAA/GrmRW5SOw9s
aadp2MbOrMiFZoMB7VX0z0eTNmdRx7PxHPF24Ou75D/f4YdRoBWkbznK+iuQLjkyo38PSJPWNZtV
ihm+Jz9c4Lt3IaELwp+DL++xOPVI8tMrlwxw3EevzgsfueW67n5pR8KzeALbvE3YWGQO+jdnGH0A
GkCTKDJrDB+DbSEjCg+n6NLoNRYvSazkbDs8HS9wn1lSUE7FHMUAG+UNOclEx4OwneUAuBVNpzNw
URUhvHSBZq56n/harOB6lKOy9YhkREuDz6UvloekZo2JR8r6YEabQX3rGimg/GjnA0PdJ8SqXNuF
h27duPNI0CTds3bNzVjmm4OUQPkW20H1pwFyTwpFTjFiexgD3ghtw+SaNjiQK6QaTLid830TDZ9O
k+tj+stzPkFyXkA4FhQPRIAiu6rVxF/q/WabSum4/0ABgnkTMK2zHQgycoLT7HBDCyULHBpEhymY
wl32qEqxeMdLTgF7wk2hSoNalNHesbia7ch8GTjT9P+7RLtkE0qazUxmHpzHR9Iwg5ovqWa4paUJ
L8XGJkZPZxHPCwUI5UPBtHhufdFx+2bfCCItFVGCYFcejuG/Rqun+Xug7SyrbL++OIPjhDE/9ytY
u7ofVE9PGjeZuyJI0PEkTdDfMK8VqlY76NzQw2n7YLuyR8kJWa9W7dof+N2DKI5+vBpkDAdi2+CR
G31nBKaisZ5sgiU34Pv+ziGiVhGJ7Zkc9p6QhFZpHZQos94XbvG+UyXl/7Rx0o1KZqitiyFmQWey
7TAi/pCXzh9VeNwUbekeTZwRRL7mm4/6zSX/dbM4iiO8x5mzdDz5x7AG2lE2/bgUQZ2Sz63Frn7j
rbFWWUFj9oPSm6B+vqASAdE7L3lcM3OhagibMxLcwLylaviuJqsla/fK+nLEsxDvSaU6idNables
tIQHrFQd4SKcTFPFzu77jzK8MaYH5q3bH/wDIEqAY7LR4g1TBHUpLyBhnJU0uur5taLyoo5kAfEJ
yoesiywof1cBphAxrdhVDBlnysiHYSLcwHUPx2qnAhs+ZNdNBeYVrWW8CYbD/L28icrlu2AzzvJD
towVqE9uAW7v7uLGLHxTdRKlz1IP9zG0hLbqPOqDXtMyYga4pMOgBCw31CmbzqE692Zgsa9LTgUl
mbTaeq30jCVf1q2H4Oy0Fh5CZLasZANeFFbh0a6UVYF3+kgAqn4+3ZMqzOx+PPP00S07XjiZaDsi
L5kr+YCYamunPzRMhrQVe0p7gKKrn23qF45ssuobrOkZKcYrZ7Jt9RZD4uvQkmcd2M68u5LJ3xCY
aMeXMc+zZHs9VHn1tTQgoyzlNd/4eQbBeF1uX364PpErLcdURCbj8Xgz6VpG+g+64JBsQqOyU/zJ
2qLkVr8+fpXDAObMEeTtUCBshO/Ov/vV8A2j5jEYM47VQti3p1moQUvC+MBtzEQroGVQNSLuLpdz
QtE0fSA1pY8hA5a86UR9beJG7c8TGUox7DGH8LECKQm+MC52bOf9k87wihQ60pYFLCvEzhAwu5Sw
Wi3jjPE27n0YMqKtc2IbwBtBkUsyL9zt5xycALbWX8mn5Pq6/WX4RSCVA6N4wlBQamq46ER+plN2
g1zaLgC/EGUTZPxIeFAQ8vxuflbMT17wSENcBsUCC8mg9JNvatYYxzvDKtt72N+oGTRhege5RfC3
eyqhezSlKmFiu+VJhMT5lk3i0WECqiPf1dXd3Y84gKircmHWxN2co49jFwVq+IKihef/HilJYFH0
VlxZe+GA5NjeuedVP/m4GHI1kYfa0naO8dSb9MatBzWNx1kmKik2nDfufZPEo/TAsvvKLgow8Ixs
fin0yNAu6TIlkzOhEVm4d1TuosGnr7lQp4JCi/de678d9qr7mFa7Y1GkbEmxPPFaNe5S5lW7GEmM
w/fOd06bpnQTYALjpldrV7kTkvZR2VOdJVWB32jf5JfVumpKbXKSDDGOcakH6uXTZdEJWyLv+r6p
E0i5hCxPiCWeWYsPMr742QXUBf9AdDWrP/LmcoqDaXFQxGCNDXLL/DIO0xcVU6T5bOIB4Q2I62EA
xm0FIfA5DVsvOBs9PRZjGBMC14tX8oHItKnchd/cxVqJreKGp55I8MDxQ7+sNKs23xcefMQdFdx1
b59WznpkrwXFzatfYo+DJdSqOtJiYbw7lYauXWq9ec8IqPayzpFJUE49s/TIUtUA14PIzbQHtbKM
+XOOFmhcCh2/YpE4p9Od113YL8CWVZNdMi+kIRPGspD7CxgJ0XbkMxBZhrr6yWfFm0Y11mQcozAQ
MCBEnrUGg50UiKg3yw9oglisRF8goHXwODKuRASRaCEPVvqEVnFvAmyMX6EEnyP3p4+wfY9JRnwb
IYZBLsNA3fELHZSHwNxBB2JENd/9wiRt2qbex3qLnefwpq55FqkA3k+z0LPpjbjg/rKVRfBeVn/W
ajADfLEFvnaloth0dxVHxA3YTwEn2OVIq6LDR0uNHR/128AXklRaD8kG+nITDb8gpM1XM4vAsDpB
+KnBXEcPhqV02dRjdPwXXgfhGRXVBAi3k9iwwjk2MBtZeTqjUpoV9xJ2u8Vd8Tp8soRpdnYtC7ge
KyvrRe47ZiUj8KHdcGHeSjGbXnYOzpPEjYI9M+r02s0dvQibwW2VdBmP4KgGoh9eGO301ggbSXKm
lLDmttbFVEtp2Pk2kO99qGgFZX0XOMh5HCyBx5C45wUbiaWPnuS5GJguLvzUH58FzDFoY/Qtjgn1
igvb0NdeeiPJ8wV/ML1XqbrxOa4xq+FHcWVoiv6A3nsuOtlhNQGekrhfl73RWrxX8eJ+Eqejd2hT
r3RDP02+q5ZUyWRDBGWrfVvKjKIUmSKiGpekXAYq7Ijf3FQcNSq03umEwiNqrW1Y12+xmvxVEyA/
qJeNoM7nPXN1YSTiWhGE1j/CYzRlH8jq3Hw1jWWN4svsegU/QhpDvZGgzo8l6oxJkl6JMI9G7d3O
voXI+1jpfVI94MMAHSr62mNrBXC2D0top6kwpFxwFF8cZ7BHFL6o1rhKTSn6g4jdp6vQGcNc30ol
N9YylrWJyyYVUNqAhRlGcitswgH5qzesOXJelMoDSRaiVlHWhIPurv3KdwRcDpVdpsclf9oKfV/6
eaJGYA/J2Ei3qPRgjkuBSFIlr+A43YZ4jYlho5nh4fgqAxc0P1M1s5tiWi7PCM53aeWgpGiKZpp1
vHby7eosI6NP177so98TCKAjxyDyvS2uY+C/GN7dpDc/indnGZIfGjsHtZRWxtAtnZO/Qh1Z5hos
A8mKX+q4U+bxiraoivLfNMQVuDUPMOoL+ZcFD3d+ZUepiorseceiVd8q1qVF3II2vmtL5QmZWBFW
D8cH9I+KoYzSJE3iQwmqyZ9DD7vFCNjsD7SzD9aa7w0iddr8sG/uO8o/imM+LGnMQ2wNyMk5gNAY
K0m1vA68UYOeRaZYp07JbE2CFw3nvuyIKJx5OFLbMs/qonGnlCHD4YesNPEQ8sr6cAEuLIYP9i8j
Gm7t/0Qra8aH733G/m2I+OmbOn+MoAo8UCOsjjuvkRwZeAvjhn5iTrM3fODOu66IYk7OKKTHQ6OP
nwpetEFNvBzfqeKboPLb51kdxCW+iuAl5IPqglc7/PaeL6mq+zW8zuV25AHZWOwMtGdEXiGpSZCE
gCDKU98JbH0snpxEvArRimJ3dqaZd4CA0PgP2z0MQULL9iA73yiHg9C94cZzbZSscmJsZzviIyRK
x+H2wD8lDiJIfj4TeZBt4vRLLuHLcApPK/pYq+ROYTKSf3/KltIFicA91uW+zWgF9muKw/Uke4dl
1bpiTIdOm/EpSR9ixi/DDS8mJXrywe5VJqG8z7wZWxNP9adH883cRLa+wHBDpFgyByZlNRjoZ76x
Wn/ApLMSZQXrhNVJDuXNoW3mKpQwnLuVz72Kxra5xe9XjaXzPcYdlpLpLdGzgqFIT0LBMkV/JXQL
A8C8gV8Epmaiv7G8lQwiwH24xUOcJe1OUlrMjOI+inikrB+4eipTh1XRQ5ShLSv+0h7ukMK2CtI4
yhzk5pZw7k068QAlQQJG+5zYjbDHtHAX+Rs4NX0UUBZYxWUO0bl5OcxTI4cyDlj5QWmPAJ4bBykn
vApt9kKOkuNmuGgXj5LT4ZYlT7xuf88hVopZabv+ibLREWE7TngKkKoBUfhQLrMNYGYoJ8GvXJFP
I2+JxpSFBzVS89ExB7za3BD8nfV3Il+qs7X1iy4VpgLhr44kDi/cZ9hmsMUD6fuwhoEKQ378+3CP
bZN7/rfEke7+zAMa2lAHvL4TArvp8ZaRlyXarFcT89yL1gerJIt5qvMku4QAWjjX87pcSR/f8cUc
PtUhRVpmGMLU8szLk6Fmlt5+2uIgiKpVut2B6othDgH0/wc1i+zZHTqFc56WMm7wY1STSouQmyD1
bg6uGbaLTPv17h0WjzutLkNd/KgGvgAQZdG+QVo6+3qLlLkWs8lkJX9JeWB+vXOEd+QR5zHpKzJR
QdkOPkUFC3C1FkhxDkxEcDVub1v6K1LqbEiZw8Y5VjG8jUUw9k0mkmCbZoJ4Du0U/ATByK52db60
RuOyhHMNs86uVD9xyjFJvOBEVmOkLSm3Q/x2M7u1rRohOdvPfIN1Js+Bu0kKO5wReIaNB/tD7uFt
WjSFa1bL7+FmIjmNtt0vms+z5t5sjU0ox/oOlnHLyA9U7PTexTYd4+BpS6QBefsxMhdvqDsCI0XC
qEbkUOxIOByxjUx2O20SbyFdkrh4G+PuXb+0yOqhytn63Dpo6NGdZKzOoLdPNVpki+PW3p7I+qrT
pdIJuzg49O3fK69w6WcM5EVNPc7z/vZn+qrB2XZkdg+6NVH2TUYw1iXBpyv+Xwx4lDgpaA1UU/rv
dV8G5js+2CmyaVOr+K2PFyffBVoz5TmXHAJmtFt2bKtmRoX8xNaMt/mDBorfP8mE/etcWVT2doeC
6xIBkKWDYJwrrLn6uU+Y3CaPn0MK8YTUuIx/rpzZCbPiqXsV6fMNNg6wWSfi2aoh2qwjPcm/qrlL
ME6vZt/fYBvr4ngHnNTPdxQkGZM/oQjTOLFW3DgHGHX12/Y32t+3klQf+xPpCSEZaiAphO+Aihim
dhjCmz3mgDyl1obuyWcAVByA4ey6WVzXu+gO1iOS1GoXzPs0tHzoWj1c8+7Sf5i+Nr3DdmJWCI7n
ER9p/pXh0vA8ft+uO0eMTDH6P9Xw6LZhg9YKcUXhuMywWgTsg6KHfTA/xx6HflVi3JrcDlQxGOwM
6S4ryjojoi0XLzKQQzYYGeYgSu3xwS5+otluNZCnSftaySVhn3wfSEtmD8LnqfigBuKK41wNIIER
sV9wLOI6X/Mef+z/+qGIHm5kNW9rXL5qDyk1rISjGblaA5qQthLAhjBRl+nF/1fud9fqtJaP5emS
t6iHu8KUb6a5X15L+vezbjSJURsq/oKPbj3RUsnPAgTf3c1mRljYbGhJommeiikdkwe4WV3NARvZ
NNfxbG1Y6jYpPCB9nIcoCY2jhnpbILRoZeshHdg8CsHmaI4IoRLhY5o6YbMbLsHiEH8i2OczqKOa
hgjSqmJBMYFZeRz3O2sSyeHedqT9qvTEdtVweR9tHBgKyt0txd3+dQqPzSg5eQDaGuJue+iIOEQE
FMNTo3CyXMNXFkyZDkhjVaYnEnUBRpPSJtuZNeK5LSWFexZOEtxNX5bxg1GsSLdbSWPU++jFm1tY
o7K6wqSPgdTsh8QYZQD0nlQO+bIRM2wOibx9Kj9ANTHfIP3xjkT1Lom1WjCc3SuEP2UjKEHmQCi5
upeJkdlaoJJ4Q5ocFPjk/v3HoJqBq/jbH/bCLSuJ8cGXBUUEbftZ6UT5UV9lNb/Hgbf/JLNkXMjR
MkHdNcIL42nualUXmzHQurViflTC8DRwhKWsTtyYLtukNBDjYflw97tUS/apDW7ffeoIxieH/ckJ
D0qbEOTn4G9atQQe5zUDKmQZamCUB4kjhKTQv4jDX607IoX6DyJOtZZLbeiTo/TdaosqjaQ87pTm
j3/Fvp0c/a+8uex0anS9gW+2POMC7xc/0UIsFGZQYySg0ilEqKJQD4IksnNOpM8oZhSyWzw1a/qW
cNb8TuPmdQImMcqwZA8NufQeIqivlBwiR5fYCiSoEUrXgrwqSUzH/pxktczE3n4D8yfZSH8gVpoz
VKiCLnsKrWPLTWOE+89euEP/LiwyLbBEPvZKBR9pfT79aRlmkiJVIYy79jBjETCkKMil/HFreJ6k
7VN16a1cZWayp1ixzrQkFpVmhZCwfrKQBjlDjO7E/oOfDcyMgqW9xXP6giWlDCH8VAa/TWXncDgm
2CpvMU1dbPqFgGHrbky0S2/IyayZEK1pvOWaXGIBsEmxM8VClSnMm8GNspx+Y0vwHIE642LnZJyu
c7ggzrCdrqNGx/HVsQUBGQDJCyK3i9X4E+fmE5bZ3cvWz1O9UOnrjDTRkKAmJ1hC0a6BeJcLYDiF
ufmCslfMG4eO0rE1OaZWrohFS2Z4jY413yLHaNR7xwpN+W8/++y9YKT7t7V/S99B3xWJPXKR+cKI
Tkq9aW7NixYeJhSXR/N16y9Xcjfpi8nopqPJkQqvm7b8s8JawbIEaiBs3aU+5RPhSvsbWix6+KfE
HarDnLgfrIBUf/jrOQRAckq7jlQ5ovFsgh7chIfAbMr4x+JMgQB+0kAzWIS9aVSt0hOo28uBvObC
dFRfhiT0SiHf6vOWIVj3z7FHD3p0mLoN9Wao2nDbaBeie3FsRJwCmSbyzRBulJJlpTU+5ibyD6tS
VwCAPbrZJYfae24z6x9zYDTRD0MNAYmj2PVqUsTyaS8xSJ6QxoNtoF8O8u382R9biowD2CcokxWs
Lr88nEcKsLf0bYEDrI0IX0A14fKmDf2bCP/vU0qLdBVXrqmWmSCuoEPpriXGRyF67qzrD09Yi8xJ
SUr1AQWuTF20JPix/sEbjhyUZOnSB3a+Xop29mMIPCOUQU+29IAuPrqeQ/YpSTLZ5P+VQQA87TUD
tQjTre9j8qk8x6ZOz+3XARI3lNABfssTWRbCD7JO9qVHN/czMuF7hkwEN8TR2BmlWrPHCnS2Zihz
OCTdSaPFHWPUY73rfMsjnbcn9oQ1xD3tMEpJwi96i8sO9eQ+In5/aX15B65g19R609lEYB6WXGoe
LTAVM/bZV5KTw2VDQywkj4vMThscmuyBMu6fSVDkzj8sRJeynLUr6MQKINDx6QVKFu9NxOvanGXX
ZcYbFZw+KaUH6xJZhd5J9SPBcyW5kJw6opLVR8gKrqBhwJDmsFw0AGwrmnQ3qp0tFJx6EqPc6eeJ
1FbsOaRy+m2qHrIBZzPLeVqqgilyHnVAMYAtKzajC7kxo7gvmz3EPT5BJk0C00jndahJWtQ1M7P7
NjfDb+fhtC5QWJkiKhTylH1am2xXrYybsG3pUYj165M9oMX3WImvnCZTvkW5iY1ndzK9osQy3en9
onVY5NEUUF8ZEN9SK7dzumcOcq6+32GJHb5qLASbLek5hQlH+uAbAOSDEwjpC9cCnmj2XsxjFdZc
LYZpZcJHjWjvECzMWeGb7izCR6pm+1I607fqmkVtSafzH6RWzKpKzX8/T2gyLMdsjPJJp/2+OGNh
pnky3f9UalNAL09HniAZwj38/cpo/7kauT/Ls4sqoiMR9fotmcpXQ117iPTirqcIHpQWmnpZqYom
b/QKMc4+qNaqtDLx0i1+ajedYoeuXkwXlBVB/9rtWQ7qGOnZiZmmF/9Jfs2/6KBu3Z3fzDeNZ/mK
1tSdSmS9vS174pbqeFojdtAV1P77jS/+X/on9GMeUk8AHOxDx+QudRamOhrkrp18BZmwuGw4wPnp
SLWmtHn10DTCjS2PpV3z7QG3aL7p5vB+dGcUtzyWJsrjrEX52NMkiNtp249UKeVGypf8uPwpuvvU
bwAS/FRkpn8BZAeQ/UCh5WZ4YFikKCv365O+82IF5zN/pf+ISnUEPQIGPEmcVpmHFSv1yteDU60F
Rc8DJfw34oJlhlO8vSgWFTX8ZLfEYRswkpTWN5QJr3VjHF6sIoGc/aM3of/IAP99jA4bWKEuxAvk
0sFUrjIPRwS8wJ60IhXCVYVLvLhtHIzEcFAmZSNZoZMTAcgB9HU+dsppzY0lwt06m51U6OlWEK7I
YRriLbRjM95vSZdkIvr65K6GMtcmpMTNM5ZCBP+71nABb90yLXzE/1XX1c6dzUZp3Y+NFSDoEgBJ
scyMXT+TEJK0USJ/8qEW6xyYD/BFobBe0GeKoFbOQTgwsf+FltNSAndAGAO3qtn6EE0gsjVBy3kn
uTunXeA0G/bMbTejJMhF7xrjUSowqqpW8A/SNV/UZdeQPL13/lwEZ2f0JYRlfox5fGfX45COUbzq
aO9CV+F7l6DfiBMWAZk+5ONG8g9vZ2qjg7Fr75KzOLvEh/HQF/Zd9QK9+0DpWLUEJVXcPHu9A8yT
TZ8DVu6j9DBAu1nLART4qKs+BzcyKF4vB5z6UuG6/M8PkNnIsFTwtlvH6AZmsSa2F6w5gZGhP03+
KB60jqgMARfOWPUuCb/FxL0nDed0nBxmVqsBG1izH5QkrlxB0iS7FCgTAQhczR1HpDwKgrdgJlz3
kGID8aXICOjDN9MDhcUD56aKM+arurVknD+7LBzA6mduyDSbZjdJ+9vuqdGV8mycDxvZbzioFLpO
p0ZtrClBlo9I4DUeC8abf4CwiGzbkJJR4gKbpKxGxkvB71hEUcBg5jvD3YJCS14eiku6+ptRVQJO
wGyv70vAaBPa0bCob22Lt2vzjXPTfoaOKoSr4h69Xf3S0P7AclqP3bCKgRohcSVxwEOyfdnjP4k5
W/AGke1yjCyWhDnHMUNnVahwgxpWKXFrVlxS7r6/ENc0Zg9GCWLCstIITXY6+9y6cK2nM8BfT1rV
QjT2k7CTFU6/EcY2vnwCwlswrWTN4/1L/CxpprqTlm2iGCRrBfque41aCtL1mjLdVWQ0D0/i+q6r
Ur21cOa7uG7ElHs1BRHHT/rEXT9lrun3TZ4uPHsAWYc+i4N2BaPTE+J3mgho1FnQtxEjyJYTM9fX
O4da9Q24kKBK61oyaKts7j/C2aFdQOS+YF5DwcbAC5kaN179fwt1mawiTbBtEhSK0ez/xPQSDWn7
8wiYpzSRz/IMlnR0WgDoOnnsou4qGlnF8TW1lzHDTgXEwFbbq6FG2C3sQDX9MFIJmwOAFnzhiZ+5
yrV6e34nRUmhupdjAkoN+4qEpbrFCRoPxavikbN8+DK4fmEenrTGtlVQ0AqXaa5YgTcInQTT1H8g
9AyUCso22ra8923vpFceISwqiHasi/tFY/M9y+m2QNveDjH0koZOVMOT0UK2w4NuIBFCTrp7dGZL
B5izf0buKCbo+EWRIb5u51MBGo7KwSkhh4a98haod1InZ9UkJMK7uXZjFgGxS5M5Gxeje6/QOlMQ
vldYOqVO7Y32RN9Gz0ypxHdX6z2yBCOU6kf+gbjYs9mTeaJZCo/0qIsROftZ1o9yHUqfwSlnY4YR
9Z/yIx+ftdIV0xAQS6AC3ME7BmCdG+vc1UUvEoDhLaTsT2fIUq5CwGDMK6YHoqb8Tp73NFbdHgG6
0uK2/DERM9FRk+ERy3Zi1ENrhGhbegOvpkK78UlFUglkGNnS4RaQBqhVhNLX/AyH+arQLWE7sIwl
WQBPHuRc98tepLDIzIsdSas3rSQ624jyLLByXK+Bp86QIgYpLUXOsUv3NOCyrsVU3LVrllV6PVHH
ztZ3EceYVTUn3R651zD7vEMCw7evyokMSTdUoRHUdzOYgGcEF8SoLhQ0NCR7I1SKeaCMNKDheD62
3A9emQYvrtFX97nV4yl0ouQnP3HZaCxFHscNqbcP/qTtBcdo6YPig+qGmQ7180Hr8uAFwGbtI7HP
7iES8U8tcBKr+4LVHnQOXAORDHCDdtlt4DtUhTUjLBTIajgGoehI4Xjl1wMMvjur/HV/0RA4+zqF
xKP+la1BB4hjnS7dAOnXiE8ocwFbRdSMZE4lqNZAUUXvNsFt3z60oSYi8776YN9qdAigHDM2fHuE
H2thE8rkHyfEtMeigo+e55AKB0QyFzuUrB4CWdYW7LBziAiwTIc5qrIqPzGR7venS9LDfyziAS9F
wAXuCoWEN/4kQLhSyTz2yVevqw32Yaxmd11Pr5vPFvk7UBKMNRI1PTpizqKpQtRE1jtxI9vqV9vt
w/gpIHNOp8FBT+zFENJSydHqWoYB4yBBgsaJAHpvyAfVXgVUnou32BbHxStqjBInPMQ1VLbiuddG
h2Bc/5eVlr/76HjdkWBEktcaNXB1dIVfInVbZ9JSJ5hdGN/0Hum1wtFy8C7DxU5uTU1ualOzf652
OE3R8aJMommn9YKDqldoKa4QUJ0wMzy+NPtlJwRtMN/C8aJQblWiUZ06A3DHlo3UHtjaq81gBF7f
ydgunAcFSLBYX3JOndxPO0EtUJxXa0WrWhgbHv6SBdmNXOwMBA5mfskmByGd1eMwDJ693cxSZG13
Y0muQ4r0AtSuP0EANWQEYzAFQnjdwhuqOLwcyABDzYkoNJnRzIhgOeEkmiPqO7Xqa4qZdttlGVxI
vWkolQGRthMyc3Iae1dduxpQXnHLLtCZDWTxd4OCtRqop3vr5DVrcc+9cIi6jM6gYbDg3wxIqym7
/LvrMCcB0RrbA7btYDPgIWJAAXY6tvUrKbOyEmotqK6hEPCpnpPuEJlqOY2D0z+x1GN8iwj8T63n
S0tCtlsTnCmK0fE6Uch5koq1RCfSQHLni6yD5t0i3dM4agd38VIjrtUAQ6rme2ZtNU5rTh8OV9UD
FBPAgx4rY0dh5C8mvQvVj8RzT6E3d1vt0ygQRBxm9XWjjgcd9nVzhOsl5yf40tSJIJWMN0bW838v
dtDejWo2wHCk6Z0Bme7Wsi6tIJ0J9BqegxQewasaXcQ1BwWxhM3+UUbYpS0zqicFE7RVGWFgbVdV
I+LtPl6nrvSRMZjpyufghY+/5cuGJsU30xHgBlzEUu+rjbCoftFtarSjyQ0KTsSgdKXzKJ9uYWF9
dWNENxTI23PeT6GCo0FttgNPS6xiEwa+5oF1acMELZ2vo7Fz0O5qsaNBrelKmSkOJQlq6ahSNiPA
D2qv42h0S6Cnjhvst014mstn9tYMfOg8MrpcoKcAC8StXUJ1xIdRpNBFLhZAuVYowA0OXf+Bw0xT
vIDEvTjA5Zwb/29f40MAuW6Nria06qi9Sne+EnT6eX50wkA+8SXfKQW19RLOAVTCPct6geZNRsnx
20zG/fOMe9Lm7U2KRRqdK4TknQ0ixUNxN0bIwBaQs07M/mODn7YZ+V7PLWvqTWWntbjt+WQ5DJd3
w2GNc1eEe1IiHjJj+laF7f/a5EUK+9M+Tq5y13KM7nVPj6M1TiopRRjCu3sX5pJVuT9Z4a8h62+k
dmvcOF13ILP+Mcx9a1F+lVsUujkg7EPovJreWTo2k1e3ajXuRySt8huxjJXf3GkcCg06zh37pBfk
1y4NhRfAEYhSboOpQl2L1uMoz64X5fk0UXaSy5JR0+lZY+o0HFIm2b/G2WX+GrtEjAkmngSO+o++
JmIb19+e08EfDUC+TSBW1d23nafrPl6s6iRKAqYHpLzfEKUu6VgCxk7CDYtAXOvHrL9pWMRPt7Kx
5Cq7iN1tAjJ6uDhSiYxPH4UqS0e3BA6WgZhf6CJCxC1gevJ+yMd3iVrSAwc7xBRv3scWVyus5gVb
OQkkwxMNdh5SfwTrdDkKN2F6j/BtQYA6Ep/qK2PEPtF4vm4ul8x98pbWwL+4ARxNUIqL/7BUKBD/
HtiGwVj7O8sjA4KrTDyiicuDmR1Vquai9lcWUdpvnDA1Nqaum8TOb6NFY76k67MPpZeLQ+AEHGWO
Ez7CKsM2VfqOGNM0HwDUp0CGOCR6Ca0sCNcBWeiGYFoTzDB3qUSgUxLz9BvwxSygu5SN66UKxAWg
+VDEMMmI2P2GdFhnrVs3nVeSpYuup9fyqUr4yLzpZwKezHNIM29nadbrZftLTuOBFbfbzZOzg3dR
uxR5zBQDTF6Jax8cnIrw6Ywk1iT8bOVb56XkAwRsJOPkSwJog8g1A38Gor1ZkVFVUZiE6xRGuxnp
qAhap24qeCZEq7v6PxD5Alct5QyVzHzts994MZuFqhp2T/XPeMOLWEYLzHfHicvLHg6x0a75MoDj
RIbF9aV1HBgngHGcC6buO2prY3S1NqLBB46/TqWxs2SNR6oqaPBH2n8Cak5z+LxK6ITEDFpSV94c
YY/r4dND3NwG21ENJ7XY+BauWSlcUKaeBNsz3ax5Sbu4tXDEeNqhoG2vzsio0wQ7dqBsZr1Er7B1
34K4KO7o/ePnf7XCDmX/l+Poraqbzo/RrPryeSO8NpfaHLTSN6dYHewCsfRkN9idMMWgnxFIgkvE
iu5Mh657AxbVZRDr3ub/qPVxle1IIOj6dTc6r4LPFFgkztV4qQvYk8XClmAeC8wwVVArx29yvGGx
m7oNamM7MDJzUH8hw5K16UZNtIp9ahb17LlJKf2ksJ4O2RUh+3vdFRK7l3orlkBGNrIKu2K/TuTk
uhkaw87By5uPQ52Ti4DHGRK2oox09nX30GEQR6DAW5GDqfPS+V6snrk4Ley2sMGbQPjFtFZroUzz
D96LX0W7H6Hy1LXdtyUeULgqCEfxjTT1IEEBxsImXYPBwIo+72WUcOtBFvkLct8vxTmRjGqe9nRV
m/Emc1sJe3PhKqLz5dNCVijSRACl+ewLeAt6NQJLLZ1mtUuk26FLKC5ULGtxPryYBRdpKMffSq0T
jY+2SbGJyY4nUnI47vHgjIaf64iqWdCogCrdqVFHBiYlgMQOS6oGMegxDPaGKsbShSe5K57cWqrl
lxrLR2y0mQLHpqtGy7cDk/KpIxDlXUAttdkUZQ188ItdRuMfxRzCpGth6Cz5wgWjIyFqY5rgkgPB
JkuPH7Up+3jyY5GaMq5eXtWwjsEqsf1N8MDdGhdqhAKA5rDlUcf7t+rv6Gl29NG7lGEq30N1PuLM
AB011eaYHzOYNwwOEFLqjXnCJ0Y36x1EMFGvPWu3/qCX/Z4x1eU3Jg/nCAc7gbw8FAYzGAJgqRMc
o9rQ9u+aUD5GSpV+w4XoG2J3GtvGxywXO2w/9FFR9csimojCPImLVCacsAZavy4+1iKg5wMToP8L
tJO9WK4i6CYW/k08Odd1oV18GwwYxC7AndL+dnt/Hual7+kYb0VwOSuIj4jkpv514JGiNbSXeBd5
oclL00EMDNw5WUq7o7y+ZEdLtH66YStOhWQpkOZT1xCAbMFZJTevUQfwz2UUnAh6nLJK/swpNoEd
i7eMUIYmr8SZrHH9Y3Nz00UISjef4DBVZteVq0YBYt1IKNYsvcH/K7ZzbW0ooK+dgOpYvrXLVqez
ZSjyRzZsKK9wJPSZ9Hy6HORAYvEU33Kk3bepnN9NlWiOYlbaY6GYoYC4TuFY+ckhP0rG4Ceua47W
V5LPaAn7DA7G3m37ts+/kNGFJ6HagcZf5Lxg9vn/eh0Tc/m1gAuAHAuWyG1T+p8ukrqlqlDMTH4P
fZ21u52JE7Rc4wuv8kPbqLFgOyZSfAX/zuduEu8pxKQ9LQDr+xQdC2MJTjLhADcNm1eq15+iFZ4w
6W1d/zaeKcdnDtKxOBOqFhZSYYcGFPiXPf9/pYI9LprY785RMs/k1CCR8Vv/tqYTHygnq6CbKKm+
icL9pe6k/ThMHsD7uTUUtBget69Wb4fLVgr1WznaWHZfrsDnOkyME65FdXYc+GzvPDddBSyHiboi
CLcGO55pKSJHhp6HC9b39kM4q9O5Wql20xx2Hk2LN/Xs01MSelPZFGxDBEt197xDzBf0F+DuwUiz
g857xN/aQ0n72L8V1/nbuTj+YwKCoC26Kd5FcdMh5aiLxexMuflIAnvhhSUBCRGkY3Xg9d8cAXrM
/6qEMOS4NEsfrA5Vn7vA3sQpWnViKDm0E19b+IskSWFRgjT1d4I8ltzcfqxpfOKkW2WOlnDBEfk+
2qLnDUxVW+bmBJcjdi23UXSkrPHlXxWuOyeI0VXUg/uy8kPtGYa1mL761XHmRvXl87omqt5ZWghm
RF9BfSUnbtKiKnyGUETLbqSyA3EtKkOhznWK5ILY+3Dj+mToap3CY+StC6ZFAiul4/72AJpb4awy
bwgMi8wy9eOmwAfADxX0/VZwBfj/u7jx6uNIeFbfpu3LcisHUBF8s+txqWxBfsZTV4qAGxNb7KyA
D1cIvGe/Jwb3vbqoA+aCzgV+GtxuKIt7XmXzPAkvyyAHo4addo076CSOFdHHCj4gJDZ/MBdDE3T0
gpiqGfI69u9nIXUwDLHr2Yo9awZt0bxcM3zScJCSy4p8Nxhj82At6CLox9O63kYTKAqkN6TswWlS
RchXz2EaGUBYLzx62uv8QBVxOdzEty3g0oDVthnozuwphwx4Lwetmtp3YCYpebPxdgRwMtEORMsR
1vti+X+HOqZBOLZ7hywChoEJ5ju/LtTNi7tgiknZIGlWhNIFAq/WVip5tRyYMrtpfcD1xA9iGifJ
At0BYusN4VcC0t9M9TdBUl/nf4oy4T3lWxKdr3F4SkIeTudpOiKXvWAO/B1MQclfkBd62+kXxqWh
JpHMTK3DPYBr0gcCE8cDD/Dr0jVJ9Q6L8gIFFeHZmGj+9v+Gyx1CgYeyDb/AMEYHRDzvRlDubkFb
BkOMAolY6OvEFKX2rACXO96b3jZd6y3ZJuhVwVrCHxTF8+joYck45OrXkSlz3rYvv4Egkb8HNkUy
9rnhSLVh6BbXLjyA0xIWDNhRS1WPPGrjam8EnL7bbxvh8byJiTQJSGPJfoW/AZsEpXXiDRT/y7Zb
KLoYQN7AW3s+aemum9vGOrotSVj+VX8251AGA+jnPcQoqLh6pzdFPbPXTYAjBAnPKuimlgDbIVy2
z0oFqbYamiAMMMG/GUL+LQ1oBZVk1kclAkkVo/2s95EycloVi21C9tULVhuLnYhGAMAbjjZTBUEy
G+K6qInZajXKhVo0d290GipRO0TuGPPGoU2WE7LxD4h582A/Io4NifTAYAtfTIDT3e0HreER2A5M
evg6oRXAQrxgnWLGQsN2BOb/dlvrK/QI6VL2Y8P5YceGVv30QgQPUwse5p2q3YlAunCjYzaC55m2
qgRIbu8O7Uiv8vuNEbbdN51mSsNGm7kF+qzK4bKgp0qxxVTHm/hBpiHzsD2tJAw/H/l7caODZPfv
4ZQNsGtzEl35JWMalIMW8c1HYwHYuj6Q5TSTRSu+5Tc6+wYyZEMvD3pQotaxHdCIYrwzi5uyD5KU
O09sIG8iVMpUwl9PdzN+9ypdlPD+9FlWFlfbGgiEsqklcOg2d+OqNuarBfQNpE8L7tKM0HuzDsLZ
6noBl5D6T8hqK8gDtN2gFxPHopTsquz4t3VNKcbSZRD0yg7mi8446XPLndyELcu5PgTMSs6Gr809
0eRdz/+ZnlvDJNogBSTB9P9UlzTQwSSlDY2bICRbLtFWVDbAXGhXOZsuI3KOyfhVO7Uhel1Kzn6o
p+ADG8Xp+S/ocsQSNmB2kXo2AlFDxi1vraX1NN3HUcEHKy09Q2XuoUToimMWE2rFzRjEhHDGpDBe
7+dVmVnIfIiJHnPlHah4G/yda7FHAlacEwoXHdxo9UEAcpagb3m4cc2auNnpxtzjZVOBVY4Rcijw
xkq/ApVqEv5S/yvccgthEi1GFu/8tyAMJ1GCTDS83Wcg/nbIN/9H8Wk+51wR37RCixx8ZUMxb+8l
HGx6sAO0Q2K1aSpk3TV5AzTGwdPzykxj1ITImmocJ4fFkB/DfD3dpG3TrWEUMTtXnIsJZmn6F3W4
PpfKvbQSz+Sw1RqxmCN1KaMCCd5iC/hckKW8Yl4h/ehI4ctN3acBJLbUc8aeBNLsoz/miUWa4kUl
Uf5F5qKyxTFza1mTMXLH6tzIG2BXKbgBGapoOM9CWmnuRp5y575wFt48SeuftA8sZY5FSDgrcuYJ
H9pqNVCkkSE1E0NWpRlNK8f6jm0LsSetcApwNiZSfJuSagmpYo350it2ZhwW3GOlBENb1wTaUkMP
fRdRdanr+4SIWDv+HJobUUHOtHX2utKmEUtgizNE4i23RPLxwIjhYuOIVqZC3Brh3LJEbQPZMGKy
qjdHhJHAj4sdQGqLC/cJzWrtgUB1rmsyG1ipO8Vslp7A9ukLy4lnFlQ3fiPRWiuAddmcFIp1m2pC
blOJ34WUJX7dWRPOp0kCJnEwxo/VqoH/1mMd2cQqX5SlUM1nnvO3Q3DjfPN9d7bLxA1rtzESPbwh
eMdy5MtOyIcOkF9RT9kY0Y4AoAoAyjZKELYuHw77ioEmumjRPV0S1oAAmZxPwDrDBMGK9SHRQOt/
1T8k1IKYEHAjbh44pwtE1YpncfXuS6ZIbA7TeG36uZbUiDP4AHav9nEqm5fd0fzWXvFx1H8OhG9Y
9pEiL/6RshaoI0WKRod4ltUyZnSV/w3av5PW33lKXrguYmk82CFo1hysb98zYtVlCAEstC64ObGF
Z+rB1pbIO4qylQIQCFxZyR2SytvhCM6i7r/HaAHXYgeRZH/yWtYugQSKWavddRvlnO34wy1R0B+c
HOTnuuEalvEK3SfgyesO5H/aE1pG8QSQ8qEuEMf9be20XqXYH2G+hsDrYL/riFk4TQjipPrLW4RC
BmkUySqgYlgAX0BKzIRaFXbCvJwWMSapRl3g/ylz3LMeqyWR6y9T4EWJ07slbdNSkch/p3SoBA0s
JZxTqVhuoeBhBOdo0LCpDYo0kjEateObDek8FVKYf6XvcbENQSW7TNO7er4jzWvmTUJJwAwVgJ3z
edYDvv2WfJW3o0FhRClzCDwwqQCVq+mpbYz+5l/um4PVPFoXTW8L1vzbVtx4kko05inO+5Q1l04a
8h/ApMSj0vgVTwejrIB+PZbFPzU8RQSZW9TgDWYPuGlq+ueolN7LHRNgDzKL6R4nNRvCgs9TFdik
gNFygMBY40tv0ZqCgXH9zmTqJvbHxjcZ1uxxGt2Rt03+HSbGijCLs3xPWWQAsqvWSV41RGeLb2av
zktJs3XhwlUVfI/JzI6uWjSQ5AioilVb6SLcNQo0cwGkjwwWl31Vnj1Q+CsC5WmeM2v15Dqu2RCB
m5kro70tf/2oYaO5NESlJm/PXxR4JDVNTEKi4x1FTiG0w4/wa6okvvTw1o6jnArhz9uqgVr2itTi
+KBAwkGR0f//42XUchtoPYSbOQgq7U9e3sAu0Y7Fb6ABHdyZ+OUa+P6HGg43pRTDUN3maCUQFWny
EGZ4BWuual3RizbCTJLk0eAjGJ6GCkZs1s9Udqs2orsyRedhiPqqtXR/vbFzGh083Ou61UL6Y2cr
8lWC1Xps9ybC2A2fXVKhTJ/DDdvTciy2auwdbgG/Epo+bn0xKu4d/Q5OyBywFz73BD3TLIi7a528
sD5XmD32Ix8/Db4G4g1HHG9Wnd/ZewOjPsZSAJ7fS/1+p+y9mCseqikC5HN9WipTGuxN4IsQSOTm
WP8mTSg72Uk2Wu13b+W50WofH6QohIB2JZognlpS4pm+tqeV9EG2y1Ef3qn2Bsl8wLzfoUTzBYV3
JRnBVxqZK75k1cp2yea/FwZuTb7pBCCIgf9FH1TcphDo5Eo0YLexTMXw2XgHszZJkThHq6m3pgeM
YWn+zFzzcNXSgZdDTp5Zfvl2z45aMB6qiN4ne0eKVFMAlMQYAXfXB4JwayCQkRCaufl0uBydBrZ7
GggfhP09urCoZ2xVNKHJBFsGahZmXpY9l+xMXUTgFl2tjZtrjqDxdgHYISCLt5CJGyqjBg7WpY5H
NUCvLJz/lAyDoysjUfVa2MAEBrdTFkUc5wOPjkZclVSlecLvK1d8dRlXHVVfETbT+2Jgj0w7BbyI
16tWcUcmOST2w8yuoBe5Eejyt/PH9WcBcntZ9md9YdHRUG2P6HE+5ZkmJ4N3D9nJACObBIR9tsrk
J0SCvXjFOQRJnEpdc/n1Av+lLXoclzUCXSZVviTelJHAjmRqIb5p4PjmKRnkj7ddlP1KERVC1CsA
OsDvaqPqYznMDfnVMpyqTk/NaEYPx1gQzVI7zZjAJq/u2Sj+64Bw42jjU9ZFn5XgX40PgWZyq8Ft
cxTRH29K+vEX281igGWp9PArbKU5NTSCu2U+712NSXd0Wf2gIzRxO0yNJggAnIaYaPBnV/86wPv7
lZ+fHRtjvoApUnO422Klati/pBMqlccWb+qAg+owvyCqBpoK4txQq1eBfUj3dS16hqvJBNeESvYe
hj1H7HirCwxLKawwFQJ7seejYm7i3cTT2eJ7jGV8bvl1gn0iPKoUJuOSmOIicS0ArYkFig8+qIJA
nbcCVdxy/pMQpRDSmco3RP9UNMwMKrpL42WOyN+T8UBYm+UkxEs59Oy+MCasSb3G7YtpOBrGuXW8
Q63S+ZmLM81K61+reKnBSAnw1XekQmLGyfhpfPiJCy24NpINbCvfldhBBrFmQe5b9w2gMlrgN1OO
7ERE8wMFGslkB5IKTG/XifHrmcxoYJBRCG70Hv9IDPGXukedIGNbBbMMfX4hW7pdxZcVq2ruh84d
GZM3j+SFAIT/Hs/j9VFLqcKT+0UEMoJItNM0pKU8emDRvh1LZEo0PBe4liaV/i/xPUJHByy8mSeU
6Y9ucLCvNRSywYi9jn6uIn+3khr2yD2Fx6i6wXFQuRtlJOXYyzkPHxEahw7z/8j1XpxYvS9kkhdU
VVmcBBgp0SZovrIURBuUZKcU3lF+DEq9z7KyUKlAVxYtzyaC0jLNY9MObG1Yp6tnSb2x1zCkxXFP
YIdj9AgwxUk/BlUzxdqAIsd/z1gDxT0cRSbrYt887VkY20S/wanI4ldRFR00CbCENBtUzL+VUE6v
u1jzldL+PjiF5XeNzMxYpIx3V2rQTLvWahCA3MZVqJu1amTqjohugNJz+S+5ZXQvfDyYjVAHnEfU
hD0awfqJptCV6M2pZZi8BEShR1jJrcsgdp8lBeKeUSinaiHVQzSSW68jinFbBWJYra/igcXSLIo1
j1YQdckOqyqFzCF3ubR4jrTMkq5hBiwnFx6g/rjFkHKMU79CE9/5eX5heX4kqck9JDsPY6pAJmMZ
ttD6Yfufr7CCCWyuXaO4zXZ60Hws9wUs4/aMKKTRae45YG71KLkt6g08VOdlwq5NifssjIIXIyyG
gKeXd6fUTHkdLbPTC1qDpUBeVjvRDEtdev7soz2UaiSbGz2oEX4oxL2yNDStkyxmx1ygFNMcHbHh
yhhA3HLB/rM+QE33fcObHtwxFnTuvpSgJ1QafoieHee6qBb9jl/BiGkHhbZ9J6KGb/xITgK457b5
D74z32U774zceJ16RlrHpGO08+zM/L4WBw2Q3ezzi65vPZf5sBSi0nr2YmceuwnFFZPcnjtWmEFZ
3KWyv2bfH9P5oPMeLApV76XSNGLkPyoHLwlV2YYHaeygygi9+fb5iaHmymbujw38mp+TT6tcYmSl
cFUKQ05R5Yz3pwoWiRitVINpxlPEoRxe72Un3Ugvmuyu/db6mSvYwI6lA+wleuCeSaz57zo8n5kP
bhhS5rBXVtvH91ik6UAtC0x9Als36EJU9Wyjoyc0ageOLHehu7GOnhGx/f7HvhWdUGhtjIPij/1/
cJ+Z3kjQBPNcb8WInKiP7ll+zN4ZFHDbgDRw8I2kj6szY0/oMUkQAIIFQymCl+hiEmIhUkauMCVM
Cz6TkrAP4Rtt3F67pwoKxsaY7gDACUgQyWhTb4Org2NSC3z/+JCeqBh8gSDlsMZGMSJHNswC+/ba
A58JkZDQ8P5OGZwVJhXm+80o5t9gU0Ss63EWcIS5nqSX8xCX9H6zmQkqdesmjG6shf70aeFvvFYf
rYRdQb+Oqi1q6KnLvBGF2GoT3EloFP4PhujOAC3XFEWWBGQyjyOF3nyzUoKUvtvWTF6gPHJBMMW9
8/rsUgAjhWn7FyIakZFbT1J6No2uVK3bhcM0nUgbmfdZ+haCL6BMHfeQ+XCO7S8eqa8ENoWagI5X
JxZ0gDDd52wdlxjfAOhto1Hbu3lJCL2hzIeh+GgjSv92CSu+Irn0wUnh+JmO7kKI4VP+CavYwJcn
CGx7ENJqp3aTBS7TMR2rQ4r4VJfJoaxq9FTCq39nCpWCHaS9HjCcL5OIDNMTjUO1r5fTZsYTRydc
+f8y2jhJJpc3Eem/zlkBYh1Ctn3UEERguY5CtUa7ngZHDYSV+2Uy0qdOGi4OD9hC1yGDhZ2rGU9E
Tx1uTlodF3D4rSC3YCqX9Ik5R7eOZqqqE39WXT6vwaLcanYoxxI3dUhttKRm8JkVAAVyYvqr2MpV
eMeGkNSE/6BscLW5MIEYb+j/JuY7YzCj7LTQFXzwurzVIsyPNgUb2247pjkU1Gt9dgqwGEoHRV2R
WmlKQbYf0kaWWki3bBmPn4QIaaoDYaHZ9C5u8aAggdbw2QzbLv0ikftx4PPywAcLnLWVojjK5BHl
vuVv3sB02nWWWI9vaDxGFLsA5LrWF6r5KPQwYVl4xmJNoqzF6uAWRuLdJmq3sb+GHBeukRo/cc+p
gsHBNvcNqORrmpadO5L/78muMmUpp9USiMTreR+JqMI6bevoUg107Yjcf84mYxyLXFdRMlPptBDG
T2RBjDw4UBZbVlF5b224fsN/ceYBF1HGZRK+GuXABOe+0csHmh0+zW+xsoOoBuwRm3zT8fneaV0x
LvdGm/e+ElYPnMchMttoRqXOujkv12nMDVVO1rVNUZTl2ZGZCimfQmqNquRQQAxGqFXYaPh3oOu2
utofw+qv2ThdWQpmpKotjB4wUiAatxjTd7Mv7J/d5dQHWddWFVIGfed1/PTV0FfqS1t/sB+VZhxp
Q7QAYq2b9My6B9yEVSq1pdFuzLuIkzoixn7XZs1aG/G/DbhjoeuvuCFEARqtarGcSsT7s8jeaXLn
kiYiHvEjO41+V5LPmmBGucvl2wggF91yjqnGPx40KA5UpKf4q8jdJlWYa7UKcWF54tLP9a8W7rrT
LoEvPnh251zqyfpoCSsuFnkKDGOrLVqd08fWIEluGIAlBgTeQhpAlM/LNBAKVXbbAzRfKVQtxs+i
aNRs71P7gXoGA9b39F67HJwj3bT5+j7aBaG4Jd3o+pXWyT2j4b0G+SaRN8Vk8tK9YAwXoImMgvoq
k0SxLXqOdZH4jka4Yqrkm3UmoRnT9S5TSgN2du9HuljX50mrBIngifTzSExoGMJoi9xxnWAVpalt
LidCohYrpWGFr0c8enjX4Ent48yKoV6GBDLWmzMGT6wusXtin41Z6Q8JIHNeib3bQszbKwnHeaSX
zA57wy7g9XrBjLp64qnfHEFr37uORP65gTig4vkwHmB1dLKhkwLIkCgI7AYRuKICyP/0olsZBTc+
0fPfAQGSKgwsW2fJ1eI/6Bogndw9rGzxOtv4tJJEHjHiGAzcQ8OsbMNJ4VgpYZiLXL8A+wwWEDG/
HeUPf0OhIf2ynMKSnfvgVZzXe/cKNotesVu0FXkbvFk7q1D+Xtitk2As/E3yHB9u2vZZ7L6PgzwU
xDTRhFZhdaPmpYwbBHgNxLa3lK+ltqiXQ16P4ez2DAKoMObAL0xI01EoUVPyAA0/v9gu+fcxUVAv
5ZS4E6awIJzUbZdItQlG1IARDE+4SpAg1R9aIwOf5Ico5fs3wBL0ao9y0eKwyLC9rKETrLwPYYv0
btokrnT8z0D8nbv0HsyKSupHcllhqIaxjfEG8KvtW+oec/J4sDgQC8byPY45wscJNoj/HYNXYWez
Od93Anp6MLqIDN/HR4d/EHzRNod2/mrbP50gnmuVAPJ0fHPjUs3+XSIlz9xGM8OpLH0KLQ92Utbx
ULvFfnUGuZ1UznL4sX2M9CvuUO9WE9NjScexxBdfVyW4DoCKGA1LbtidSYEs79gF7mm1ywXtWmVs
SDOvfY4PMt6qsWJZ4pmbS2iZNN86Rsy4YhVLYtXk8+3+KZE4fhK+/nHfucFMq3HWxgjIthXzFksF
/RRZHbC+2ksAT7bqwWKjOnRDXVEuWWJHAybGV81XDgZuB9sUXVuiVLoTZGIUsV0g8O6pJ7eVnlZE
Zeda2Oz4Jnelr51qbDBpiBnbibpah5cv6MmVOWRIogOXTZCzm6HKjpP92eyDlnFaVAn1O7ILw9DM
crJ7P7dOv+SeZtqLYgyaeVqu+9qCEfgAOaxtXEStlZpODZM0r7vPTazhS5XPlecmOpRa4EjZgrta
7BRhlNeDJgl/ToRMFXtDXkPA4thpJFQbuDAepwSC5XW7+IyI1EZqaIKvFhhbBAABshsBk9THHKXl
EddMFvwcdfED+khtMDxKDRi/xxKrly4G4XDJwW3Gt83ZDZLGv3fO73CG9FOLIhwt73vS34wk4MLi
g5ETS0iilXuQ2AO8ktEEcRXIRnhcml8kQxF63VH0VbPgJFV5H0OmDUvNXeld621qio9KMebGvxkN
mLbTtM5xUfabBVcVtN8TEAJlWpqt02GrmEi8O20l6M1TdPJMO3R9uO8nBKq+rpFbSzdfy/Xg99Df
jVH/zhcs71+GLrjYKs+pG0eIPdGjp7x0hDkuum+ge2Sl0750popVSS8x1a1fpLoXxUo6ZX0Ulo8S
bq8pyCwnI6t2taZCtDmhgGcAI2gog91XvWhGxQNCdMy37BbC19kZJ4i6ssqqFOdDj9h3ME4tdCbM
CFvSKHT1tJl1ytyuOEuF05r1TQIOWkblVstyshe01bDw52DAA5PhnsHc72juJsUFJK2pxe98k2cA
6x8MPwJmKt5924MFyjtUDwFbU3DBIFuB/8M6/T5z53JmY+n4CZS4QLHbL3XL2ycvR5eAVswrmkHd
DV359z0dTdnB6FWUGqlX1cWdsPKrjF+aKgayvB2/zgtkR2kVEEqUEii9iqFRG+zCHzq4sNgv22gW
obBTxAfF1vxcaqJMJqTULOi4RegEms/dntcfmkMEn4/DTENm1iZPqjPBED+zELirVhiQ/1aqC7sJ
9uV+XKVPihD3qHVw21DJKX8H89tTCpdokFDF3cWfD1voVARMsOeHzn5RsJMWqiCp58Clznqfwkac
84itn9xy4tZXysp8AVhnXDy/mHBC93zE2w9gxwyJx3lmT4HvmKSqAKPz2Uno18x/tLi+hwByneuG
/iVcFa8IKdBtxkYCWPukOHCsWny+dWa3q+6tUlBA1dGKpQiawTtoVJiBHejyO/F+bw2eMemeeQc+
jMsjH1sJLn5LMbaHy9CagpQrrd7BJyobx5LcEAKCYeFOkUbeJUl/nmzf47QhnwAwTAR7xd0/9GiC
SKQNV/TUAxjTKY47rC8shZ/bIatubrDxVHctjS8ssWuHxEVNMSrZ/mLhkeFPSyfTjBfqHfj+6oZ0
Zb1J4QBEd54/djBHsQVPUnTdaelkBkROpxj2vC2hZfKbjS2TBRZK+m86GGB3Bjr4iOyDWVg42Qyi
3zjHOLmNePijuUpR2HSf1e7Btg3F4fIWl/htVw/mcf2CmqidsUsLsH88do8Dr1SOYkZMMw8qfYuG
J0dN3sbVzLYZDe+wfBqej2XhEsPx0BsnFygTBg7C8UY6NrauFPh1M2PzMY/uS7I9vA9el80WNxt+
P7j8ZdX5Ja5XstSO0++PDc973ap8T318odxjIH4nYBQPNeHF3YwAlG8X6UDMz5+aFVvS4KF2cF69
fFUPdxUJOzseVEqk7LkA+VyjUf2O73ergCF6h+P9rOr4nwbO7SRfgVBrpk+LCDrJ589ivVetBn/b
wJWC2CPTRiEjNppRo+gkI2HxcpvTmZZUNNONYck7gH50o6hT68HTZ0ku0+QX0votiFm9b46RWbPV
4JbPebD+vXNnfQJP9im9VmEvUL9s/2u6U34TQH51PZCfgStCT5cqvlgyDhCxHGwVLNTrNbRU/jYQ
4SF5j4rWvwnxqEU8oVVC8tqs0rKdGJ3tjeQ3nuu5PzCKEheLpN4cyPoprQomodzdbX+pgJbnl4Fp
5Te67q9ccTvC0HBxYmqYpMOTh/Rr1VAAlmQiFJoGuTt0W8GU4q5/pPYk7x0r+cbtqfWLfofWCnS4
/X+/6i27caolhRbFHivvvpkVQu8Ac3ETjTV8dfZba6iILvQ+QEafCArbAx1+lHz8iosaozSN51aM
eJwzhl4iUGoL2aaTHgwKfBf8i3vvGRf82XLBHugCTF7REHcOXHLsAKb0oe5iE07V2KuScjUql5pY
rk/EqH8zqIBppr1hKPeKX3f8AatBhGhyMpWJSBVmlkdaIaTIreaBUObAeN+fLq/hpcPHHzJ/1NRb
U5Hoy9QuwSRVXCM2DKNGJU1zHm1rxx7HftL981OYbCowQGH6E2F1QN7Oh2yX4YxLe9yG1hRR9I37
7hv/0QvIRGqfXK0JsvoNCivxwwfwo4W+QemK694t4/f/p1hSa5VezjtFWQ68w30TPnqpFi2LnuaC
89KomF4RxFeMVFfiapq80nHx0qadtqr8DMhKezOniqT875rcltSl95PNyUmIh7GCUvej/lmyj/rB
W4zx20x9/I/agWacR3Fnmbvib/NGZDf1JTz0lJYgnU5MMSmKdXpW7IEx8xMLe56vdzpzdwJwI6QJ
DSiaMKFigcnhbvVJfBzPPvEMCyG81/m37KP3WU7k1bSfqc5ggfX6q2NbN+gEgqzOpSyRfmZdgMUm
OldM7j9q3bI4GJQJDloR0ttcpSU1060Ont/XqK9Rz89qoy3jLnJ7x7j+J4p/KKzzsbj3vPgWbp5T
bvTB2Yd+No10tOdlB3ZIXq7Tv2L6Ky1TEVFheRPTpw3PlEIEv17a6TUnYSC1Ul96WS3ANtPa8usx
ElWoQNkdCLXuOm7lf5FoX2Mc2tP8FSlGf1PH08WLI87QfDqY02ktfIxLaaUmgZlpz3ZAP7JnY5qX
8JVPYRLiCxUdvOMKkMHlJLuLmfb2i8oAad76JfXBR6hSdUoyks3Jxyiuoxy4hSsvVjrVwJHmXrBG
c7NLTfqbedeF/KHEAr8MKwRczOHwnpg4OaEzEE7OuIe+FQeBQH+y40xCONze29GgsBFXOkK3zD32
iOSlVv9PubnZbUNKFkqb3lsQMJ6qbbtWvMWLXbTYBfyYlxAZ4LsolwnmoV9voL/IsSKYHy3WCEKR
A3j1fmeO2CQ94DcBOftvfXHDzmkiA34RhP62YZvI83X8II/CL/ekbOuBWnwLJ1iyqlIgu3D/b7xI
s0EjjZgE1PqejXQBUk81RaJnX9M3uBL3m7zGLgyMs7JzaoUQ5JOv97poNKvt2D1gvlltJ+mAA9I4
VhnOv7Vl8cclqSpEtMaZX25a4MphWX3fIVNvOH28R69S1D/KC6opbgaR1wAkFcRSwP/mqE9qvKR1
vGdkCU75wwp/oP48csyDrkg2KmMreOpn9r1SDN3X6ejSnUHtsz5PZQD3e7q/bS8IIFwAw47CWjY3
xp5UVE8JylCCIo8a7EkfI1lhBIx761bp/uEyGXVRrTHXsd7HFPAe5Cf4r5TRCnpv1zlFkYGOb+3j
xUMGkCahlkN6khef14x3D/IxxWqcWH4JqwL7QqLCJ4HuTBc09u96nchYrYmKF8gHG6u5UsXjD0s8
QQiFwukSKjHXcGCXEw1ETDi/w+h+SgjNWnX04sowt5L3fmgkd4iMn9mKax1fjnChIWPBmKMFlakj
ZjuIJtzFKtbuk0hxU4Z51ZjRzlPzn4vcPGTge2U84puwqbhLexhjCVU+ioLpUKshqxCPXXX7+o5B
TtatsCSZCWLm6PIn1ZKwB84TPlVf1UY/MD0QIVfHp2aF+70XCtQ/HekFFcnqUQQ+w/dw0adE/d5m
03TzFRuAJIIo9fpEAETraL0vPIfqf4ODmjrn/FoBwg8dJKwMt5lt6TdyebmjRi1O++PtieNpqCGC
cxcpPEGhhPC7Pa5G4MxpvLjq56LpF3kWjbS6hFrKBH3EwYrmXuH5v8USkdubboAir5MK1XiRVbe7
7ytEAzHX3CCrP2v4z6wat/+N7zdAB41h/cxNoqL2s+AdTUjrRs2tp3qahkhvXf16lbUqk+VdOiHV
VPlPKtUuVrrlo99ogwv10hG7YSEvC3eO5IJT+U4m5uh7EUwo4ZKsXIUQcpnfZW4ioduKK6QBd2XO
w+zyoiu98/39CR7xppb6JMdoOi2myGun5cYNN8+m0HqDHPvjm9rrE+rpN+k+Az9m8TfKJA/34s2i
LL5b1xDyp6PyFzoJ4LkI7LhhjaLR1andzESnPWV0aWyrHgDgEA56q0GS+ka3JCVXFek+0hFrL2qt
0hjQETrbK7lkGZ5oEn5Idhpju3tg3KPam/w/WKzAnleOTuXJ0NmZ+iWvcPFCjPeQmPw+4VJfAYWm
4/zoFKOVamPbLRFhDgQcUDWg1+1P7VUUINRBiugS7lNgDWdHsxBaDc3kgxOECWtZx0oWNzxQ5+VI
K881N6DZml9Ne8u222aKUF6bA8NFARnLN4nDHx9r1//59j+4uyePrq04Rk0M51FiA+XE8L/DOTtG
OtbVCgOY5pKxdD3PID6F9bO3RBJbNWI+wsDW7yuv+50KB1k/X8O6R9JrIK49HdPrZSCQ1YKBo22z
jhsIHlsCx/XLmDq1M+2PdjRdzlCvc3Nxcg4h47jiF1qhgFk/Rzon/Vx1PlQjF8WjlSuqoqCkX1K1
yLQYWhZgwC0w/ROr54jbC3q99GcyCP7viAZaCV9xXG218mbZEMtLOdARwHKmUuyK+CenpJrXR8R+
UDGn7jTzCM9ErH6rHo5JG/ykRA7V5ZbJSQsP5PBS+5v6RPpt0YNdggrX2CtTn16D9wPQC4vqAD4E
pvIDYCpHnTKgjUgpqxkcA5xxHkZt1siMQKFNi1KduzD7bly0N32d2mVCm/LBMSQNAQYLzFrNoks3
MiZTCC36L6b/u5H9dhv1Cv/vj4f5ozAkz4S5l5smNi0hSNqEpmRLTt6iIJeUnK01PzUm1cug/cYH
cTAr9wHTv1m7gb2hU/hjPOVWFVortOK0si/bTnoavgK0h1UH3sOFjNXMwerJPRrw4alI0TrEW+Nf
qJeiUNY8ZSbsF7Ya5LhtZMXJme/xI3OHUo8L6+Xtajlo0Pj9ZgCjH5tqYvJbPRvtSyb+l0oDKqPG
pXA+F8UkieF4qm+mLUW2dnsiklHo+QICl/I3FYMsD7MmrD2BiCHTmLYlU8VbGBzaR2ACVZ524As+
nw7ECX/a7wH8TdKnnpQYqp3VUcuco5f1J5fS4+oYsONA8UAIiqrYFi1HE+tupaAEUywqlU829OhU
ikzGtg+fmqgfjCQ2VdVY++bLFVjzwbSqX94hb1HbqDMBp6Pl9n2r/32zxeiuTCNKxRFWGNup//Vf
if0vv2zga0wIJvvXxjkEz3m9ZmbuRTFa17eG0f/oVtT+hXF433Zivv+3A5KnTjF8UdiK99Yb+z4A
UL9/rJU9wcNLwVpTbnr6KpEeqf+DsIWcrPEy/8OjxZlK6xPBAkeTYwgLBYMaE0/yv7yO+o55Q4cW
lw8D7f3zUP2CIxlp3NS17c90BYsBzQ6tODlP9WpLCK4m6TwXeKHRJi7Fd9i2+Hlmaevn99l/jb8m
d8HljAMoLBKuOXEBBSpkBgkOACuqnqxtHssM8gR6NxQYJsac8T+jwEoViSwhkEAx/la9DcjISkUR
67lyrBdi+aLn/Va37AM5AUqE7wIkJjLNJ/uW3n5afHqgwCHkqwGzvr4K3CyAXChyWiQ2S1nvsIIo
KRRKEk1YRXrDWHgw6VyfIB8J2tfFf/6qC8iaP1qyoFjomlC/GinO1tOU2ugxmeb0jlnF6Fp1Qd//
NGRgj/d89YDv6C85/ZQIlM4pTeRKaM2dBJE8fa2p/1Zsg81mcFFWIlNrJ8Q/PPm8YfY7jHc6gN7K
i/vBJ4NhVLJaDc19TJFuZhGqfo40+rk4Qsie0pPlyLVnPhnZqhkO0N1qDLic7dLbz82OrzdMBF8g
Txdbks+lNIV009o5TKPiUyTLuC1pKSYZfTVubrOCx+4/0tgXnTAVIodOh/QIRcs44DAultA00GTG
gvsb6G6naBdKmCg2qGBCApvMwIRHLgOFAW1vI/u1If9XTzPW0QNB/QMkH+io036lQ7ewNC2wrCOi
WC0GOXNmVUIUl3TgJGgnsh4ISJ6eHz44q778H1lAV1wWq9jR8Lwht/HRhMBWsIv92OHR3wMQvl9o
S+bovoZ/IJdjDVzaZj73vS4Qh6NLWiXiykyP1F6NmZBqRE1urrVYC3jhwMKC5zmir1fktMBBEGwn
5dkvvxFQ6ErwN/YB9TMbR/xFI56GWQukprOk4N81DFnwoGq341DaTbcRMtVDXZC00OnLCEXG8/ac
gEPwHyGv5MjoZkU4YtHMMDrPOFEfESRu4neDXOXOccNsLH0D+FK6l3+Goqg9HWn+HCvMBG4kYgr9
EpYGFRBc+Tp1Ue0yRECYVg2uKCdsCS8XrQBa8I8ReJQA+YWzpWEgcmsGwsPPGg6yhD8lIu+5kUZb
VOPx3jOUVkbfRMvTUGtvMAqRL/v1+CMakDbFBsd07yHaFfaU2Dmq6s7Sw0Mjt7AdRXNBhdPMjvzI
vY2aOB3n3Aen0fplt1O9jSBnpqtJQjcNM9Gz9lMD/o58V9IZv1ZV5vBCoBCuQJK/s1mUfdMpEW6+
Mew9EoTakqDcOc8Dh93KmNVlQxiGiwvfk7B+t0Q/Sc00fqJt5FuSpas16qbySg2IXwLklBpfNoLb
gCCyCR220hnUFxxTv/IyXfzifi19ttvqGS2o/Bht+au4MNRaGMhFDPgD0p8QB7tZEEeZhb/UF8t+
naRsJ1z3RjDmB8JZmsQxaaI8IFFUkc/ZL8Nfb/5Alfs+8w0ZuxKS/4I1n6aiwBS6mig2L0BX0P+N
Cdxez9OWYD5OvIv2lqN88ruShxhMMoUQilomAxty28kVUknTioRHzhaPUq0udyFtLhkdDQMpnwEd
KxqoaTThYEQJjF4TmrfXIagIzcbf7MeG1cRhqeqm5SNhJPC2MeR3LCq6TPiO/jj9eoDGRq3s/c5S
WyRLIvkRbZ9GT42ypxGcQgY+nZLADxtupYDaYxpm/p6LgPM6ubzVPA3Y8t5wLTyMPrbTxcgy7JiP
0b27dacRVgii5r/ASM2eri6IPDFu99Cg5s8K22pcmdLaHQjcjkpv40tJmJl6By04RYihZg7Ueyur
qinFMQS4t79aO/uWAO2EkIh9+5E7CG0zo76g1nWsTy9rytcvKHFNR8mpXeqqxUzmd4v5m4dolVl6
DUvq41EqA8i68qDl11mtk0eeCUcG0up549u6A6hX9uHjRuER1H/U6H8MpE/gcDF629yf2Cc4TrUP
WCOmhI4ivLchVLbP9fFTl/e5ZUMXcd3yeQmMX5ww5kG/KybJ7r6Rnc8A37rPprK2xHIPlS+Vhmqk
RwwPpuUhx5kH0/eF5N79dy9cviJ5N1DOpVOc6t9v6rhYme388gVke7ixWX4lfv6jcWGM92m4QOL+
864Seru3T4Ub7W6CbDQDpnWE3JKkZBH5tZj9RDcYjpnzOAcgE/hAw+f7YI5HY3lo8x/u2kLk6/kc
BUZn64EczGx3SZX/IiuOPvyfwjVxmXLK4mtQRS9bIx17eSPLR88dbp5E5iXoVcXv92RA/DjkbMnW
EscX4E146en+zCKWLhohRP+Hc2SnHmdbzbx2Oeh7ihKRGsP244/Ero2cWBjQ7sedUVtoe5eUvRwn
FInfMhEbzNpWD35uJ0WHk769NBveHjS4RUAXWMHiMA5Kr14Tc4azlZqy1w8NaSHHkRb8Hi1/Cq/J
Wznhblt0dR/h1izhSszeEj95FvAWcM/2iQtISKWVUY/+1ENrKa9Fb9+V6oWCHJNl2vdgrs/F/PZz
t7VFhkDUkBHAjZN79+Ql7HdrrgPLA1yRFZhmCeGjbPoFmNG7FKDzdUWMjiFFdp1Y/aF/2NHkjxTU
VtYeWfThIZiEjQvhSiUfUSMUvmkYlI4F7LTxfRLtu1WO3CFrrVlhYaplCLl25TJCuHMeBAMujzIq
1fUFurOle0XmSyWN7JcuzM3IkgAx+/EAjQ0a0fc4dWtm6c4gYpVZWqpfMUfT+mG6ZRbLrRpMTFYq
akdQZYemcgrvU57Du42HQzYSGxqqi0MygWyxbF3bptV7HzfFeJuY8kT+/ZNlFEmynFpP5+aZcfB0
eQwMiRKQFW+L+4fCuO3YeLWhfuVGGoeg+VcTTu88YqG+XXRuNQbyyqRMUtWrKq+tsTz0BNt2x9aJ
RgFzGXadZHLxrYa8beHiLId253gnEpD+wjJGR4dNJyACVlz8wWYZRErnSWZ0S05RiSuDJcw9K7+b
6rDCo69Oapa3L6d/OxD5yMiDAAKYpeNPemUrajew980bi2m2yeaFlf4114VzGnjUVn7PiQf6kqsY
oa+doz7kz55taS9cwPZi7egoudkm9A4Zp7gQ64PxYTTyTdJLMaIVmNgkc80MsFxq2wUtRFuY6bE8
FzhvK4DntASqdpLfkWdNSgw+8lcrHKurLDgt+lab7tcLgTx9RP+4ypNzvna+QqXYUhc4GnjcD1a9
9SllkPH6cOmA/ynzdL7WZSPnNxzIQvZGvXY3yz23jumKcQMoBx1m3R8X1zkyEdRIXoQKOYi8EkDy
ZIM1y1dEDXMjhj8Wq9c8fr8ep/T9iIvGlLrBH/Uif/AeH6BjNr+Dwg8C5sqT27DM62t+Tanr5FiL
E7D7qnVAIpwzlzJZfouRS+a9mgbSP3/zyWuJ7eCuZXLwGACkZTMBoQm7k4CA96LA+JgvNLcENWzF
4s9rJlxdsPfkkCZcKjwKGQRaX5kfVbYgeEQIKEZlbIn/AIERkKYOJSSsgSVGD7xVJe3C0QZFsKzc
VQVMIJQ8P89Lxci2v8rZTTn5xjlyRnp+zK8+UDAa91eMx3pwSARQA6LSTGACYEHLqF+lBn7k69DZ
uWa7+JB6mfWtq83P4YzdBLD9MAEQVGX30BmnV9pZwGDUti+OAxYqGncO/7l3A2Wo3qk5tuEAZml+
cRGC4ukDfx7fOiOWNZvdzxSCKkL/Q7kLegynDjtX8z6QgvtaFPRBnzYRjkG4B8ji/7W1lFHHGoMO
WZpibgdcG1I8E+k62jEkUZ7w0tiuNSG/Y+pNf32HWb3a6bZWkrEMkeTSlwB8Gp8KzsjK1Kua7eOr
jWwf4b+YAZjbT/91LCRTaySck2fbdCbpoTXZgC227MSOjLWPd2IIn/hXTlaxgS7Tx4JJ99ARKyAQ
2fmfz3ZAlt+Fen0dG4t/KvPgyKN9DRt+r6pOXvLXtGVtDNDbcfCNMLV60FlYdOQpzaiOmTaD5GC1
Cm3sinaE5S4LceTRKiY4N7ujOY/fXAdDkSL4R9XHbcDc7wDETkTiACAB1Wmaq87tHwErUlnbANo4
01h6vGb0xKTwp6GEmlvGOP/nG3j1/CeZaleO7j4RUV7XAErwLaZwY4qMWvvcyyo+tRjNDHEABEkE
Lyr+L/6I4+/UNfwVjAeIGXytkpl+6ErlNrAzhuSxFAm6ZxN7eTDiTt+jWEkmGcg04PCxYeCZMLkO
/ra2VA5N8TkDuSTaQqk7gHA2w8TbPO4M57t/bOsHjKHlKsxWIzuLT2gOaOotQ+/yTSa1ugK7P3e0
Grhbn1FuJ6rmgdN8Bd1+w1355q2xzKeXHuylxjDTFBR4uSlTmauQNVLAKXTcmYd7/k83jL/+m5d2
W0aALSbPVlxXabAii0nsM3Dp868Akn3T2J4ZxIzZN+GNCVB1xOE4MHtEELthwYMkrEToBG7gR9PI
JeitnuRsYSHR9cbeonr9ROizAAAv/yX9b21B6kfbap801JnFn46zh9sdn/Rts7o+0gZuHhWQosNq
6Ze1M4k/goBDR0YKjrfv/cMRbDxUOPLiGsOrfRPzhpznjcsaTRomxp6Af70DPLKmjgA047daqJ23
inkiH4vg8Ast1UM5LlAGInKZfonDAWSJl37RNrCPBMzWQFdi03eZlbFwFBX5mym84mz+O6OdKM49
f1Zld6DUiK1ZCmg9QYjZnWUe3M+8RsolVaFY5fXHFZO8WOPETCnvxTdF1XHL918BfdyMeTu3jkwn
oKNY/ig7+7LDUjBtmYvBiKDVN9sDv6NNtujZTGOAxV99GC52YxZwtEw3DGvJl1+nBrXfBxQZbsrM
vgzcAWAyOGWEkwTeaX/mstFiaYXEN9reDfvgWI8DhXv/C6VWSsD3fKuksvncHXVySopHDaFXVXpF
TTmdlUWTjx7OjRgtE1ErckYf2g4OHC2/Du20IuYrEjJgSe+tG7qo9jdf+yWrsp+6TQrr7IhwiRWR
OXho8GbVnGe6pceCSuwieC6u53yBQj8+T1DjdnoCAJjL32UTmE70uqANKCRmsAtb8DToxo5B3CAX
RYY/F7vucfwpk+xGSlpSSbFnE7SMa5kh6r5FtZDJZrjtOWc13hxmXdN9TYXh+cU+xJuHiRmxQPFz
Q/AQM4i04Ru2AXL1ZNAI72QmrXaHXbn9helpYzMrtlCW3uRIatpnUOaal8KAbz3c2XH0SzRP/+v4
JlBTMQiWc/AjJGQHaC48RA3Suf0+M6nTYXrewfSx9VTZR62NjaeJ21KZ/1KuSDby6cjxTnSVcA2q
1vtjlZfnTTwtmZyYHFHPy4S1dpMyzbIIoze0ubx7HJ/TQJwHy3G50ftzyT3G6g2v4D/2T9vnYQWW
6IJZ8F5sLcdinybP9iy2wC06u7QnsSGHgJt23AOPT6RIF90I1BXQ8924HLQ6DpDxzOSN74U9H9Lo
/i9SK/ybbbTzSeocvomxuwj2d8NfBXUMYMjHDUsLahLdHDmE4JAse01I5FH7bRlCRiA4nFoCTzDK
/kkVDLW+phm8jUPuvak+KNq8exQvXWUO2q8ZOcp1omc+XoPp6V5K7JKe04r2XPsl3LGJFAH9yCO1
JD7MYWf0rwbV8TbTlcDjZFBrq6CL2m9yhx85lLXuhvjSE7wH2MnM79EECEvkyw2WTettUnEAzzJB
LgEMmkhL+dwxG4vsunXnrkxR4kDEAtw2Dhbp9gO95otvU1MoFkr6lc1rZZXsITLTGV2NLLK6hGRW
zYLDFhBgmjJcQoLgmCBewCsyMhWxvHVg31As6zAd59ljoXqdkK9/MIAM2z7aDvCqKSZf3p6o4mCP
8Rm1tqloN+Au1EB7EZu3zsTqppr4ndbQgzuOf3/7o13VTvrSlu4PMnT1QQv18RdBq1Th0eyM6UhK
jPFpDF7faUlDnsl/YlwIVwmIqMf8BlaZJmUfJ0JhIWZ0q1P133vVOIdrXMkRE4ns6oApCoeNNs5R
zsGkTiPJdEp3dUXUsJteyxrDSoPL+SJu1wXH2KndcP6XLx7juh24WnsjI1OhMqcXP7ih6RBXSjQp
ec6TxPosfJoV4YKWLU0gl0BPX+oXMAssCiJC8X6xat4w82Ncq8LKIh4152/j2hRf+ETF/1XFLFdQ
20vAtsZo1eteVDVJMuxqdzEwk7XauQ3yqGnKXkG+jebJdbGN+5ALa80Se7wD8DweUJdIkIavGHbR
c/zIdmGbH05cYUyGeu2gQsjpjYYBEAXPgPGBoOjXJ0lks5a/eRU8a7e+s5l8R+QvyPg4/4152Njt
fPmvelUpPTLqyvgwhkXdhRuXI5IxiEUqN1hC6JnPnO0hAokTx8IsX/gkCM0KcBjdu1Fpywf64h+I
6AXtoDxloEXtWXrVcGewLWYsZNSwvb8FGX+/SRCDN+JwpCJ74qznz7rwGoBvijlKcLsDE4DvMe8F
X0DBiqWWCzklmcz7ncUz78/VLcVn6BN0gvB02wqA4I9/3ejeej2huNxRG7omodskY4J5Jds8Sp7y
BjyvyG8NfGmkGnRjjrNmi+O7vMopNeWbcLmjap2vW5ISYMBL//7tILZMdSlfSRuwM97eOspXYJNN
wRX8NXZeTS6M2yYpmvxT/KnHnRWZQrVpSuebX6093bBI22+wTXixdd0DNyEIQJNsrjMdxdEnDACm
FaL8rcxfzY87fXTTDPDIy0dC0uEbP+obn23gwPNJhEAFY+YeVQ3X0/4dZgSamJwuIGf+ICr9u47u
0fu5t3b1HPyawiX82mA8J4RUP0At3kIVIvuLSnWfkxBy8dGAh2eQXni8zfnlmt/ZsEMppAARlXnq
oZRE07QUf3sQFZ7qEnoHW8xUC4zCUtSs6y/FIj2CFrzyQ2tFVTY5VwWQG372/IVHt0/sflsHFXQI
ACme/kd0Tj01FpI0pRj1RxEpoIY3C0qU/Hw4mM3eZLK0O303mG7ZigEGG7EdphEIGbI9gjdgLIcz
j9a49o8JrZx3zmfi219vGZ99CZece/s2EuzWEko2apOKemMZKGnX5kuOgeoTBpGtYpdOfZ0OOOMc
w796jj2IyMtL7NVB4Dbc5I6RmDnfXM0IRVgOfKyhoeiOI6HiPDxkBcBMV6WHsJ7yn52Qtvrf8e/b
ylWFT+Qi0L6msBjSA6JlD5I78Cph+cBkQ1e3GL78QLIA0ln1Y5fmpNk9Ce9JSzXAhuQM2+ldtYkN
M/6PE0Y71EHRUCRVQYMP+RcnMU1NpyEDVfRa/mUhjSQ6DsVNA7h4W6Ayc0+C4quqi2h4cQSq6nWz
Zrsz4UQl+0CIkSx5iiDKIfvZo6urz9k6hI2A6vc22Db8XAkMRsjGv+feLsfXA6GtESJc1Br4IxSS
a9+rIDxmFV76xZlTTm35P0HCxQ9T5eeqqsA962p9A7zWVZiY5E3BwmPJZ8HkHCVUHNdOQ62VK6jg
c0w9i3OMBQiBYyozV+efPzhKpAYBwEr9X4d/cz0fNTaNWpCCiy7dUF2RTm2OAM/J+w0YaNOwwMAU
Rm/OzLetlq/+K1rKEFd9DCiRZgs+hr1upwBSRaj9AttaMkcYOPJj1dXfCCrk8lg7vBobLSu6QC/M
hyYQX+qZ5XYys83XdZh+dLM39N25u/Ej5Qi9k6r6jWq4/sM4x9n22FmPUvmH6wSmPwKCK4vT8ZG0
vXvH8ttHxRTRIiFy07/FlXAeHe/jasMRPSZmlpyUpbGj67uxq7VmI+NDK2qyIwEe236VwTgwndho
7Y1C10cbGbvZUZT2OV1mZME5OJX+IhkYvIIeCQvPBvKbIj4qw+psopzZ+XoznMS7q46tQG4oIk49
ynPkHZVtJhXC1EnNcbNaSNe+eNp5jvgloFtsuFsD/mD9VByiEfsByAxRHF4ukaz6YhhNYyHkAgcR
AePSzYyzseFX48YyM03j84QLuJwN1g7RRikxYhEq1DTPrSK9blWnY1dNl83InorgXQ6ayjbr8H3d
zOlrwEowu2H99evLbcLwAapSpGjqs9osIl9ZDGtCS63sRVnPh+vWM95cA9UwqRPpsUknXzkj9oAx
Fjetw2ammJ9jdRTp89gzS0x4k2s95jfD30JGZ+CkPPNoxJjjmZv9QkpSxLBLd9j3zOI1gIq2I55R
gSo89lw/tGwD48/MWHG3K+aDwLuWdqMYFcWOJUJvEEHKM8aQX166QrP/8ipP7IgrwVbOsvBQIq4r
iBhKqxzuUMGl0e1LkWml6cu4C+q62boFrP+dti9hhlvQmL5v0Odmlltl4HQ8ChDKhF0uEeLIptXc
60mX90UYWmDUJ5CYRZa7RynK556wGQFF/rWJaz7Ix/YTCYgFmEb9mDAhtVaeEHTDBIWLBP4AxKMx
89dgytxv54IQK/PBH5oIBCE4Qsk7n3vEqLlwd4HberOPduFD5DIWcR6XnOV19dJpn0UVAmDEZhoZ
CWqIjSKU4iabUHWyh4INLYXdt3kRq+sPKDNi3yBWCYnFG3buKvtHQLuwd/xVcZoSjqel0FZAw3Bs
X59rkfx3ENMLfuYiZxpmQT8WcNYxhv/STmj/oi5snQXDbwI0pmzYrHoSmPmgjfNxLCkh0lXDdQw7
axhl6Z7+zZymRe496DdFh8+vQHUn2SzrYGjJL5Zf0rWLls35lut0MkXRWtSDG0zInXpKYQO0/rd9
ywFHuoTR8WYNUlWNsdppo+CTXFQ1sBO7zGvxDHlMfhbj+huTp2qK0xTbN9LLinp6iONg2YgZTT8w
ce2ovUhtAwHyoXtxM6W49KB8tv9Fym5QILPNnya9MMFPvZMW25AxCiZmL41AOXgFcxMxFZkpQzze
XOywQ/dBIALce8dy7kItvaBf0Y7DzTsqYZV+t5EA6ehHwgHyKuE0l+atQDp04ITFmzDZDdYFrvnt
BrA6YZmJ+GLeHGzf61ST7ZR2DMTiSNgmlVEmNmCIkicVnaX5yGDd/B1zxYFJ/0w9tgwhnI4ellC2
179jf5e6wjjJxfiK+gA31ehRJ+xrhXfx35dCHGtbBtAPmKLlGUdZTbp4fzpKBUF42gxDK0P5oVBp
E62kry2jvUxJEOwSEOvU5DiiPTCVm4MoazfuBu1xigsAoZ6VonhV8fXbTHJTl9ghlwcrIJXPFnYZ
S/IJV92m6sfGcU808pmbKMlNRzhJsIyCYcWAaLYUZPAVzX6CpJeO7KsvJND5sAPsmHVqepjIYPLd
6GbUqwg98S4IXi4xe+I0hGucpG4N1OyXoD/VE1fm53qB/32q2gvhWgS+6Oa68EsBhPEnmXNKZJRe
+qllTSgc/ZQH0B0Tkbw4E7DTgPQORoS8GjhlnuZdqWtngWi9DfwlCmKbTiCBWgdSjqxSGqEjpZhB
5pX7yEXErwhavS/V7jyEUDfdPHE/JF187LOSDjxJQCrJhaR8OBl3ERwiPbhHAeKLLVYuG/pitiPd
Xz2RTUCERJDZnVNb9ufmkuXmfo8zSJFp4PrBku28SmNk7vp1gx1b1dfs2YFIjD35laYzdaNlVeD+
qgdvJ9lhOe0w/B2HPnE5nyd6vjz1Y34rCSa/ij4uS9FBMGunAV1wMkcw8k52Ml4P4cCc1gT269yU
y2hnYatmEqjA9bh2SuPPVm1isECQoI14fTqbAYqJFkKTEx8ThkIblK+v51kcM/K1IdBhQn/6YHjh
h+clv+Wp8mq1T3igYJxHxJLK+fkvRXMewjUa49L4KVG4/i1PHUdhIsRFmziwMFTygt1d2TitCS8+
6ddc9lrH2gvky2xA80/mhuFRuTU8//9AFObaCE6Z6UPO0PlBWe4KyveNKitmbqSJc+0KvsWhzQHa
+CRBfM1HccDWvLkv3n1I2XVfPZjG5OqnFExSI8PFCxiP/Djv1NWYNvSWIZ14cnKdunNO/DGL38Rp
rJMyozIWnMJXcBg3xUAKqWnKmcbIB8NpB4GqzClvq0lOoRZy0gfmehJhNTxzE4zBzS/7vg1rcgKY
VrWA4weDNFG41SpU4Pggaq7PmGJ3MaupnVcFKwJUhFNDPoIedrX3zJuGWKzakFhHigB09BSE6pQF
tqSTZQ/r4RuzAh9u/M8/Jt2ZkAejnu3nQ2OLkBQJUO7AEi7aMZi76g5+4lCnKjT4iUoWNUhUHy9H
aIlJ7PFo9cuLkCafuvJbQ80oDvrmLlIKm9fx4XGugHbu/FLNOAjWKdvHiBuMCRzkumlnt9E2FMlI
KA/7DxG+qj00oW81kLCPNjkvKEdqnPVeaQW+VUriifzJbP3fgCAiA1Jt+sdkb9uG4nlKD+z64j5Y
OUOI/6buM01FYOWma0YzCN+GoHcYll2yWS6u2r/bqHvcxdQN2htoTLyKuxVGeTIkvRV51/YUmSpW
vEtgW2F2HRzIty7DTQzivU3DN+zFarVK2u/VGiIB7yZ7MRZcEqsmm+Th52XEWM52ItxI1XoMAHco
BddsRB6jRvQLsQPNqyg+q2Ivk+t3PjLXhJ7PUINaYetV8Kl2UV8GTks3NFN1gGFHHV3zhPDVZaau
X0ppxtOnh01vMFNmQiH4emrV0kziZ5bfbHKM6FdPV3svCKnjYFCotYmynvKs4/mpwsYE4WtElBpL
kDjN9ojuwMj46wKplIotWVBcWrzSDlqu1hypzXsfwcMGY0zQ6CnL0Kny3xG9OPj/9+VNMqhkNJd9
Z3M1tBGz8bLXMvfIdM8Qxaglg7OXksrZCZV1MU8v24g1oyLx8jlkX9JiOnoicJDi6k+LTWrExKiQ
YBEa3RmYpWGQ5Srpm/trwKIoQXUIIi00sAhHycBP8owgX5Z5hTRd6expKocuctB8wL9cyKfw8oVA
k9Ynn/kwYDHa/TnihRn3otPAfmXNfZF7NC2icLpVfOcit0nU8jcVjho4TNW87byX746RKqaBOa9Y
fdiGoi0M+IyjqUUZ2HQ8kIVh/PwhAXc972jTF0DnbUc0shHswjv2tdR38ZiIse6LUnr/tdYIy5Ab
wZcD7U0QKnLFvNyxreFTYp2xzU1iEpkaWKiYou3yRG1JwVrhmzJlwcbXDXJ+E7ylIJufNusCZA1G
HxfLm5tgU8ANCS7oMKgTjga8KJnFPMwR8zbPHTnbI7Jn1yIQ764XscDe6Un3Qgp8K6uFIr2+dcnN
bKVeaExydSCu7jCi0TpUdXaZ45ilHwSVNOm0nHRUeXL31GyhwSmZIU0ETlr5yeyEVPd3+Rphb7XO
1kDWCjHFSimeNzt+sYePs6qTW1NB8eGTBFPCLKk7CZTjONysDuHryFNoxF0UQKulvYc6LgklFxoO
cdn8R4NTs4ClGihHtM00epuXVOm5Fra2KlRtHH8/VKr17fLI1DSE6C5vAYRYt3Qsdi6/3wLYQEqP
FDI2WtjOCA1B4+nT0bORq2CbflKac7Yvd90scSZAPHGLV63v7WedQP/Hv/Uyo/1w6VDMPI4i5pPV
PP1KFNAn3CQKSCsw2cClgfOz7YZ56it4uQ9PzyMU0ZAkYKdjso1Ypeg3d2iTetV+BMY/A/8ZyC7P
5cWdsUtYkiwtdQhu66gFbl421qVqD8lN87T5yUBKwFUg2FQiEZuJAxLBFxguxUKvESxGdpg7MS+H
eB845rf2ly2m2WU8Oc5dmHK5DJzGJNAetb0PUDTO+ggypyWhCo/EtnDqDgJYJRc6IGrgMeLeS/JQ
y4Kq2nR/XdlkuhvdbpodlypAYEakuhFknQFGEN3BOYNv12ubWUrP6Vxwf2xbCqoXmlXWQSE3PKTR
R65t1sV9M5JVIaJ0aXPXb2NWMpVZkzRvM6Yv1eAXjDGRtsw7hdHNgKEusRitEGC+LLBpy2XAQepP
Rn4FwvJIkb2BQucdCKup02kTbpNcj56/BlkHi1c19c5xeMgMVp8LHmskfd4KnhxmyjP1BfLbAwst
+5+w9On1ieDU1jIipYjBTu8jsHQnYAYheuWEcsSJrLDaOrCaymJDIMpkD3r2ebIBET+nifK0hqlu
cTIszeOjgJN9knAFki3o8OG7pbZ7cTPxt0U2E4vg9GCedOziuREdk5EqAHFuLS1dVTixwOnpP/iM
4UAb8jslUgz+jceh4qAAAz4IZEGK4sFc2ehmxwc8kNkrnWDXheUrJAcDtWqugH96YzTD9afxKgq8
GW9sDgNzqFVQjxapua8xUeZLfeX+EUpY4oq3D7htea9Wd703I/go1TnP78r1DC/DpKYMxUnNBCMK
7hPcom8mEOiOsUQE632iux5qDZ2aXaNjTHpSZoKuc1WeNb47AJ9QSazaTmqSiNRjARu2MwJ0I2uY
zK29ahiY6QCk8zEQFr/efXUnwCPCX4KgNKvTtY09RsxqIioOVHUwU7w2IRINTWiGp9vWQMowE7fn
H98M9lPWaCniDMsbYw4G645+Y6OdcRXW7Nc4S3AA6tDyTH/uKn/pfy06NHOaZTeHzeMGRxIupyBn
yep6Mv1KG7LksmXf3i8V0nr/HoqHtzS99gmJ/v5fbSqo3CfBXjzciGgOTMegih/ooCthRsGmEl8f
ni6buPnTOo/ZZ72d+lhtQ3Cg4AnmsT7oHVUQaftL2yZO5a8k++OR8Xqd7Q2Nt4Ebr88dpYXEkPCT
2mllYHXUnD97ouYwAD+XdxTICK+MuybJUfm0xkpApGcsGTHLUk9+txi464BHahOZqsUc0M8jXsYM
mgloE7aJHNy8Jph1h6KHykv7R8eOnoo6goPOVsWdihDHOd+t1WfH69ZyUMTx+0VguVrpaH2rj98o
dBeQp0YX/IbzlBbzCuHpG4/EwAk8nDhD/KtH3VmM/LfelUpKpa3WB41jCEXpbCh6GEpbBLi30Boy
VwPLCsYDfyN6RESv/RhsznQ78+bgbvibC3/Rngqec4B+jkJMExp2LIB9Jxj9ItMTxhb8TMPQ2vHT
UsLEesv2Ptn1xPALr7Jbh3VDQyDEv3Wsuy1B0JTJRGVwxKsWGmbhGotkvB+24YvluWqSZq08COhc
6Bj3PhGpCj7MghGfCeVRSZtsmpkZzwITTtvWvVnpJtOGj0uiEPC3jP+d9cC0k1IBMqlowEF3vZXA
G5mXXGaSCpB7ovL8vRaWIy+6O3BML4SbdEqjijpRKpeATZC9Zv/Vz5wBfVUu9Eqp0o7aht9orNIx
wOznk+VvX848hpL44+Lt3ZTTK4mNw1CA3t8jdKHWxrAwHqwszvQV/tYrJPHv/TukY3WyUeItW+5v
GxZXu6v6GtnUx3dUHsV/DCNnBbZKjUR2/nB6h39Y3+opIfKfjyq/chNHHNwhtQp3YpVkbj4irHeR
XmKPF0FkjEY3XnrASdGQwF03eRkAdjPSx4UF64pF59K/sgywef2WmEKwbujN1w7nYqutTxt8C3/I
ZlcXXuF8sgquRHTD+jLSEVUTELudCEyB7RoYh4mxivm3uKxnf62ICePoz/kMd5kvp67r9K4YEGMd
VBIRjs3ZpszJ/7Jo/vYiIXZ8xd59dtTTRPi6NrA2S06TQ12c2C4U0s5Es+SLsKXdtKrZP1G8dfKi
7zG3yvdeiCy0MOQbOun6T591i5+9k/AJVvPtE+xsMHrpgvG9ipcOk2cU75HPm9WYiNehWw/LBJuP
7+BNsEMTH+suZ8C/BSY9H6qEQTMoBULXcR1C3/125LKCmD8/jlZbxlm9L7V0kkGRbRxQ3e3HkDCN
Ehpd2H/G8nhte0RearEXFgyZim2gI2ZjLi6NXrHOUc6CoZPufcRVQ2wLty5jSwwIE3N8L27p24Ja
X2g+bflggG3aYsVC3+fpPIXJl0MiDo0Mpyetleq1n9TQAJA8A0dTIdjVhgpdXWRn6hHkpGjUPhxg
sUpBhSDwAdp+fqqHYzmXTeaGVdwGFvt23rmsmQ52bBlUingO0MjbkuzoPxLFrAuRpGmKDHUrFeOW
94EeeZBfhinUkJBrpFYXdILrpEdxPibcokW3indkajQBU2W3faw7WHLIcI5S3OyqklOHylyQrqE/
7B3PFWMAdOLNSUPVOkgSl95Us8oD1N9vGB1/yTRGdWQKK3OwDcwiTxFciZIMLdjGpQeuArocI2A+
vcA2ZOjlc8Zxna2pNG5FbYIesbJMSOYaFluw2IhaD6AtZFKo5fa7VxrpVYFqiKPAMi9ukazJF+6C
9ZV61eo83wNWnYKSlhZfNhVMnM4uJfRVd+qvrRLVdQBfA4HSmr6IcORbkg3+og1cq0SsVrHVzsbw
8coKR86xtlxVlZJ1Sz3xkkGgtOqvQmvYnPgnpWg6H04T7JHNieZ0+tSQ7eXBCy3EhnWUSOuKYRPV
jiO95yJRP0mPL4ZB3LSleebuJirhUDOaUbuOQPedNpd/BVvGsnyU4gCoJScZSlgKAvnKkvTqNvCI
YLfnbLgK5dtqZRkh6ige89wCRZgJbIecjCrrrS1Qd6503h60b31nv/r0theVcfQpKc1rZq2ocqXk
5aJu/DcPrMwt6c2PpKU8nJLyw31XCOBL0AwwI5rzVuqaRfBDMRCYzj5ShPdPrEg5W27S+qVsshXA
Y1Kxr2mufZEObkXDwWnvISjR8S/pG937L79RMzVPqIgvZkTZPrNpuZdmyn02NDX27LvWNsdn8CqA
HipINNF2xxMwq6WveOEltXw1fjiwREr8MkXuMK3gsncIbQ1wXgQWs4t2iDjVgYinUORB5R4wsTuv
HYEr1IvELV1HUG6j56t/XFWRbTYJYsNqEkczI32rTk2rrdcQiqtfFNromKJCz9v48wEijX75zilP
9ZJt4I0ZnV1YMbu5KRMEvon4lpzpox/zQ1ydewTJ8z/AQNsXdjEriIgIZmN5DsYGJLjZyNaRj7vk
+TUqKy8X5riddkv7XwCEiwhG6lsUkSrE2hAd4+GJP2Xm6yNODuJkJikI+VyffoI4MqTrDsGK+5tj
JLlsaJWdHYVqC2+GKnepLonRr8vu7JxvthoAQH6dV1d8kBSSHBEHkmjXIwba5MfD/X066lDVm188
0KW9bkpEpvJOA1lAgIjSUC/mf5/aquQDUqEIGzfOemw/wksDC0CCuT9HJvXHAte5frL3AFNv7pt2
aG0B8orP9j8X+2TTub8WfhfQYZ0LAwipBwvmj9gTBOxE0/dYCem1Yyo0BBQlYSxPPCJt6fAcb0ka
hKzdOr3Z5q4vzwb2utYnLXP4JtBld+KgEmwCPAZJF94yUEKdR241tAWR5e7ea6D/233Sf7U5ziS1
sQJE/m2Anrfk7MBYW6Wil32lvaBfuH36hNjojOTP9t+QAzmiSel/MfZJsWSN5/JsrWDe6uerSafH
NTcGkDxXT7EK0ncFzZyOPpqtE8LRJidXbZ8sy0v4blr0kUMCTag9Y1qRmKA9b4/eCNrn+Po4qPkp
vMMyiIMgf07o6NqeoidMHO0hZs81PdvoxtqpHFFNBXrmAo+J7geNyPHT25WzkRwV3D12VL+FISEK
EunSJW40hIBCoOieuIpH1C46ySfDG73wAcvwwUrFNoNrmMdMQBWONeZMGA8UG3L2Y9cFltsJJ8sj
hAR13vHq6qwWpi+lb+mhEt0qrsdO/AOekLtorkeg6SmXlS8g/mg7weFLvK4FL0tfSlTo9xX3ykoh
rRwIyg1IZ3A77a1Yw+7Px5i4SM91wJ4I668BMGwmcZXoFBQPGYGoqB3ZQ1kVSZ63YtgLqclegPus
XMOUCHgbv+oBhOJ/bC2eHdaOWLHuzB2qmjqZRvYYwYsUOoVr3VT1ibV/1Fe4dmPYAEuqJCWr9bc8
FWpC4UFebTXYNhab6Ulw0lx4Tyf1yFqhayhC/Wt+V1fh+F7zKUXVh5tpvrTmy3ZklDfiIQUzKHwG
0SfAgZFphT89sjb+qyjohwzNGhMRhhI6D9i6AWoj9cUQWUhyWBqcq5Z+8mi6bTXSqjyl3PxPzRl9
sZiGJ/U81zvMNaW0qxQ7mH93V6qmeLIvMUMgxLxxWXiHONZyNEyH1iFJi6QUX+5SrJDu9hMDYQt8
osbZZZ1C6s7dVzvNnxyMb2LCJ5yn09rwVaRl10Dpm4zmYZg19HFRty3UQpxXd64aEPgf22Q2U5eP
223Boj6lTJECDuYznjJXpJR9KYjLg+pb2YitsTYatMM9VtC+Hn+oZjHX+u/pvk5kUDXnd/5wy1SR
xLj6a7oT590vADSURRjwzrrnzg/LwuXlFPWO+nkrXPcv1IDmAxIUX0UITy+bM8Z8TgxdBBKQYv5y
F6g+AnvsEBGXghvxa7DCuNYwlwQWDWEbweFfcb0/0WDXbbS7Blf0ecQo/WtAK3ip6e6wzt2MSEXe
r88YPKKgKAancVzyOCLgpo9bW1aj9MIU1p7IcRQ3RrDknZPfy6/o4IXcCot8JOY3bfcHO7L0RYQ2
hdSSVahVGB6QPZwJ52gquS/IdGdAdd/zz3Sm8dfmX+u42ybkbro9iL8uuLDY8Tpex3krCNJFFSWG
Z01zvGAWU6BnjMYSOAGurSxfiZglgZyuM3/IIQZaNG0WdWtSQuL9AHbr0b5aLpKLYe4JiHhiB59l
RJiLwEjfe+KgRSnGpsYb8bkJxvRwHBZE+g6OM+DNEC632IQw3r/zKBzgB65gJxUyAqMS6x+kHUSB
ckk9wlviZgmxRAIDju7DMEm2k7ts9Pls/a48vKCHsI8gsFm1VPlAlbcQkxvzaNfxY5sU6SB5i2sh
GSutJASVaFujyowb7VPODNWrjoGZJK/ZIm0FMF7K4Yd1x9swFkwImMrLixEmaiXYqHV10m0ixUck
vb5PkvaQla3B+qtM4nki6OtpWek9NeSvp5HEvopDVNEuTobhHGv15sr2gmiYV9LpqlgSyPdm/KaJ
G9+yVFewHRWSY1Z2nG9LmDSOTP3kGDNaOiur6w0qybZ88mB5vpJYvj9uj/QyGSXv45raHQ1pbgwM
lTBaHXcdzYDhmRU+ldVaVS/0XoRt4cY8iGj0mc5D7UJ3coCMlXqPwVCMtCgwFIYC462TsZ4ppcFU
ijxD4bOCYZvGRoIUzp5Hf2o2KrSy9L3x6+JU7/sC6c68LMnN1wnnR00NRQDwARSrOAwf438/7Iqy
T/d0WKAIgBpOtQJgUPRuC4Z0IRGEO0lX1mIq1HjJHwBRu+HV0F/udFH//Hdjr2sv2E7k+N+Mglae
eHNZlv/MuL4bIvw0X4xLGc9wIf8a5AsaMO9CU0D7vx9iKnoKQGPcYAk0WvtMkinme4Kv19dUFGuM
4kBIfUV8hSi0/Uipzq5/A/zD/5c12Ivr07ujFnMykseADe79d7hGUwkQVYp9AaNv93Tgd9kEhU3l
C8NksbL1ckFxHprHlGKVLxSRgZR8aJSH/BwHn3oOObWl93SGZIMbdY+RGjxdaHPqLrpWiPPUeE0C
qunbBFSF2rWW4j+ZH++QlXGD8oBvAcdtNu0LlpQKvkrRrGK5OpGq+mdS1vqDtNP2P1MecBSyBHay
Ewqr6QRPNMwaT+253R6UpqxRChRTCYYrBvUEEZAgaWSYyAyadmoxxbsjPfPIYYWuWXLCQx2gUhpl
8rJ2qBTuNJ7Ahcv43I38FKN4NVOHmnNaA+baaO6gR2amksa3AecVDJLvvkcY7J+eLfH3ZrVbeP9R
UaepFgvt+3twdfakaB533TAAlvBlxGrBwjtwgHA5NLhQjtHHT74VFcLpl9/aN2H/r3HnkLEY+Q0l
X3YDq3I77VpHd74W8Phf36Tg1yQtQI+y5GUoMHNjwchQaa+GHEJP9gX9GPI9o/xghN3ihF24lbPX
DeYR6WaaNWO2N4qn2RVSNaUC1EV/bhyHbiBapGjnFExbXnaK3B1pX6Kvi0/Wl/rUxQGYtxOzxkA2
BgWxoiykUh9SIQs/syZHjXc2hpXGAU60B+pBRbvly0FBThtP0wgE8pKt6kAlxx042tjH+c9UmssQ
XG5HxgR9XCtbNcdK1IhQQuKjZ4Jn/88DvqfSwmmzJf/CRjlh2GMqAZLPfn01N/RfCodtx+h7WzHP
BB9XeTD+k1L00BkTLOXNfbE4l/7Or2+0otnEfNqXeWd+8aLjrQiXkkS8B3o5qKzsO9TagbA7fYiZ
qtGtqGuYVrD5ZVUFINDOdbMdAcZ3Id/4Y0oacrMeZTxTrHvZOMzYWT+1kodlcZyN7kOJpAApKjvB
pGqwFZ474+WHVzS4UULmnstYGrnm5mMDbgv9Dr94raHArEL8tHqDc80973MyffrMDW+b+DKNhouA
zv+TlWKuKzZjsnTR/PVLt50t0/9tlPxdluQnuKyRFkKpHo9dzL4OpAdEvsQdhTdfV6puqo4iu0ym
bbbWSU34XA+M2HpIMk5bw0jKQygCX3CH3GpxxfKjfiFIE6BFPNP8yia4fGDjLjZ67ve/O8Y3kZ0N
V1bXZgTsR8K0MFb/+CE5WkgjFmc2wCLuiIkWOYl2aMhfEAv1rIaMiHMkVaWVrOkgXZTLDV734teX
qY2aqh+gB+9mDW60qLEClzAjO95WTOUFGddlHlyTQcykUC8OKhkYgqyjj/g9KxHsE2jI8gjj8g5f
sy++at7mDxvZH8QlI2f6gAG3+mRWaGDws387gp37i096D5xqOQAL3BfLWjKEw39Xxx5h8LfLv6M6
VofNDUdEaqkRxXOwVYn2VF19sKoP5hzaZfsCEos0ihA8Plz29zQF9EnfihVtZ3owsayZvkrK8Qyt
+TLtVLUjqjxyc131YlcF1+5fkgI490MXOpapxvkSZ2hGbduYwNfKq8LxlFMn516aZOKWy5RR7NSC
WIwq5nquEFz6nCzIYlw/Z89CJbCSDEkA62Eovl5ftUl1koZMOl1irp3Hg2ZPpmtYI+KdC/GKMBPo
fIKaVZyAh2IRDHirrBQ0y4OMYbImqC0q3HcftaiTzgMrg6Myw887cNBFcGAaMhXtrPlh1IQswDn0
sOwo3bG4JvwdmVv7QOq1aLkG1aiXW6kF7VdE4Hvv8OtK4aodpLa/kLyugepfXbxOhCSdrwIinC4u
IkaHcaBe1AuMiWrtLyP7i36SCkTimxnWAH7ECd4KkFy1g9EuTa/iDqV7FbF5IdEKppZSv0/0geYk
meN5/GUirwCETWr01wR2Dhw0af/D6hVgVyRiEpJNc4fotZU6pbL56Jb1GtmR43l449+q9YLHiaXr
yD/Xf+CG+stglaumGk61k24TBJevNO8OPT8lL26ejXknI5WU+swu5CVnqDVDLn6M1P0GjNuGOdfw
qHawfIV1De4QHxhXTdw7Jf9Tiu9JDbkF/Skz3SOOapO6I4nJ3icsHrZLQKPAMhsTcxCFNBnFE/Od
ahanH9hjvtmwCOXLVcB3n2WWycF9XQOp2PrCDtf5DSFEqSkES04pxDfEe7n6sfhKEicx0yMPVyMD
YKNs1I1/wRQt4O0FHGT6V0JWR2sEiYLFTqBOHEKSPpKTvBgKqOuIgSZJzkHC8GGiGCtlMqaUtXAi
XC7VK4Ti7xBtWjUFbnyDk8lPqr85F7lsx6/Ec8gm+1HoWaPPfW8zqJ0v7xSffz6vIYLhGixwKRej
jYciIIgyQwkYQ4di3rc44yNgXO9jrjVORje5vT8uShhFRZqe2zdN7Fg+kIukqnMfIDtluw6tOnQd
DoOXbmeqwnj6w6Q6h7BQwVPHWJsvKn7VRffIOQ7FtLdK9QY9JsaoAFUvSoEn4p/EI68X4MKNOp88
TkDVrrStyNSV1X082LvLUC7WhEuNPvthvdlbWpGcqn04h8TsMJWfforPQ4UdXJqxNpoCkbK7AiN3
5xFeLcTAVYnJhMXk5m3UvMmbfInwRh6VEFf0f1+BY8hJ6siA2htO/qa0vutWy3ug5kHjm1u/dM4Z
tSjrQyG8VndIRMGJDPNPW3R1gPMS4DdN95afWYI1iFWoNPzSEKvpFSyINKJx58ZbP8HYatBBPc+H
3y0t6ipsizTOTVIDublmj2UxLq9LGLSGWloJUZ3qk1Xsq81tC4voMH2rSC3CazIh81xBW6slgtsb
/a632ZACmMJV5MbYhf07yiMDtut6+2sP2uxzrn5OVRn7ajiK5Y1tfA8v4k0U/+GdwSMWSWY4CMA3
CuMP+WVpgh3edTL8t8PTkKYTaIKtNz3340ptwP6HBS3xZvFX2C13jzTMQQm8C5cG0Mlwm9fZBZ5k
kTNPoQC9mCW8gH5V49X+yqCD3B/DbeEPM12vyicvRREUqk7IfG9hD2IQfQcbmpl1JFXlVhIp+BNC
ga44Fu/NlkCEZMcqxpIIzAgwZXg1nMqYDGdkoXK52dHojO8bcEzkHaeurl51+M7ZgXSWYp1tZgLf
V3Pe+pU/71Q7jaciCiwM7A3FA3O+XRPpG/9a14w2jgnXxRytzXjrZhvKjhg1+4kL+FIcRxjZuJIN
neMSQ48foFButFsIhUEGMvgHfaemRHXzubSxmlshglYoLoTigGM1B+w7ufnEW5WBqwGDlg+lAVYO
pIlGODebRlLUWvCjnrBTNIJSEDUxmVHsw2kH1q1YLUs3FzuFrrfh71LiOwpO+zmzJX/x5m1Ca3CH
9pPMhCgi9fDq66cGSDxwa1/vazwWuEgNI4Y8sLAEW4P8n/j11/e/PJwUdz5QX5jMGJkSgaPR0mVV
lAJC3/oA8GzzjLO1iYUU4vXUMB5dIrvyZxew/NrBMOKC424Q0FUmTtD/jb9FD7y9Tz/gzksE+mmd
QLVUOGh8YqX7Z4JSfUY68IPSqn3f6Tmz5k6FsJCkx/1Hs2sK8qwdwkTltN3dpqyWaeC7FG6/+/VN
7lkI0A5suodv56q/eGvHLbPKR5ts69oSAHdf4Y/03D2mwi/ybxBKqY5g/SrgpsTfdMl3BMp+u/d7
RtutTnMgNfn9ADAXC98yKpwqFhx08WpkP3LQcSUYi5qSxDBBgz+n7VPIUJC74A525BOsuuAcmcic
6IfwFiTAP8W0IO9UDExeP9XtpIIW+CD9htGTOVtWQG5PsQQ87mp8Gm1IyKF++DRu2QXajhdjvGd+
BHkqnU4+1WLJUAmXrwxX7Tpw3KNqwIbAOzNEmQ39BshcsnjG3yT+3hDDdT76uBq7mKt+Nn88p3Fq
x1utBUMS4kpXsqK6uMNVVd7uoXcSkAQB4+MCewuqhgSV62pyx5BA0Qs9Kt/GVTKm1ZWrNB6mhevr
STkJUqkRCzD1jWcVAT6JqITVOjAFOjpMfCxMEZIam5+NzNOSv/eVdoQ8A6lZk4zjmH/rHKoIAYvC
+mntq4+ux0rtdGGGIgZw4IDwprnOZzzbbt4Zg44FEj1I1ok3spk4vZa1pqIdLDzwxlzH68gxu4bs
PCI8wO2kQowKiMp1UU/a14n9D9iLcZf75ha4fkkyDQB+5Km0YxDJHBVfPrmxQLd+0fn7jmBSGIuY
cA2D9pVUrMymIK8HZbEPMMTAZySySUDLmyHd3QcgWuduCagYV/mnvB9HUlkOjjG91i0U0dNV29p9
AV5FJ87ltmd1TvSN0iO0BQMarZ60AFz7NZh9Wv3r127msPxHPZJ1XH7dDpJwyu484UuPNKdLGhha
b702rpaAl7xZG5yeEKMnIfpB5b9BN0WL3PtKR3jqe+OnI2ovp7rXnboadoz7Zd4gTxfhOHS1aYAb
d5YusP3PgxgXZmEyGTJkGxzItgkuqW9IhECRfh05EKaeDwfdsdDZVLPZcCf0khnFh41apNNxOKlp
s+4lsIdcOU8XmIuhrtwxj/O55KAu9Qa+qypLggo1N4xCMfqQmUAsGC/dy1RgPx19hiK4VyT3bBys
WBS0LsEqdmwkKNbbp+HreEqpByABvsopeQ0gKOhatKXdtDhaW1NgpTLldjZ6Mcqzt3lW9+uTAuJA
bGCi6uCFw1niRQ0M+goNEwAe3vEJsaoYLxGW5qeNRQ2mJjbWc9hOTRJL3NIZ/JR13I+eEKb/v/E5
eUhei9N0MK9K+33KGXXH+UuckZq+EcldXgiqvhRZrWwNZ39Rn4O77C8kucA1iWOlL9lg5v5/PIqw
rLa3AsFmTKpBG7/HryNmFZDuOKMgY4Al0mqR6sU3JphJOgA83u6AVftHmkctQNfCOwYzogB98Z4I
PgDyzT+ueERBswP6Rnp4yUKw1S8bXJXC21T30qX4417SxmP5+xJdgUiwGysy4SdSF04HUWz46wOV
KX2ZeA21UbfpznxhYXZFAd+gdi0eEdp7JBAqg02XNdFmdcReTKvF7tbZeDZMSMN7ANdeGTlLSnAb
8DxjgXEvdoXAd7zhH+blxoth4Jx8qn23TMLP8pwCVlOrrGpdVcT8nwBxaG0ZjoW4jagbyAFR5DIW
8gmyKKMijlWnSWV+m2KMd5jNnO1A088FfhNeVRY3hE+lZjPdmj+HdV3COcT/9gVcTxyEbFd5axDd
4F6y6pWD9TcNopozuIFxAJfG+sRn1Va1Y4SKOoZgyLpvB9fevLSehT829UQwUsKABhWbUuKiVDbv
7ilnd4KXeWE0NlIQssMbIstIf953zeDsudgdIBh41h9kSOI+75nlHtc8ZCJo0+ainWaeDwHb61fM
1Poo3//IYDFm1dXyG0ua/5VjVIInRKdJjXXnBtcvlO2uCVMDr191upoJmyIA5vWvwvSo0mjj7Y/G
C5Era/9N4qri2Zqt7IkBVaIEAKYxkRVqDmqycZHec7b/10VSzZ3h4+cvoekqW/1WtPlC+UVr8Y3I
HpP9E9R5Gc/UqRHd1djibyKYUuc2i9boiYhgOH2W4mcmNv8FheU5YntmdOLCaf3iHIDcvGHQsiJQ
zax0bT4Oemg/clLFD50Ljyy9x56Uv3yTK89d+T4Rf4gCF6m450IGJxzhHW6bZSYYY3w10DYc1aG2
H61IYK6zPMkMUPNqc+bO0hZE1Gv6Hoi6rKi1zgsFEEIXVUa2F/SstqA/onNv8QscN1DNekyv+71S
6eVzH3pI9a2HMtyL3pS6k2jHaQZD94OBPrj0b85QszWb8Ilttvf4PEwO79Fyp8oFQxg++/iSApiJ
j9b7Ddr780Y+kRERqCjnbaJdpcaTW+HjrIO8C4me+tVS+CjzP4S6E2px7hyCJFbyqtFIuu9ygpk2
mtNGR877+Gn7dQTd+qM5B6V8Nzq50kflOXx3axjTwXwFUppbaQ4tfiSPeSsSdpgwd392U44mDWpH
2okxkTQXbHoLhrsDb06uGVERzN6/XxbFtPeI7C6KKXpvA1fGcc21m3LYeds6NUgFOUVvMoDhZGLN
TbX4JEP9H/vI/n59nTYl1YvMuq3IFOXqFgmZOsqIprGYKZZBb8qyM7VUgpkebFWE4IOMmgaF3/cU
ctg2QjUryRWmQmli+T29+G1bn5neQq+PehUkH4TfDYeRWE5qqurF26rvnkJTk979kD3gMDmmABf3
V5SlpeAtknwLk1zXYnY71VrTRHzOOZTQaRhdY3QEYFEF3hN/fZJvD+dd2qj+pl9bRSrmpiffR9v0
vfnj9gbcXBks8+XNmYf8w0+obNiJQjvOoN4pHnze/Q4uzKRBjZAV95a4owFENq/oqijUEoqK+SLB
jhAB1h4iUfwBGQZ0aIiHE/YFCJhviVsl4J7hKOepa3NNKamUYFAu/TFj2AHN8aOh4aXtLF+H3sCi
FYQ+YHnhC3HDw0ZV3o0osXdeVPMtzcsH62B+F93XvhkbuuiXSmMSOsUqB/KN9Em10F+ISvqx8Ini
OD1eWfmhxQPZxvO0E3HQ/ZsY3vXS7Ok041MidCG+R4/39J9Jk48QsvyRHyDzCymo84zNjNQAduf9
v4SsN0iwN/Kqn3/Lt+a7mlxWOmbU5SKvv8hpUGzoExUjzmVByWjf2uwrdK1biSuSklCDTVzueEFY
1pS1DtURyygsOqpwYw1WXS6DRy+VasbWRWwsjiYugK+Gz1UcLzBPs9MYuienrqrkuV7w33mn6KN1
mEWDOWF+p/qC+vJ3CSw+skTaggkVS5ovqVgFQ4ZZ7k5iH6SC9kf/ReNrku9VQiPCud6JfQcPdlPU
eaG45BZdgAP5ZTz3UxIpVj3gWaQIMaoNIgl6F4wtSfafMglXi+TDdFkip9s6E4lwPsraLeBBldf3
QOYNtW6WP9fwwzGHvh+Yxc2cOQQHdlZ08SYVrEhV7XptniJQFpWzkvA8RFzieRK5r9FOO4gy6f7L
s7J2eiIAIannafJJQUud18LA5Ol4QBvjJkpxuLzB5CHPvhO1VtaCJ5KP4/GOlvKtiMcc41G2U5/V
AQNny0MuNXBRGYkvwWlLZbOugDpGORtUmlvmQoOzR+hRYb2dM7u7thcTwdp1RTwWxoX+7MlRmyJq
VMqp/NLExHKXSQczjhFVfwM1uKqYVjg3JIC2Ha86wng6fob5Jo0pbs1WFDEdAn8HTb6iJ6Fh9Eri
D18qBftgiezUydPzMKoNWSJFguJCIwmfVHgZnC6QHjSxxZjRFbJ18NpNtrDtQMUMClLYkK66fRBv
MrW9HrMu1ZpjwgVWNtZ5geJ7UxDUq/NAl4dl8DHa+U+lQnnc+y9kT9OnKfD8qYdkzJmoaERDRekJ
Q7VmdNvKpHWDkllCdGnhmIGHVbqdDsPvq6mHHJbQK9nLMmJ+rffQky+78LBneM9jQzbnje9BWz2r
6d6vYB6XIseDJ2Ee1P+8Fs7zW3bMIAWJ8yk6/sJIJxoGMO3Jt9yF+PAzBKUFsGbv/JN9vQ9iQkg5
st5TK8u9m7uA87W5xoflxQ0zCFhlCKQwCtgg36MtLbou2Y8WQPzq65s5XXkgBFr3RJr9L6gAsrYY
ykhGsAJRQ5H8kkJ6EYqFKksJ3DMCLbR7O1WnNVj/EMWMpUFHAmAGLKbDGLTWN8mrwMtwTogVoqq2
c25KSZhUXz8l6CxsvrJGq0TKAa9NxRKy1oigh43fNkRkU9sYB47jXmhL5aRYdZ/LUsqRltJBhvxX
WMV51+G1QfbwbXloK1flPotDxYsGOE2PO4ePJqQa5iTTW3slwdJUQ5488IXb2m6AOy/4bFz9u/5z
xqbMiLM0GS5pV7IzNA0vy5p0GalPpkY60vH0BKGK3AOQYQtg1uK5lB879mvoLZ01eIUxD9Z6rkt6
WDbPuPJT88DcerPhhJGPZl26/8HKXGL33lAEihHDAe9iE0GLXfY+Kf6Si5wsf2xOsFyGdnrR8Y6G
b9euUiJnSYdPRU7GlUFBBR/A/Ehh6PW2LxPKIUs3/xwcpBiTb8NKwYtqkTV0ZVbZQS/V6aB3u4K7
OH3LN87uBplG48VtnmztzTOU3g41/IQyd2WJWSQbkbv95wesihEDLkKhp3zYuZkZ2R8nduPPr6+/
GTjRL9wabQp7ThyMuHMq5CJPdRdSfbKHVKqFsG2owQpMc4WuO5I0L2MZbJsATIqFsLJUM4E0xThm
bOIfokBd9n+uXPRfU0XzXVgdx40w/OLva5xtXvdlBJkPQWg5YZBXGPVIZGDI/+RHVRSK8m+rMtJG
vthWVLqt68WZHNx2DcEJhKgCoPCTznYU53EABQBZqpx8otTz0aLl9RgWaK2rVFNBVv34H+i/FHmz
FRANupo82AOBaYB2vXBay5tC1mbt0inugBFSkSwMWnG7KZIcyInuJ2zUM6dhjwVJpZMk7eBSnD2k
c4U/qR49esQ7nhC0wH0z4U/M2G1xXp2xvl4O6Iqzp3f5CzSvikFoJZ/SrY/40p9sC3slu7dkHYNv
SShFbyhYNrq9RhXRTSnCF8d+7xqPciEQFNsSWarZCDdyl1JhwFzgMWlSmBnXvPCvbBLhrSMVWyww
nUT7Z1XZTTHAx1GP2l594uK1No+swXL49kmj40oGJYvAhwbGTL6wwg57d72ZZdlQMhZJVciM8G+o
c9tLQBv7Rn2whDzWBoTFf2zisXSDSdbFgtwu00KUZ00Eld0KAexsWZvLAm5MOgAEPD1QopW+Vk8u
Dg/RAMjX198OunkQ06r5KZlydCzlWcc6I2pQEmlTysGB9TInAzMzMiTa+2jjvUl4i0YOgMnVeVxB
XpuZWY8UmzFLhgywZDrurgr0T8UT2BHTiXXvp8TKIT5tkyyS/FeGi+jt5cBGIoGgJD/WZ60eXdcK
HHH6GV6PW9Lx84TtiLcOT+Obddlk7jkMoT672TG0S/xgFKosjUE44nF5HcU7hFeHbyTQaLZd/Cyg
VfT5x48vvwde5CAgSKyplHClGMveVhPtfe5XZ+Ap5/E9YM6zttr27a6jLTrkla0GqTJa0R5988rT
NM2nl4QwnQpFQjWw/J7GjFK59jW6HSCJMwY7ZM/BN/y5OEWOLPIMkglzBwP+QP/gupK269+EPdcX
JsSZok83QFuM4wmuVAH8hj8hSv7u4tMpuc4j4n+cpoDG1bsrTv9UnWCKR2hg4H0EcptxFR29kOYi
UOnF88Uu1G6iipPrLq3c/vKwCC0vC/93REILpVMk5QPeAyJJVnAQpWfncfzP3Y4djjIw4Ni9bWOD
XLSM28kYp1PENgVqeINbG4SGU34byp2KOeMdMFjLLftmNCfn3mmq8MOcxr22eili3NH9PXuBV/KA
QrY+W5frOCP/IEam5ucsrj1kJtnWnyK3cBfUIAqGlTgqT6tVu4mvr5u3O2+3FnnQzTiB3hZjxGmG
/FofoHyy5gZKCgTobIrK8xnhP43dGkg5/k2UtkHaCHscRfdD6rJOy5fgAA5qkMp+jLacOtJ538Df
qgG+Gh10KvQNuJlv/XzikQ6TYz7VXvCVqdEM4FisBbV3itZcJl+q0DSL8Igr6pPqVT/NcY2R8YAC
zI1zk8ud6f3sXFjViXW9mlAvwTXXNxr+MVH4rw561R5pRwLZUWTygQPGqFSH0HtKPAC43Zw0Cdl0
lCA6NnNjAMaEQpvH2p0XhbRkdYw/DjI/rA8TSDtqUbSbj6VYPANDhsFweiZrq+kFi0oSziA35lVi
iBSPu/8afVoN3/T3L9yWChfhWbc2ZNm2iPEx7VbUUs+mUN+6W42iyCRC/71/D+r/U045/HhBFiIE
SAsyo5grmO9PfANmQEkld0XU+2/hHkSu0bXu0c0FoWktt9WReaGN9OxkDpt2GP7SJ2iYoleCmYI6
4Es29dP4LEM8hLjKfnLaXXpbAYLjO8JIw/MCFo5NXSbNx8WWLmDqJ7kEXoRyRavyuccr0ob42tbf
ROWIY12nmSD8WLVBl5B/Rg9hCA0o076O3L2uy8rCcsP47QBg+9j4rVVxg/f79SsvHpK+ra8bU+WQ
TCmcrS/2GIgLwQwXEos8OMpNCLOhdVEjfBMQTGuhjQyMBezOyHEWzAhDQTk8+4Nu9KOPKNh1omhT
J8JDNMWnkHiHL/wQFZ5snpi0PeMQpGxsORiNEMMDLjEdr5DvWaGwyx4Mhd6nidFObYID2rAKircp
dS2hcoRlZjYsSicjQRZHQdxi1t5bQP31uxC/SR1RxrV4hRUx4NBi7YhylSN6CLGONo4yLMwyvdg7
BzxXSgQwXf5kecV0D1ARVCq2y1vo9FDjTRvb3Q1t1Ubh19GH3UUsObbXXa22xb3hfqwq76t0WbRN
fiCJHZjl3sX0WTmdKWjfAwLK1d212QIPe4NTBGxBN4Os5pPsxJe1mz7R0NY7ldX9CGj/0pwsiC5c
rCMmdTlaKhpNA+QAUXu2rjm40xHw1lWSBhERLjgvdvw2qBd9Gr5ECmbC7GsIAHKdqIjVr0rPVscf
YTpNGAqJdP7c47NbwF2kQTAzmpiEtAYpmCk/9U1FOsTOkXs0c8GJ9YZ4CnnC/O69pXbErfBovIh5
f2YG6CfaP1bAqJsbUMJfjMZKrtK/mKLYobBaIXzD6ywf1eencMWcUokHftljGvTAdKdM8YBsrNLF
krxdxllNfo5bcrQvadmrPciZUNAsheywdYXaNpP0gTYNhkU6dFj3KOiU2b1BPF4jWvmNra9bdDJ1
GqKpC7XYf6as+VrwaX2iIMNwsQ8koTIwAISUl4GXs9J8xyN47jkgWNDmI9DHU6nQjfhaaxU96/OL
PDL42wY3u6K3a5RnRNNTmBqw6UlW1HH3+VSbTR+sCz8KwDejxkuCGtLuq1O6wl02WmuMrpfZXbH2
2ipRfYfAM2gMFDYb1p9eAEOGp14Y9Of5kmzI/EROdZ+Eh/JsTB9dQRJaqExZzEUHWer0rRwyRSbK
D7/e5dwx6ZgoQlYn7bHdT8XP0MlXtIwIFEllf0sJiN8o1k0w82O9OUxnfzXarPrtM8ReUH2E3J+O
s19oaL00uTrRipG2rRHmZvf2rXnE/c1Y4+q4uZWEsMvu+w1gVBhK96AFb95MYBHpfV3z2gaRaBF2
Z8dErKrFaIIPKtx+xYTEtD11kSFk0Y7tGaFw2UBMSV5E2zeN2GwwtDhZxxu5cZbmuCc0oeomr5yZ
tZAoDw/Wh8zXd9rj4o4HIGmxxh3NbqAOc6Xg6RWZHJXjb8Xhs1MVoPQRWXrMDKvvNy7VLdIW4/Lg
Dv0Xq+8Tf+6m546vOh0ipmaEn1fjvEohiu79Mq/gNBx9BEA2vnfbfxmua5TTCLHuemIfY1wEKoLZ
azKszssacV/6sJFfmWpCl2UPls+XpexcEuCt3gbi2pUSZUch7FSUgy9Vys2Dz0NeeD0cIeNXRas7
u8AxCPgUupsjW0/hG7FIdwtgUzcJX841W8I2No2gtKVkvk1dxgFj394BeB0Wgtpcnrw5Nn16O3w3
SZQkezrJa/mj+YiOmkosur084wu5alvInTQCCwLr/QjiBEpfc4jCaAplnUwWqcnhRjbrXk2lkCYX
wBRQS7yqsp8mA0QvorHj/1T60OHrgHZ7QeCSQOPqwuC6bKa9bqHWSFfKqlY0WGwMOx0DjXj+iQT1
1tN5U3/2pv12pgK5HY/kCgriYX1HK23uNsNE6EqSinFY1z/A0sJpfwRktsZBdWoKqimBxhHTy0Bd
idAmTmN87VhAf5iY3fzPe+tkBEzkqQjddEh4vXAGTA2R+GjEej0efxkUP2+XxdFAHkky3JgDplxR
sQhmeSXeum/kBeVgD4TUUFX7RftID4puOJTs6qlDHGsLnyctfgRQ/HFE5YRpcTZ5m3vduefy7QUQ
2C80cIn9c1PwSW/tAiqfOiUb5RXV7GfTS5iE2KktoGE7LBgL4LkpvPwXs3dwX+Ik7lun837P0K+u
144retJWtdqOcQ97t2AbINu0Tx5dKu+7YGQBemKigpp2V8pivl4VCfejwLv0uRzhQlNFV2tqkUQ4
9LgNUkC0k+8AXHG2BXFRAs5kIWwq0C0rOmPI2NY8txZOPUZ22Y2Qo3n9B4YmHtYE5UVfMqb8yBWz
mmZSmd87ZuyIC0eUmPOHzDThE8N7tMjUyZRAXvNACTibv+gH/jQ1Jwnw9Cxi7PkAUjoiNSr0WQed
c4RHyiUeHdyjQIEW2iCtCilNJVtVH4tBnzwyAbKbvOWamkEZ9roSOLfaUJWWKPQ4NbrkOtDOr1rL
jMdi9m2EvctEVLfjZoOYlySsClkX/gAbyGulAQfWXEz12C7SUGXNyieimcNofFAuyWPEvmmsy141
jYDq8mReYmy92xeAfcA4gkrgZ9Ti8Uf0NXSTAqm0qmo2wOOgJFf9NAP05yGUrDxTi+E4tDFWqw29
cgxAQ+tqq4wEsieJjHcbvFgKBoh/+Gii18YGJ2WJ+ISqBa0wYwMINvzKvWOs9JSiy85Fa4UZ64xN
PzSu5JzbzidHBvLCQs0rT3Eh4rrm1jITiu0JGq1Y3lrlPuRsZmhtU5kxFjMvDGKTPbEAph61yRCw
MMMepDWRFZEyXlXgrUEcCirCFawquGXQVeeqFejFDBDz1JRpbgG4I4l8SZVVL3Qqla90XjH3gZIP
83aXrtkXGLAH9ftYjOnCHfR+AbxPEitPsa3/7gU4sAKTFu8L6Ae+dBUNW/5Uw9j20s50U1Xuc8qO
vh5ieSk/uMyFN1uyG8/2pzT9vaJSTAsveBEjx67DoYzNndJ7199ZTcnz1F+lVm5WDtEU9zzvvJCw
+iRTrYYHwK222IKyWFS+UpkuOp+1XsN0g2eEtVNGGqTrFprbueJQ6TtmeQAQHkKy5PNMb1/8C6F9
+9PuvQGWiXH/OCBK9rT59cN+ADLGuV4aV8z9JbMrKfNcyRO0y56RujeIzouzPlAH7hSIo9GMqW6a
Fu54hcYMsHp/GAhaV6r9Isf+XFBiX+aY9XxTwUEpeZb0hUpI9CISfhFiao1y5VlEL9P4zwbBUt2B
2ILQPzKxmNfnZixzo46R9eC2V5NF2cvnf70WYrEA0+QTUyfoF3IjLaKyquTZbdszDOaE00/KwyBh
drj0yFZZrR7fEve9WTawJs10Sh9kusmaHeotVQf5LDN/LxxvFBcj1U36zu7EZinEN0Fl2PQSru4q
miEPdlhhCPagPr0AGgsSG9pctUUKnqTfooP1gIQ5UdU5Ic+A0I+MkQaWK26gzRJn0AjHacuhKoj6
CaJuEPy2H8gEufxPzXXhVcNSZFFL0tx5/OtOF7JXJzgIbcZ+RyOROkuuC29OMKvTDcNtg++Wlqun
UIu7+0iN0tf6wgoWfJ31eqRupnSRCifLySBrnRFx+mzqnMSsC6Bmc/yBd78Fj+MBd8a3LN7vkpq/
yUAV06iVfUgDZo0oNx+Tan8eYDe0hpbfe3TlDy4Qtxs53+dgnQGimSRJWyT1OJKzpmxPYoEGZ3W8
hezcE4llbX0cnij5ABokfRnd7sSu6RdMh8jNCiYzIqY6Vhd2EV7Kg7G49MkeStnTrL6tzazn559d
Bk2m+vaD4QRxJQxXZquDYesNKpLdjjlzKF3gNsbgRPkrG30oYxmwUg7pctI4/tPz6epQ8IYXu/us
mUif1+osr3xKvYljTJI66sR8GVTty05yqpLI5Pkjq/vZGZgWM2eAo+BXdZGbjL9ybu/UeHHat5Ob
yK5B263k5kKM0FGE1maQUsZuODWE7andubJkqYq9JhO2Snl3zIaR46SOdQSqkzg/ezsVLWMEgWvN
zGYJwEInS8m9vQAVFd1mpLfdIvwpHzY1ltrFkYvXyw+ZLj7me+3nfrQZ3ppd7ZEMZo/ba+RZPaCx
z+7R8eH0UQHvbloQbU9fkmWFjY8rX+BeNF/eenkXj8HzFCP2CH2HySEaySZE1lEsrB/t8Q4ihxgI
KBc5OwrwHR13nBJV4PBqeWSk9vmTp+wHb1MjPK1Db469WGrwbd9Zewzc793r8Ojj9tqEi/SxCIDY
2ufVb9iwu/IbfBxlnSRI2cSvPeRvDphvmt9eAdkCKOaEZvwEmgNpwS2K6J+rHbue2rXUp0m5vwyb
eEYKijVXlrvoKSjVCeL376hnbl8xHOv3uzqAYZsXAKfQG7zaYxJYEE5p5tZQ28Vh085ToDptGfNG
DfZXKUVTeZXGRbGunK2TcVIs6TsGsvJnrDrY/iy3RVszD/n60xkv6B+gVqfIXyTMxBPnuCRznoba
8hf1MMcmMEDcEqUuCwPKnip9WIZOaAFcSdKXQg1jaUWYByPrGhd8PljF+WF3E03kggfdeaYf8dee
j+u+m2PykcBsJSDmOyLC6lo6zzQS6Yma/HsRgpHz051a5iLdQVeGCQU9knyhuFgz/FlJeJVdo29F
HDfkRoLKW0RehQP5h1bn9TRGmC9YgtdRi/gkRSrdkF52OVnntz1pdrLHeYqU7v8+yf65YL13Q4bN
Sg64SopZ4GiyrxhB2Mz7n1Ih+veYVXSijcFMNhu3Zd5NkIEcPcQWMctlK9Gbv22q2I0DVtjcXdE/
eZeOrANSoA/Mfs7rH6IXS+f93qswmzG97ZQwmbj3vgKzVfWwFXxMj9yoIx8e/0R3BNMQLh9E3oEn
H0k+AeRO9GR00XOmKWuGNsH3Q8jb4FdXrgFOx8FrNqNwxjrilFHr1v2JcUmmV4a5ieIhYlhqiuNn
v6KwJ1oEixOs+dzW83+PSj4PSQwflnSvLt2eiHpquXz86OGuMhMGaTWOVbRoWhh05bK8rg42C4aK
S08ru5CZmiLyHmokvqD4YLuILDOZ/vqMjF9V3W16d9dnTUyoJed2W/NGYjq+y30yqeqTk+R7QSrg
CqoS4uzOqZcqTHb44XJI71YUCa0sqDcCiFYYMWEA4tkzWNK692lLpAFkTLBIOjdTodmWc4bn1Qei
zt7KQWlA96pWbDUTrAMx3+gF7A/bF+f/inkWTEhGbVKEn0tReV9I8/7zvlPlL/6rq6LxU6vbneZs
dxhcCWcM21x7nspU5jSeOf7AYoIkgwLWysHm1/4yeN0dnSS0pmYNc0C5NvinypwBVKBlStle0UII
o495tjl6EFxQNTDQRiFUvuCD0VRoa7jHHg8ulPdtxyYgfn2Hn76gt68YD+13399pRT3+pc/miHC+
IT5C/XHBEHm3k8cMEOjvh6MwiVcIt1dFXMEyUDwLjyW7fMCCQVC3tge1EUqwiVDtraVS7e9rQePm
NqUh7WvGqOOQwrwe51TqcAb6eWdig4D9YZfv9lXZcWHdww+eEo7qtkLLBfgjX8RhPVUrgCEcpsJ/
Kb5l0UGMetNXfEhZ1Mu69LW/yJv/eDfh7jHhdyve50QkUdmbgvqz7YMucYiD4ImuHnMUMvOg/q+J
2Ef6y+sXd6YRS0evugcTnLD7AUPnJXKqQPwAxQnrhrDgqYsP7BL7+Kb3lJxLiGcX3xM181ozH+IQ
TZCZeZq4Owqna0V6zaaxFSwSgteYXpN9x/iidPGZagoo+dT7ti6aIpBEPM37mbtbWr6/WZxPqIWE
z8Mv2JllOCu+UsYnlflULwAfToPu96j6jzZSL3YEh5TeKqgj2/AwkHHZ6Ch6Sk++v4R/cfq4/khY
YS/oh90bpRrDzQuzuL8+oqwl6r2SlksZNiMOtKM062C4hRG+S3O8IzKbHzUFDAMZk4Lk/w/tF1bJ
IiS4k8UbUlI4Ojmb4iUR6a42+8+DCd960zY5gk2o61ZiGzOGKb6+y1Q/rWYPmOgSXPklICV7GUyz
O6dQHfXdvAmhRRzp9aJz1FeAuPTJmRU3iVWXzWy4aFKPtXON9VG07RnEVPMlS/vCBPsfWOesTCVm
VbwCJaT9doHLcyeHPwtrjB8AKXFfd50EYnWYiy/ozQeK+MOyGn9R1zDtYQ4wifKjuMzohm3LXrbd
UB4a5nxDS3M2CodupRQ/JVWpXVNkNPoikYasjplYAf8l9HSvHdfpMtkx7Vux7Z/cGSeo3qpVPNny
D7vBrkXmq+FBtCn3GAVAQmV3eKrkWe7h5wQFZy2j6UuV/cNsnFsWE++r8GGno06VNn00AsoqBvIC
nCV6Szhfu+5jfaEBD/2mIc3xYOR5cvmgqzjHKff8MVJ7G4KRDeQeK8U6q+TrGLHjZKTbPOALjgnD
csaShr2pWv7/LK0Ccy5EpufuWvSr0Fcltdh9kjs4SK9xLIc/MwUd3+2ns7IlBasIm+snco9jfNH/
OnpCiaiTiy+vVFZpxPrlH9iIcr+6Emkj+z/aMtF6B6YaBl9KpCNLN1ZUfYT/MDXpiLc5sCG3ln4x
yye4hBFef26s/FpOPvNhccBtd5yF0o56Ue518BwvqDjC5CuyKUMl+1oRfK8/uRTo0TdAk5RsM2Df
EzWyMWO3E4nmd6C8IG1tf0kqDs/piYswCAYcADPtnKUSduf0m+DiRgPb+n8hSIRALdGDxj1JBwWh
2ZlFZOAezpnUYNpfv5TYiN5ECK9Ru4WwhWzt1WWtBdnURbH/cNtZeKiDGqftGoEFPxdE86kHl12M
0KsZ4mNbOrtez9qxwqapWae32WkSIpHAhUfvUxLtAqfF3VlPrqo9V/W/FTkQIDUo4lAkcUpgnxAu
4tJRz2v/RMWfgtuf/vemm1rWntyuzRydApaXV47D5WM8hwfY6g8nJuS+zlKLehsVFvVfvPKKrTiW
OH3O5V0WSnOJPmhTQyl7E4ebT2ulPTxRMXyjc3rbVykaEMPpUT0FZWI7pKuwU0RGAousx1oUPsg9
HFkSaQv0fSUEjhJ/a7f/q5bjq40JC5N09l09rfGXT4K0CX4zd14hdQISCnG+jBrcBtFSXxK/dj9J
rDooAcHoSaMDlbiw72q7dz/SI53ny9Ebso88X0xEiRYfEeuwKWI2kQpWKvvlDkuoWtK5TCpHWcon
VTXPyVqjdtIWTmrJNPqW6Fl4iuvc54+jQ4g2BwFt1LkQG7DAkA2xXHsC3hGs29o5Dt5dNRjFqLno
7yGlxlUXSCW2mvFrLl+BntjcjxSNaBrlZgFM2u7NXh44nJl2buZ7GS38N7/3DLb+ZGePOBNelRgv
x4GiH6ItzoSsP5Y0ldMH/IZWVQjuN2epIu+YoU7vUMPUJsbcJTkzXrGsQnSaxQy2YvP+Ox7hYyuO
8FHH46BNPqA9oXk6hcgMcplzACYsl9IQBFVXdbpNZG68zgbksG0Qy6Ui89BwUy+B0WbNwYronTNr
IHieWYSjUgs7aJAP+E/mIW1b+K6GpRMPs0B1Bc3SrA8GfhkHvv1vw60n50LDw+8AtJTwro8d4kqF
XFD1RfEAABXmQwevH1gm0DW6kWzkAcf6tmiuCl9t/cWhv7pRj7gSy6ftMDdD7zBJBF4Dyvs3Fu5W
m+Cpq2/sYDwg7i3v4rVVpC53ZS2IQ6gaOIBiFcI4BIClI8bYuzyZ6oUNePmJUgiSACLmuePpVViE
jrWpScbhzpQRig7bWHFHf19xyFSNDgC/lpLKTmPeF9t03huBFJVqSyA1NZuxG667g33F/G2iH2Kd
0byaQnh9KXgkvcHTPd/esOrR2KSWyfxGO2QwPmTxnNPWHuArPcLuNEgnzQXIATz+aLsQEWYZD/OY
jyvn5qTRh7CRcSZoCh7RhkXbhrWz1OjFIR1I90BxdYMN9wa721MW3gCrci4pLws6k0YWp7bj7dir
I9hY0QMyyGe/WOWakswQGyVWsSc1nBLRylkNJ7Aem0JY6xTZBqLg1hdPuV45HXmnWwnZltZCrCvf
+x69QHwuui3AcQR/OpVW6rm6QQ3UvxxkvGSfqSndNSsJ603sxAi+6a10x39orUnk54tBmgfc8Mm4
43FQGUYfvZXdeazfx2ilFraBYrFxXx8ODfphtYhoeuY7xapJ2ZsaO+A5u7Dsi8E9b//9eq6wKyC9
RqNOdFWBQeP1Z/IPZAnujHVtz9HbmnltkVJKqdKyFBI1nvh4hDzA5HYKAug2hwyyAPVJLlXtDFMW
B8Ob1zj61ohDLvSC+SacyHi6EckblrUN2EAEC9JyRksWl0te9gB8seK6EVxH20g1ZOyNDRJt7h1M
0pM1Af4G92IxDAf24gNxb+6POf7Q2eE6+GzX1CT02a31qCAxcKAVCfKAt6vtzR6BzZo+mRIVOuS5
zbZUFTbYBJCcEFlDmNuG0SWzzExDEmjfEBWTUUL2QlK7hWzrl4+yJn0JoUPxv0FTJnqZnYYLFTeM
f7npL5rg7FFLpkUREVnPoKO8hCTnfSQX6s6Ti7M0JoahVwTPDwgbsJZmRAt86bXMPk0D3/+81TFv
/pTrlOZTccjkTD0DrkflhA/HNhTNGRIFrAUyHhvn+4NwYVq3ixL2ffLHLvv6CmZyMGA/hrHdfJkz
E6iwBsEPEiBhtBO/LBcc4t6y6lvfgkNej7E69Xwra6bRHVSHV6A0xgoCcy0yh8MCbC9wUujx+1iL
bb/+zif3+kxwmVylyaz2PbsN1b2O29EqPINEM/pLTUErd88NT6FpfITElJfWHxAGdteyMUTgDPr8
r29DI4JW97v+YlC1STWdkQZZOsFTo5FzQ494zguFcLzHy6NrQi5p3JEdo6xVTAflM3E7O3xObZnU
GoyH+dHjQt0QdXDAm+lc4blTDjrlvMHXBhHs2iwdomCkVeXwk3Sw1R113AfEAjWbTUkzsCX7zeBY
kxDRZEQwE+3N7cFqAIuP4glYpnLsux/SpXj1BcAmQQl3juIZSLEk3F56lupyvtEW+IJyOI6U9JuH
FMdBjoLQ05Cc+z/8muAqAga5Q8N07+eD9HKcxumOp3vWG+rh9FXXcLNdDjHn2LxLg86N/4sZ8kOF
wRP3lAoN/XcFt8sZDByikbOEoMm0BU8qrmicK81PXEhMPIn/iJ9HUgXxy8xiE2xKFEDJjrLEt1oL
PDyTySpC3MBRq1FH3yKiDQIpCIoUQbk2+9rE2PSgCA6+5+BNPS4FiLWfacLOSiMEIXeYTFWaRJLS
pFVLaZotmLoIZlT39lQz+PehbVBbygepmLI8p7q7uMRmshxXOgvEMd+KEq+47kXG7Y4I3savyuKr
+m514VcDpO++x68zIXo2FWgUfpiDKxBTgazQOtYs/pz6MRLqvLCKXvrCus7vIgKYaLWm8g/PGPaO
eV+O0GzgULgOLCwesQVrp9smxWu9KJA/m9oyc1VZsRoQ79X0RrIVRgapWJ1CuRDtwcwl6FwKOHUp
S4mf9tZXNe+viezScCBG9NE68716UdYBlzx4jWkjqgaURyZpF/8l3WdtIwjkmX7x/y21bcYV4CMM
5mHDY/5p5V6MhKh4C2YpNCL9WK1Z+g2QPAb707y0W780/zQiI84hEtyUJ/EnHkCNuVCETDJYhsTf
jzlgf9fM7rYFp8jV+3uGXrTBsBqlC48RqiNJsQTRHDNMFkIMIJJGwGADN4yoD5/+rMRH3ZznwohD
tymCGn5bXN5I9Af0iY5qxOMkjG762Tzrxi5/YUJtv/9uhMljpgnAnB14n7PPHaEcY8c2q8QTcrXU
r+CKZd+6OhVNXE1ovi1GHPioIuByWLzI/xGJpZxrYZFL9X+KTDmqShU+sZm6xgyU5PeyXVIuOeeS
HdkITtxLvCKdBtG5OS4ugq4XmZ7pVWkMVF8Ur791GzaSD4+M05D+rFu7lAobCjr7ydR9Ds1A0BAk
UGAExckUu7xng90Wii1aEctBttYGY3fDjwVLqRQhxt0nTBrRd1SFHVa8EUNkaVu+9ZxBVn0x+65i
gp6i1P2MNggcsPUALUtYhpVpGYkYzbyVikIOcwQN0hw2LIA5K5H2jDQAjJ6LEfBVxlo8dCkigbft
6SYvVFcX9HXl3arhtQt9JjV6reB5Mn6h9wngJl9xKF2pro/2FAdlBw4KPONvyMV9NGg8Vyejyj49
uUPai5Ak2qy44/2vITC5O9FdpxyKiMqQXhcKJv9JlIN243ZtoVw/IZ/RshbB92AGqfmf4JUt9bQG
R7To29UZGpGidi5XGj7aM4aCVsd0hql92Bd4V6coOVpDxB4or9YVF2mF0ZbgX8Ba91Ow1TEH4OpE
Tz6VSuVqHVQCIFNtw1JtjsXeLxjjddR9sGGFwYJS158luPooGslq4EgIyAYPYN2Sjsa6LOL5+sYJ
azO6QrzXs6wfZKTUD67HHDpYIv5FovkZ854lg80M+9ZpeNUxiV9Ix1xOYdia3t6RUSlhxZQ9tiJC
1dw83Xw6dTG1llkuur9Azg5yhUk7jAJsEZkIlYcvDSritkBnuCg/i8KNDU/irsNalVrt59LcnV6X
vS7C25tkqA9JIBVs9G8Z3/tfalirt1I7a9mwr6BEMmuZWOP/S0YNfMpukcV6sHYwg1797capfW6B
nbzU2zBrtWNoaD3ACnSd6lBTHD+70CRyn0gHBLfqy3s+7/oFl80+U2J+S7wgmOzYHxXu3pfIOEBH
9zQW+06sbq5zWKNSNwGV8/wZsMarlGRj1sRAspLeyg3cN446rd0agbAEDNM6FX3RbtG6j2VSGoWR
XELFJrVqH+9H9VcnR2USriazZqBqNpZIk5DOhr8wJv92OwdM8MwVuRif4YwhCbYnGbpvmdfNkADH
fFUO2i/OLaq6rrfPE+yiCFgOf0l6VN0JZZPIWM+Z9UrLrmqRBoAi/R9W1j+4VHSyQIF6rUw8Qc10
BnDuxJ8dQWqTavlcZ2IQkFYAD3iErdt7Jn0YkYklG1VL9Gl0Fv9q8PaF50D0CKGzo2mzHYrms+N9
9R47uo1z8hxuKAhZrvYHEmJG/nbRuP1V9/NW3Moet3kdoTiJfRSltM024kN4LO1bHZnivZpQnR7s
N0HJ37CmiUDc2lqu4dcPhJHh1A3aWB8OcdB0gGebwG27DF2Lw6edPNjBD0bqmsJ32UKwSVcvPZZH
0FF/tzrddhbNAkVoA2t40StDWrkARrdZLN41M6tPHdkkEkdW2AFBi5cv1Hh36rafk4jIPwFJyw3o
UBgoZFaEbX+sVIOfH3NHa/jl6gZUwkshL7uY52LaZI+22MSfykqz7jnHQRtVaK7WumVO6Y/jS/HA
+Wj1tsdnw26t/J9fbmdfKGAFEQKnsSLeS/tlCGQQI7mqhzt5hB0fizGckRvlhmZDCgPn/UAHkMck
lX/aXIvLiPG8PWFETxAEZBnLTc0/sIoyIyNGqfWweymJBC6c5hd9o3PCG2+G1nOdvxQ4cANAb0sg
1UK5eMlND8FmRlZn9z79LyCIsvyFxldJpEDm3liT3CmYmw06O8j7r5wajrgdZJ4jpjxM3W0+uw6I
X+Mr6/6UcVPxe8MkxZsef+ftWhmMOT1/YVHX5Pu1nsA6OQjTPN0G5SYwYiHxLb7baIdk96mcIdSW
aL0qKdaqT8adniuZU/rIjBZrz7YH7DGTjabXNk1WuFostLPYobX49q6z/agZIWSlYxp8bOujWx+f
4vfib4UBb5qck5Mo5fZJqsDV40rob1dfhUumxXqpYIxWTMbbOamvOmXmL8lKD3/zOsbe2D4tCFk9
v/ZZ+gaWlrDKKGxQEKmfNMiJsOktkjtITxJyqbE5ONS2aHcJnBNBNr0BiMjY/8zI3A9eE9PnDQOJ
y5kr25PZBiu0x7hPa/FSvpb8IFPI74UsnVS12wj3cdNwzr2cHujIc2BWGkNPmOfQjnP4umy3Fial
ktBSAwzm4uqXCJ+g8k/4B9Wd5Jom8DPQxR6DalZI9KU44bjHH3OUNyaIbzjXPYrZlcx7KqmFSFhI
KG+y2MR22eW0XvGND3XvOtF/In5Ai9ffgIJvpeD2YQmioqnoLsQkbtrsBmlA7JKAXHtZRFtL9lEZ
4hjCdVgzewYpOEHlxxKLOFGoiKvx73THL2PPY9eFnvBHn2SlfGvEPC8RHgcwRijy4gdJ7YeBEHN1
igJS98OixeW3t4EpkCDLQYPYX6AZ1KRFYbZkDjiRSbz+4+r69LsFkgF17DBfXckZiSKVyecCdJjV
2n/ZQFaMSpGMgrTbCFML5ago5zI4dVlD+b8xKRO21WaXKq10keYnZqcR3DNAx0HE3GgQ32dA9ZN5
rnRpxFgxZy/NofZ4sRPMnIjq7kS+mA1PqUlHchIyLsWiZKLSAEUpDyoF22fKw/clvxL4ix7wAqSV
khR9pbiAZxglte1K6THPooIDuKMPVHh0fkVWu5mNFEEEl6S8q+j6ObxUlxDa2PskE+C+LFnN2QaD
jdmNdVzlTe6eh1dSaelFLIy4sAqLjMA7UZvE01d/RwdCaFifbgn369YoFkTK8/WDqkRWATht1DmP
JAUi628CUrpatkHr7TnlOTpO1HUfHKopHiKgeV/r2fgLruA6ec4sxImqTyU0LXEBotMcvGCeDgAs
uoIuPOTm7bv0m5vvqXXWBL8APHtTWcztjb9XAPKdrErVOnEE8pdWux2Y0Rm6P+4pBzZNcsrUWx1w
5h+5l4sKkrlRPKPKG7Ngz0x7flehMgObu/5x+RXU4VlsoCv193vAcRLxzh46CmqjtzGkBokoxVnu
UCYO+6EdDHrkfaOVzoLak27CxP5L3YEdrQX4uZ7q9VDE8mGAQJxydNEqa5XsbPiGntm1UR5qsP0M
oJCp0xhqsd4wY1lfX09714Evy3m6MRQyFCGN6JN+kZXvJe64TVqFcPZVhktKz1vxcJmcK3sUoUlJ
b37Iz8xiqvU8+Z5AohnZ1StvqCdqMKNS25MWKAzX751w1HHzqW5RajP39M8yhGkij3lz2Atv/Q/k
RI5Ndw++gsGES5kY9ALplxXY4bRSt0YhyAKr87F8KCuTTwTw3FGMOnwwYjRl3/0zDizVh+J2bcsB
QxvnE5gl9F12jMNWvKoS4c6jBp3n6SiMTxsEK9l/uCy7rAhRo3RQOZM7BWxdl4VYHhkJiT/il+Hz
yS4dgd4tpwARU7M9PoAY5SPUwY8Ei3tX5vWTmIIiEAEoB0/wQfbUYRBRvj6LWq9oB7GEJxRBvjTO
P0wS9xvh/e2cpsngSzfh54SRz6kgoelX4zoZdKkDs5oXWGwLodsXAGaZ+AT26ql+jlR2DiRd/vbC
80WDT2zmG3qutScwlX1Zhhtw3umAjTX6vcPt5TL9Jds8/cTMIbgyrVrZQSigjUxdjTiVU8Wcme2X
zLUpyxOtWgFRLmYCnnwgBKIhjw/wIYZkxr+FLDz2H8it9QTDtbAT0xNVCX04r0m06NA09EAuEFko
xwxEDdtNe+p+qax2FooUqQ/dstEF2glRVgk8AAOGmwM3ev1/8oxuhs8P0S4c9bUjhzl/xzTNgWkF
77uzdb+1W2fFjgtnkcbUfeOqKzWPx4/0KpfuS9jObNADyInJ65DelQziv7NwKgyEUCqpmazf0g27
H579NFJTJZ8hpaCTkxt9plzr7iK+t5tk69a1kaQuicJAtwqcFIJlPalC8SMA/OpNsB29RumY0Lc0
DJH9cPoN6fgEYRBIKEm35Eg6bK+1UwGqlL+LlRZ9wT6JfCDoR0s55wlmHjMJxE38JOhFVhF63vHo
Tf/xgRWLQkKcrbZbVEtz24RtyqYr8uupuTKEADWJmVYfysagf6JKPu8pjaq+uFvwuPH7w+zZQxdB
KmOf78g2gUCskwIKEMPpO3XGng4h1kvKTH0M8frI8fmOtDZ+9SuNgi5DZVXCfv3/ofcML2f+sMML
biaIJ65Jkr3kAaMKzfHM9l7AM5ylqRf6FH/QF8b7P0yGX+8p8ffN/Kg7yWLRvVvCtBqlP7PnlPnA
xut3nLEks1tlbJ9QJI/P0K+8EJU3kRZ/f/gUT1CGMftRlqlgmLtNsjnAedv16hsqu6SrO5Cvvufr
wjdFXmSwxQhCfARVvS6aZJIwVMSQZVDRFWpF6T7SXWg7V2KJr1JjLDbAuMO20qIgM6RKqPpaLe8f
fP92w0aOKUQ5/ywYWCCoqwwylLfHkHZrK81EsekpvYTUWpDTI7Y73fqvsnt5u5IqfCxm1m0kHW/O
Zu0leer/f4qtwkm/x1Vd3TEt6CvATz5NEMrKE+A/4d+2ePw8RMBQkrlyTZjy+NMo0XUMUmDnDFl5
wWV6C5f8dqUs15vg8SBI4TgO1oWTNukUdD+JpUTTzH80tXyyC/GgkhlQbFYyZtus+qe63ifvKTeE
Wvw6aAciqgP99eNbU/OICqd2tN2HVNYlMUpqAU7Oel3fEUgpQ+IrUdlB45MMAeexXC4jWr0XJP5l
I+yHUsju/js1LZwZr3rlKFG+D3oMSpVC+7R8zXAN2njMCacvWubz7ZLJ1NAt3WhiQZHU1uY1vujn
xkEfbPcYHYDb1fRl/Vuxxqkc12vuDdM1fHF6MMXmZPIx26nJJ/7he07rV75szw+2W1J1biJfgtCa
wH4YEjpt0BMWhZPGX6jG4p332/lGbp/YOMCqz5V/yjnHDTG0FUIlzACOYEebcLQxdw5hK4mO4S91
523rX3VK2Qgvg4MTy45BdH6fiG4bvBQnzzMJeuHhdb/zCmpa6Pi/fPn/uzFqqyDqT4kQrK/Tj/cw
l3+8i94SeEaZCBLkOiocL9U2lMO5WhHvhL5g0uSva0o3k9+deULbw9uZiRNpxmZWUmMxfwd76u2e
t6vpmvoiqF7hrbYfHGaK+uh61nhB2WpDJ4FsNAX5VlhGCxzWAT8oxcsR6dAj4vVAhc5xA4qAj6k+
V7QvHy5/Qox1EqzOexlgtxwxvOSBfzLVS1o5JNdSnZwQVRW52GsdTpRLcJZ0E5a13EuCY6+YrdQ7
a/MJGB7ZZWSbVo4w0iVKZSBcy4w+VFqghspeJEO1wPmvMpALSqiuVmLSYcKkkn3U8PX7OvovPdav
dfuJsndM3pmFFysilxoHF0U2+6yb2poV6Q/SBVcZwTXLRPQBUae9pOE5EBWOgbHZ/TFzuWROPRsY
lhs6V3Ol9CBouA2lBGoBee9h/J7JxlGkcp9kXEQgSRlu+6b7KO9lvxA+jdvklhpPkdNAFd/nTMht
ItHjTj2D66oIT/TSVupvWW+Gfp4U5llE6hNPtezilO2rLjq1FMICDn0KNuj2fPrEzmRAcS6xPHCV
iR4a8DCzmBtlZgXdqo6knrEcmf+BrUicqAQpQLnRI4pmT21vdUXoEf2xIyyT46FFEYF+sQI/UK3w
HN9OifbDu+j5xFuF/YLzGb6Gb0fr1v89HupJbghV1O6nx4IrmsX2vL0oIiwB8QQD8gQk9lRuoP8A
R0lTNqUVK1FGTztnkkmMQcAqxtf/qH3Z6Rijraw1GQwPV1xDjx3e3DD954Lx6fe4pxRvwLQZLOZO
CPYIKjfx3ngRmnev3+9dYErQ66QSLkUwdyhI9D9cCFDgxhzdNd8egM+0aSv2I1crdTfJ0mOzt0hw
1afr9Svop7b/RR6y6Bo25dVUQGXtsKPbKzWb8OPyFVAAghU3eogo4PnZWILr7MEO7qb8VKWxWZgF
5bie4x3rC71XmKuHmEOlX/Wa3eZLwehz70e8UeMbmmnrodGz46BedY2l9tf4HAoYzPUjV4oPIUSU
th8174tgMh7cMKZXRJzEcC5L36Ztnz61Mm7GFgQCM40rRf+7kWVfLPbxrw+M45vApoflzSWw7Pdr
UvaZ9VJRRwc8TR/3oR5Nh7r1azozcb+o3FL8smZQtBlzFtf8HcFKecDo6kOcspRvjOQq4pjKEdXq
8jQ2390JZvvXIVLtxbJ8whTR1/AztL6k7wZv/74+WHzJdUQ6uLHlziMHbbF8h5f2QWkFgANlbMrr
QyBxXvpCiecI7qeWex/pXjNc2CP3Bsz2Nl6gGrMbED7zzhZLCxeCTGgUibjUi7/bh5gMk6lR0b9K
17VNLZkEMtMCog6rJYD4Q11SC4+ZT+aKJ48vqYEN8jhirRGw+apIqsQWb3WyETK4z/Imx99ofeD8
hzaF5zXOcJvtR6MRvy7v1DJzHKZ+Mw3z0iNGQn8DiGY9TL5lTEBHRLcU3mrslkH7q6YRaH2vC2wI
Uv9tjIzIWM2tSrieIBVA+FJRcREykUzj8r+UFSbBojQDsqwsky13gZ1deaWaeCSKucH02bUOZoWW
Z0G2glURzD+8tJ6VTEo2BUT3D3U842lO0I6llXII4pqAO9G63r3vFmVCkBkjyB7QnYMfD44XT35i
HGG4E7Eji5ZItCSZ8dicpz4nxFYYMKkLwbqPJrzU5il04QOqz0rD7u9ZEu5J8Zlpj+gYFnlFZFrn
MBlm5+O84/iP8PMsdNKX9jxgBL1OkkeWB9eXeIZYJbBrHUDdz1qROEjraMc0Ovta4BwGtOaHCUnc
oE4lbTnWKJSNc7fLD+Gn4+3+GLr2N/EEtNE0+udmwKETuN1AYQiyTINDQmMPe3/Bug3IAvjELBqp
wCMdK07E8vNtubPXq5P5z99OwC2y0U2fZMkOkpO8oarSHY7juK2DANnfcOXXPv+2rs0lLywK41zw
id3i3X12ENa4mcgi/dZh2pR9ItRK/PQkOyduKvSLaXvQpy7OBWGhzLH9apZjbPVjc+8DOydrHh88
vfjpNl/EI+vgkR5q16crL9yiMcoEG2OTWuoJtGsK98ZJGYQ48DT7cBcPFN5XkKsIvuHaqjnDzbH2
Au9ohiej+CSCC08iJ5cc+nj8OfZM5+MSwTr2OK2tHB/Hfmbc1ZFLenzlIJfLZZREAIGORAm4KS9q
olQ1q5nWOSGOMFlxTJXiOaCALUtkUwj+NtojQDScgZPVy+pVo0cfH1hEHoYZI7E4g51+gzNguFtq
08lLCboO8P1PASCnvO8/G3nqVZEmZJiDAT9HGBwLTJZY4JRUGXxi6DXSEX+nFu0yBpAg0IpNqDbU
0TvWU3bTDlfw/hHiB8t7MSt8OQ4yA49P5AOl5taxpyPxPRSAloo4qsd+W5AZShQ9U+LLwVwtnDf8
iC5EMO1OrZBnaMugCSRwgy/oooC8t2V3aTSSFqzaHANVbTpqBSAjb/3AFdlewM2rEe3PtDrbMpvu
T33QoQAbvjLpK3bjT0lhLX/D3klvTIY8EVIvusLWXgdrvBCKcSYcgQUOiaMdHevz6Voex2490M+8
87CtCnEyEDOE07sSYuvhfhlE5K0zpJ38N9kzze7C+zDzvcJLUCCmVBbkBlZ8hef1T84MBUosf8l/
HM+6Vtg/mmDMqn3fOskz2Qibwv4iFBE3hzqgMuA4n2l3GtAUNHOdTQOD+a9Lkew/JdgU/KfEVz3Y
q3Lo88dQmGuW63bq/9OOE50F2oD/agnaNOP0IHP3JwQiWmoxrnAqOEOWRnh0paO+4pZTiShO2QW3
F3dR7CCsqbGfPGmcgTlOVyX9BNWHMgjBmMil4/8mFDSnRjOQ1AZiFFsKbHf0XUDWYfqdhlWo8BVv
f7eS/OOCDo36ueuhbKumhCCYSnK3ymAmfVuU81LdCTrp8XZS2VsPpiZ4psa5liSt8Rcpj7HfTcPp
EGsydvYb+MXvrwUnZrvlDXks6v4RBBeyukPLesb+7ieTrxKoqlzQOrNK+qnLiBRu7X7kInYAy8n9
GmXSPPpC2hCSMJ/nAKjOnGdGP12qpy+gZBtz10cnNvOCtR9KseKF6iXM/VV0TcsITqvJbWsXcJwJ
s6fDPWfLvXZVGd4CePap61ICzmBNFCkJPODte98EZAe0oEAm2btGEs04nFrblycHOH/iQYNaTf+4
pMCRelKBQsAhMguX6xkP8drtx0She3yK7Ebsd1kmPEuvXZIw3/l+FHXHIJj2Tx668iEg/9Ubng8Z
IZAWbzaI44iu7DIRdIgbXCzJClZcQ7Ajwk4IguWsFw2O00Ud8K8/trtfnxv8NVPGLPp+wgJpXzxp
TzR2T9WvlBmhoSOoTyFRz0AlpLirJSQg0Nwg4uhuLF/CYcwT+hUHG4uL6H2qDSyibd2SZRngypZw
FRwPJXBr4Drjrl3S2R7HMecriK6B1P/AqVOb6LRIKxw0aJMG7zJe9NHv9FHxGvPH4ZUpGY8scBMb
ti54OGRhcf30YMG0pIiZe3U1BzrZknCqXt45PEPhL2pmTcJiYjIYSOpaL7rlulvJX+K4504GGGZz
MSxYsS/XGfQLI7lZ1bhsu3uZzdbTTXYEVKjo7m4echl9ML9UNH4QcO+ZIRR4uuNvuUcWhoizSIhD
LcI/vfVmPXKMQvwVyR3Bj0h9dDxMAT2kumFUgDwUZV5bJSac9RIY7ZV7FZkDWPK42r5j0PXEm0Rx
sEtQSEcPo7OIJjKT8+1JVr+2cFbvYrxQjki2f/bNnA6gS45cuAgl1+NL+Af/NqCuWxC5ke+vLZ/4
w0069jlOA6enbvy+X4trwJZWilfpntbjYQe4upgMp+msEfFExS7+ZS8i9pIrGAX+x2k9lDK/JfSG
WoG4EeZHSfFSLTUc3tCXDJOxY8pUpChmAUqesBsUX6B7pHE+fDR28rjbqP0qf/GjhlSqQBt7QgZh
TqjGVxf97m/fqBf5m2VBAX9GD4h7qIegMvDuhu7BtvvgTcbUKHqGSiPicDhEZsicY48EMIzWIUDo
yzai6YKYVOuRr2NwC/sOjWBoPy3h5Ox1POtYeCgSfLiVnulquEyjaWjCWftIHafB0bYxzWxZMCWB
PwUDCmyd6b2IMD+miWO75+ksvi21GtsRIQeh7ey5i2zAjQ4dnDGG/1OB7wYVtiD2Nfz+wzY3fqb9
Nh7fGLZkpTgSjvF+N85CPe9wNti/wZjy/00dVhHWSPKc7MhNxloQ3vGnXneENOYymGWpAK8tXq1h
X8AF16yi4B8GDPvCivsGlwFP5fbbkK3TcYNlqvKHnI+piBXhblRQh7twXsIYY4qXuNE7de741M7L
CkcRftqiYYXOD7mHKjRjhPurg54WgonHxxV2AdwOcWXH/zQBGyVGdUxEDoRNVjHErKX2TYQaHr72
cuMCLmQsvQGQgKKFkiiwtvYVJZGBYjVAohEfer3S6cfQYFbTagKwJdScZ0rk/9QFVUXM1mAYEWPr
7CnRE7VcBI/XvXhE00KQz9lgkEOwekBRDcZMofmWX913Ia/HfNCA8JM8lFYCt0novCOvMxz/rfHv
pMaiFNfUZxziPx5ODI0jr0sxz/4X9IzvRbSh1Iup6g7HyhSi7wxlzcfuzPUOkoyiDn94e4JbQJot
R59jakULdWCFET8BwH8XMU5of3ptQzZiFksL3pHr0eKO9iKRTQgLbUvUePLUzMkd9YR4fS32xDRG
WcyQZ6WeEyu3cf1Xg7gTgQOmTWQraPquKMMT5iscn8OsNdNqcbnRowKa2/1SAhJt94lEp52ZKwCi
HaTRyLiawfalT7+Alcq94QseQ3NgQ4h2JW3KgMIeCL3hrTgE2YnC0dBakCrg+1mvTZYzzMCurOjR
c/G+o+yPE2YKGD+TWdzIA2YVxZ7DJQ9b+kgiFw9BUuVpu1/wpcu4JBTZlaAOFGfOGqicnn8GpYmx
obAS4uSVU+GVVqvgi5Gb5h2/l4Q7AaabHz/lXj+SWotnnN/d9ZP0KdDgKG2HH3T4rIDuoSihdoX8
3Gi2YHyOYGvUyP6RI76JuS+cdxzJRyylAJQnt6egV73ZOa7+CRCC0HHe9lT4hk+2PBkUAAdqF6Mv
ep4o3i0aLm2Nmf1pxP+KSvIPCUBeOwucWsmfzniLrU6lpqLyUhAJ/Hm+ikvm+XQqw2z0IZt0Y5o6
tBEIYWEjYBFnMOvt4ElqHNWHoh1VGheP42sHMSDUtXPV60elaCQulYilqk6gGGR/xqs9vAfYdMwI
hoSdoTlAO+0J2kMn40q3uOcrfG8fBf3b9r9TcatuD37gkml/a5kOx0XykIYTSM64AunHpx49sn/r
ZOCqrCS9K24NieHs8QPaWgKlAuz/CF4GvhLIS+xkRcA7orCnoZL55bN+uirOaj6k1NLvxy+3SbTM
UsSllU1TN6UwPHnkmBJnbawsXdI7m0CcO//jDsJju0Pn3wktGEGbRPMoNOzKD+LSAWVO8P6UM0J5
Vp/F1jxvMvq5FSynHFpMBx7Wxqm0jUkhHKMxVSR57K1x/SEqzSl3UAnVvtmFqZOJEB9LnExQPNHd
8m9RS12R4Y7+QnulnZ9INS+IKe5x90RKtsJcpJHwliWRH8PJRD02WqyajBmxxYuBvcPQXruPHzMK
3L9AEW3s4UzCTTGlIhujm6vF7fSgJEJBhsPVSHpWXpifRMfaCpPtR9IESDoOku0U31Ts9wVdgJkz
yS13P5OgBVNFktuQwDIPOCMs2aZ8HXKZ9fl1XAtucr4h6ZkrpY06xGBbGovVkCEsiNH8S3O6zhrr
9uNIggNflFuyJDpHOd1xAsaui680d7Zbqr94/P2XZ08O0lZH3tjErqGEVgn82zYSS5rnGBXOONG0
CzF0ZWG16HlWiArvJxJo4USfc9XuMwpPM+3CrZ/LX0CaOq4ezGATkphyi58LzbZ7fPz5q+5D4TyE
+A2KmARcM8X6fhQnIvW6aBgdUOtudfFVpAnzmTByPAQ+zcov+goKY3qEwlFVhGrrCypSuqYK332W
dTc+AT1hyDJQP1wJydkemZO87vW3tqG0yyt9Ycx2BpT46odnXseduXRCFhVmwj4cc4LL+Kg3eoge
wqda1vsfmDxLcnPxfL5IOxrXlg+nTbbsCekUR3C+dlvT41Kfc5FCMaGeVnz+7YPXgRZJ8LdB7Cgk
sAPtZisYGh8wPOFyWVkm0nvL/rOc1Mp4S8j5z4Dxo6zM7jZjjMfRIvSIAtTIGOS4djE1bmUIBOSF
BGT9b6BQPBugn27Yj0Bv5D8MD7fCYoE9N5kekI4uLY/exftaG7s9ZnS5JZ3Nl9pXjN2Cq68lXPUf
UTgCnF0fX1kpfSGCP2ugdiJUgsxmWjPyIyfTZ6ob8L0HkO3jQ3ZYOwTtBWELLyVsBFmlDfaU6lIv
NBIJ9PLhc1/KpZQlBobxPydBnx7F3y9aFD5A5Pu8tQsEhPqp8W9aYz+qdZll3CBOf7yv8Q+ANVi4
huy21/YzcKQQxDEWH0WbhcYTkSCVqQflw8J1a+JvU3g14tV9gPVKyJKdvajEFJ3qm+pK/UpcMCvu
d30U1TGm7OmyPKUdFIgC+ZUFohPipv7yWTJinDpVjwbT8lNfYzVEBPse6fFn4TkxA++c88aDgMoU
uT6PB2vS/ReQNKSqZ350ZogkTDq8Jlh6P1TaXw4+CJH1MgwmQjA1eA+Dm0q6dZXU41oyQ+s60iEQ
GQajFyTjx5k3P0zUGm9f/lGfbIqT0jzDr6dpoZp8IwRM4B4p+siBU3pOAMEPEwjzEwTc/1tTVfNe
bW73wBw3DQWYvyeTXblNDRA4nIh7OxMKJdytGT0Qgg/7vcKgqw7iwvL2iH6JK7LagBYypAs8g9xI
8x5cYBMfkSG4lgeHsSVVqa73rrhMWNqReHev3XuIVZjgxaBcvHvHQB7eY5+QlXSA/nbT7RQPRQRT
lHTy/wxC0kDi5UVS4CENSZMTjnug2WN87mgwe9ZzhgIYYJS/AMLcR3nxaVj1l3X7sWnf7YwB12vF
GkD3jko0onsmhKaG9L3NGtTDMQJGUH4E+xj2CHTBii4CNNvn2kuBMr0YkVjD0ZiV13cIt3pf7Sjd
QQg12LfE1+evJVmsAAlfk0zBi8Dvl9T4aJuK8gbK7qUSZ1LTLDPh8sRF8L9MHkS9PfuitQ3Spt/N
MW74HBh157JtjnCbRzoFWTXBQM+yW6xrRTJvl2rthMs0lZ44gFj9vT80B5NLb5ENMM8o36Gvhb6p
BEXnM8mj3k9NUbcX7SzLn3ujhwkM4rGbKydSRbkVRh4hZZwLCWQZmWaU01zKOW7L5XmCbrXwlkg4
3sCFuQTJ/I0z0zaHedlF2HIYPyJLT4Nf9ZqdzetdgCqHHoUo2g/lbBBci2RiT/DIYAcqltuNJKf+
uWHdhBjHp/HIyV5UlHFg8QiKK+/ejU5SmJReEC8Llj2GdEA9Rh5h+I+/6iBGu+aBQTSQH9lm1o4Z
2qt7rTQm0qOiE5rAEKBTz6H4pfiNzPeHjbSJlY6VZvHdxBZEkZ7WUr58IHqRLnAIyXISKeWwzNUu
vc4IEbcxf/6gOYvEuDQ4Qk4T7ASG4AQ4rRjlyrqb9UticmSEf6mSMERLgrx7yfLDOKXuHGyr6jeH
lO7e5W5a1T8WZww547rBTSqTouJ2q6N4PdjAOf9NMNB69BEToOnN5hUtK7DQtgb2eN/O3F9XRQP4
0OgQOd++fTbj0+jYB26obaESf+rNQx3eqrDhxTg7dtB7ATlJlv0Lx4dIPru2mmuaucOV+a0rlI75
jGLBu6oMW7Tgwep6J5ZJyqryKYoxYkHkhVbFq3sxS0hWMmLTgnlsI0lxQXVqjGEBNWGN06cuPCKX
n2bW0wCrVW+LAVb68K8Xv536drOhvgU4QsdqWhsdMsUTHV+h8DPbSb2pbtO9Q6lcbtzbWxR9x7cX
u8snfjoVzpi6/mVtcfBAswLMfgTBX3jxnCBw2iAoV5nw2qJuH6pMmE0dJc+weu4TiS7ARcHjZ9Rn
6J+O0PjrU4IoQR/oYelQFkzxfFjbrfDUu/O3x40OV/3P1EnntfSpxqCyhTbUwHQN7HWqem7tNukH
20kKHgXAee0/5nVMg04/Ey8pMlb2qjRBmMWBMK+bJKaw9JYV0X8Rcdqyz3Dyl7K4Soq3Buw27Tj2
1Wa81sfch4kppEifmyRv3pP0kDenFTOVFyZ16DNE6GV5OTZGLU4VqZ0dZw9K12tAUtn9P6yghenm
LeRKqTh9gPTjCdnoJHn8UeTHUNdzgCNESG+B7IE1TxxMZhRUzbrekMNB92xQmYlBy/HOsmQsimqk
AAyLA5DKq+vSsl4N+Yu6JBIejJCxKZjuSGaQlTogDl2n3V2W2UrvFRCK5w/0GV+af9Xe6nX1wM1O
FXqRjIfv3yXnV67rM1OC6SOaB6J7T3syHO2K1pF3Tj8deKUp022vWDiQz64MB5coPYWYWgwgl94f
/yH+lkiKpYbkMOHMf/miaYZBgW5/xeOGkbifk8YfcHbQzwm6+wQAkx009+YsNXAaxfkCDeXLq3Ij
BpijLBpEgbeLcRT6pNAwkw25bhpiHQx14/M1L97z5nOBISU4MrzynT7wUT31yIfIZRc+5/5/CCgc
UkuSRBJNbP4ifeA6UHtqx50kv78BnQtd/ixvG21lkH002oSlQh0EtSBrP4Z5v2wuqhwvu0q0AZk/
Ng7XYx7U2AoJ/IlxmMGt3ZtLJlUPzYmhLrJkpmbL3puRzSfQZO35OGwKP1NaPQMrrNZpas0iY2jq
gT0rTUopmiGxCNreKA3hrOu/0L7alze0XKxWFOY3WZiTNb5lTjV2Iv17zVTQPb5WHAemWqYZNDQa
SiBaSN6c71UjAYP7AToN/MHknitrRkqlTue2MiBR8OJSuBOWjqRbFtS614VK3aJ3Gdu0kOiaXTx3
pr52JKim9djWYgS4hen1l7twMr0FC00Zu2gQK5dhJFdkKMXxP1RBz19P9/urQkIQLGulRliOFSLn
63VeJ4wZAp9k46KJHcGeIakQ2CBV8D/X8WtL8INWcvEk7ShHQcB6JlqftoUqxaLqgFpdlVOlCM7J
XynL868CYo8RB9Gz93g4Hv78AyvYlFAEELRP/hY8l0QCxjq9fISpNsqfYhRQUrVEmZ5RpwnOPRHt
yPJIE5rWqJrxMcFi5uTGXYn/tWdDnM2yTD0MGrlxoMMfJ75SvudC5XrUb7GtxmO+pQjQEwmZP6rB
aP20BYJqkA1ywZoTKczIX9W7X2l3qBbM8sUeWSEiAgMtqFoVXXhbmRPXm2vp26VzbxKd9AvOGfI2
qSRVhjZh9qldJJEm5sq06WTJZFReWfnCI5UJN0IRxQV4SixOgrdV+bY58XqWVrs5LWhORCenVIov
GnMAj1N4Kx2Q2I1PRznOnJIeZTtLH55IC/HpS6SWdaFwbPNT5yMddsQByIThVJPHAq33NLN0fU7w
vTXWCRT81+G0lj/E7iQXUEphtQ+YpgAAVZGfeXh7ka5g0DOB9r99p+hqKuAjHbMawm65JyLp++ZL
xP6zq5IcVOrrJGvuzdfA+r1+NOwffuE36rCzwVKpsuMUfSEjltzBBRHBJvrlfmvNYfPl4arQRc4p
lmnxmNXg+tLGxjQETffnB/H2SnA7oSWB7Bx8u0vsQ+VbFNoK7LoE+Yu/KmisW5tbymsSoyDulRti
YqfWsnWf9k9cHpYoufOvcgj1tti4fOAqxaf2hdB6r0WOMVpW0zW2qtdw2KizYhPCmcskitbO77Ge
+kF+EiUjGZ8trjdYnI4fpk9piJU3M8tfcAuWC3o1TJji1s6rmgcMfWCR75pnk4TFra0dv2wlLrhB
GzeU6G3aiE/+aT/GmuOTCx3EzbaQ879e6IqUjF4mn+hsTYMRiQc7lBH8FRyamOCDLbHTvkSO9Bmj
FAmxpIDcQfymepUW7DYcCBhxp9CWcaRVw+ZIUsJ6v+TMg8VTAqIfUkg+Wk+hMkry959WNVtWdGk2
hwLfqN9+zrYp7R85s3A9Zaig2zLryE0zsxIX6mAiYg6JHYv7bqtgnHX9E2DalFHkBYKLNS5RaLUk
Ws0oRqp7VJFE03pGfhYvPWDB5d7A17diyM1+bjWcHdcXy283VNqB/sbq50dH32LBQoXQTdjH2e9Q
vk+UAN0IpJ8vxE2FvSEkawitDA4EwEh3y4wV8o6t21cIWsxgZ8bJQ40eTyMxxDueXyv5V+sWODCH
RAw5MQyTMpRY10zUrgoB7tum4UZ7V4nb3HMoGaPgvTYTeHHL5mwha1uY0vnt3yiVxXiUvx7bQmbh
v8PEMosHvXHvpKsHyuM5U0PNb61QOc7jKsK89ZOo0pKN3wtTByMzJ+GnbYI5KJapsRBVXXG/0a7j
XkWzW4IjJYPC71O4u4lqcWtFVBGBRavL3g70xZpU3l1umEjZns8gCEBCgObwAdLUHSfLTOrzV3ik
JyzkOZ79n75DqGYzyeyob8DO1Le2a6KWZUQp3KsPC1fXyT3DSUTg81wo0mqLqkq6moK7YVNItcpX
SOYw7EAkYKqcDuJNiuznSWZDagLW4KUrkfG4X81yMmQ6iiVmdPO7mSY6RXVzHJJciNP4AreiCzXm
B2BBI48o1U2Rv2YgMJwlql3QRl4tzmJL2UwNOYh/gn/k5Sm9/JoNGJ6VT60aBxQqs+6hFJSvKacI
p86s/7lBdU7rzZsVRsNEgFbSH3RCHppDSMzHynJsXELS7FjkkCbrTkTXnku8v6mGzXXePBBjXYT9
R3OWmMEsnpwoeYSnTDGc0iSUboTdz1rZkaMkQQDC2zbRwr9J47HtBjeVxgEql+L1ZwEsg5iFi48g
o3Aqzhezax0xkBkljBBbWqKe+dtx6+sUDnpl3b+lcO9yaB6wcrUxd9maE/KtDO/ZT6gq2aZKj7de
Su31ksC+BEAGb85p8aycxcGa14UwFFHgYVbiu9N2wx38Gzkkg94HevtQAYnC9iTH3fnbSopJ5lr/
Str7zkp0RC22vp1mbhnfADoEOUNNTctolB9ZP6JR9bwjzTC97Khw4Cr1mhZbgkKyU1hLbCsygEsK
iP0OD0TZYZDlVr+F9HhfVlmAxG/OPptTge8fn4hN+f0Rm0A9mE0zF7vafinpHReQi9Rv3lZSTOlY
cL7cdWN1sAL6MrSwOu6rOiwQ2tLrt5Lysr+RWpWB+GeZeTARoZ42Ep5REPjw07LCmspnjS30FMAy
o6tI5rxMsqyBDRGT07azc3P45HWkw/iAVnx7g59iTFFPJbSpAYfMvEmdttVzTjjIdgDXsWODXyD1
Nilxw2uSPXBSIcHvuSUWnx6Z+udZk5ifVqZ+x16VFqxXt4HMBBXaHNBOvMpgPLlOe4CW9G+OyJMt
nEmv9+lfsRVL9x7/DXQF7H5dKwyU7u/Pb44nLAEdpRhgFj7VKQp9xELM0Kck7MBdcwUdfCoLYnd2
iItHiXHdlhSffwkWIu2A0i/H7HT14PezuDxqIlhvw2Rr/+dDm9QhEkCULvI9M4UWvKDaAkVU1ZUW
mtnA2cDuCN0zt/3CKDCry5ANrTnlK35Nvg+KkN/Ca6O2isvoVN0uD7wl7nG1UoUBKlXlVweS6YVl
fhpd2TGDsiOPvMo8M630tZ10Cnh9Bq53ujP26o82nypMrJlssikcTAb2HU10OBYPAUFTu2fIhZpk
t0RcrrSg/Hov9CnavPdaCSss5uJ9cGU8HKPJ093o63veL9lba0DpSOVWoz0vVyp3+T7z/Dwa28su
keEwSdCTOqEK+hYLZ6SIjN7A+awZrl674iTY2lpSiPZT8MqNdGUg6z0Ez4y+Vych/uz9Kxezx42c
QWYJh8lvfhPcBrvgQlJ4EvWbw6+84bqC55M4NSdsjUsknMETO6RhQpEGIEzouNgzZDPaVW0E7CsV
mxiJ4IJHJpeY0PxQwnwEGyuc8uN+aJ5tYpfQDhunfeCjUwDvYXrDsEo9u/2vkmoD0qjuvFjxEqkR
edJ0dhcf/tvlNz0Mc5AOh/GEb5e+Y51NZVxTHhee2boFgmRwTimdnMZNVxfgubfrQKwGndtCREXA
ejsbdEYqcBCAgxic8Jk6sJWfDx7fp7OveVWlaQGQWZBLSyVvDF+CVNB9i0jPPQ9QYu2MNHTBX20o
RNgrRpYWDLofLVDrEhJPFA/Vdq6B9DfMrFXV813m8R5qv7NAKoFM6VQMT42G/Dl61N4b5DJB9WHq
wQhrbW/o4PUVBoBkbYn2ydO2jolJR36ODnysRcnmoPeHb5DlppgOsOHnQHQEPFzpK3uwsnD4H7rJ
9vriRInGw9dV4UBGR6OmRVyvwrhPnAzWm1BictjNsTeRpeTgZgZbjIt5IVVmRtqk54onwW0GtNkH
AmkWVAskdxEHJe1ju94rqtZad+Iml+AJWKzc8nfdDRo/dop1kgMl9u2jDluJ33Aj/K8bdo0OF7vv
mRuO4x7+8RLaIJaNwcJykPWzCFsxdtBzz5DZUYDYPt54tsvUzk4JSXW4mqUvJl0tecJkS6f6+sJ0
sMKFru/H2pu1kw3tqR77+L+qTAN/2C2YexE6wi6V1ZIWoe5qsKLgaKbqGVkor9CrtlHvHnT6vtZS
MQJlfzJ1VQ+w6/o/f8KEI8IIHLNokfp3xbx+YPmvFXqqqEGOgW45OzqezkCc6KRxrhmEG990naPf
VYDOkNfkPdLFMD5+ZeMOdt3syqmz/hFxHxV2INjSvQDJhK5TyEMZypVevDY61klIVdelujoAMKLY
WQ7VwiGzPXqCrhyTF7hYJgGpvWouf4M75COfncY41TJBo448iRVTuQziBbmYhSkOHzdS5M91LPkF
DefKadUP+XwnQ8v+qXuxTOQAR7plOQZsexSbjam5gvEkf1BYpFyCZ1qXLLaLiNG36RfORdZi/a9B
tihPQD2t1WXFyKfBp13pX9v6X5B7EDfub03FC0DEUSpCnWe06l3ZGa5u4k6iN1Sfe4sUwmA1kSGG
SaVPj5rQiqXBup2kMxg/KQwyZ1c3PimJgXPi87hcf37l96Wt7fq1RNI4pPw7gTowEvb1hxweRpye
gE2rTAwFmp7JtSM0mfvZeU+Ltzx3ElAdhxHpeCoc35ZtRUGXF47TUo/Zr+eBuaaaM6Z39eh7bDy8
SP9dXJROItBV1Yh+U6r69XLq9Md8Mus6mB7taCzzyVX2zaj3z34xqXBdAAjQo46z1qYXvTxGE1dP
CphOgUsHDITjCI5wfN87ccu9sercJmH8je5B6FRJmDATWps86Lon5XdTuGLxmb++BrbWr/yK3iFw
oi4een3PRuNd8y+NH4vjYZU5qghivXmTdM/Fzpu2dx5lQWm1k8mLpttEU/JUYFPliW141oxt8FLj
L5eRc8SWyvScid3CjCn+n1GEhPZV4TTGxNlPXcC9+i2uC2S4ZzFwTIWMmw/IxfcXv0cwFgq+jFA+
Jblh4unax5E4Mu507Zh2XhXNIk0recm7T8Ejr5/BAkgsAqcDJ5g2KGwZmJFzvQj4z4WdWj+f+SDH
FSKCmOorDRdxsXT7yCxmnZAsdl/LYLlgXTRmcHjzTs1ZUvi6bZ0Ut7qdU+07GFoMxDSEpBU0nt90
5+dPCgNPMc2DROd8hjgRYx5DAsQyvHlXbenznhoOzxK/W7iggSzJpazdZGgTURLkJd/W4YxVMUwY
Trd5rOfPghqP8nlQWUpDeCHgqiTPlFLkwrMQ+U3TIVTkwRBYQQye6Oje91i+ym6VHPfCJKwpcu/K
ji4YI6BvM+ktMWBjK64KkR4Gk21TBV+zauK09OHtwYwO1iKaHByswtw+Z67f4o998t3zpPbY0L3d
UJVr801vB5v1Xle9QMnt+q2WOM/uRgUhJLuyX7qOvrMCt5QOUJfC5xOkbkaoRFoxv/KOBwd6TZkX
HgxsPDEDGONTh1dgANhB/sbSLuOCnD31fWWxOXJXaxG6Ft3uija8BYeGaM83YcDXo1ignlnS5mk5
F0iKp6TiOEyjwUIX2V1Ne1O1OaH02IgncuQH00NSJhZVpsmTBL5OEJmfj9YbwCsWJyAwXf2Y3Iac
hBhf1jj20dhpY6lh7BOnEECsEEHCXdKbvhfrscDULs/vLGqpeEq1WtOlF1KffcpNwlPtTxYoKrzU
Jmt2P/MylJ5MALDgO7Z+wgrXXG4d58YgkmS13oeearX13XFvkRsWwkL8KKfzHBU8JwY07aiy6FHY
uQlLcOW6YonLjPjbwiZiDaILVe0cH+v5rFjCNcY6g8sRroPJuVURJIue3ZNOTYIzFErBTPspvCN0
gYkd1jlNp+lO+3qFM9BDMG7pyA8b9CxRkCvF1SccilnbS+v/ogGTLkM/vU+NhmA35l7QfjBQb5XZ
xEouIRh44NYj6NQiZah/Pa83qVwLbv2dPopJYA849glKdTEVxWb+7hcx/prQEzBE0rXGdM/qV0oF
lxLtq/7csIJFbN0185Q8mIqTIys7pglsEwHoKlwbG0ft0L5/4dGCr54bcMCbD0v9VICsURgejK8g
jRwgZI6DmwYo7Rlvunn8SBcDPK3VjKV408Bgf2rUFKdS3gl2viJnmHJ1djBniER1LcUUDHUPrBQX
4pmi0d5iml4ZfN1tEXB6u46zXbHle3D3EtAdK6rR3/LusmancfuUMzMvQ9Auii40IQQZNQIXeTbf
JLYLWi4z+7jDWcZKFa+8GAS+0JPLLy3D2VIZzc2n2K5fhfOqUmweh5aNVQF/2b3F0VSHBRSZuUV9
jkcF1k3cg9w7tVn4Wd2h+Ytb7AwX5HWS1YIPktjXWFUPBtAhXpL5eSfk8l/Y/hkSsuHjwo7wtwXy
4ZA6LRiA14ULdTA6/TE1WkN5EIyBzhqHHAAvztZbYF93FG+H7eTLfujv5pebVZrIi5EFkems0sYG
XEX24zbLQEut/m5bc0A3l4NN9Qmp9LS3XOzIzdZD0DswAkDLgM9rnivThIiKBiHqblZhzi4GdSzG
PMasrUGgavWaLh5ZjR53VHi6atBsk1pNahZ+jKAlflr7Rdd9kj0H8pkzMXdc8kO3urhyjLTXRxnV
IDsLndQF9wJrMIr8KD/BBGrYqF0rYmkR8zLGE4sCY/ediZlNHDwHqC4sL9juB5UuSHGWe1jNJ/KB
tDQBlR0wY5qLfJAPG51i1zkqOXkq0jIl/OLqcwoDkaWAtmhEOw3vFv0ffGTfb6Olue/Qpaxm1yJd
qb80DWQgfNY+ZYbCbRKhMaF3SEph7FamPncDjVUY9X2UIuEqEwou3syRsKYMK43k0OrbtrJ4YK6W
XMe4QG1OKKYHxGnsbxi1N9BMXmsXPUc9WpUnbvL5PGrcRqlR6We12VwBonGQRWpeJsvC5IHqkxKK
6QBtxM6rWi9YXp0PJBgnrDDaMYl5jRcZV7ubFXnER1yGbGPDqLnWnUuIFVz2T9km099GvDHZ+Z3o
T1a5APCyQUNBOn9O9Gx2px9WMyUs11KKxooxApaNJY3nfc4J59zUYbxr0lcfbuXsMonsO6xZDp5w
cRxSBWCdjYHR1r9c9Bx+oyhIC0IGR+KEHNblOtRAimge2/BbpfEWuAlMaxOc+iOXrUuCx0Zm933Q
+CRASL09crC+Obyki4UOUnP2qu1owJvgfitosrHnclnzBWSBkhx5sqLDMZBPODb65AiJwI14b65l
VSRm9GdPyZz1LSRt5obptm+XGvHNJHw4QRaAX92j0qqcFcpSPI+Y6L+W7fS2y4IdkA5LNn6xZxNS
GW+Iw+6TN4F3jHD/rhkmbllDYcPwSzO7oIfUyCMK9x/rNSgshFWRY5MDAz5WhZU503+xy1xHaWUa
uNiiKdXqvQ5AB6xpNTK4LtrVlYt1c55/0wvYvdR7MaOn+LrLNgeg/DUomh9ZWS0/3GAknFHof9qX
A4fpzkjnVf4Q6DQgGd6paGww1KU8MACxNEJyajIqkoCQVc2eTzmIAUsxEALMPC527Uig8uE30iH4
5Au+S5BFOaOOdM3XvySGZG67J05DjE9xuNlSImOHn27YTzi9yXtEGLrwL3FqB6tcRGlyCCBJUXKy
woTUVdyfHqdl5l3Tnygpp81v7kVVgS0ZhGSvUOu8hGMu4583Cg/R5kDSe97FnaRTnXABttUlD+TW
14zpVOPR61m4nRg8uDtGiEXTXFRUw8sU+TfkMrOmC9mbs7mE87aYQm6M9ZK3YbILllZ2ljnNMa7u
vUNujMCIxzZQX7cH7NeARjUg4leoY6s7OD23yRZrYNeKP8M1pvrFvRWSN3cxMsu7WG4y35XhCqW0
e4K6QZy9NTDzxH08oAgMzzr+1/qI4CoVz+Jm8XIou8AepDskM0zQ2wtgxQWMpBGFGPeOYgTxG6Bk
InjcjwqqSq82JHESXvauTOnK6ZMq1mlTvhvWTIHthoB4Z3afQ7ltEW8b1EolZLJiMrffVNcG1+Ye
JGKgpd8CLiRZSw0CMTtYRkghNcL++vYLm+C6c8BPXMsLkHAiKf/Cel4L1xe7BEoQQiuw8aYVVdjM
lSroHX1SDnt9iMqW892n/6mdUezLcwUtG0MDRQTdsMbXeAUyP7ZsTqESHNt8BVD2OAXhog0u6uKc
Ks/sqMKixlrxdmTc34mxRD5xWk0jH2lG/YduGVxmRUuhGecYWSoVuPj5wWO2MNVwrr2TXZixkHb8
kHYsbGV4dYdRLKzcEncmgJ8HfWIP8IulJ0Pi/ZS2wpx9TOKjVklZzlNTfpukXyCtlWTJwLjVYbTk
HNpYFdG37ODa6Wcbz052MLxvE5LGWe9UCEANqy9LUWYjg/aSobmdpzjfP22f2gPD1zRSVfJ+ouRx
NOqwAbIssS/1X867rSsbj9bmuzSTVtdlhoEZ7ZzFDsS3IqJQjKLjaLPnDisoyZNAGw416Wsi7fKa
m+e4Kzhy7XEfYZ5Pg1zBoYJESuQZ78kuNOY2D9+mzN1Ln/6e7MxDCTvz769sXqYJZPWOncFn2X4m
521SMsOw0QcAElnya9ufJQdwXqSIJy2NPydZckxm8vO+Bkpn2QNgUz1c/3znAEsz3H8NI01ei67Q
gDtEIdbgmn487re6aRFng2u35vyAoumr+6fI41DLEMJjuI2SSQmzAgbnvDl5hZJulZ0o6W224SPG
enhfSC1KGki7D0WSUgT8dE8XZyMRWv1AGXwQEPGqNMMlfT1+/EmNsyeRX/hleJll2RwAzLSj0HXA
qhLRe0BDjUyHTqK3vwkcJAVXQkV1UmQ5APHv9/3PtgQmomnRImb5NoQLICMeNccydyTyZdOylZw2
IWkX4YTINSD3yisBq/2tdvZ1lOiTNds6Qx4IKMq+2i2wLGkoXPph+oa4EHTzJ3yt/6Vigonl9Boe
Ka4d+l1xWCmiIVi8k/8qDVKOilkHBvHqN38nTRSp87ec+6AiRlQMHRf9IfSaNKYnDhQGBJgEnbhu
3zp/6h/J/jlv2gCVaCSDj8ebwwD53lpgzYd1MvtN9NtJmWf4B+IciczQh+ETX8Sw2wKY19b2fMnR
Iuk/gqGaA1lVWi8UBiH3/hxgWBenm7BlP50G+aw+ds4te8hrzwx5TeoxnrCnATtaCw4iRnUFi1Ui
6gOMoCmZJ5pyQsRSNqNFBSlovLiPZhLjZoQ1RM3ONeoN1PMGK7tuy+KqzYrl2Ty6JjJjGlv6SqUW
RrUCHqhxChyKF30hNQy/5oXU0GbMtVvl9O5kwnTZ5EUu/qA3uqoM31V38Mz6+/6fHEn/0HuBjRay
qkh2e5rLwk5/vtr9c5apVwayhtMsHe4C7lsqHoBSJq2Akhv7wrx9aiC2c8vuY6fqKPcOoJhCEMC0
qA+mFyO+AdRyOxscDorHCLNYRBOG941Fzy5bsjVWHjPIlttNQelWQHEOW2PKL0XZPusyjZenoH8H
1jtHCzwhjei+msVz7r7xNW+xEfSOrQwnPNePLoo81RN+MdcVORflChG2zfePsDoecktvWb/+3AO9
NxlfFDBp3OdkpvJQhw/q6CARExEgXbhNezVXIntL3yZyW026hTpV/3QHzJWYfOEDWBs/pN6qOZ3C
Dp+exisO0ODNjGP7DChGTuBFTE0hML/gYT43wOW/NEUmp8kPEHhOCHa7Juesyr1buQ1kv845IEID
Vxs4+pzt4AFqgoTudxPNbgrRplDt2/8COX0ZjOEfSNrQGISdKQFfoYHiP7UV+psiboF35NTw0XDT
nsYBEYpPGatIs4KCm+huUTQXldOvq5EUB3oUAMHHQn/ImtZs0lBMHfhGX1863gjKJcR6+WeKELMl
dFMiclU7nUpPKnd0q/Xf0oSNjE3gTyYhCx7OjxrEU0MBn8vxnB4kAQ8sABOflgvaqhdd2WP7cJsA
1fO/+G4JjOtXxdNyZKw0cRAWIQ/klPycQB/6RSTITaxL0jYh6llOGnrKShKoGcj6ACRUCgTW9zTU
fkCLhh1Gmg4DvWpi0w1ZU5Nj6y33iB28sE+CIMpONGtu51CGIfDuB5yDLneDLezMRzwWaRKTEmCW
z28QVBYMj3fHKd/SnxUmxU+C5uNVCAExZKoST0bKOC20mxC+ZsZOkjSoRyX6bjlDGUoeJDwvidF7
GVrwM73iyhiqrXB4Nui6PYfxaLlX9zwcoVL/inlY6JwPS8RbZ7wZHzhby8R9PBIYGDD5rLDtJOBy
jJ/vrIlBA1OH1o61JoI/l8LZPwcpidvpWbtTdMq3D4E1rY3y7IcafSWC/mQ4Bh9HTA6B8LY71X+V
oB1u/D8B0jVwYx+wtLkR4rawqu3spwD22L9Wt5CQUw51IeEbZJeXZwdFLrUiijDm0BBsIX9BYISF
ygNNjF1J2uTko2vKNEb8Dy+W5oQ2coq7FJzN39N17SUTYZJmRzAlTzeGtL23Tqp3BCKhPuOgzHfn
1TjREJUGRXFm6ebf23lalmXt/fReQUQsJNrI6TGkHFJleZGrKlDa0SM45qkH+fEOioZ5jHHVfUmC
SHE6tcBcD8lqHP/RBzqkl9itpgjaKz1Nkvcy67afquFw0fqlOqIK2ITNgiR1PPRcxNDGWtER3vFS
/bjtD+DQXv/sf7docc7mIoU3GDu4LmTMHN9V+ibcQ39kfarSSUhf9inAX172urXLJqeshmG0IPkV
eGS8epSs6SrNnhcpLstq0l8VnsJxZIytzNKX+egNn+jOvrvlxQhmZTCM722+jsyJR6mCT4kmbi7w
Fsrd1IbhiLAQ+RJo8JF/X2CJiTAtn0hGvDNew5dw4YVweG/IsqDVDJsLQQH2jqFLjVpSJR3wC+1P
2EOMQewn5fy1jijg2MoVpg5LjuMJx/aV86xeSJsyujJ8O+5wP1gtxtD5kuMq1MLyLaazSkioGbhy
J5290Z+O8Ls67cMLxGzZN709t84VJq7QAzFwAioGeLWE1enn9h7e1LoDvECwO+4omVD4isiDIZuX
IXnCOgN3eNIjucS+tbLZRMXgivYuI7z9ELMsLNvk3ZujsgVz4HDQzxTRb1IWPFbYuUE5pRR5Awhv
DJcaVec5c7BZxS1Hnp11vB++2PsTBRcA1F6MlikBr3h9J6UFG7OLNPPlY7m1RMxFhenhaI88ssxg
X4z+Hyglp0TaQISUqAn6FyRqmU8nT4Z0g33rf2NjmDiHJuFKYOo6PG01brTzVsVgIbwCM1COEemT
MDbVPPy3H/dbX37BgcYZyUd5T7chru5U62CkWsrb9PEzilUmg+mqxyCVmX3ruKJ1AXpg7F9/xcsO
vQDPxWF7s1T8gNIyc2hF16DBN701UTg6Z2sDkjVKn62uSzUA6FK7W7kq66BUfJoufzZDPRGHg1TH
HNdBOtFjX/thE4/q7bju3us9b8WPR7gJGIjYIsvq5KHR9JcprnhPLmN3i0wwcv/lP1iyTdDhOHyf
Otvf+5rH26tT+NlBb/QUDj4FmZF6Om99zrD07EDaJHze6d2x8HBvgoeXj/vFoDaYWOBKQRxmDto4
ZkAhjsXQGBsOqT0wnLfdZSVJ0BZhf02n8+F2C/zjATg5ahJtkgWf0G8yJVkGNpIgeeRgf6J690aF
LHEDKsKu1qBDYQ1oMrxie9zvgJnpxr5Lbr1ETH7swnmGTcuYPEr0jpF1daHuY5U71YJQRkN1dGSN
XGZe5G/00n5CKMmpmuGkuqWoSolJBfdYX1593QIGtyUbHUW+OM2BymtuUNZZwkcTGgVzgvcaJWIo
aV82uEYJ1QjXrj90ZNDNl9KdmrtCeuVvHb6mw85sYz3CLMh30MrU3w3sf3ronO2C7jGtzH6Ek32K
csnVNopeG44yWwp+57VmFiIAOpRWEHfr9rptVG+TeiQoFpGhsgP5JJTa8BwqzUn3yk4P7+3ZDbpT
7nls6G2i18lgPewye12rTiXXOC+l9R0+mUZiclKntvgeO/7hd/x514bcSBXj1bRP9g/fuzE9JBD4
5sJwdVIvRzmvlCKnyalUGWoSmPaecXD61vQrfBFcWbfZPQcDOHvVIdTBrKdoPXrlBNoLnyTHHtSp
V316QI4ohb405MmozVYtH0NCxSkYo8AgFkjQJ/czGEWoH9H4/Cl5Lo0j4+HU1CT3odFjatHJkzXv
KyqKMzPT3+lw+88XfSMot44TbqAceyieLlrIV2DYEFcxwf8O7jO4tIcFeD7es/0om3xzIa4px2rf
5ZeNylF+bqM3kIs8RFe/eSR+HaTcIiunFa9SjeEAmKpShrGlbkN0K2++/i8Nibgp0JDT7geJquSv
xBsFD6Ot7luTe1p3CmjXGMI2oBNIGCd/ghWmkN6U0bVw18f43r5cVwHoxcMuTJhdnZLuFc3j9BPR
rkzdwmCaWtCBq+CYTvu3msnQxwbEEbvfDirmrJzNbmNYhUass3KJkid9d26IOHhJmwf0dG+wh6Ne
KCcAD5sjpWfM4TSo7VOvQiKlFIFAQ3exPph67J0spPxAP2Z+CZRxO+JC7JaAuYiU7QWz8Lzs88Gg
8SXAfgVtJua1Ymc0IxFwCunqCXBhllAWWtO3HjDDUl95pzil+QQ+gqpRq1deWjWc2HSXUMGkWDUt
CdsjJJEPWCtYVHzDO5sgj2eTfz/7CPxt10So4OzyXVwXp3y930hrhnoJ1sVbiEOhSGpt/CGuOupG
Zc19HJ5DVgjZ528tx9waqUeO117Srst41rHufUe8atGiSXyDlUo4KIv7iXrZdi76aFirtgRjGtyQ
YDV8hLYX/mqBHxzmIT4SZCr6ozbQ7BRNpyMHmqEUu5huW8izvrR3jIt4G3VtFwCpfiOQIevpe/85
vPjOytYobON4AJ08OhgnIZ2DULvy405MNy5tcYoK78h9XvcfsUdSggO7V5BVaog6jBGLMTOT+yHZ
A/fBzyLBoAs9HH4l0HrpIiDjBUuRp/ED2mAvHR83c1IghMSTouAV8t2gciNa7eHAPnasLDk6Znm3
+bIPNvvnpWGnqk4SCdGL84NKoD7MW9x7HhqpOfmQeDpzBkWRbIgLKhhycMPnjubtea/dd4gi9tvO
SRL6kvpsBgiiOugBwsa0aDZ7mOCnp3E/YRPXkmKI/rTlGR26f9S2eEhRRgtW1m6LoPLNoAB5+tHX
WgzsiWwLiKsG5Yn99a1IHW6rJhnvnhgqgTvsFEak2wh5JNtk625lNMds+tfyqEpzMcKNwfc4H6jm
MSoK3j70rctt6CRQmtGmq5+0P4dt2cS0BlsMdsOcRFy3G2OV6vfV/yOZQKK+Q6QH5Xqaxy13zf/g
AYTXuHSxzJotCohyqaOWvuAWKWymXZA1tRaWdXQhWLR9aLyOgW9AExQFuet+WCGEkfltvuQQ8QZe
yfBG/cxjO+bmfcR3GQVmfDrJnmW8A9cGqnhQh9CfaywJkxlYkN6+SF2NCwAFGTh/rBBi9GqJT2Bq
zBhStSqd3hL9m2DprDqqoJnFqyPUfflSdtLBri8yOks1NA7XFp/mf0CGeePIcAu+cRyvvcUc12MV
vB8TJfh9akvqpN2KwZdPFz0umCyDtddF1aOKCoOsOK0HulnVKIU0s81O+e8NQDO/rpETyzoZA0qc
XD31/jg1+HBPwx7sqkI48Yf3quCc6F643AP26/TpLGmwnabu/ZAJj7sCT+mJ32BcV84cU2ZBqzwV
TgPZtdIA8OfomMa2hwZyrCI+Mcqf9xhnww0A3qncepheTFqGLwXb43qfJBaRRes1nyyWAXJi9Sn+
9QQYlRs6YjfHixOUpgj4CBVDt81Gbh1WnMajXB1ZvcZGud1gE3UyTK6470KRKXkllhA4/L5EuRD0
UhG6OccJjEbSA9SZCOyyQc3GlaafmpNIOjw45w8dA0tLHfSn1elt8VwIeVEqBsFoDjzLRA9vpkVn
2s/RXJBPom3xLXAbSlz5kpgJdYoOJz8LZNpqlEymS4wR2rGLO3OgzgCR8cKlnEaHnBgmkiKE/Cxc
iYHTNM2C3byel6HpSNgzWoJ0q0ZpcNRE7QSPbLw6twTSeG9cefoZ2y6jprUjO0sxk08wnngdBxeu
Z1+QTDtPhH82OtaUI/Xiajn9GMDxE51a/kXRENttoapAHNtxGhJncKhMuI4t+LZnXaAbgMBTxo3i
o7UzRatS+r/oICiaLjJemy+IItreQzitcUzCuwwd3A4AWBSrBWNhPyV9BGqN/eVPjWkIqBA6iFI8
KBW6PnG/+8ms/zigwWRa4Q+zcA4P0aC9VxHiNQUragYkWS6D9vVXVBqzlF+Q5FtpRZ0R363yafzh
MCykFJ5P7ZtQZGetfJIE0BGvquLpJIiWGv4sEYZNXH0MT+8np0VznNwmy4agdG2FGdBI5cG0babB
+csezJPgABovKdLLTzDLWy/qpNxDwa+KGwrxXlFbwOw6AVp0ZPw8zfOGZDVYijIN2SnDiZPAms4u
+YKf9qBCRg1ICMYtfOTSC/heUXiI8Hc22vqSGtF/89z0F2nXguWYb7ygV0+Qb13msqUkoa4HvIzI
31ZlhnQn0rAd4aDBaKRng6Dq5wO0Rcl4uR6ANgYx0Ukvg0HxdcPuCjOOk+NlJTvzvupBMNA00dOm
Vrm7f47NIazdNQp0KEBh+yCd+0dwsV2qVJoKSMyCjGKzp4ywgWp8tQsOCrDlAU6dK+ywfDvi0Hxd
aBFNtPHco1/Qlr1A/RYOv6Ho/AweOdR3+Tr6e+APmblB395qupoxYiUMLYy97FAkiZPewHZOEjat
jASM4wyO6eOqT9+QTuZQ+nd1qZg5Nq/YbalVLNmhQGbN7TMeIo6DpQv1uP6XAVdPz3qsN+g1sjoa
ZqxpW8AEXiwKFwRk5ZkB31wDg1XLeW2s7T8HK2KvQN5IyQgXsPsvSa6iItl5+FtE663G/6nhsbNx
Y3NaQ/s+UYG/z0IfiFoQ//tlblFGOSr5FCkoPEEz9BHdlu2osnUbT9bam2sJf1N+z2PHk2tc+m0j
66Q1iLZiG2qTwUtg/xGhf4pcVhC+jZdZCANAwJI+rfeRcoz2QFvsMY0XEixG4hwSn5zvF81VY+xv
GSUDDhiQrPFwIQx4Y1v7dCTaCKCzB/S7fAyBo+AXxPWy9nxfP8MV+QqjzAWcqamGdaedL1yx8iO3
c2wU6VcKnZe6QIll0zIiNN1Fp4lvymG3BiRDBOqpfX7lRHS/mrG92qOj9QwHXKht/IqsKMnRN7zD
QESNuatnrIgBYtpEOxqhpEwNvwX5e3E298Sr846gyTvSmVXAFaUW9kVx22Yw++tntvsv8doqzQ94
Tl/vtqnxwv6EGCMg7AsQPh8AbemAwPM5CVVqxY4/K+kQbDYqRZZCFlGq1RlHEGIfVY44I2T07nts
vFfpX8Wzaf1bQ033uUc+1qkZl0vO1hSeXADB8PwxPfqrgtR1NBhnaqqpwrFf/qNBFuWUjiZW9TF/
fNFlujy17Yae92gGmYv/GmvrtoEVDweBQRDiQJFFBKE4OunpyQ4IS7RYLJhFiE1iPtgaiYLlibsA
gVL2rcF8Axf7qN17jjfszED5QIhD91Xvtxv+r4UMGemToj32CHSHXF5l2ILajh5v3knNCG2za5sR
zgDi51OsvIAI7cC/RFeOL6k7lTBBMtpgGy2kdfziPyJDLYn03DhJkY5JUPhAi8j4qk14skoE7JPd
/KorjIWqGXGGfbfUZs/VjCUHNG0dvWdh5Ux923hNrrrFr9b4UprCE9ecHkH/XjQ4c3dw4NCuTLeu
9maQJ7ndWyxJQQTcHIoXlzK2RVYPrtr11Yyw4vpT3OUXMgkOYMrl38omFWbFN20VFAktpWLXmYfq
irFy7jRMJx7XL+53Ahabl4EnCr9UXWF4QRT4GrecDnqrVIOcR2naOTzwWwLMgAhvoJjiZVjLsB7e
HStjp6bmG7TRvBuHPVJhNN8CVDCLd6QC1oH/sHFjPuVi0imHipRfIb1jlaHoAZCeol5mtOHqAmeS
g68IiwHqhNgKmPk9+xoBattE06LZyzrbDm6ryZuUZ76TXFlI8fwNcR43XB/S4gvjImdopQds4WUv
9bt4WNXJFg21sBVVhytvE/rpOv4Q6sYbGlt3eGFcLrjSFgbz/168UYltIYLAlVrTSdCVEDW839LG
nNdA25i8e6ATkFOcPFzulDGwhUTj/A8RPaDrtzGPCiuI4OxHK9u4ziMyQLzMHPvhCJPrzjvCE7a5
gVGs9VWo9Gl56XoMcTGZz/QSbORYfAzwgd4SiG9DcqIcVkB5hifl5g7Yn6RRTSb/0uOHeNy1r4O8
skI09HvnA1x7sACHDyHPsb+UmTi6v2rh6lbi/2OLwjWwEcLr54HwxftHy86DSy3DLWwrCMZC0Qfs
yYkel/iXfHMu3Y0emc5fHmDrUsRlZ+fft48x12cNT7m9/CiuWHUEl5ozi0rl/8uPrH7qJcUl/2Yh
mrINmE4U6X34shdJAdUVODjivgZYg/A8vrhY+0yuCtNRmkwlPN7ZOE0O5YwubbX7MIf13gHwXQ+c
WHi2lDAtY9r7bNwQxR9dBgY8KEnRgwlx2u7m1pMYj9lmSmtBS9nsPKVGC6okiuCj5DiSVD63mLAZ
vQWrBSWJ/orJ+OEhwmS6fpIYsUQe6eeFLBlh6jJxboICiLfEZVAU1kDj9rarNZRlpjA6wpFfSM4B
oxkRfuqPHogQQU/Ashgp5v9aS3k5vWsdq/vKgDzN916lj1jPtEcVc+Ux4W8LVg0nch71F/RQF1ha
aUUlCANzK7ln1cFnMPpaWD8EDMgRJoWz56f/msz+IZxX++gRcU68VlDBpnfJxDBbwFzE6dk+D2fl
ey6D5ZTyEJ72zEuGj5wWq8zCvLc579+7UARzm8xr/Cu56o2q7n5HiomUczbHeIosV/bmI270BP6E
51VOS4tKvuyPmEItBj52mbeI9PaaPvow6iunSmfWaHFwOCnqAHZe+lxfQIXRh3rO4y1h8jAzxsbQ
uwQjGfEkmwPQIqvB7FJ34B0M0rLyol9i4c8SCtAe+ojF5G05LtoIp383oZbKk1dWd6pUIBPeJMbs
zJfKLBHsWRg5UvQl69ULf+QfWTRep1tcHvV4J+SD4Cz37KPluE7FBXQuE1Mtaa8QP1pME4IU1Y3U
gfOjugaW84BJaJVau1/V7sv+NO6y/CQ1VffYTuLdPOnIeo1mpozpIo6J4TB/WQQiG4n0qpPeOaJP
c1SIauh+wUQ7k3jSDOJp1l5KIj257C++I5PN5Hak1uzgRBm+4nw4+l7Ic5e4lMeaR73kPMJoZnAc
txAqY4JS9TWYLqxUMlzyH9N2c0H9f31eyUyThJNE6ndEoZzJE0ta1uxgXCDLHYpoGY9PY8tYGQxR
dWNVjiCgeU74/olwh4WmxvYo+QONViFbf+wimzACr0NHnEk6hOBq530HcMYh+VkPvwdPHr8DH4FV
tObBFbjhZnivqpb+v4n62/sfDsFj1OB1hIRT6ulZhY7ad+WHW6ipFXbTratA3J7t62jpbboLprcP
zNJeSACbtsxW/zai3YHd0nO/GhYogRrm3fmB5AaYNgwzrC5UmBWt/bNizfn2xWlKdGEQsOCTprGd
trYur3/IqBKHYHXxLM+Lw5Rb9hIpjVt5NXpy03Bz2aQHslfdTHoJkSjv3MK1KaXYPVKLZqMZIr58
/kQsHEj2NB4M3FW0r6DBYFqu+vdROAolTxrBx/VMiPqOk65oqhyj9niiRgKa1G2HGMdz2S8wl00h
R7rtzYqfSTaJ9166Ht4Z/ddgQeh44MyM7MeukUOcPMAqIDIuWr7Ny7IPA9vrJcSsN8py4/nFAH+Y
Njf6wE2gFOlO4YJqNUaXugKP+NqnBrLPM1VtLwpGGs6enmuDTR5GJkkZC3ZcqWQkFEp1+CRqRr1L
vrnW2Etnr96+Rwxse+OT+PJhmG6ev2R/WhebIOibTH4uPoV11477Wm8ayvxPA5kQ/13IfIrPjngc
SxiJ/RCfz53/expZIWXswkQuqgE0joN1aVqZI1WwGFIxPjtEjbwYYcySPk411Ya9nAY8LqWvTjnR
Nac5zl/nua1Zw/tYEnmMCNK9yUvtENYTR0MzWJHq5wGD3Zpl9928I2ytkU16SBEqaJI8nP39RPuC
rmUJml81oysEvHFSt4l4U/PLAnl7qvewgAI4wHgTGM2Y+UDcHY8G+tx3/0mqyyhnAudu56el2QTV
EWr9YoMtts/mxBkaLWAOwW3OYIrQypx9qaRff28y+P+apALumVIJBa7GQnSfIBHRI9509N9Q/2LM
xAGYWWvZVpajaeg/k0Mc2YLDZdQoWBSvPoh/Vex7/Bv6Y4tQ/7Pu5lGpQz29HrsRcdAzrsvSRvPk
jWNItX66vdhGHAx7yqbXUlBo3ngmB4FjkG0E0eN+iXGsBsihvXq2jgtbzhBaDyeREdqUeYKT8gUy
uvhg89W0eAoM/z4GVPOy/9idTJ1PCshLx5t8+GolZElErs0Oi/M8gPcgHMMZICcsfzExfSgbRCcV
yZLZ6YaNIPGmzUsJDh+/oWY/y17Ail+t/ZNIvtsKPsk/pUGw3k+w03+9C7WgJe2iGzyOAuiVx0SJ
POYpvkazcgaSvOhETtoDUM7iyQHgJvDdvzvrqlDLmv96cBXqD2+kJ2A0UEttxoLaPOFUDA32FzqW
wJKfL54/CpWt3llFVeslNtHX0Mf4o2DAAwuDJXmSDj0MjXrzEWSG2vQEggYd4gdkoMLF1d7VDb3t
kL5U0c0BJJ8baGNOr2dG9jO1U/iR6qTmvOyEzL2hPrYaNrtmzN+IVMjBdEQN5yRxHfn5BLXt8Jbc
3hi0Tn19ugPNd8DIZii/Kh/0cYpdKtEHCCBIiDRsZJHlXTVwBPFAs6nRmjxgvVpqeTB3RCXy1Kev
KMMPlPoIEVOMfzD/DNzamco/P9jkPp2pHYBsAiWBM+PdgJca73xFIa1OXNH6skZC94nA38whHYeq
OhjmzA9IEs4/1rsDGko7Ozg5zaXuwUNl5q+2N0eVG0ovZPYARDhP4C7pu7Dt8Zx1x1xjvEqkU+Y3
RkWJImgPWiSg6w7foci7OelPTwOWdRk6OkSp1tDT0J9dBpLwfSnqvydR+42cunDjV+BeUzJxmIhU
S1cqSGDERCurAnwPILaChq7T2bnBzyFTKfCjkdDT7K/uTdE0AP1gOtNrN2uQuk05X/O2KrNyc/4x
45PVwQ5G3N+MowQi2CYb7OA0B137ydKgKnrKCBxdCs86lvtPvITZPUsNVMJySsy/4UHQHyrBzxXd
gQpbX+kZ4WpE8uf6pINIjnsahyGkdnHgFsDgCuiXgWd2s6wzBhqDRtuaS0am4DzOdVe02Md/enmd
HO6CYrc4XAU4O7s/BYmpyOVMj8Iq69UeKCIX3ao4A45xgelqlyqx5pLqiLOB3hIsBCxAeAzwebAJ
OTm0XOQI2JkXaRF/KrJknmBz6b/5GP/wlHXh/MqFiv9Wn66q88n3Hve3NIamg60d6YfDcO9J4/Mw
SH99i92dYbARxYPS1mUB7CLf4tt0VrWwqHoSb4lbu9TLhmiiNDmgUq9W8Qe3K+2yNJGIWgWRycR6
F1Z6+i/q4li7nYV10OgYyEkAnnpMtDbvC7pTsgFdL+vIxAuNevQpD/t0j7ZgWLipB/t/A+vGtiqy
ICnyPTadN2FHlrUuthEs2hYj5ZaogFDqWdfnAhaWhWXfDmH9Wed14mjsnLqyCa59REVGanGmZgz+
6OJTIFnSFNh0cCNq+xK/Ja9rKBF5J1ZjYVzDI0Jr4uCMVMNT4RIyKzgU3Z4xfyIHjJnrikt4LXfL
zVvSOs0ByFZJMfrfQnbP8tpBp5o0OHIjsboQIt+GVaPbO30mbQCP0EIuZ1TRqu+xqBhpfUciD044
vpkJJ95L7F5MWMoQOr1PhW0oZ4fuTabgbcgeXRuKggwrJf4pFCL0DAEElQxp1EQMtkv0ikefil8J
Y79UyP1nYEvlFR5r9TLIlUl1UsxtZZjwxC/fZAclMjdTy8CMLz2KAWRhmv/FnqB8U8IgWjK8VvJ6
B0MYm1oh5gZ04GRMAgEomYKCe7S+R56aua1ruGv+LCfIOAOuHPAXQN7A60bGs3z6XTn7txIe+3R4
Oq5MTSJGgqv47IvJjizv2+b78fNqEvY6DkyBIBTNIV4jlOujZsdKwPkuSl2dwITc3b5Pr6el0szY
MGxRH8ApdmiSC9Mt1E6UgKnf2En4g7Hi3/z6wAr8ULe6BNdEVKvsRrSsTi1x4CQQTpnm08JHjan9
GueApcyGhzIFT53vgwcVWL941FSgJ1qmXtAazqAH9+XiuKwQZhO6U64V3+2boXRvXhAEEiK/x8Cc
RIsS1wE6tcsVdINuVusZxHVuX9KuPyjCjsTb9JLD9YbkRyhZRQf3MSdJqg68KZ5lRVhDi/yMmEjm
bH3tkYQ6PTt34s9vaJ4wmc7smzCTGsj9X8IpNZt9ZvpU/CSEoVeBg8KREmyCpr9YOODPR+ZlfP+C
FMHxP0YlevBW6WAZZXDcNj8RkOzA3xPt9VKgu6/0XQKOa8FaMY2EWnxasLqqWEfY+9N/KnNc7QnU
9L2C4EJwgU1AMgx7ojFYXMm5thkptqMq0m+4dlR9LAF7PGNGqLhVq70o5DMqXYrupfVMd7sGR2ir
R/waoxzucUykEhDglr58e0dGTW3TIaoCBfSkMsFNdLvldMifO+h9J7exkdJH3JFrAFHIoXT6usP5
JDfYfI0aCyvGy4unTqxk8O0LQzAagMg48jktk5/LQlf9HYJXY/sVYMz6pBG9zLE+TsWX/DgKi+yC
ueLjJJQBJCQ6+wFGIpmtMwvaQpG7s85cQSIaEZSsARJc8zFd7Ki6aIQMe2+uhScUs6CTSJsWZkmU
NKqCoQawdVIGQrb6XYm/hygscM0VNCxnzpOQtywUdtaoKtg0lZVB/bU9MCjXvW/K1igxZpb0PRq+
0UP7ulTGP10iYsDEgMdW+pEy3NR+huQjDmJQojhwnSocAZSH8rMdoRQFO/oDHp30BvTMaTX7mZ7t
l4ce9XyxLLpEUl21GbbPsk0OJkVZZHZ3bKR1KMAO9EiovOOSUBMJaH/ChPdMJAzlNuksJSBO7FDK
kC08V7A+O5PQm3a8AN14oo6dHjm6WSjGrcUWNx5Kn1R7pLA3ofHBGOcuYUmCX7Opbj1HvUGmNoHu
twV60zFAMoBTCIi5AX5Y2nL05uUEPYzVL2hsAaD2DGOSS43MgfuySPunLan7XqQx7cZM/NgZbPj8
LCwcnQt2Uf7kaMN0H6+7BuE+bzzWqDNyxp5hFOg5nnao8fTHVKkRI3X1eeYAwP7PsRwvd/OxUcCM
COOWBXJAwqkPc3c41OfzRm/lqohxUpDUzC6ZnJ1B5TTaNQk0aUTd4OZ4d+4QGqgbTLHtKNyswF78
cheuyi2s/Z22RuLiuAhX0mi9q0p1qJej7KVksqog6OZn+xzvEyi74gF9PnOBXyjuq79hfiMOVtnD
J63zUh7qr+KXg00vwoKohzgr0/+s3h3i/+1X+z/bZVuWYKnfMRoXKrInnvvOjbDiLaKzldAAWO3S
2FfsNqBIEZOqhpfVly5DltZnfN2wY0OwgC3mRANw5eUPqwPjuf6vq7+7wmMib5EBUvW0+PcyFE7g
LYB7GSN+3e1fjpUpA+6BMiNkl9X7VPaW97AmVOJLp+MSZUXK3aH/GtY+gc98XVw5VtSiarLOYHEA
tb7C2D6L5I9B+VECITEYfbBF9prK2lTmAtObQxFPjxwRFCh/RO1XsBpBS2nJyHhLjXg4p/8HO9bG
1IU9qCGGsY/+y7RfGiuKKd2A1Fnw7WJ+VB6t36au0UejrRFQIm84PLtDVz08TLqNt1gMXq3HDL36
x24bF1V1L0TNniVRJcGkrP6X8J4UvfCMVcNqxjtm5NKThVQtiAINx9ydY4z4+OZp+/lDMZq2K7Aq
AtMaU+C53gC6nIXWGXo7p6bczwLKfaOg/kqN+jjxCkWUmxzqPYHDynoatj5LCwIHIFiy+7QUWbtn
/81sfNE+jME2puSI2X99MXZtJdF8oXrVCEl1hZdeWO4QPzLN7Sv+vwpQ2pUH5A7upHNB7ng4mAml
rkJFuqoDur+TY/9IGv/vlx1vYgag6x2jqRZUI6bEYSuDsPWhkJES8UZE/gMp6eRr7mPJgflQI5Qm
+QPQDoyapYBCcxoHDuLmMh1m9a67Lj8ypHEAL5ffmWHdLoaO5cbeh1zdTaNswB6M64UGtD49J/0t
h5Z9rZ550LjhdrpvY/7B2XwBWqD5Qt41Sjh1aKfMOc5Tc13GSpvt8cJuhVu/HCJ553nmeClGSlnX
huvv51f8HaXSfHYHIYalBi3dY3uvP18It7+U6nxqETDcZp0tDejBQDh2c8W5AoI8RZEbw4AX9V58
p93tZgtoT9OZcmgl4C4W6F7O/c/g2FzID6mWYPTih06dAxMr889lz4ojBuWG3npOxW5HRQv26+L4
fvo8LoxwU6EEwMA7PNXBLCkaGpwcvXr/tsGkkWYuTV0jCQt/KbPffqlcPxGltOzOkQCCQqt5icj8
38VIv/pcxxe08PT31iF2qeGhQsS+2OUc8zBj9xmV+sZ3BSlPXAeSGRHDZF/nodhbSFJUj/ZKIHpo
+OGMJ1p7wRmXHtut/k3Ydogq8oFLY6csJfyZk4JcaDVvz4HizvANPZOMBV7rGqTZeBWZ9BFDeIcp
ntWIpXg5RDKYxGdNcccmf7qr6rwo4hMt6/M9IPvNhZMJ/UY+ptNmzmCgXC++btwmPjXf7MHLFLtA
CQoL9wz/0xxEq2exjh7YCRpFABC9etN9+Xv6ZczOp0d3ReH5xrz0hYrQhHzJhpSrsH8FEuyjRfrX
GtFQb6X9xu8iervTcWyoFXKGBiIwmIFXAF1/4rKrdYSYOoVzJmW80ZTHT9y4mFaOM0YIJADVNDU1
wrZeIxBM6xXBaRzseOjMqoHXQC2A04GPWI+Z+crSKWd4a51JOn+vIkcCBW6PI3laJp7qFljrPQkz
2ZsRJBaCAV5ZXTZbQHJtPpabP0B631av4ye1omnOZxj9eRQhdOXygPkC9GUQ6VazFS2LNxfvlW8j
7uoCHPGYCEK7FMqOD7oVRyGl0vTldFQ5hzhLfizsOKMPdWwVMfn17mf/QkBThA70yCFfVkYsoHPf
vDRKDM6QT/a0yXoM3zche8O4FIoS/sj/e5iDA4qrLjyH+3yAqpIyUBLViGI1OSbFikMOBwn3o6nY
BmNfh4wF/GyIB2zJAXwShI0Q/twgiMTNpA/IsIaIvXNbl/s2L6RYDREgdsBFfL+FmOYmzgOyXu5E
kQ17Zq59egZxzXgfda40t6E02Oas1SwJ4/o/7XILjd25A7ZKxWWDXFkoQUknlFPCYfQddoKfTlJJ
omPM16uchVhazX91rTUb+jNqOhS7i5UOZbCVeSq3CnQY96K6Ga2+lnIr2mMH1SyaJZQVbF3pyOx7
hD6vEPaijDaxi4QGdnXitrz7kEmZfE4zcqKKk/3znPPyrUGRYJjLOSJ1BuordjGTYN/55tUGqRZw
7bk8cChM16Ilup3QHpFMW48D9TSnfavZjbDar+AkxpKElzjFOpX/NbPB2BGMSE9ZSON03ZtQo6uc
bHi6AgGa+KH311QI3D+EhewSF7Mh7CWxWRp8CPleKrrUrkCCPl1mMxClQwBHnh3oj5REXZF8PeZw
JYpLypPl8qpCLZk72nXFmOCXcJYltECrfjEZ82P6T3miAdtpKmYX0PiqGGrDg6sfm9yEU2//p684
9STeBux0k8QrWO8JK1uINgW9ZPaA8uuSOYBYa1IiUyBwfy00R1RiswZgyIXu7V1r/fnZIgqg55LZ
vILdvrjTQ249J3ic5DnER1O0lYd4J//h0PZCMdWUjAp9HbMHCn7dRunBzI4C6UqRutFnGtJWof4B
WAWY75bFSdB8SK0jY0B36HsUAcUPdzBIhTNewxLQ08kmT/k9LIlSBzgWYIcnD5YilEgenxvT6+kO
bShx5cgbiLwLdPmb57ON1kLdMRYShsES/oCSHjRyFvDw00uxG30H1npEMRRzgWw3wvAsMSLfInPY
vkqFK/yZij0Z/eQqEsNfjXYt36JRKQ+J0Z1/Y0nZrdPkVyRd98owKHUhbokPHrMBnSeYziG4dGeE
vtKrBIdUqqlyYHhHi0Z3X+1Npk3grc/5Jn4cUc0ttE1kEa04TkOFlXUyPJtq+YomFYR4BDZ9lmOG
ADnotnDlwLv1RVbfKkmtLD832r37cFVmsey73q3vopCf5a9nwT3mHX7mlpWXHDrYKZlvw9O81p2Q
mKqRYnvWAU4UBpCF6LANFvrmwu4MNBEhuAwWJs2qBPj1wCnlYqJ56u+hYeTQlVkRbdngyBNIVGPP
ZCE55VTn5Zqf2XXmwBmsAd2OjxLbwFUWuM9Zjio5mDg7QEE9RaYfOLSP0H4Tr0OqONVB1o2n5GIL
bU1IYiBu8CGP/w6a33vDcwoj2p+FJICHaxx+VMePJNgH8PQvLnjDagJ10m6SDLvHiJaNlJJvET+E
5UR3e+aO3Muo+OQ/kmL+5/sHThkxRkTShn5+rpW8b0b5KDrrwXyNtt3TUAcedDhjxj63N9QoWAfy
BV0m2I8ZZ8liUfkWhaZFja3ygVxgOnpxvMLi7kWviwqKuwWEU8W75s50lNYdgvvVLYJ/VEl8QeN8
Mx8Gs/pMWSTplXsrD2eMerKbQW3mAyfYkxXcacpjO56asKGerni52WIBOtQ2igX2M/Rw5tDax21E
fkmd9+K2axr1PDqhzyididBrQvbsJlUzwIk4Yxc5WPP3RJmGKXRhNsW5AfoeXwrvC5gy7dVGYl8T
djhS2ODF+aW2XwRyhKxLdEr48cu4a9/uOeRg9RM5DvG7lhOI5gQz/2m8itlOgZz7ey5d7FVkq+DQ
zK0BwVtERm4oHY/A/Th5dk+ONrzOog5zn/Fqpm9f4wxfU23xvUxC8r3ZSxqpyY4mrsMQZ/i8oVco
kTooyoLoAg0SV3dfIAILWxnAe3CGZeAnfE+Kun3KHUTXfIduoxzzPNQGhq9IZ2clGu3VMngGXYJa
lpE4deFcAXB3t4131LPrLJDIwDZy2nYyt8G83HmijaNacJ5aPIpbu6iALvxaA/6hEccK7p/znVpK
SebY1dM7ptWLSWD/18wTMgLmyI2tN/+wntDAEHLo/hek2GrVfFRnuoPZ4O4AFXpqXWLXGdFYcZY3
mQ8Q4rNmy3FY8qSXTHRxS3bt6LNj9uUwaoPaxhBv31WKmPMtsF7SYBAeMGaK0snvgknNqWE0EB+q
kW4hRxyotAFbeiiJo2rhUfhRddIN/twjC6J2Z9Td4T5ej9tiUW15+D7jbf8mv1G0FNQNRXX57bk2
wLlTWkiW3aWJ8Kacu99bMeYE8nL7hVJoFgUlt4jut5Lb9GvzzbUNNyP+zJOzRc5tWwuvyJKMQOX5
DCPWMU80nXg9zm7nGKB/csz0YeJ6x1sg9ZoSuRwTo8zRd4yn9jahLABz3n6Ts6Onugh0LIll8g7e
mS9I8J9wtK6bi+dUuUoANwVXS1bU3igTpycXP3wWiZ3NYrR1q5Xlpuw7b3+ZtJ3UAQr5iHp4Fo/3
wPUSn4OlaYb3fXXAk81YsMh22cfWxIz2j/g8ZOTUqg/vzpFb8OLn8TE4+V7l6Cmeh0dkVI7Y9wVJ
SROPfRI/2ScjV8HTRmBa9IZZOCSfO2YrX6Xc6LIoAWkBl/YhG5KBmZTtN5OTWXyhelcwvhBv7o0X
AmXZDDfmbdVZB+39uHrYng4xvBreyrjnRgdphSkx+xzE4oBUbh8RXgZeFtf47u/ScOZcTCeZiaRF
wJd6Ia763FzO5Uj7Z5KFjRspuamuOT5Hmeb46EoEw4pBChghEKcTEFq6gRM7HyTcdZLBvuaKz6ay
2AMIy5MXXTKXn75BA5cUxvZCKaihXurxaxMA83WK6UvjrQdlVq+CbsWyz2yXdNO9RnkRtN9z6T9X
k27qm20Fd8ZGUuAS4vvHPt6VcxuOLRzOL8S9hnWNmSTUKaKalvLTBMIjjDkvzwt0YFa6DL69hEbV
9ogHuRTCpEKDT8Hhnie2FhJO1Rrjp0C5ZR2Aw0HrjVd1LIY+EcPN09txC/zBreOSTo6qMQJc6/hB
xVABhu57hlrQFjLCTNHrrKvG2FKlyxK+WC8MH8Z9uvy8c43dKD7QpyNiHk+rUa2g+5qdGaRsM8JQ
VYqhD9VEIa75BjIulyQikkh/KfNGaI2BGGcKDyWE5zCSMTIWZZIPccPGm6mSjsNUQ82Gj/M4H2wL
PtIm/ESNalOpELrTNa4AAotTKRGtbvoDJFlimP/QRV7TVclwcoO7Udmjwb7MboZ/yYgQniH2J4Is
ckblC5dMGJtV939tfZflRvFpn/mkDp02cBT0IJa4V5PkCKfYNHkwCiYqsWtoLHZponmYTpBvMJ1r
7spStNSx+mhPpKBCWo2Ej5f9Jr45nKal/wqnyR16J9BjKoI0l3z40QBYrGR2k+FzN6xuOVzpxTH1
QjQkyaCEkH5E1tDdoozLB1aT238GiimhtksuGoRtAX7aZwXpyLv6PKMKNW/arRZRY3pJD1m2jAlC
m5w4ZwjuU7QO/JgbHj2RP6YDP8XUAD84HHWt67yg+QZLAHLZS/1+FyEGjCrwrt0lRCf9SWda+P/t
8OOoTKsCUJZw+6bBNTF98giyy2NaFauA1Dp29nMBXP4X54fHgfLWtx+bf7FC0e//nsVkwSS1hCPY
WKYfFG3vXrpPLYU0V3myF3lICBsc5VKiP7c3MRzO0EEHHO2XqXh7KP087vF/R5RoMOIqTXvuLl00
K+lgGZrCrGscZppFb0YUZgmhteybzJjVaayLGhQuXzNvFgNzKc9MfJk1gFxK7+eCljmDCUrzFUv7
Im/20RCbAxsxtVBNmpiC/FZygYPFUtjnIqoi+k0wrM7vqsctcw4As6o3RURqEDXkBEeksqBO7q4T
c291bJdu9SasQgjeiVsxNvbJwp61luyaiV6kR+OoOqEeuF+D7AlpdwmEsAo1ZsdyMaP7ncek3ZIv
SblAMIJSV7WNVWr7Y6ngkFTi3SJsy99EFU4Wdn+ZLD7MC8rUDVTQ+mfMCEBuH1VrvC97o24xJrGE
Dx37ipWGIr/PL3rhuJr4WbAf2x2L/hculMeCt2a9xomGpi8uzEMCcWAifrJHaT6EKRfMFdeD0fMK
9AEN2FYq7KUs44tcFwW3Yi4kOIM0FVDx76mHXxGuVuDBuZWBPlkqWfGIX0jB4lLT9pZ9HgwzFdbv
fj9+/vfNiDl1Lvk6xofs70D9Ux/9BuJbiBKWg87F3dKMBXOm8wDKeDGAUZSYseVBEhv2kDOeB3rx
ofgxB2yBwir0FcPpbV/OoY+G8hAp3aReEo1xH82VYfEhY9fSj4Ux5FBoEtrIPjWLLCcYHaiaed+d
BkW8HKor4GqD2JLHunTwDxIvp41OSGBHsLNU0G4a/0nKIh1pF90CXjfsWGNhGXBvawKY+sJiOegD
nRU9+sosr2eXy6iXqkDAcBZATonE1wclfCDMoGk1nhU1Dc9FoxjCiKn2SL35y/2pFNeOdNHlziJx
7Z44vyM4A96p04EpwlKjsm/3nJLJnKmcpmwx+ZU37rwot15oN7p6r+Ovf7hbAX6iR4Hq1sc56AtP
bGBpkPk4Ed75ZM+wAZzqbecGcRgdaJNC1OQiIQKAhqPLRGwLJbYO/jdpYeNLM0GVgcxk+f/2Hy5J
WiqFHueWnoC8HJwaATZksrk+dMCXtRt0g9idCyAr+xNDkfKm7z8G8sniPjTthEqStJpd4nE9PP5O
h86kIFVTklVaTERKeDagd3Z+R8Job9fTYxUusH9WiNqxsap7c/Oz4qwO/suMFBPTQVkyH9P/euP8
jXIy9AXkAJEa53GRfJUl9wpRHPPoVpTF3sanx7t4C2frcTKq3eLnX4e3Lr1kflTO1KPsdYFSUpBi
QW2ulYe8c9opDmPExltuBW1hOVZQ5VY7IYDjUwHVC7/a5IyXkpkd/lfisrVusSnEiZKq+WWM6hbH
V2xqlp7GMYUAGtLIdB0zHxvd6pOVk8Vew04TGZ1frTd94vEyeT0Rgu/xItkVbgywNNvOxPpoqPIK
pXAHmjQvuRqMvOrVFuU/ikvUYg+fbQBfrO7nt65c4z2+K6sAN65DWZEzjppguZAVja5EwNKCoj+a
v5PuyqjLDl3QBL8TVpjPSy3u67InRLrzOyehmmqc4PKZ1ZZtWR8SLJqTUp6ddlcgaUktQUROs6Av
9n+wvHE+xksmqjhYwaYs4BHTqxkKvLdyz0T5hbAQe4TDsrcqbUDJAVNsZgfGv1UQT840Cpcm8Swa
B5z6RsNceja70P3kis3QQF20OWRqMs/ZmPGARUJcUG1Uc8j9gkNfQLroL8FgxzHUOALTUsA0lxn+
lEtdXWdtvhUnKlYVi4sbBLRNbirW5Ou6G00d+g5aAsd8wWFROewxgSybV4H6R+XI14Ytiyg3hNSd
6GdTvG+lJC11XlmceamyIs8FjXH4MRnILAKg5XbD2COsiktumoU3tenBa/7yn+lpmUMrXV8/U1QZ
ySRHzRaR3pvZTDYML35A+nmttUMYNzrm6GMLdwWmMfUb1rvcQI+C/cjCBoHi6NNOmMqvGpY+Rutn
pUs7lgEjFhc8QGhooKwcHNUcfUxxds3EtiQnx4TmV8568Zhdq6/wgHNXD+CkjiN5Haasmbm9K4JB
yXdebFQ+/vqLO87t8tstHATdZScHYuJLpQqlqpgZNW/OTHlT71w79gfmBkO3sP8idLWsLTtflej6
ki38oPi5CAA23rfRLCFkz1rpQ1wJEN6tvP8eFnTQaQyIbfP/cLlDZQv9IhbX8cQsq8nEkojyIu8V
Mu3hanicxB0UG9IDMY05fjIYc16Sq0afir4w8md86fjie80+b1ZKwrGdCU08krmYIpDK09bGrRET
9I6A4ZBiBus8ReCNqEe1Cgamf3TtC2ram2HVW7DYTmUaFDupiGTQXYkUMaR7/lK6giIx570ubGtN
EYaxLzF32wG+Y9bX2oAoRugGhtrd8ubw9nbD6jSnyAsVC2BR2JhUSrfgBpndjReqDTli7R/iwsqq
icNdTcWIU7nF6JYiMXg8UYlsIryefYT+Zszki/hlFSxOAak947ssnLz7TzpYEXuaFbxS8FAHSgGG
2/w7b5AimnB9S3/gt+X4CmdJxlTV6ogZMqehwhTjFz7MQmexTbQG7tCEvFPP8mFiknsaDm0M4HEb
Ac4eojxVUCUfRQaapI/ZWaPPvt+XSOK/5jOziK3Ui9tosG4YkV3EcCmHq8cL1JU1Ve7UrVFA6lq5
c+t0GU5+ainVrIJ/sJ/Ya6XRgwx1PvO2yHY9E+W43sVOGxlyRFYTnbTakQukJJFz3ZBRYP4a7KJh
ez3OqrcD0ZKLBxRjtYEgVEArGVmtKlyYVIiXAiTZFJh5WJD9n7mZYmMoKTDHyKX55aSFYj4UZvGv
mvh1kAXHvLrYbvr5U4hTbU82qOa9xQlcu+oDY6JR0c3vmRis59dpW9i6VAdo2LqR0uhwNIVJUAjx
3uUQJ6k+mUZb8hdet0J0Ei5C248dEcN9FNNv5keuW0FV9u/deVplzqYEJ1oaoA46SxLDIuuvpABZ
GSoutAPogRBfsgXj98CVSNaFwguHh0t7mmmC9/k/10G5HIPh2v9QjQYvCgFR7sPhuPtvYAG+o34H
YefWIDGFVt6aR+uGaGn8nxPsRLCEtiGb9vu8lgHDlbH0XeHAnSn39KGiZ3um0Cl02hLsgS/iT4VW
79cGUBif8Gm39OOZnTtBWJgnjy1kJe/3lSjcsZgKFRzy4/Vencl9qTi88gHv1dYhwcoi8oOm4j0R
61tQ5Ly3qqskgNbVp5ratv18c2aZG1To/n255fiqWDw3uZV0oqeipgOUi5xMgfLnAAa28X7E6HKa
fDjzrg7Sqc3rVrRag5ZquU2V9twwCiR/Hk49kk/49FIfwbDJmH2RV3mhWzTDFIrJ7SrFXeJDza+F
puQieuJ/+mPH2BORobup2m9o8xNfwNbmgZgOAgL38KA1jwec7TZ1NJ8Ie+PFfMl1LSTHpYccExqB
6oD1iSfWDKhYcmGtkob9sofZv4j2/rt2sQBABrfojRROG3hRgjsrt/vZISBrrV5uJhq/7aGX9e3y
KHLfbl0WZZiq1BUwQFFomKpxtFiWcjqFzEPbkoBYVusqxaNQ3o9Oc1KUquVa62KkIRQlocivpkD7
QVWzedkLY5TiVqYGYUU3nydGVT7EP6O3JcdFCytuqVbJ3zIyDKDjQkouX4LKYW6BqMHozo4L/eV2
wtwT0l/y1/eQtJQhk7Gj0HjNUTIGJFW59l7V+i+QdGGwgsde2JFrlmC4S5mMyNq3cbvHoRiWPVkU
x1IaYPWqB+VWx2Pmumw+iK2iz/8PRwiNAVEUZYYOPuSahGblxhjpA3amcnTsJgw3adEJq/bXawYe
TxKzPphsxXkMFj9gp1LW2gVx6GGym4ZHEWJ5/rt4MCmC+z5UhH9zjbWiqsik3w/RtbcM2qLyXRIQ
5jiwHoAZRG/UzrsgpNIkoJ6N4dPBTU5TWKtQHogRFDi0j6VDLZvJg3w3fsAvllIeCqz98CivILPk
haE6duUSpBu4wpZJxVc68BAMsVdXSvJ8kwqMzuV7tRxeOzrUX866l/nPhN0BJpmoYQwEtHSQrJEN
XwJuh6/DJ0370ifOwcN611TDC7dy4nyEj6QG/l39QsmWaG7WJaqHoyb1t8CU6BwMGBr0PZNrrnU7
CW08IG8IJNPaArtRF4+Kpubvc9SdEbYDqTQF9BrW3vnIi1Jil7s0MjALCT7vuAFq1g7wOxfdwdmR
iXC4EpL3/42mcBrPYqLKoYeJkIyUsT5i0pwpknsWSyqVvEpbDyaI3Cdlr8lC1lBX5+4nAFb2miiG
whbPwII+eKl9gvSCPCxL9MKsJfQyN7nx3wofxo1vx9bUuWlBGVsZcNtUpMfDBITWOokd/gupdo2v
I0P98x9O9axf0sTB4p0KM8KViMZJxMyY5vwBZtItOunNSf8/B49r7m3QLoNWGNooRN0WnVOLqKE1
5QDwUYEWEnSplbDLRArMbgnhpCA7Olugaad4QmD6JgRkUG19oObekHqcdX51nb6g1NGVKRrmAAcW
YsGvOdehRSjmEzSZdeBddAHnzd8rkhjs0Q+niXibHl5O5KR0SdOb2hnsd26vSELHrxGHLUquuVlt
33cZK56EErAuuTcvLRT9xnq1GBsb00uu6/oyUWflj93tNk//KcSkfBThfVznscaTJPUHp3I15Aux
RjqXpydd2Fg7y97g2xMIgSgTNynd7vFd0EADW5xe2+zxi8IsGfREfwB8rPruVi39oE1oRg9+wTiK
GGjaGVbo1znGA4o7Yfo5jKEafhLKoe9t8Vq5OsF5KRftuiET1R5FePEua0l9mT7EqfXDO6fsYNzV
d91jw17W2YjLnCrCfxwPEgibXYYLG37D2IjXG6HqgU/U0wML8nXDI11T/RZ23j3H40o0ChMJmFqc
VBkeJNCCeHm12lPKVnysTPW9+VRZz+0lMamvSKQq+tIqonPyuahzbRw0/MMcf0YJVXtjRYy+5Fhu
bvk+BFPawjWQCvmMsVKVQsInCTbNAtH0pbYN6HIyeBLCKSK2FW6blU7oxz7gHgTmpnc8cZgGh/xO
1oZBdvIU5jWfPswE97kIgxe4iF2RDywe87FU+BOEknZYaD/3kcngcdVodEM7LDC7t211pFhL6awW
7kmshYXnLDha7kG06qzqdudsg3Xn+z1kz8jMrEw9NSM0ohvsSVTWlRbRk14Bar8tJ8gQpfRYKZ5o
hhvh0+Cx/q2VWuXA17iqExxLDET1E2tff4peHa6XquW0V13cJa5Ylsfjv1qzASh0xrOBGAt2Ovme
o8GOllA+5GB1OH0GXNir0z+RVY9A4YcVngfIREP9HkfAtFZ2HUdCUzweqJO5IVfvZau1wBXaLSiP
xE5NxinDNf5Qp03xcAPl0t0hMrl3BKMGqARwzKcAUD7kmmHMjV64pP1pLi13+rAwvXS/lQz9oM7/
85s4KQhtent7EZgmvA8WtR4DizhVractI0U59NYKcZNste3eunJrNBzggejHOmEMqL/Cg9ajTrIz
HIHRQLbQwZUUMRMEbZJg183sZz7qRn53wMhwx2xJ1zhCasL2TXMuUG3tYTSeMm6Kp9V8WQ/ckjQe
D+PDP1+6+7Ceot5f25DJvhpRWj5fQyYnKf+1qVB37UKhCPaptE8KuufzIHCNMvIMiGQPtzOBlbwF
j28jCItOn27w4eZVTeKtjqyBF7eSwKi/3VWMqMhfhVEWCqtc+qje7eQlo/isGHk37l33V9i8m6eg
sBjFOsHdHzw/lg/Na6LhlUPfUuJGW/NqxAP3L+K/n3kfmxz4RmPsxDt3axo1wTCQmbdfvM6paDAW
O+/8OtD/O7ShVooLIa1wfh5HswlUqx3Jh4sGF443SWg/uRj6F34o3ZtR6sO2zwJwc87LtUXsyAcw
p0S3qM3hSYs/2XhWFQMLCOp4kJgm94JIm8n1Jr+dP2Mgj57gHabPtvirb/EjYiD2mUAsbIdYisWm
ESrwBA3GTk0cDIwKIhH+aZz+awGYJkLdm64+QnUJelzKsouUOIu1DvateRuWaO71eVGzJtgXQENU
JS1ALoXY/MOyBYAYTYl694E6dziBntGgngP2OLZE0K3qoXiZeTwBUVGh4Xu3HTrX170pbouQl9yo
l9UyeTQm+943sRsSKQIbY8g9RYBYNiM1daWb44eFwnfaq/S2osXjy2zp4X1rzqY0Jy3vsiW0vodA
bgML1IkPGI3ch08qdUPJLTW2P9ZyWfsuAd/6KKUVR6/oa50O4+l7DLcTpxBPDo6qVLyZKAmGOa9z
zNTsNJDtsFPtlF/mytomWNI3/OwQmGXd3SH8mxiRe4vEYtTzBrDsLsgNpFmsGhhH7BE7C3yrPJdk
g8zcakPPYG87qjl19A584KstTTvGjpiLvcj+qKwS9rZ2aQRkdaX8Jct1Zeab8dqSMuRmYeb7alAS
tH1Dinq+19wccIseeaHFhyW3Xzanil1fXvoyvOcfbgvO9b/sjfFCIM+iyR/IuuzWbZyv5CPVAng4
oA1er2VDr1hAAS44SdvPhmAOIsx0Pl7FNyYHaG2IjFo5+q2Tu4zH69VtmVmgFCSa1Fe/SdpX+fv8
0uy8AoTCZZchnBagt1t3EVo4KS0UD4hfmgBEJzKpTq5CTOMENM9AXnFKRZlMJd8BnQMKZbBgMuHH
KdEb/qT97sPWMV8a3+8kzC+2Ql05qTaZ22v8rUMScAniVD5g5YaNdI14egd1pbIEsTILDoy7z/L8
3xKEemhBUBV41AFAJDHq1Jq4w9WZkjx60eg1tKPsDsmsfvlVPbozD7BHVg4ZfdQfELtrK4HwRM/T
UdkJbKWq3//+JAe8l2hBgTvg+UUVa+LdNNwRTb1XejfOk579Z+gVo1DBtb7MyndCkPfu+eD8/fkz
UCYeVyDsLz3HwIUxJOPt/oJIsKkDGV3Ibpft65WxDRBBMv7s7YKyUopEe+b7G9r0PDWfBdeh8yCU
ZGEyOEyYweNh7mFJphSzC+1wwm6ZcVL1dydP9oYSGndm8OLgXmqlEBblTkJeuuzxwdnp0NqWCZmg
RShrtF59wUbRQ48wE49JUd1iTx2UZ3B4fHX/5t2+NpDxiTgANx2PMzSxcGth/Gw8eFvkZlCy5KxQ
g35FJdfnCC7FHIUlVDdxqkrM4Ak4mOzyDTljckgnEC1EKj9FpbM2DeXkAHBz803rjzzuMS7cWDIn
CV0o5ol3hfmGBcxA6s8PLlqEcWM42J11wx+gBRCTXJLHusoG5QHSiFZJiGvegEM8uGlqZP+OTQU4
s3cS+dFxK80VhPpD/ecQZZjky8f9icf45A6PxibXgVUKSmSpPSXhEKgt5C3flCKez5pltExoN40y
Hd3n18fvxK3Pgrc91W/V7J1VyTdjAAQhjZDUltMliTVR/Y/VfBHho7TUHGbMlf19f5Rs4HDgFwSI
zbzi8Gq5eAdlZ9XsTOypbS03hJ1nyTxcSNPXow9MJRPXGlywNA4jw2oub+aOV/CnILPiUIwa+kum
T/xnIJXSJVfEJkAOlb3XotYK2EuWCWOPvbkpwvhW6l2Ufj1CAlFJCOGNl74hrIQfd5TjLxzAIeb6
tCvAb65rHITe6XkIqQTAIIlenPQD2Nsv5tXika+KqbNytZLrUDwxZwzMRnwM8vsxd7rSlIh3iI0t
iKwej3mgLAW17PkOPaTf/XqcACU8ROtlzvVX/oHO/Dpn9lGSN9I5scv2d4lKpp6QnH+ro+twfEAa
2JqFGUbZqk8nMeJLBHg6fBZhgpUQrZDSzcg6X4h2AHt34ZQ5lJ9htUHHZwJEEKUy+goMFZcUCWuB
Z9hn0VYRna0NAluO9oLdl73LZK3vyqfMY502inMu4HZyYeu4/SJLhA6OP1KEEmWYYsnfuftVEtEB
ckVXpZtdVPWW+IO4U6er+ksojTqOgk1K2WKAkHe+xBZegp6eRxd7GMb/OYhczetErtZB/uVctTbH
AaDXlwozOkbyhWkGGQX28uK+Qsd22efk1+//u+MFPG7Dnn/9wYu+dATa6YHZfNg751adXmnqDCDj
0ZqMT8giVcMP2C1j4XNOzQ8xeNPkQGSk2auDlhXJvVjYrgswpqToETdgO3UdjmbjuuzEnEOPR5Hq
/cSV0baMqvjf5LjutihxVSbOTsHc/48FL0n3xE8qV59E4wjuoF/6/QQZ9bDutgmGpyI/OtkQ2j31
9hNga6FQ29pNX2EHVMHszWkBjNEizg+l+4o3eWwmZxoWemhKdxyi5yL5psnfTJGw31e9eo/cowrS
pGXJdZ+5VfRS9vfM+MNEVyQBQdD43vlRBvvqn8ecWsL3zEbin8uC0OAfje1XNQWQO6hshS9KYVES
2bkKhOYuAlESVBxCK7PI4VC1iOQtLvGqKhauzJ8oUGw6hhKSGPAiRtsMkh1Ew1EF7rQyMJ0oNmc6
UwCD3CYvny+Cb3LNsWJWVewwoKVS1j3l03UdfIAex7YUZSiCnzfuXziCExwrI4OE1nXPKkGI9Lua
CR7JPKwzjsv8kvWFSwF/wl4x8upxBTxv/WpkH0GALT+EQ8EsJ8IIrCXxVhwcSf8WXQDMeboJ6+73
UTwKFrB/BUC8hC6F+r6mR4l33PFM19sCXkMKeXf0cMBwLkNktqGWQgI2pbw+/gtByoFAMdWQRhYz
z0NgnWxQVUxNbzGXNX1r2JvUAjXccmIwt22dDgurVBfKNPIkKSWSXWg6XGD8UmRbLj6iBBlf+9zK
XxE6UPPWRQi32unSMyTqVUDWWAM5NlupTB2aBG9rm4NzGc6cZ1xrDgpTvHivTt5UaGuUOdKoOz4e
4aD9P1YDMeaQskUwtXIj0gdPp39/v56hIf/piG1TskCbpvuLABzn+iKc1HJKc+RvyJaoOGH1AXAI
NXgKl9gM7VA5UXQ9i73Ii+AtUygsDpd/RWUa2FR0jXLAqqvKCavCG+I+Cvk86FzKu/80sAE6rGtp
vVWhBr0Hk+ab2IV1kHvfMJnCWV9hYee/no7OVMn0fbzOdj9uawFbu2q4DkA/C1AMcsWuFsAVZ8FP
tgYGszeEQ/igMDvHitbNNEJsqqimc2NEZXPtEZnl7kHdcb6EAh/JFJlNikomq9AjjkZ0aydLW+7s
IlEOO3WCc1Wcm6xcOTpFL+i9OTRY1chziFCqoY5sRk6aYI08zlx69RuwYQHCd6rugrp+yve1iRlE
AC9tg2ikhZFf7DtXtBi7kpOPrtI+ezQGRlttJ+biE32bLMdXwRUnM4oYeRmjsaBylnGw81IeL1z6
WSQLfXyXcU+zlizFMxHzxba9pyys6kuP/G25vFz+/9xWmt2Vgx2UjqGbT3KBI2ScU3dBpS+jw9gL
TvZtyvbbJPy0zb2lPiGUskRaSJsGV6Sj9rfHb35+J9cADIp25UIMod9Rz4KcMlaaxaJ9SD0/oq74
kSFbZH8G1tc5GClKIZC8IdQvlUVmyeGKT7Xl0IXbQot6XP2XiaApSexE2mZvSfb5vrfDkYmcSLVJ
y2GahfjZIqWCa2bB8octM12kLlS3vGBErhGBq2i+Ze/7tY6w/w77AY/yQ1UDWNzT6lxd5XzfsWeI
AnmEtrW2VkuWRsBxWZTLn6ypTpAMii2hgpVRQnuzwsv4uqGA5VLT7ZraNe537hN0zZgxzgpFOrV8
rBtPbR/fHw6WtD54C4Ooi3kHct8q8p74GuQsYi0TXr92CCFL8Bi3OsENVj3WPiztzZ+CH6ve49EH
MjSEK77lQQwdAnZVDkD8JlQoPgCTAz4d8bqdZk81R8vVDdA/OMR7n3y7JRApgfHTOufS8GxQfF4+
4aYsoyc4TL+a7uZjl7MZ0rOpqOenBGWZ8xF9vWqaJjBS0G5DhrkHF0Bd1VjnrkGvkhEDIwsbJNA2
QWfiwlC+m4En66fhjfnB27aI/g/SZgHRX6Tvh+WaSBQmALDMLfF0/VD68O4txT9NCgChz6zlCOkh
iLt2+nB/vIy3MnmS+TWhu17q+Jlb2LIsy1rgsMt2Ys9XbVsN+LLftjtoaXjw2xRAxxfbHv0/3w81
1qIpZy2PumVZvWJmd7kIDepPWvczWj1Oi0Q2ct3C0u2WqpXWCHErhRGuxbnGJHpU7iFwxMxjsA2C
ih4jYlQKQi6+87cPXkN5v+tZoiprPlLbVqabtU75/2f2BgVIOmQULSD5VyOGIE40nzQPd2xSsisQ
HNrPBBm2mg3/5KG/HSYms7O/Ky61IToz/LNDPfpCOY+CJjGkTJ3PwS/toS7vjQyZNUEcrNxNLBvC
72/TaPgTMz+/v89Gav6FHz0VVGirVkoYuWswnr5mJZ1H1SIiQ3u4MJhRHze5LHP/VixwnygMUfnU
0wyqMs6mmOQcOl8FA5RRG5IK0/wIh1HWfVUr4iBJmoIw834sYoEOHUk20phW5qFet1dJXkFo85uI
6phrum0z7VSwLtGQLO0iKeVjW3AQKE9L0+SXLXiuUOhvJ9BQyxdIAttQtV7DDRvAMAw3RKDZBi4F
OejNEmgtXmdrvO8WSlXV9n2qoNBGDsq8gbiT5ueLg9zb52TuGGPmcmouHheaAO0a4F7Y7qDZYpyM
yMAGRqYDiK+SzweDsfZmj2gLiSg5tymx57G1ATQBEW1HEkwuWDYxyPEDIy0G7ZtFjGv/Nlr/0SAM
Ynwcu2wF7OlNh6sglS4zl8fBt9zyGS8uQPqlUll6cGcHYd1s10EWvOVH2cV54Z8q8Vm/yPCiNQ6T
nuWjA0LpH+Je7TPVGQjU/Pf37XlUh2JWKfsoY7F28WYTQaGTtZqn8FRuM9RCUpSer7zsYSqYgB9j
Vo5XXLatcDR1eETKOn1gEuOt+W9Rpu1DhyaWTtPkjMKYUqAaNXuNWkxeEsYWcBnvpFe6xVSXpl6q
NvU/FgLW0jj6gtNVEkkjqyplUwdiHVsJTge/VHraXY3MpcjyxNY0sm4b6Zv9CnqzO6m2aeGId8R2
LUKF/Gz1iJwmiEmy5fp2gci/uWC1dThVG3cos2F+VEl7sILdgA+UCfGaziNMWrtHmVEnozXxw0Qb
pfvVwJsKifkozby7SyMGN4FfrJ8/ZP5xoojM3lhAWX3WhjKqm8h5L8LAFGHN5rIBn10x/Mx8Uc06
ZMLj6ao+bldJr1K3n++kazKfn0und70osy4fM8nSfqXQoiD07gSSCpUKVKcdag19y0HPyyXL00KR
aaow9ckyNT9ngckOlmgHK2/JFc83GogY0eyTYSF++J1BPdEAjrAF9lzW0V1k7qere4eX/g9nsS/R
qIb7JntIPD84wWXTgfA92WuJmdk9uc1LQTvFoacnh0faSg1yOwC4tZEeiW0wItkPrdlqCfxgjwvT
QRiL2J9cIQm5hvaEBn8jefPXxezJ6kFPR/wcHfs/qqH2y1cf/m5KNYRpCwSHhTgwBTbz4n2LIWpV
PHoIQJIozfIVsv+J3Elz4RX/mDdyFvAusb4Z9IrSAzeozwCI23160fUyPPV3eGAy7cJPCDKdAOmS
tt9hQbsVOXbhsokG4JZzYbeHZV69uyHN61D87H9jqSLLOfgXr0MSjf1cq61RC1ukv+Nhfh2dIQPK
EuhQ/WOztjXFpzoWKTVar1WfIlIbrHEY6urHu410o8RT3jeVMk3OwqxJYOkUufCWbF0cdUEFxNd7
MvCj2rnNJ2aVhV69l9bcAy/5jrvpabRbzR4D+N0xHRht7mIvQ/QADc+JEyt0kpjnNcu4GoE1iGUY
weOactGJl/c0+aw3XBorB4CjtUvONiESWqnBP9iQgsa9EqOWxteYDdy8ZobqpulvXaQPHo6VDGUy
tXtqUVp1v84KA/pkyWxDsXVFoB/nKSFg00OtmWehxjR3Byd5ao/1xPqSVyR34Q/0vuzH2MTUanpK
XItinpfgfz0U8+FZ5MVhUd65HHs0RlBTSmz5oB6KzBo6oJvFo9xMLK6sj/iIVCm9HsG6rCbGXdEX
523BaCDwqwqcDDvc1DJwnY6p6+H7zPt7A4Zp4kCadz2baOJfbj+Dx9vKLLpqv0HAuGxHXa7UB7et
Arxo2XV6dWeKoFDfFFUf/Cgdc4sZIhxx2jT5Dabeyj/qvDp7TPSmbkz/97mEuaLY36LnNQnjRwYL
KuTCjtDBJUo8n16pgunA6Zq9Sv/J9L0STtmRQJoIzGBGQm21ickET9xzY7I67LmbOURD00qVbPo3
fuk6s7jZJDzI81jMBdURjhOnwnpwXnfELNIaL+SPJ3JrYNFPaeUNJLb0VP8w72zms2Y3p5O4VL31
0Yqi7dUSmA9i9d4Y/H1P71ZJihj0b/gorx6oF2aDAnos5F5V9Rm8YUsArS5vz619hTWplPg3n7+L
sOC8vzeUKe+ZSsKsX6TVBdMc9D8uAZM3tOizCHGJJLvNoqRNZlTPDYbE/7ZhKPQzKxxX4FSIsY0v
OSktZyoD5CqISDLnfU4YaaaXLUcXz0JQVTEIocZXoIUCRpr9VtOp3GUA2oO1w0vBIhP31+FTOE/P
JGUFWokfbzdSYQm0VMyWLIR0T1QKTfutf+M1iDw69Df//pjvgdfoT2geuPRI4pkxkJcYcxU79Hrr
SSiXcOK+QZpvRmDHB8Tlv+btPGl8xldwYQBlLhRSxDEmD3+0BYDR9PzygSpCl/IwK9NOfL9rJaeW
GTZomPBj5QSQJu18V88/Z14JFkzMlYG1r/f0JCnsghxSfV4/QI3mM17ehvyYnCSyrNulLkZvRMVJ
VvLVm8jeONJDqmd0SvlVZD0VGZvK+I/E7ueFHEOHuT/NnBOcZXW3wXw4qQwxyXldQfwLAecGbx4y
HSPy2Al4GYEYx8ZtOvjE5G3O+3P44YGuIHXAfQFCpfD6/ldu4cvCB0k93S6MkcAfKtzuaivIjcd+
525WX10KwYaZ0pVMM9VcXkrhjRXH+mH06uj6rbYMHCE6V6BnpGB0QDlkbhhAnIpENqdP9mZujlAg
918eRyPrxwttiRzILEwS3WCziuld7TwFuvIBbR3GntVr9Ys1fJw7AuwUU+TE7lifG4pHMv5oNq0k
F/q6tv4ae47+hl1CifPuRwLIeOIuyeOD3vxDqomWIIE+S/S+o5ZXrMrvoXh8HnxQHfeVLWsWUrPu
zGJpG5nUeteZIpl0dJJyXtDuNimyKh7SWcirn/N6PXotcbSBbhf8Sw+hIgnSunRXaQiZdhEJVxob
TZYABciu4EOgQ89VrOvIFVEHeErfncmTrhG1V8PdAM0COSBb7J+ssUyeUajh98YAT0jZKFi4I43y
cSqoucNdVxsgMtUK8keqPZWGbWooLhB8DwuyCrQeo4E1koDigqfPm09JwxJfCd7ZCfv9Vr1ntn1L
f3oasTO1G54jIPH7qJ8JbqAe8KupEkSzWTKevTJ9CjyhRc2WVVlxPSbNsbK5rzIfOccz2bCZBKpw
UXovfnQf9bBQULDaiEf4RNybRKUCDizwiKgYC9rXaOogDdClYbkarBCkk8b+uSC07qCz8Q4EHy9h
16t5DMdM60d/dca6idxCGxjc8nIC2RVUnCfQxQN2e8WOLfNh91n17YHWUjHbo6AhZ+ghpFrJ48Ta
F3AfZeA8ahi8CT7geR/MGpsUiMLFvW5zd+6lu97Rjx8xdeVg4zilIMgMNjisdHu6KwoO5TZuD6Q5
YCrfIoF8NAyYkLSnrS01XvT8sRNAEKtwFpZKl0WaUAwv0CCgLMId+dcsUiHypdrNEie63qpSXdrP
StM2AaXZyM8F05JQJBLQKZ4E7EkYrnfyKUcavgAXEwXUmiAGQ8mQec07d64PZHiAUgcZCvfdVd0d
ckX+ZJmIWW92vpYJLtVRdfmO1wXTl2sc80uTtkNUaJJBt6MYS0UPY2zViG9R2yDp16YL8CvNNVNe
H4PTRVLbcjdmbcT6zuGdGQ5WNtxut8hkK3la7VU7ubWPYj2OrdjTJ+bxswl2BZyCcaPxKEcKZfFC
f2NtijIeWVr7kK+airnNnDW07vuBotmpZno3WG4NW35sf+zzN7e8mmctv2C8FV/GtbOYM8S0+PAd
vCbDUEAwMj9hMOqT5+atEWOi3Gn5Jz4HuxMJP4nmvn/Pg4Bh4Z2oivt+xlGe00qd5PDvC7QI12lU
XfdpKVYDg3QhBpW4nbSGcnx4GpUWcG6FAXNewP1z+llYmyv80TFEDFWMDlTzCEPfx72o4p70o2H0
6L/MsYpy9fi8mE1rOAGE+3nsE/CQFa2av2YYIgTyBpkGL+Q0Xvby/lq9f10UIcTx8IZ9iAbw2X2m
6WnA9K1ACrgKfpIOmXGg6ME3yKy0RJlz9PohjAh/V8gHJ+6Mi3Txuj1WmKYAcgkHdAn/hBPtl+yU
qDkflg4QsTF8QxfOREz2XVgI1AzLE/6HgSzbHaLRv1UjQUSrcY3AQrO/BVzV8uXkw0huyyYvYa9M
mX7aGzanNgcatGkm+ZJDD6f7ZCb1gU8raRIYLe3C4oj7eQKhF3FLCcvdS1tWk6RTz1d2+KFGm3QT
tWe81G81zfw3kt2G+ph4UWxC54t1PSzHaddVYhh3zNIhdnMMcDX3+SgaZLZpVq87+BBYYZsUlAhC
3RodncbgaBRPCtp2rZQnSVs57V63xQ9GG3Pf/mOJClsIrbImZqKfIuR2hYy/R8oyIVipNHl9OuOh
bHz25h94ioJ2gzywjhkogomln+DL47amBRIXDJMGnwoncVPkvtXwie3k+beG0NoICM6c/hDedN9/
rnyy1ucr+NEFQdWPY36P3BjLFlM0HCfjDkhQwjbF2cLUeADRKJFBpRqnbMLxZfJP+LhQTUjVjNXQ
tQbRs+UZnIsCHGI1cLYnOkyujOEpgFP+gWj+0D8EL4f/HRhusugKct/955PoNiwdDRH/C3qUzWSP
U+B2Ep+KkDAiHCjPfnknpXAMpWfQQWMfyOI6tOfvl/a5hf4aIA2dcWUSrmFnu9laqb0UunoJ2P/X
X0LQpuFh0s8BcwTh/Pt5h8Ndp1dB23mCRkc8dtrsC1VbPGAqdHgtWU93IW2BqJczWro77Ur40tFc
A7aBUwqYchbhLJ/+5H53fYGDtupJT/5kjSu27a+I/i8jspsQElxZ0AQKUXxGAevpXPXgvi+6pjO+
vECSNwt0IDpWMhw5OcQ7/BMdXqOsRPz0qfqxZOaK348V0SBX+EOeHzfPhurDxVoBHbUx+FUw2t73
9ME6r5gL+geCx8w6kh0sJ4fP8w7Kj7wiTI+hSMvFNIxjMgxCD4gNZzm1F4nWx3paRWprzhdAuZ7b
A0XLkM7QWQxCKUUJd4bPnd5IhNoIGcI/X37oRoYAHNG3/H6eEUdEhxOM9kiG5wIpaLCp984SuqcP
ozwhqNXY6wZwN+EUFLcucPFHvI7kbUj7q5gHLeOilnecdrqfRj9Le5n3haoC+ObUJljgExuGhCPz
HK2YbqeokWujHg+Ae5aivqRjZVZtInD+4JyCzk0LjgME14QVjmB31d/nhkNhCyPM2pZm1m1MluaG
yYi57u1hHaaawb/fX/Fk0CY7Nw6Oo40qraN3lXlTpJtf7tPxTIGr46R7VDgzCc9h2afdkVTIrp8I
zkajDy9zet1RGlp3KhFA5xk+XZX9CB9pBa8Zdo5MhxSbD47lsmKwdb1Ch87tNpMKph7c1pjM7D6v
3NIUmNIjKCylQAsr7pQdga7p2yYGZvj3tzYQXnea6nDdrrYEjiO+NcUsWErl4WsktI6/pL32xxmh
ryWVkVGWmFbbXhy22K9u1A1CRS1d7IQFSiA+qM6662fHrkbbLt1Nc5aRPTAKeC2cHaGoGVqduXFS
pefgR22+UtKa0kslYbAUlVwIPnXBYVWdhwXZJsuXw52Ax0JCJTZ7HoDIsKp+VY7Yf9Q6u69fJuhk
zBKKiWLo9K9+8Qge0uOjA0No4tPoUtl/w7rfdFs/1SMIT4d/6G0kQMxAZLnGfryUZl4ylnoz8178
v9ib7YQGYGWolDEAYLyVpgamcaLQMiD58kqSPLSxLPJtQ01yIjs5hi3ujrZTDxY2SFP2ygceiEqt
2csu+M0Sgzq36yi3sz+9SwphhEGcbVus3IruNJnP4mPs3BV6AMlQa0ubfuuH2RnbHny/SeICKxEI
E73UaSu6XFvKoHYtf2BVX+BjRhcK3eIf0w5qOgZ8R/2H6lXmO18MUGczG0TNi9BmJes3z12RIm9K
5O4Dm9XaXMsyL3TBmDWAt4SirLY2MPrYP4JIPEltzMnENS/FrkfsHWiV8ugNVkAtiqcmZgxe8iXi
QGxbL73tsfWSHmA5up0V+/+jpUZmdhEmtSXXPSb51n0PiaDyFn8YuswgUCd/LShBfKR05PjbFz7X
va0O/md0BdFWVnTvjK/k66qc7jGR0GtUIXD5+e3Axas5SR2eY/INeeKFMuOa5+FrgPb8TFIRr6MI
tesJDfxBe975aNBYaqjH/x/5KJoE8gfUcKkrSnkSHKf9RzJ51ZNJvfPPofrJNa8KoakSj7FUsdOH
svHgcwasJM5+fHnKTFDnbXb3t9Z8Eqf3rRHf6iwd0fp3iyWWpiLAQ9Sti43DKQe1A+PT0kf69ocZ
2CfDzoAi2w+oC0RgmhsXWvkmjlo6GHl+eu9xIYUKcAGF6s2PSqzRLDQfY/1KjKhUJurXODrzP9sS
hhNaz91QlBIm4WIUGQp9lxzVDNpq8q2E7pdpqxnJ1joCRs7GxW1SjwwVJAM/LMnG4IwMo3M8FCkQ
o3i7k4V1ltxPzGqkdkVHDMOxIX4lqbKA+wYi1tBtNj6yMA6LxNtkP9i41l9qfPXTuwIPM4Js75F3
4jPnJWvqIEICnGqYC4O1mdIdT1+gK3YPFpy1lLKS1665eowH6g+PgKEY6lsxNxjiIkQqkoTaGnvj
l3lG4gEeT5S7Tibmc08QU849EqSGDMW1lJQSoz/q5EjdXOGsTbqXUVITBS7A6ZWjwaSm1S/zdlr3
7yfN1aP3Qe25MzS1/PMIsFNjMIFBoxuqyQkOkr95a+xVfGkbYArmvKqFUTvp3+yI3XrfLYVtcWtp
piuwm57P/tbDYjZmzjez5kL8LbIvKSS9n63ZMYy7SLnF+H8C/BM14ish+3TtSqAoQUNEtKaqbgIu
ySnMfMPtTQxvT9Sc2CraDOcmwHKhXsny9Mg9eOUU34wwn5+oWRpj7uJ8Cm64kCuDEJ/QHabpQwj3
yvP5m3cgpLITmPzeagLIOh6IcHMYM0SK5GhorBnPHtrPpt997uU+aX9torrn7senkw49m1BoWLbL
tRv4cBW0ik0izGsaeK8j5BBfbBuHmj0X50ANBadH1gZsp0sKKm3GKP31d1oTd9QSKV8cWrVqd9lj
XngEhFBtg/yVQJfFbicfj63A0k2LornSshWeeowJP9DjpgkAKIoDSMhIvTvugIZKqAcLNktELCXR
/A4h1LdEAppqwVupOoeFHaXxI3ckJ5YBqKVMbtAUckXpMjO4YfDZxHUjjEwvzhhQ5gFr4P73c1Kf
GV4B2Ib+jjd1OokvUr7rfAvP62aLjVfEdI5FerURC3AH52ZvxeTuPC2EbNBOjXQoEjVdL4W5SFjL
OdRCFBj8NQfN7w2oWqguyUGN+lA5xr+69Q55zhgMlC+MuZ0ZCe9rYLJ0MPrKPZYjcDz324erjIYs
YnxIwMqjVr3eqcvh81D3uVjGdZJ4XOGI+TUMqh6P9VIJi27nxFsQ1wB6mdDX0SNIidiIufOGnN9A
yDO2Twes/YpJDI+wfXv77mtD6Hf6aVAdmpu70nFPAcY/GarP8/InczdOP8HV1Y3doY7uZmj/lXpa
AUFaG4wohRr3cgZMoB11ANEObXPJ4M20aYz1itiVzG3Snw4JLzn58YtfBgfukXj+90ZG6RoaH1kP
KBmI+rwCR948Wji34iM4KxtAFkDYSD8Mi2VRPpGZUbwUEZEKeTP4469uro2/Nd8HPN2c60EngrKQ
RbPlQUumCAnm5+2evpxC9J9bodnEQ9l7+smySecACEYHkyCM8/4sKcKsgwXxWDvKWBx0DzPAO62H
WQZXTXsSBOZiv0CHsg9YtGu4tow9z8aWwVq34av/pHUXWhiuudCrQCS4+6qXvOzz2Z4ZDWpkJvws
YXbV/3tgh9QxvK/F7AlXsrlMkQZZlEuoLzKWGys4mAAN76JLDmLqTiUBfcEluqTb5KRgYRUr4U0B
2jl80CbNe5L8m7ObpV2s2LCv5tbbBpy/OLAm4+dg89iWmaLrMWJniSM4CSPhB0Lits6YcWmO+3pV
BC7ogdmuFOjjqgcM5+E2AVwNGu5PXYtA6sxUz6qeL/ZZN8/Hzz8b2X7lj1z/X7QpVz6JwYvxHPGo
8KqCUUoUOFLahZmpqGqBdq2r3jfPgiBd7goEcZQoqFmsJB3zUYFBcJebOkE5PMwDTq1/nTeZNxcH
TFc6te4wtbL9I9PyGbdQrHsrFyJyelscl5kIWLNwwYdVn8sfzuKpgTIGnpfSa/8AufIV5ulqpR4W
gIcc1PLonSAaEaebl0KVnTjU4CC+pVW7KMR00wZg8BlPlQu7E5psoQGJyiK3GtB5eEVnPcG0IVXk
kK8LDuu0pNGzGnt8bnyAfa0bWrDiVrduA4EV06gM1xs+aYed8sdHeQhR3x/xwCEvofyGVmZznLcW
T32vkainGDJWOlTTdeqRqG9I2c2Vfc71TCT18TCz0k3MKvVYErBneLZHH210KGKqOmIWbSREbV2q
tQFHHjy4rxZ6Sv2CXQlxp1pKVaK8aLe2CG6LBf9u/G9Rp43fTcQytmCr6TuTRG6FfWQFEZRCXXTY
bDZ4Bq9TxYBa1EEmpy1wBgEOaGZfBGYDpzKO1gRGpOIj4Rl7Uo2pRiRNg4v5nNsw5Zc7yDwd/1xC
AbslQ0lc5QqUhZuO1JHb2kRvwr67TVRyAcimbvxuRYXsYbhYHhd6n7cqlrNwWLEKbmw9WFH7bPEd
YhOssvnUJEQEqUpAID/x5YNPWLPNv/7RgiD2GQO+fgB+/ETp6T/xy2gPKbX80fYvXapcbYIUDtzK
VSkuJK1+RPC0OmwYL39xdH4xg9EsOwRQjUgO1PRUMW18Q31h/Ft88At0JT9cT3iICJ85PLHZGPQs
VEQOz556O52OJRk2GwUhJPbca5cKQpmWXCJzHZScc+ausmIkpEShzvswiF2L8XoTdOhJy0PLif5m
B9I4yTsEhGfKt6Ca1L/LvclJ0tl0Y8xT5Yt9yCVjM0BpmAjZzgPTTSrsMklF9o7ZvVBJbg4Wd3BP
HAkbUINIQlRagjlDrv2KADrwz/ndr/iLWl6C/T2rwx04MrjyIu7sxs3U5xtWLYfi0OWGl4AgqwVF
Q/JlkidqnTWyFW9lZ6YKq11qcSXA/DikQj1CcMVtyJc1ZHiDAlSVKNaZYTq9pQb/nM3/sJu8WS8i
gIwN0jWc/NqHujwaSnKjF1Iz7a4ykKM0H6vnoySRE5lPiu8H4sUlmIzs0BK6mUuOpGZxjglpoX3O
ApzYdm8JFwAILzJnyjJpSFYVNXNF6Zv6RNFZ19cooXWa5P2gKjSdjSqvG/vkshGRmiZh3Mb6in3O
J574M/bQM/OWOsFP+8eSTiTZzLXKRzaKkZJPqLMPlOeVbzdlgLUgvsGOUJyjyRE+zTsA0ucGo6bX
TTbxzuI/lj6PBEBIQLdmYdJw3DnJtwMNWKGchP6OdKuQH2IdVwi5HpC1p/LEX1gkpwy+0pd6tZMN
TfpyqfGvFr71uv8H8p6I5Bsh7r4dPB+/TF1q6hK/NT5L6HYoeoscrPAQGWXBT9vxsmGSnIy5thYi
CPxU4rMcggWBmn+rFkMbtIXypkT8tW9b9JPcXeFi08rrPPhgIXC3VAdHkpMIf41ahDTsQEBR2WnW
0BkqOuyow40QQvWCByoeG3fimwKTpgYGl7PqJLrVIBs7mrJUmuzlCQhzSTlfhpbwhZgakoZd9Ba1
ObjE3+jIzDHz4qH+SY2U3BJ7mo0fWlbkzn0ipRFd4fSiiTecpUPhmoE3Vyy1wMI54VswyQNTMVXh
33JhgilzBfrj2rG+uxpWgZilS35ql/AOul/zH8MTdAClQzPUOr58TtXRBD+LzN+QnyqqC7fSId1O
PFHmSHvLCkXSQdWhjiOnEBlIe70ibGlQWovGFpW5vRhxZguQNnsj6DrXXDWAIrcnUQYemAZ1Z/7C
i9U6gW3Ue8FqU5C75zWx7/DjeBap2p+PzIgLmxK+6AyFK07HwoHj8pTXWAdU5HVc4cEG3L7LCukq
zZaVsif9fqTjO0yiskThzrA59yf4k9qsTVd6Z8qGXo53Ij8lsWtYz33rSILrszgS6joNXTBWUmSQ
lEA17oRYGB5GW5K2kb1nJzI29wclgfuhc/9atLBBX74KLeoFKMICGjhY7mBjeZVvoGV3D2Kup3rd
thMTFune3pwtO22M0UWMyCaSnML8w5iYPeJCS1GaxidtOcjNnXiJw6Bjn4A5XxLkmhFL5xOKn8ZF
vm3DolbXrm3maFTXQpuiT6RXVfnINGft1ZbYH8em8o0J0v4WHFj4Eta4BtulJqg6lqrNNxAEfbFb
TtWspox4nTVt3m8ZuXm0dGA3dVDfVVSPkzZbTIfz91IFJd8GQWRnITuvvFnKBgN4vp3oyWnAIJOi
HPr7QkOPzwjlrEWqPrWr5mV8HQACm0wIovsAFt4Yba+mici+KCIah0cWNrjxlHF7wLPbfD/JJ3/y
RFBTXQy3jrGWpr0A1d1yrulE9iXxfU5Nug8cgaic5uPZoK751hWi1v9554vAJOZfaL1yqJ0dIMN8
tSuQ55MUdAy5guIlf3q2cgj3PWAQ1vi1wJuQ90PBLeo34c0mUA/TdbZw0XxXhgModa0r/F/dd3kh
E9H1C+7HnKNmrwYITAOLm5KYUxJ55mX77Sx7SvKQvrUgb7lDuxjsGgdvqbpH8kHjUYkuMcKv6rqV
QmjO/oqFIvO8JyKMOsdbiZa6AKIC+r6DyhUqcjqQ4IoD7eAy3oT7XQtgKlopR62fMNk40YFcNhQN
i3Up1WrIsgW6AOAFOFEs8zc42BdnHoOYrCfG/5RfE/lTCO7xGXH7gPnIvYol9+HmDDclSYXY33uv
rr9JMaDs/OMwLLB+wu2UlpSPEf7koZwl0yZyIfasjcBrFeyOBLOY/8XFoDfCDCBMTQy0Y2xYhPoH
aToPb+iHZIBFVdU+z9KKJa7JDgGKYznBt7Qy5mDacRJk60tOlFtaNDEstLyKL8f5nf1cOQPZSx+d
dnPF3gu2vdBkNfi7W7gSkYnUjSl+JlbmK4414YTttc/grKox5Hbw5yhc+uWpMUJQr0fAhzJJ3hPP
kAvGtY50yW89L9GjGBeyzEskuk22OOdn7TA8eYlKrqIcLzEtSLwimKyPoJpw45+TkK1hFEOyzHke
NQTgXWeUKVQHwjjKCwIX6NjemxpQjo/iNyQ/kecWs3CS06JieSF1tSUkeEV6bXE9GxvjtZUbq796
9MC6nEGn/8wmxhrVqGdIoX5ybmWVqEoESqp1jdGob4aagVefLpiTS39iBd7juMFCbghy2D+WMh+u
bqJMwwsIqtaar9Q4Dd8w34rHMOAvp9qPfnX/MIF+Q2+6TofNSeiOweym/oi7pzA2Qe265PhccRxb
HAtagSjJnLUyZwP74wHkiOF7Dw/2H2knmNAnU91720Ly5SDOkfAUw/Fred+6zyBGs+nHWL7J4iDH
/bPdSRVZv9VRGWLQI9notT4z9O7QDZIwanqSioGTP/E3aL1KRMBVObkutRCy5doYnYEQTi2Brbu4
M17q5/cUUHkzCSyfKT/c+8s4TVPfZSNUS61uHocPcmGP9dUdoadeLGNNkvn0ylYiZGd3VN6WoeiI
iF0XQEFWvMDN8XKIOuRAGeE4g5XQaH/3qT17S88/VzJRzdyDtfWr2rT62fMcKGovaTBQuwAfXENk
MtT2bLo8dBrF/3Js70KiltXxOKe/4riROX+bw6XoD0wtsHgMzXavgIubzkaRc7pNs/37ZWFnJ34Y
k0uxtDpTWdXjxfH5yJJ+Ozv0SlHHr8NvcX0LIkys2ELVi1W9bEQWAOcMnOuiramonncrvcCWQybo
X0I809G25NX9m30HuBVkaoLPQf8A+PZKoKBfV19h8aALITvRSN1dT5rqNVGMLUdY8B1J5D2t3xk0
WAYEgQlXw/XM9f8HEcu58DPPpShI99FA1k8/NqortuZfMWApvr9tQQElzdWa7fLQ4n3YnHzqRLQs
hHGdEUnM0XGOJ/jvJVCPfwDpZrZyC7UCbM++k23j1VWRFznF1qNaflPYHs1IKG9lvwKjgS4lL7qE
tI4Y6k5bdxnOEiMXOg5GlrFct4Keea43RNFk8+Bq3yPkjHPJ2lvWfNYrpucZWGEytAYa2L3iDckb
2z8Eu8bEmzzh9sqLP2IMAS6hraNpWRy9PuW8Olys0LupPOtGLkybcHPPX6tEr3MbSgkSh0uGgD+S
nwBpq48iLabHc8bbeSOTa0vGHxdm/93ihnOUlNPCTQMSW/T7Vr7KdDevyE3J+KZLH8kuqB+Rcu6a
Tf9665YvKrV5htR5tOJ4R2Tr5KAlCrls4ZpZEnXnj+kp7Qu9oDRibChmh9wYWKTOn9WDxjSth4fQ
RCxrrWiNhAmTDoJTaX/sylwt8zh4zU+vHVDqPL6GA2xgtKXYltSRLdhrGuVguoeOm2wVm5kvJ3uR
jNHcDSTg5inQkfpg3Ylc8+uq698XGuILYfBnFFJxFBQqO3HKgRAWBg0ZKhozRLOUvXWUEiiQBqAH
vZFFJt11P1wbs2OzocQW522Q4HDwf2R1l5fwfgqH+28UqFz8/CUNsjfDP2QGDcW3pgOBdXN5QuQw
0tcNeiCPZolIUQsmDesIOCBcBlW/6ZKPjYv81/s/a0WVbhPvv4k6CJv1MO8RkCVBJNY0xY7+fTMF
bppld+vtz2TrfIe4+RqpF6LbggHyolRqQqzfsS6hCOzyOGS3pRvOnbkS9dJtx4pOggsMwrMoQyZp
M4v1nSDuV9sVn1Sp/wQR0qTn6eVLGUWz+Idi8Fewf+WLwCy6qNpet5WUtK59bSsGZ8TXLn4sN1s0
C1GMprFTQApDxLFQ7Y/P9qNOOTCJqz9Wwtxo6YC0rzLLJmWPJ28az5qtIoYyQEg3QoVHzdqoOhQw
o5qEC/k4Bv5YjekVSj26mFhEUdO6SESqiyDXZkUUQNwHkq6KbbbE+bZIAYeCRU+fTN9QCELhxR+u
oWcvcRpYIM7pSbpTZYWoLThqss+sGAlRc11/phtkurokiDWQ+tkqNeVJ/tK4OWnR0bRBOUiriQeL
BFY3fabSwOqjn9fgu8yUBdeEmvFgMjqJ2vNrezvBzDOKhnzARr9DRd9rImmVsogl/ek3KVqZZprE
7iJFKwxUFuZ5/gUomLjT/wnw0TVeQ4duZP7P9Am4//b5JG8CPPlY/eXevQH9jrbvL7Nlj1zXocjj
08gUV8UvECxR3sOa0usPVEufDTQdkScFAX7tTlCHp9gUv4AYK7U6vwlqhzSdCQcoQSvUNgoSQxsb
tOwNHmvf38ucf3yXv85wxIUMnjOS5ZuzaUmifDRVHxzKL5LkJpUP8jSHZUEaHq0OqNsQgauEFtBG
TXQb0uXZEyGDBaC2iZ1fG/mciwXKu/1wQdjBSghSSDISz52I7Se/R5t5znWiu85XCrC5d9sOMZ7L
2y8C50VhVjpFZM0r0GdGGcp499KoRTWbO/MYPIdf/zyBjyr1lHhPczMU+mh1pJ//c91BT2PGbKOJ
WzUtoDvSSVw8YS9iYuSi6SvvkbtEPrXoxqIhBDHH8FB+Ag5oc9i/rAjD+GLuaUzwDebWN+73KcBx
xFgxMW/zXjS0P0LLQgJjDVAtbPhZjwhgE3k3pRCRPpLfRaflowy0BN06VVVjrFZH5yaUJBcW5X2E
drtMfZ8Onxpt9DpgsbC4M4v3GuGM2KgxeZ+1Apih0H9/s6g/+wcdkcxNQ8M/W6ObrUj4FrID5QlC
C+JoRK4rPFahfSppYQtSwaGgQBnLOaoLDVVgLdtqICdNC6CM0XhbZQu2plJlWErZznA2/0EZC5/z
ZqM/S3WdU8MoeBFK3JKlRZCFec8S59Kw7hlL0tAt2ATR2KehqtVctV+2i2ylzJQn7GP8o7yE1s0M
4wHxLFYMs/vbYmVxAsRlShQeaylKU3swhqrJg62vglpjjD2kO9f22f7ZDj88WpFJir8QgdNV1JlZ
wYkbiDIVr7REqcfVZQUah3cMDANGekAulWC4N3XB5b7v0U1hJs9cLd2MiQ5EXP9H+93kfoCk27l7
cWssHPw9EHTHTYyB7CqURCoWKpzl8RBS5+tEjpedMY10lMDX8LnkL22U0EDeP//dL/nRSF/ea6D1
wZ5VCdg2wwvFTMr1r03TmHQbCjCR7VwroPkjTPdnvYtWi55+elImbv/E6cSrGNumPAzBfF1v1OqK
TzL0JaCEezZEwO4G1fKgo7FQsBJv+xIWA5G3VCB9S/uEEixqdBh0JW0a/mrGjBzRNFkaRs9x66RR
2mQFJzHYTelpBj5E6eoK8J1Wu88q1Sh/gL/LtQs8SQjrz5sjPv8l+hgyPME1GGgFmdcJFjVYRK3U
2JQJXg8qZi4pyy8JR/te2JNg+fvchtSQpioCdMWBNh/l8RBIm/n8iqksnxhkYaInLk6xyhnJDuqC
RuZ/gDxJg4b91RPXhxtUqjIF7iS9ZLFDuAZTzjsB1nM7w+ErCE518JhiZkJq2AGFRwvPanV6ADpb
m13faakQKxcwVZs2EsCWwDLqqhbZA+8Rv+cHwGua+RoDGXo1moydWQ4fQC/Inv3pm0KA+7yj6sE6
W1QOyI9QBuGojrIZuPq40e3hnSz5Zh3zoKDYhe4rqoBXk1DUvNv3h1m/9srSnbJZjgQOV0Gd/xux
m4gas9Db/n11D4RhHP+ma76IIQdkbqxHj5tu6/S5vWZK7RKTuT+TIFvG8fzkJvjVLEwg7sqPsjKj
MVynkZU9NZx79pdwVaNNaUsTrImhYRVZsoHBwVu4+DMuiefwAIxTPp/u44CQyCk7gcbpVNafjEPf
sV89wQJJuQc5BQ8Ssl9SArJiUZR+7QnXROF0Humk72ktXJ3mxIzHh8U/3nyDurHfSNiZ2fhG4bsA
Kv4yhmCTYx087/Km+xWgxMuHvvXG89ha32cZeaEUpXlPAzhlXzaXLekBnKmfE0bvLn7BYB9nH3sw
6htJtoC7zIqr0SZV/4YfEu4hOc/MAJBQHeiQVMjZ3qdpoXcqM7ix7rV/0jR2ZJW9vRxfLOv8yzog
V6mOKHsXsVOQ2gfVTYNhu5Mmg7chM3nZIsXlDFE5kZa8jyaQHy9sk99KZXTuPECC/BWYL+nI5JZe
pfeYm2smgy9aV5vcp7lTWV1E7fkR6+p3WoK2I9toxDkwwILdoiHuuFg4R+Cx7mIBAH3cEsJBrjma
mc0i8Nv34rl+yIc4bEGisG0Zda66EJXxQuSYto5/+fBugzU//vQTvSXotT6GAmrFCWIhRi/W9JME
f9uivtu7WL61C+r9V5Ow6zpkCGIQF4XTwf9ujgrNWi63ypwaABEYYeOkB7b/vxZS3UQlIkbFpRa5
s7hT2A8Y6DdEYDW/+7ZcABPl4c9Nk7WK6DfjGsP5hFZvwdTi8B1be6aKnjt5R73VfcM9CwI6r8CZ
S1gupcm5pO9SNcbyi5zDgf13RPq+jX3JDHBi669ebJLEKSjgBTUVFSPgiKSdoA1NFJyBk/DCQRna
3v2Jgamp2IveEkzxh+P9cDiDK98FSEm/LvDZBX8cOWuOhICD9jv85TVS39A0sM/Nfi/39PI9pjTa
sw7VdDTP80z60+RXEp+VttLjNY7wZoOy/sdYQ6Q8eUYjmIRuGPlV2WIKN+t2trQuhl5oqdMtJxUj
Boi4bnX2Mi2rI9Mxt/nFRVdHtX2R776tiRJVP9VaIQkwfwoWlz36jaB3ejxVLpjDbKCIt+H/jHPf
K4oejSTIGsio8omu18FTr3LZgOjbt6FJmjo8t0PWfl4WdIJU1tw/+sO0iwVPL7jT4K8/oVOG8mgD
5F8nEDEwuBhS2pXGHTyWMDfgHYm+hl/wS5jXn0VfwPVKtRdBep7vTOD/JSsUHvDs2OYWOYf1DbcQ
9i+e8BNF1wh1ISBZ/e+3/F3zzSlZO0CS00qOYuRXl+JwCwh7S4Af2RDfApDWR6v12Q0KlJekIOgR
LyPirs5u3TkRRJuUqzUks7JMV0s5ioF9R9VcmvtsUh26f6Taq07/MoyTkWkB8rbHDxkdh69FBWJH
slWUwx60r4TP8C1YGVDflmgJ7yBqELkOpMxxVt/t0lke2mw3JXh5gcRGqIBcEG7KsrgCMSnjr5+P
tths1GtZ4lt3N9FbuP4MdsmEDgaL2D1haDLItJCCg42qiee/sBZPvgmBtC+bN0d7fW+3AeK5Rcsg
Zx/hUKVJIcXRchxliZrZ7rk3caGjZ92Mqk4t7AJwS6iNU8WxWIPd+l/oeVL9rTjfIksAVQviDL1A
9rviQKi69jM10Nv4HuRPWbQHk+3OV4cfVLP/lW5PwrrUZSiz1q2iAO7DftWWefcjoz8SaOa0/YOL
xdXy1GWXp0H2+mUMrrWJFf5iVM49hj4++6H6fyPlDkwhggqRA8eblc+VdoFD36HoU/lXGlqxp0RT
qojLvY+44hBZ0M8ypzntZKtCWHqTo3YwtiFvrau4b+8AL+V0y9utRkhZo/g4ZzrhsRh7LkwHoyxP
py6NS4+Ripr62xSqhpW2J0ARkEJpiRSDEgrc+Bt+rqQAKs+4WYf3mBm075ec/hqjT3XaESmc7eb4
XAxWIKfBm3XoPCaxSUnBPhUZ8BBBs+ulwod/uYTJWnrQoaR+bNALIjDlhxvRlowMXvIdfvwtSiNC
w9VY8pDkQ+XOHAw15QHdh4iBz4ujtlEax4R0CLPqXcj7Er9cldOy6vVAXUQoCnX63XuvoZirQgfJ
4e0ez2pGHUYn1XjrTi5BJd0ekDzRzNXu6leitvRyZkXPgHVS0D2BPwRpZlkwacn0s9ZCtcxgt20L
Qw/R300DPb/mZ4Qm8Kul/rE8uKSzueWY0/IvkS7S8V5AJ8UuWa59dWo1sNecb5U6JgvR69sQ98Zg
DHxRTTaRLUXcqn4e8hvhvpxeNsvpUcNvkJHxR97h1ZidtrIk2QVZmJkZDwU+PrPuQisOQoJ2P5J+
qqZoSTeIjfdylQsgPBWi7XgFE44HZrklgnhOg4+lVIGDXoWL9zvwBh0Js7dGXnMwiAwkpPs+Ocls
i0tREwJDBzosT5jSn9yIm/e07Mne8CQf+dPtRKRSgplUOxu7F8UaeX2utWt2sc5bcXCCBFv12QyY
cLcstShfKlOCGjtP6zNsae+3PGGJdKzwCLs1MSVzkpJqQcR8Yk87xKBpD6bXrAzp3resY4hDx2UT
/Ze/mFVLGSyPThWqDUrCek0IGwaBpTRPI7v2R7nMSCdYK2ZhKIfba+C6FLXe38wF9CtM1YF6YWYV
SoTG6NHrpvWJ48+6k9n8GkWey2TaE8IKY/y1Lw5DlgzV1t2afYg8guCJC1loqyEVzjLXooVAcdVV
ZqXZMQKoLSn7tv3j14aiIbVYvnfAu9P6IFyxAUOmdZqi/UxQbIVuS0qe1GCKZwSpjbgvxeEuqhf6
WvKsevra3GhcuGqHg6skSZ09wZflRhrQJrAWcJyHMUZIgyEgPWJNsgy99iPb1264rrMXm1Fgicxr
V6CxsjjPCgF/rBCO3sOTQhspb74dPFsdr1wKQS6nQUJTeLEXmjl8HylBark1iTXyq92LxeaFtf3x
YPv4pzhcwrqVxj8sT5l8XiK8zLF+QR0gpmhezU/Sopj4VlhCeh4SpTfTolQeXIoQ5lDC4V5Gk8NS
obNiydn3uvLgkFuEid3l4bNqPqLT4UEY4XX0qyy2siPgeiVoHYKOZ6FEJczLuWQXBaXyitmrX6ap
JnyD7I7MGZIvTiktB23O+dxI46V2psC/kaGRMmmPsf/wx+U4akPze/qNmib7fw6gERDg6Q94LQZi
MuvLqT8n+JNUqiod3Ek6etYDduCW0i5mnTqbxubFw9Lh5Yzkb884FkXbyUbw0NeirSJPJsvmneh+
U2jtR/cqSYx2px9Adtp9dgNkdFXxRg1bymcGQ2hG1P+EeP10QEONJa9ZEHfz9zwjLeoHvAAMs6SI
Zbo3uLZzRCwSKneR7RXySbAFaCX0HPg2yIAEKSQ9ypn5Qig24fzHg8P3SqjiEpmAvbm0HkKNDALT
Nw/TmPqOLk+CcYTdF0Dn6xfRLOonjrOie4SQfA3+5MZPxzNFalzL2oungo71zGVjDT449v9CsTd/
nB0IHjJ2okjuFdMsje4+B7Fj137B3cWl5ofAceRqVOIz55O8NS+TNGk7gA4MYIHmFYOiXeV/iq72
rV9bCtpA/WB/60+nLJ7hcxEJ9F9hYvxZGHY1acyiC48uOU3j7a/EuvfAsMPk3sJ9ksIolrXdRhJG
jo8rcTz0vbCAJ23Boc3VuYJfn0JZpzds3mz504CX/SjKtchY2TQDawLRjNfpMRIjjzgVK7PAPzp7
nfDTOA7plZkiNea1ac8UWMlJYAs28LDVnE94s+bS59Tt8/shsMlgURe/ETQ9RlqBaz0Ee3LQRjUK
qdrBaJuppxhb36zuSYMnGyIHDnj6UJyyyfTWn7UuXBBnyyoX66DyTFyz3nYx4ZBqzTPNNChc91Ji
GnwCgcJ5bUaHg0pSziePX1lHhHm4/VLydOzrIa27fwCUYzV7TRKHL+qPY8vLBmTRmwc+cQEaWRch
4qSlswUih/V68C0BRhPgzjXNqV9oKFarc5A3v5MIGeNQW2ptlEOCgBSazx5uEgXGvAuAdfDPeZQw
w3sZzqCZrgMiZtTzGyTTWhQj48xX35cnUcDGxmHO+M4p4hhOSFW/f3+nhjQfWgkbBe7tfbRrozqr
fgW10ljoOzjomKIQRp//In0kw3D3gWJKXBygCNgrB5Jjl4e1lCsIsy0Xeg3/Tzm7u1TwtUWEQFAN
t/B/TbJeb8pSPdUP6wVinIDQI8qX1UNr57DEBZZr/oTgnrQH8aPHVt9qDuEk8JL2lzr1a824m3WL
kExZu1j/c69nFMP2e82TyAMXXZfAzYkhL0Hwf1Hp/cMIo2ZmS3R57Dns3aPFGlOugEgnoAEMAIx0
QG0BcwFfZtD9lv5MnTYMdTaAUt/OjzE48q1k2/MYW7rEPXXPV+aKwjq1xf9Q5gYA7TyPAZlMmcpc
z6qf8g35OEeJa1kswNPvv/J/KKwOxY4OpFf0SS6+KtJEvaQPqesABNMXv6qIrYVU/17s/RGJ4lu5
PyraoJpeWNYYzcXNhhU/wJyuMAezGT3boOamb7xlj7V3S9WX/1d8jBTJ0kTGhM/lX3x7H3wxICUZ
4FJOnApHG5wgaONFZG2tt/wyaCevrfL/e8VsXDFBMWh9kamgKJpLx//1F0juBG0SpG3qQYG0H4k2
xy+UV+rd6oJfssERAAK6e0E6qdEmaF2jiVl78cvHhO2W3rT1c5XfKeSEVAWCYjfQGGBSwZ/E+7ki
0xIWonMsbskaKgh/bItjEUBNfYXgzh+UWyFb8iyPgx1KyGHQPcVo++pTF1Jep9Z0oJV4RI8ETon5
GJlzbi+RLBqT75bgU3bAFkIK8h75rlvkMqatX3xUkNrOWG1sVGsW+hdz71XdDpH8Mib+D5yM/eZo
uyKsj3JPsUuG0c3iTy2IFOiDV1H6qmkS+y1Jxt4wKoSMmpVAR9xQAE/JaTQ6gkYCSORn6mVGD8I/
xnFRekdv3bEe3+VFYNUm5p+pYarMC4np66iyStXOth7ofxmWa2AZi7rOUWZRpHC5yUDAEYoz+YxN
ulqvRgD1IjPs9hFtyVU8AdVjCG3fzBJ0qKgoz1xgGYl29XYJMAz5QlvVHpvlEg3weKXWLbaNb+oy
Q5aOwcOEIGhJGL3+HavPU59osWpeXH39QyFwSvsR6i1ewOrTnF/iqEGPZEa7D8mo6iGiExRJnOjy
2+G6jzw/sNTjhT2P7TJmSVq4aV6MHYsEQz/SDbPZ94WfhGFf+Ye+w9TSeXBaJQy53suBDdmp1g0n
bR+rl23k5e8WGStFfDHQRNS7PjRsh8gA0UEVQvIb6LVOtKyHEpkkjrEjBKilYkapE828oZFyVqKp
r/36biPywcNd6P1wS51dtoUPbQxwERLj+OrYlYXBcVpq+0Zpb4EKHlHrk6ISGrY+Ibmh7nw1xij3
DnoO8A2WE4o0uBfByQ+h5Kg3I+6+39edqkbYKxIAd50pSSdpRmO18OBVELtGgAlpURTnJ3xkSG1C
ccQZP2za8yJQ3dmVI13DCqtDCvgt3TFjKzbCl2n0MocHm7eQoLXOrUdGZjrzci57kQuWe1qlT2Vx
EOtvg99iAcTnPCvpzrq8WVGxOQ6pf4YXJ4HeB80oElHxWoluSsuPGIOWcBJUKnzUoTnv+IasBWMH
VYj6CfxmK4TrKtgkdLdhE6dNhh65QrHCQYHHBGOz3qzQGpb2zg72oFULIjgHq41A572x7NQs4uuP
M2xYoyoIKsU2M04Et+npn76rKlcJxJIlqb21lvaAcrEeQWCgzbsk+ic9M/SiT2r+E71l/MX2sXtl
qwiQQpHrgHukqHHcLL8anoLv9JkE/xBTQ2Ma93j0+ldgWBR4dWn1EX7UiwP1TQn9T0QCFrwS9sCl
6VyyGXBp5geJHMNiSwPnHVhfmlzYvtzTGSyzZIn+OuL0PrXR9DRoJ1K7rKtdT7KwS6aFv8roLy7G
3AsRCwdQAbeedWh7yO59rjYVumDaKoiRVth/rEqsmr//uaKr0JGzE7P2JvZxm/8UQJyZjE6G9hvl
jsiVEaJaSGRpvBIFV3IrAAGqvxyR+ALbUXh4jeF9pTtwVV3P0bQEhvNplDGTaFylJTLFqC1yANCd
Qs8ImnJwJ1YqQEKmazlVkhRPnj3F9teoF/o9lQEOC/GfXOaqru6U7iPJTh5Uo7qn4EsMAqcQ1/nv
R/UlQ8Ratq3z65SmbZCVLHl0yL7eJcNCTIF1ZiT/dLMgG8jbSAVrYD6rVK4bw3beUU7koEUEtDNQ
fjXdvlkcmQtR/mTwzcdS0uls0AthPNN7Sg2Eb1VVgNMDPLG3n/7B9kJeVIFaFxIb3Q9YvlVeC2Tc
iQ0gsD34LYXJCfBEs7Ewj73GPPi+SC7FVPe5LnA4i3FNCrAgG+ZHfU+4DEA5hOW7EKE6MRRAQ6FZ
szltY41u/NSykEnsgB1S606t9lziagzajDLguIBatrySoIqah0INdRGQn+63YQca7/BLyGZBxxpw
+IiIoNUq8U3ViNv0SAGsX/yhgWklYfS0GhfSRQE13wZgsX9S/FKNNKJJ6odpQNBBnXhGhCzHRH4r
KdoDHrso5rhxrNNVFZu0LpsJrtLRa1okAF1/X3Jl+WPugz2/LSBQGCBy3znRh9Vr3b0cwoQfPmbl
cIsbC8KZxltmaQTDA25Xbcmw7fM8NM9jrAr4gXzu5EjEq/KmHooJeVO0WmAa8r8KP8u5071DuKaA
nJ0lw4EQbwi1H5UiewZfQ9hUYufeOSeqlX0h4WQfvHjR4xnV0GFLzvt+nprfWNUshH8S5kZf3Dxh
Y7GnRSPZf5GVmB1Dlpif69fc2yrkPXCZRRQ1P9P6BE8c0xyMuFXvpJHFmkovG+HqySvuXntNx2wl
OTnT46tvh2YqJ3KrsZdcGa/FOSXMNqZG/f4JPd7T/amnu+3am8FlLmM9Pf2WoyLPo50n0MxFMTeQ
SBFjYGeOlO+hCWH8MszKwJqfTjWR8M2iYhZ2Mge291mN0zse2d8/eePEABHtIT+uy0w7I3vin4ib
AQ4Io9Abpf3gRHrhXLRb0U83FbXmctXFF9OZz5pxrtKWvJW7q40O+1GU+C8g4134hBaOZy/6O7Y3
OetRtTT9IpGRwgF1ZBpZGhnBxh8Jc79nIi+BriOMPGzMoFti4W0io69G2NLPw8QfhvRgmSeVHuxl
cfU7JJZ2yGNM8Uvxx+i8ndvqcEYCGUo/AjuCoXTZmsiykyUbx86P1iiRuiU/QtTB8Vq0u6E0EQL3
ntzs/+YltDIz5JAKSEiK4R1Dz2j2+5XflsALdo/QSvr/CAtNsmwcEToV3cUUjoIimQr1NqM3mGN9
Y3R9ACpbSHVhTpc5KCy86LzM336d107xJWHvy68moFvMbzwksUIKbIB7f50w5Nh3sCT0o6+yMntC
o75WG0nYQ8U/zzQ7DH6lptW/D7n2wZ1NWwL9uvBf9xo16M8VVOOgs8HiGHJDRSbOkImKWHuL2tUK
uhMftPWUKGGI+N+Qi2z1fTszcC27KQmQh7A0jqLzlF7B+vvVOC1iFGlLOj9zMP+mzN6aM1bc62Iq
8ypKC6o10RIeIKhluwpZzRsd6IieCpldLgw0mTlqROcJAaTcMnhWjhD0fE7xzdUtrQgQ5hcK/tHN
5KlW9in48GESIxztZRnEgsK/HjTV/L8OomSosaF30NMvkrZVZa1m6Q9ZRc8Rba2QTw+gBjkczx1J
2T4MICll81idflGeUN1F77SEuszbZDQVvCJHIuQFY0dM8zZ5T9KHruIN8qqmOP5UjP+LhF/bqAyx
+0iP4IcOf8UDzyR4z0I8jd4bh8+UTgjmWA0ZQKekP8SxOu2Vt1cVQApRNmxx+l3J3Fas/fS6D9t0
AzO6WH6Uw3pbpJqrSeR8p6MMzRHgFw2u2NoQP9bpGE2Mek1y+k2sFwhTXy2eFm/cMJtH3tHyHDpL
UNGlIjTRSy0n+X9Z6gHcY8qNnNbcVTzIIczDvJnksbuRQNYsRxkvqw6ah1Ahi5KTGJZT3qozEb9z
ZCW78IMbhc2bKVA4QSSuZqaBoNIEKRN5ur+KBYQZ5NT6y2NPSKy/b/qdNeXb5MPWnGuz0GO679YQ
1sJD4gCCB82MxzvY3hrL6XPiF6qYqdimIMjBDj9oCOJdoc6jlMiLq8jyvnKz8lvwc7euchMR+Qg6
OKNPJLQ4DgoVUQurm6i3RLwLz8WM6HBlqC8ixK8mvXRyY/XLOH1ugK9cBI3keSOmi1aNTIVJxWUt
mh3jBSCRvYpOXPRniHNRKBicxoMlxjgpy/QdnJjMbwnkFk6AArKTiS1TFixtKJtrnzikuFosnu0n
dZFDnIg2ulmi8ZN0nwq91Y19+NpWYw1ztTJ1+pcSZMYhJ/XesTDNwd16Hk1GAwJ/5UqgG1slBnUv
zUUyNXQzQ53CYYGSbW5ROE/HOrvR0rKBr5vhRIBH2qCdV3Sy0PI1FWJF07SYmdMXL7jsGQIeCJRV
xbDk4qwrkHA3OzUpdL1h05brYgoBELcLY4PuW+bJxcYMIL12sFdUG5FQxm1+8MtJg3ErHzAZkp0x
P7EyxzWQ77+P7zdffXr+Rh+sU8a3zl9MZDYYa2hspVmLA1gl7fG6twnId1RgWQSvCU/PkoLpKrm9
L5Uh23DhF0lZ17OqzNBbQgnz3yXsEXCIT770+uKx/uesRX2vACrVMsy3ONTZju+qNkclBf3nDqUk
4EID2YzUp9vHty+8b83XWRpxXTkRDqLEAaxlUTW8KTogv7y2c7QFBjC4rUkxEmvM5Mo7bRUU94X/
sR2WNhXb3wDzjjMWvS8nsMDuzIZcNr18eqBj2/U+ZgtkQubbEHpDzuA39DsLB8Qz/Y0uBEHEtYIf
ZiZbCxs16O1goCPaAW3zlZZ2WJk4obfevOY1VeoHNP4P9rPRULKHy1gDnBcszT6xWqO7ucWzOM5V
9rPs35LtlyK4YI29ScW3Ml2dhEb0uBtbQ3Iapg0jdLTaPcLNqhCvr5vODBKQo4DYfalnJn1Z0LIy
Uz8meFzZVsXj1G7rOx4fWjHKT/l2YIFyPmXlVwU698xHjEDK625k84roBGM0wslcnr1hVEKhIaBx
z9DL1PpNDOIwUjO5EfZoyU8VAmUzsNIdNIe+F3SRiir9MtYJ2OrUdCzI1CiUvRmIOOUWPW7hqhxW
7LqQt1Ast3ZkFFpaRphhKRCIE1Q/56uhE02MWaUM0mhuz8HSea6PzbWh6siQJEP8R7K+dkjhrYZZ
XDVpDeW/6btVxDv6ZfEXbZv9+kTpDRWsO4YXH2gP92P/ArJVi0y5x7+cAIHZORJa90YRAkQwBKNp
kK8TvCmkO7KX3Sa2UEpf4VK3s7dgxqGTk+o0RLucXGWVedt/XD1bCNoL1fHKRds0i63YxJpXMelg
LwkcqPO770DDCrmvlNw/LZiPHl8tGeL0BasRY7zGJAdLySuP7Yu2W+6WQP/ffVbyaWALNfa6eLfc
PvNA2rK4QwVkij4AOdfvkbXJ9Cw/n75Q50PlgLCeKs471+qvLlUWzU/FcBhiTPUYmaYcb6O4UAPC
fTr6J+P+fs84TEgq6/6Vqx1YM/ZEBaEHlNQ7CzMvdTr1XCyY+sH7OwLONuW/Qb14rShFAqmPxrbT
2BuVnxxRLNW9826xx8rRSLjNw6H1dkAW7rkkwgptLDJfSlMLG5sT6mgjokdGERy8sASWmJ9RpYOI
LGARes+TtrwIYxX63LBreAMX6QRNV2eVM3Izlvy7OWnkuWB4NOUI5x4nFAnqJ2kE5J7GyCoTbMBa
gaO0u0bwKELtJIBdp7G0UxlzMyIEoAQV4K+pF0VNSovShpyE5WiiaybVdirI1/nb6PXlkQvoz544
kJ0xOQHeKs1SXGRHFptuga53IarmTrNUJvvD4Kd5pqjQFRgTGyD5sEf88Wur+QmDAMU9vltRcL5E
KIv6Z5txBADOcG2HJ8D0+l9XMApGZRptJQghgOiQSCz3wSwo8RcxV7h2RiD4bQAnoYWwGDoo0Srl
O/15WKG/Lv/qpSog3a+UcXmRWyJBFaob3z/LqiJee6YrjgDo9AOlkB8OO/F/gIyDVciqvZaNRB11
ZxwjB3Z7upXaipgr5+Qx3oGTyTSHgGlFj5EtneSgOLZp6E7hzy7tzt0DWuCxKriMouM7C+1CrEvu
SmC/A/InDsn87p4QqsZ6gy8Z7aC+yPgin2qYF8DUQiGFmKUb1+4msMfdiQZ+lpeLW7uPcYLq13kZ
g2cDMh55uLNazt0E4exe8F+CScpbaAZr3jf0ix7KQdEQzo9/IWxDA/x2nAD9TUUKRjmYLa3/9CLF
NoOhQe57aMSUj+3aQ/lQ6MP5C1nRZeAEBNATAxSF8LEcxIF2PXuFljTIFyENSYrQwiRetsn93V7G
8PoHwaeOLfaTeCdkBQrCYH5buFvL3NK7gVVXM2Br1godaZoRvb/vw7/7t+ViYTTvl8wJHEU7sdYz
S6iwXLbHxj51jvYjBHcTXIEQZMjqmuvfT8pxj4ctE2HwUfFvhEogjbPfjJIXHR+hbu0UtC/442z0
Fe5YFQ/5JGFskLEB5bz5lVYrUFWA4bh8Gn+NFRs0BU9h3vt7ghMSvLEiwYBxKojNofGS3uDlXlGd
9Ki9RBBoMWQxQvsSgKiogCm8WHKbLQ59F+wxEtkzmU1RHuwlFjEVVpGgG4NYYGT/whKj/Vzv4anP
ZpDbhejFQFd4JNeybf0aKuGtyp6UoEtj5nv5UaLWbV72kvRrs+XOGOhI2axQT7zvmDANg0vzZZOv
xvqxontzfA2A+nxiTlIVyKq1KLeZgtMiqNKhrPY72mnldXD6kzYhP3d6zgYxbS63jD7Ag/6HAA1m
AxpUAMklNNLqJ4yMGMGKKpx8UixPgHn7nkA2gD88TsxZv6Bykw9dVP05jhoWSD3YzLgl0NHGdEpN
2cf2RFzC0L9XE2IAqPPNKPQC6D7U3XlK0edIeqN4hhN0UIi/UDWFUx8EoTjTBcUb608fTjWG1/2b
47AMo5XVFEXjHKjP0zElWcyyIDnzXPRYwWyP259Qz++VnlyRFf6yiCOa8skffPSpX+9GbOfjiq+H
nnM2ybjNGl7wjtQ7UBaBuNd4CH+VzWSH7ynY+XeRc0T7rm1zz+Bv/o5+a9fs+4KxniHAuIEOwVbk
bf+T86o7vWJrzHFDsSWnUkz05eYny/LrMYiKMmfTikDPov7LDv0VIdPVysjZzzrYj+8cAez6zzSx
IHp81oHlguxU7kjQa8JJPE+VhdpHLDN8llqlkDC0CnmkmQjYYiD5nAV/i2+o9IgVcZYLLDKiExZo
xKNElv2EGzFoeuTbvhDoMu022KAs6OJ4DY1uEYXggkVSGKFbDLxxncVGCk9SOOrnGSDa8uXxjiWA
9pz/5vqzUhjCul4Qh+ghk6JYflyYMkNCdHufnYcLORa2EfzypI6uLutBiYCDYETFwbHyQ+OOvfmS
YzDDLWTzYHBcp6UOXBb6JsKHS/H2Aor1ppBe3+GCqVsccZtvHxGlQhbg3gUZO5cKp/o/D5JNP5+N
yuMq4nPR3B98t5Cb812Ak/1Vjtph0kZZnCJxsYQCpi+cfxZ91wFpKZr7nZmsRFm4ew1olS9W4331
cLG8NF6LOnxg/J0TPQVg4rTpP7oMnj9IcQYf+PAINO1kXCDJXzEzAjlD8PLz6MdAZqbls6aX1QFA
jEnBsRawxsZfKJhD/8Bf4f9Lr71fHVH7vbmq1Pgyy4bdMqwPv7Du4q5Fb8nLWidjolQBB1d9rEjG
LPRLrun02du/GAJ5xD/pKwch0E1NY18aVx3Hiir6x5HizAbLZAV4mcNiVc/KqR43tUqpQoSWPY5I
qcIgOBwYoblWrbqu0InwHmMJXSxxygeuQP2ichk11Z3Y45U4urVOckl3jc0BBs4kpZl9EpDfK+W7
gqdjXMlgzNJNZAFQtr6wTC7lQsl1jE6HNKvAQJpwyMkKu3p56r/Id0YS/HvresFb+5CiObtyQsIA
BdtQCr70DGWcPSLatW5UTJyxheC79dDI+GPBe7pjBCMl4KXmTyzyskr0Q0OtijUwSSqowm44q1+h
7Ln+fX5kopUXJ+M2ywJoInaSjeA1aovKSfsMynDqas4pdNdrYKlSoyioAQJN3Krduu18tg1CKghd
4tDD9Yp5W9QqLK5cBken+PyN51cfkY8gnmA+L4NUtAhVJlIKXBwAnuvVcsF7CRjkpexeIrVCGd+X
Td6LNOBxPUfkoQZ5uTaRExeMrC00SrIuMvJiAFsafDL8m963PmL87dLSDkEK+D1lnioGrHHxxDKO
zXOFdg2n8PRgoPxomiCRb3TnG0XvgwZTrPJt2ZL70UmXgk+y2WDKtxPTT/qrEh/EClYyUrNRZGTy
JlP5xAnM4wYlZXUMysvVsyCuf/NiNuJlqKHb3hcxQSaIvqwh+Nn9d92aonaPWuaRbmKuPhcMCTkm
CL+qYkJmZ/1edkHqk15GF6Tz4DZsjKCp5BmHdGzk4rAZzZzg48n3NM/NsJZq8Wv4atin8nN3CqC7
4FnXQGu0syZDDPNH8IKh8NhXJuuOt1la3bxaFQ1LKrclfnRTHoPjVP2+u+etUrBdRHueTFaWcCij
HDEf4Ob39lDagLHy1h+RukLvcyMtM/IN9xi/ClZdN84i55/az74wrKEeZ1lQ2MrxhcwBm7dokETW
7IAuh5lkSAuc56k2v8247894x8AFVxi5ENjsYO5GSy4oSeZxEjrVE7nSIObeZY1vwmAFKIz8o1Ri
BLnEG7GIbxaB+RzEO5AmGif790aBoXc0O7qb7kq58Y6V4YnE3fwpysi3/iOY3KTAK/O013P/Fj07
B6tiEcui2noRHQ/uMDCVvOotkda07HBUABQuHJQ3jqjnLaSVPRHp8AYul/xleArVKXZ2/fZ1dDhF
ATpsgAeuH5f0mJBB6yc9puq2fNtkMVGYgtOdet2LgUo2++IU0IajjCgANIu11soi4ICx0MwS6ReX
Aah/NowmqBmJQf8/Hhyg0cyDizYEi81ucc13jepweRepLN5R+ySsO/LPH95UkNvuSli25vqiQ9Jp
6nbu5erhf2kA1VW3SAwdpzpuI+yZ4jyjF19yHcWpLN3szcsrZhbvY8lwIoSXa9QHf/F8azZsFL3O
oEYVWFNhCu5s1ZN7L5t64AdZ5QSu9ko59a8hamTM5aZD47tpiaH4PWLY0bpUzVvA1frpSa4gKkaG
9sLlsOz0UyWY86B+sbyr7KmqJgcy5YY76lSBxicUbTmhqPMosXNP7SdYaj2aYaALBxlnafwGUrqg
AC3vAgvzd/yqCOXgST3SPJKZJyo6M026bUZYhbADkUsqvjeSAGph1U8/Ll55GORGZONcQH82X0mz
brnHZ7ngYcnB8EGiKHFP4pCHTjixYYZaJDB3RYaxAQKQzFIPvW7RhLyOvF40ci/5118EbdSWDH1x
qduhXTxxXqOoyg/Jnq9wcGrBEZ6UlpYBrgLYRNXHtDAFXubLQS56zpg4MGlqFtRtmFPd4dTsXoc/
CRq7lZou3WbOw/eEGIgSObE6mCghySHr0ANqHWPQeAOqv8zVqS6KA9Vw6TjTtQLoVSSRrF1In1To
CWLxRNB5+0R6rjAPW2lmeugFqyM5z9ncnI62HcWc+QCTaWgGNMzIC5TSbr4McIziSpMBJaCWB1I+
/YTGDRVaZrni7RtU6OdrcXCwONC4ldpgcIU6U6ljYCq6fhcWgppJJJamRfWP4tcLYszzdwynGJM6
J+FZdSfQSwG4DNvjNbctuFmGUxltKODoFg0/7J56mdUU0mR6tgUtbFf8mbNSKk6E0spP91KB2iRy
z1eND+1XBy2q3T1gdpGWg/8AiONUCgW8UDu8S/aGecpiy0MK4phxFm/6nhiLzqc1njV24MjEadWj
eU61EZ2ZSEnlrZRc+Z791m13QlP87WWBXvHLjcu54WR35idSpzRabm3M+MQ1RLSHMa0fyxKKSxaB
m6uejZYZ+uoUkSebKF4o4OZLCAAttHuqqG+jTdrFdNjbtDFwjQHwHANxGbmHk58RQCMqkY0/EDIr
mEvjFwpbFavxlOMpg8iOn7zyeV5sBIPY3iqCmoLc332yF4dvLulW+T/VeZOa1c7r2aKTiNZx3BG5
Wl3kc/VdmR5vG79xEfiVIjMr4KOjYuONh4mc/JXuFEseSxgUhI42p09Hnx+4reljcn2GXIONIL1g
UVO8tm8cTMK9dwRVxzCj87msp3GS+Z6tc5w0G5Cy+4QyJKRG6jdVdIP6BAVZp2yFcxvcbasVANyH
Ng+j2lAUeti5ZYJO/vGn7PHKJ5HBvpvmaY0ENzZ9soJttCqJibg4gSpXJStklNGVX0cBMxo2EHqY
Jo2uT4u9nekuPFd4+aBg0lo9PrdUCCuzPR3PWJHsf1wmpJwnqX9NqHJZ+TExRAaEj9z2MEb3vNuV
HHLUxNskLe8quU3OPLsbLcfd0Y8penBAiXnqeUn655/WW4PHq3G3xjMQtH1ukb5u7MqkWDuyzQ7n
izRPAgenrtqka4dTtRUN8/an92Y+N/B3rO1mfrENizajoSARYovG5d8bocFvlXT4UCYBMQt0ykcK
5r9YKlfFRrOitNevSRC12rs/J+bfiO3mX6/oD3G6c2/kcp0N174qHNKuqCWZxsc8ZZKwwFotruqr
BKqVfHZ4q0kPjZdGJG6vJfB+0QoZb1iCiMwB27ChSJNxTDwkEBgsLSHtPefc9DRIAA0ef9wqvRlW
kOivfueEADICbwgJJRd3M5850KDE7tafS4YWOqGlaCPRYnqOQRRx9OHm2Y+xUa0dUsY60cqnTB3H
uCDwpJL8iC0/OWXaEGlhFmaGA+Qb0SDip+c5CYF5BOTbeCTTTgSc94fIwHS1fqNaFOmtVkHMV0Hb
eEQXV1KR7DTZKTuAaFwDL0y4cZwxIEW2VbHdGnx4AoxIE2BljJX3xEbJy24ahwz5R3ULxLDMPfVW
dSfisLDkastEc4Yx/ixWeS6SuVuAfHLlGAG7p09GnBrztegvMLhuyfT+ZZcngyldfvOnPm3s2smL
gD4/aC3qwLjr2sB0Z4d4OvK5buPwKMlJ+p4OWkXLXqS5NxBaxVLjbG27MJaXxkLwp0QJOJkYbggB
bKu7HssqAFQZI1JbEkJr2AoxKhB7OsaJn4NH80CxlY5ZRGy63lnesrctQVwu8BEn2D+URtIKqT6Y
QaxBZcjuSN4qtRZprej0pU5x3Y57GOs7anLy3g1CiehKMT0I25/0DLY9Cg25RrYtv5WWm10AN1Ld
dJWQN3ex0g/0ogUzK1o4iqIY+crIOsQ7mFcCRFOSRvxf1FrvjxEkDMkiqq1yLlxD+rNKdoUAmg90
E+0gUXHbi3+Bp6z7oa7GnB0G+I2c5i8GsGiZTY54/SaJG5m54aBlhtI074CJhCVRdxAaiDn9vNWC
NVpHAr8svU54W493UPVuoysxmeKC2NPtUPjxtGFVGYOmUDv8f5LVDLs14Lgf5Fykv4XoEJdYt1P2
w398xcYk/4XujkoNPQTkfeTUg/V/4Xhuv0KmyXlPkySXoC6SCxHPsLePMPhm6FVkNPF79aZZno7C
aQHkEHQWS0D/VFQLxxA9UuilGCvGxYO7aSeX/j9HXoikt58jSlf1XFs1fKDR83Xkq1hnxndy6MfZ
purkQrwbdDtEfQ/0Cwz8c9xAjFgB3U9hL7IDwTX/T5qrKHi/ftAxShMozfxpty++GoB1NcFxgj9C
UbwzyNqn9nyIz5SMEZRp5Bpr5ROMdh6UjUR/7bsXns75/EMVBFvwiAI+9n7oq1hblHVandw04ABh
dyRuYEGUroJ6YKzW0fQPF6mClQhRhhFSsI6BrqRtdXYHwT7pX0E7o5gFET9+RK61PvoDr5XbUcNt
O1ojZKqFtVqoEd5PlUBKucHD2mRYPQNXcAMgUKnOb4q6lfCV6ZVncX2RHB1GZ/248y38Iy9XfA1U
c4xqD7AR8qo11q2SeEjBMtLYn+Wi9xXGApFUTuuFURYny7/DkVBhNWwyYEzy7G0TjOtU7agMPzbp
pPQj/AZ4/uGL/Atv9kU+wmyGpkQnIPb0t6sAN84uUIbZZEeth+8NnNgFrH1EL+QnQktsJgx7VLrB
kUJJjOzKaHvsj/ys7zQWkoK7OJv+o4BoeXbEON78vskdQ/4qvhFoGssH5KsnNlHVql3yES3GSTXD
Fg506xd2JHK8DJD3DIkOzN7RkzgfJpXbxgZQVWB41DGmNBeEMcGDMEN2ujsLh49wvalXE250SzqP
OeESyVImRKg5FpMffH0QrbFHi7G6dRH4BhgunEDFhQbXtE6MB7ntLfGUmqyXVdCClKKd7TOHllLD
XAcPskJ4+m1bEfE6LB0mdY/OQ0c/HH2bBh5VTrNaIFKCmX6/td5Hvkcgw6mkfrWIsPO46Yo/FbtJ
JfsGgORZFbUQHi6CGeBDWCif3aF3b9eCOpd7NkUg9UKJPprR4DN15OwGRkWwZfusw4nz1M0kuAe7
VUxpIMCUQ9mPVUi9a1vJnjv11u4h0dqPUJIzSBNOecTtR5Cn+ofT537vCwg5mvi9JpMAevX+GqY6
f0O78AGUZyk3WY0hdG7m0NQKwFiVt14e28vWEUqHMTls9QlJuODGHxkTjgoBkCf5LhbcBhUg2ZsM
jiNvOyUoKXIT7H1I1ZQ9bC7Ka0Txerh6UW1RhoVOWTWCqTEMmLdKFLbG5EwALGkh5jypVpIDtTEt
5Im9jwvDZEd7ifjyrLKpTz5X7qO7SdXBrYWeceR9iQNke9aBpHr/GMf7+jijokqe9MBjneJxeo9o
L/wXlN4/cKMKaWIQwJmXPpUoyZKzi+HGZbmvA8OEM8HlL0V4X7hErjqKWKFtw9bp9nsM8bHXIv53
ipE50m0XXqm8eGToGk/ILdJBINqY88Q3AcyBh1CvsK0kwvCzX84KVlNGtGTFWpvyvw78b6XMqW6E
zuoI56jnsH0MkGYHkOdakpScQdFz1Mwt4GB4DVWeuYL23UUtp232xM20Nd+mnQha277vAa9emSCF
MSQrOffcINyY8kEtYS6o6KAOshbOfG8CcUWEo36ojj87SAlV8bXyvUxKxYPc8FJKmUYAcPjJuWUm
nIWrOdaRm9/rRjXno/NrUYZf5lBpp6f7QD98tYb1/e6apGcDbp7PbthS77wM7x1/tKssC1Hv8ciF
TmJPnur5To5BmV7qBrnHtoH/zzfZMO5jFyNUf6rIlfggbKk0m/J4tNci0imiuzTACPksA1ueE5NK
dmJqxhwp/+EjCbG++K7dgb4Qi8hN9siSGEYqBaWwPgAx9EdBPVgK4nAe8gxrm46G9xi1KpiE/1u9
Wi3qkNZFp7CsavNwaNwuWyLsyKMoB3x5BUG+Hnu5JJQDzF1P6yHTNe+QX7EMzc5ZrcpwW9Q39c1/
0vrdTF4mKyjg7oXgwI1RVlI1DmLbFMpMpI9Aa24LWlsBUrKqeEhrYXmFsVKrfRMfeZR8k6riSDnf
E2gKdSJQ4u16f6fkhYwtStr+pkdNLyh4fRoieQEE3w45Qrag7v/7gZ21c9L9C90XbuJkqVF6yegt
gtljRt/m15MKdi59nck/HUYu2pwSIP8AT6i8mEMl7TMtAyLcccm2b5JETxzobVjOp+mzfXIce385
C60JPs44IAyszk8l2w3qdzbm92hGlcBx5V168j8ibnOarE+4E1J+LPYvdAnvUxGCiKqSdlCJ5i+M
hJ4dy6UGvQ9PuqkkH9WfkobDZ7g1bT+UUEyvzok+vNgURoxSKUJQva1oBPmtjrpt7XNhZ/hxOTtx
uvyMHUdzcIYehckj957RC28Imkhpt9ZEC94h/flcfyeAcBDxYKp4UJyxpOL6PjMK7TrF7+4wRAFx
ABNsfaNKSxAYvOfykUaviAujWhGjnJi116CjGk3PNi5hRgv8Up5gU2uyJIeLZwKvWlIHL6UvfRxh
Mw0XUKgfmi5EHk9gY24AMpLR1MUqWtTg9XdreTGZR7cEpXGJPBNjbPayI9t5/ClQtVeYRrgjtui+
+G8X/NesM/OROZPw4IzUjjth4EMiVEuXYQDEQQsIVIsgGmYkzwikX1d9Pgi+1pXGHFTnxq6/RH03
jjAuWadcHa1FRVh/YJ5/9obOucwYtY+/SVl+oZvGsHHI+Fa6HXDijy38aPqZw3OPiTDjhIo4Ku0L
et7NxULw91S4AwHlOwINVko6ssBkkKc8meKFKfof03qUpkn9Mq6nHCcUNiMAB9iFOxyOsO23NS18
4UYyIJrFCDrOjVkxOOv24CNaQjx0Psgy+qPJYFRgRofR3edIRS24H4SW8mGFg0GNPiKPvG9vHaWX
yJ7P01BYVEGjVgR9Fx1Cx5qTnuHbGGc6fn1qAyv6Qbb+P9RLmabntaW/32Mgt2PcJUB4oxzdksCK
jNKz79p8r5JQbtw5GyngOjiuFmT7VsZ5cLrxgoQsOo4Z/+TWoFPCECZuWu6BLPpGLz4SMswku8R7
hUj6XYhCXskmULSsI3ullRDmkrXsi6YPdu4DF/j6h0noiZM459MQTywiE6qyaVESCVioWZt4oFBc
ytCTbVlr0VDZhxZGM+UeE0YSjvp8BGGPUi0pa9lwrQe2ay49kes4DqwcKcBLqKBa/B8cC12vay2a
gw1yoGW58gVm66LI1XaHdzUulhQccNWS8QqGfnPgHn2l+LZTYLUb61QoHmoM4LYAUzdjS55jEBGk
lesLZBWWm9MhfCSLKyo46cAn3WWQcZq2rBoOpwb96fzuuUipABy/o4XeK9NRz7XmHjNQiBsWBJC1
hHs0ApizegPSoigHCpDiTRIohx9Xf10AhN4yrrIf3hyX3x8JGJ1Xc6wUiFpiH76cW6SyewPnSCzA
Gq53KfEgFGX9iKtwtq023FVmlDmIjvZWsXYZkcDxGkd6bnxnJPaIYsf1fLOIZp6/DGWLGWMiuXSv
Q3+WEfzzOnLADywWbmoSDed+2757cTKVNmMmAvcxQiGRr5eP2clt7NbqX+5cytpiADiZguAvuTEc
gSPsyhJo1UUWt2wShXtSh350hiyR+ZQZHCABL1DdmMYeFt73MaGmI28bPYFBaphjYsjuGtXLea6X
UPzC7wsQPSJLq62yk69NS4VKetmdw8k8/gZIkS5ImWT43FXA4YG1z5dVKRU8WRgaISRcHTjHa69X
jMO/yIdWuKvE7I5JYon2osHKz7n9VoFyHTer2sS46l5B97Lest9pYz439OXE2GimSPpb11rzEATy
xk6Y49+9ksxatrHEwtUrPT14ZR7NTdrWP70KJbtivTXKEhZdGNNjdTpdN3lgTu/+yZkC9Cde7L6u
aTOc6qkFcS/SkcPqIdla8E7obOBjdhCtdtv+SzK0JRIXbXoft1zSM8eciHchkggigOiUNixKSv0N
dJV1H2VL9TqSXXzLXQzFikB0bJaG0ge2IN19TyEFgefbFjVLdsWoNQ76sDa9YqVzGFsYJsMj4vWv
KGDSFoMaO/u1n1agyriPBWyC50Zk3+/0gUDsZEMDN8GOvInYR4i+a8Z9A/+FvXQuTdjgMqLwMLFo
NIrsspOlZAAfHAc0MtTcKhvX53EtSi47dLf9MvWsrwIqbG6ojqkqICXRhiwb+92NlPNdsBspZLsw
0t8B96ds/WtOGHnb+EKz+M/rEWyRNolIAVLpnqd02nGUboMUNS1amGZTTUSwzaz+SaImEakO6ggn
i67mOrCYHDGz8Ec4nKw9vId7SSemkJJ4iUtt/l1snbF4SJKN7rPvy+xYlyhEfSsCQUaZOxdOM57C
BKEBl3ISVesN1kRF5cku4xQIQZhhfyX2GMDZRHR4pHwpLVPTtG0Hr7Ik7P7dQFkGWfFbTk7nOXO/
KE5Fa+vZ9CTIHBdNER38/kQY7dDhY7Hk67g3M2qss2k0y2oF+JxBer9rO8zsVSABMShXt3JbNlGq
2CVxOVWIF/lb+xIaqgYEM+FjlT7Lc39wjvZXW1gzO4+k4VR7IyVVilRFRRYsDqZ94pZgJXX3CZHS
5e2y93P/A7O4sFykLIokKddqiGelUaiaXtMi0J4IpQGfGPbhVdphsZqS537gpz7c5b1wHHpC1Txr
Cb/b5mhnZ1rGeogPTpkzpyHwqjBqAXDjxP3Cc7awBHQ7Z9CZZ2/BdSmxnIxAFDrHj7Db2qH3HJX8
dFc2Wwzx4YepiKMZqRj4rAxIhI7ynIBOsKox5VkqCQoQc9uVp6KyM49jexJuBEY5lTBdwyXwpSBl
MXGasCVp0mDhTqfGHM0GjKKMlvX//w+jg32C64PxHVnkPVg0DRxkXIDibuuyol0CdnoKmOrDijHj
45RCX3WrHkfiWC2kAZglZASvp4pY5XmFL9e/BiduU0e48j89uZDkAgr6tmWlbL1Yx+tH4h0nf3fQ
Unjn49K4mI3t8hCU1ZmuC/kAhguni/ibNqZXjpwOhElouZNWp5Cdf7D8St8shrrTDzwtHUT/gANe
9XfHnmWxfrRuIlotdXsEqFnkxX6xuUnBMSF+/PaH7BPgEbM4QksLO1XVyfVLUCaRql74YAW8BBa/
AK8LSpD2eIU/har7wBdsQsCXiONGmckxGUsdc4fT61xipa3H4giS7uHxFjsIkzbAxqGgWoC8S0ff
LUSWyN8epmyhaf/l71EKkx4zuhYOdzNZ4hd8CdZp6aduRkMTdraJ8v8rETc4gfnc/KkwbP+hEG1u
a7ztx1XGEneTsUNAiNl7kKzWvBHg1t35DZbTwsGZ77rpf5g4Q/CtfwBKvaiCGg5M1pFCvPkUyDa6
pnPtx8GRAT200J9hbms6ObPqO/O7vo+q2fPjxhQFxc72g9fBz3oeyQFv49cwrBQTR0XWuK51qK5b
BrPpZ/i1nOXz3L5L1efPSUPY70yBY0JPqUdxsbRAQGZCKKGp5Kf4gblQ2sbo99refwZMVD1haWE7
6HADxV22P5mC0Vcb9iScgr4SaZDSq9bdWEqYWFbt+kL+PsVWRiZUWvYqgPhPHB1Js05xkEAzcR8Y
SjjoJmJSzheRsMjYgHCwKYKfdTgQYa0oe573Jp7G8Uf9TEa+GlFnEwP4GeRZRM7eh3z3hhmd1oGr
t5bVA1iZOX53L4q7tR9LnExkdVSkxKiRxkPD0ceoRzR65GRePz1HciXwUK/1AKehUgJDCb5Rt6UH
aJV1vOcKB0B38JbbTenzIH3fx3CCV6MkIcTEHI+zaL1S1+3dJBRNd8uhvg2QdQULJFIE+5IJ6TAk
qvRKEVmtjZhyf7EQlRa9l+oUqH349+FXA2+oXh6r7zYpeKM25/GBvxfy0aCYD8qZyBkEA2+2B5Va
wHKYZbo4I8dCnevIVrR/tiHrablaUkehP+kbTJsUO8hNw+eJZnFbvXnP+m7v04r9v+3qIQg6H/Rb
JS5TfHl+Tqlq8fh/BgaTurE3kQqQ8+4ju6iOuKac5DLZgn3qhTBgkKT191o1hTFB3vkf47Z7ae4N
izmO57Mr5SSCGwkGYMnUJIbTVEvc0Y3c5Zj6mSywuBJBVgeCzNjhz+C6hAuOtflp3Zaqlp6Ar/cy
jMfICAjiYhzLjX4yoqCr9Kk0JVnI42fOD9EF6m9XnsnNycVCa6FX26cI5DgFkNTOk+22++osa/vE
EJs5pJsVXZPnbjnJVtnDjLup2OTqlEOHptKv/9dOX8n6P//ai6sTmjoRZ4QNIbxz+vdWelDIsyL/
wxrmxSaBJFQcZr2qmJbjsA/lf3YjSyck9/NRtW3o84Ga8PcJ2W/UWVCngD80yLFwIgTctZEFVtEO
xJAf7qlg6nMIqQZIF1KYDDAk13Kq772Tl+vZLE/WB5qGPO29vLhAUrBvgGggjmMuGdHqkZ4ncXxg
mj1MwgkoNtYoLIuNtZ0CVf29THVOEcYnXk7BZO7d0w7/4iFnNXiV1SdsRHAq1JtoZByoAsE1YgX9
ZeHMdNtP+fjmyvpM++0j8xunRxdI0mXDEj3PZr/OvTKca11lsYzIvHa24Qzf/JmGpTN5m1YDJ2RL
g1rWB3y2T89db2r3LIyaoJiDFZlkw8FsOMPaI1kluhha1NHeVnB87ZovVgozIoCK8deOmI6CKfNA
TX+SmJrFXKceYlO8h5velpdUEcesBZRFoiwanyIhw2YuGJKNFN6OUhREmnOKT40Vttx+fU3fBQ7v
KUzxD/+NpIwZFYyjglv7egfcOuIOQunNFQc2aLPA01zUvjv/4jili9SaF7E3QoWrbYXpWV9pkoZb
RBrZvwCfcCuKc3vUur1YmL20Zh1+HRzgFI6slTvof7uF+vORnkWTm24iIVzhDua8xJFn+ajz5ZTt
VsxcRR8Ysxyk8BnZaoTYIgj5y9TppBFon1rZOfp+F5a1uha3tC1zi/r3qxwVVD/rDiKJ1LqCkZHo
x6MMt2/RL60blTZNioDFg8l2B+JCKQjXl7qI4pR9R/NjHoWvSa8ZWrtZp0RlE+sArWAu/cXSIR9a
aO7j0Zni4CnMqveZm3S8f6yxYQrUdt6WnJ993YPpgYI/oP35t5EihhkkHromOMa9ZiOrZHIUwipR
x7+MoC3ns/bRFefPJtfaoJv2Gk0SRmwuxATHukIqVhywHNsh2X2qIBNwfP6uyHS3vdibrnWEzO9w
rwuZe9UOYnafbLRxYUcjnYRc6qpBljtQDBrPRELB0OEXovGZuAljCHm3W2N+cegf4iuE73jOD8JF
SA24XyosEmKL0IbItuKBmTnLfJQzmjoLSj+tjulJVLOip6ULpKE0+6WvqBPLInAvb9UE/gWB5+Z/
LefyUcze7YBu7z1HB88mAzu/YwHo1zh6Xp1oMx96Mg/rCjY/7Jwg/lOJsKZcrKJypQmn3sxLrSTo
X0+QGbQnU5v4WoXj2INJQ4XqXt0qO9nN15+Xg6TYNNiwAHpTFM2OhJTcam9AmUGJRRIjmSKkvfDI
IQ3sbLrzKpsVaNTKLIfBCIbeT3pCzrwPU0QjtTVgf+w4Cs1nu73ZWaWBpmcHDcEfEIdr7PoMCc65
Afh5QH3KyfFp3dwIYNPjcbsm8oD6ogj7B1JCj+gUE5iOze//Jq/9IekYY0usUxuPs2VeIxymMknH
WJZ+M7Q0bJA/DhCw7VrTULbksP42Y4ckB8UrcY9JddtoXpqkh1dJuEfqAw/8kp1oMyD7QrhTLwTl
0aL/QO8DsaZ7PN51jFxGjxE+T8zehTt0lotyGgvNf12wKJhJk24pnMqE1Nx+pLUVt+kDEjbFvFY2
GqGm2V+y5CK7XaqHlmewmx9If3lcdevviymkzTF5MIyEQ/dYY78PjKZdS2sqQF9uFHzAywiL/4IL
Ni2H2BmwdQ6H2DOizgmOhkmjz5Z2RfbvGTiD8xCaQ+uK8pugpx20xAjVoxdqeLPpc7GNU/JkWmw2
mF5DV0g0LSikG+nLyE4mX5d1+ZwyOMQhomkQEyfBBP/t7avRW1DPtbpm4CcopnXoeFU8OskfUCEf
9oQSv/GCGyzpySXtmvOr9TCvf1CL82c6y4JhS8kEPTgwIfVyWOr4D7UJeDo6RzMPFWtgi0g9iCBi
1lhMDv4Wp/Par/NPUyOu5dN0cwS/Fwtp+0k7hSbN+03qhFBWMoGiAw0f8Smi/yZX1nHRxPmxzcrs
MjNEfjx0YylR/VJXJuwaG1FblPj2yD2A2VhGlt3opg50zxfFbmVInfonOkq7DGQItxX2gE2OBRt+
3fSp/19ysfp3laSCmNGnKuber/s/hftuefMYdSzVnPg5qydnt+uG/QFpyVNDgauwzK/lX5G1baQS
4rli2zzqC9pIYieud1WlyzQXbmVdVhzOEaA7zdVbFivExIQGDfWKYLVhCvIIaHzyyjsxbHo327rP
SvAkWvfkgpPoUiOYMIFahR/elsMMLZkflwSmv0ksp5pO6sG2viVZNlRlbmZTpWuXDYkdcJ4/Gc/e
/cWxtdUpL6e7IqDcLENGRQ/kvpfbfurLQTgJGTt6ACH39h5ArfrNwyxDR3QFLelNdXP53LqHs9jr
j4VQ5vYITeNStI+PiHd+jgUb6wmPCQwHmDerNJMeCJs28zLWmKHzhVr7PCelm8SGYvSS84fOWPQn
hCEjAw2KQjeRe7kxOoEPx6DJjoCH0z+OUU9PO2ZTczuhvt9fILG6sygmtbviUhhuLbP+hufvfqNC
cUsJWoN5sjiUIxR2Q2Z0ZkT0W2MZ7AOIO+m3R+no0Z4H80KXzKLr09k2enh+TTwfdcp0WAxbvw4J
4gCUBYCPZOE9NXHuxerIUvkC5te+Tauctq8rB4GL5PHfPNC65FFCDKVmvo7bop9X3beNXQnv1tjr
k+yv08t7y3bmRLQtPBh2p4P4iP0Wp4nUxYFVcU7YcJiSYezXAfD49Q+QtvDmBOSAKp4+Tag5dwsy
h8DObPud2QwqAplePQb5FfXqkwnZDeXMByTwqGBRLrzFm6YAuuO2DrTqzj6VJVQtRqqcFiokPEC1
s0bwGY34zZC8XIvfwwBDGHej9ECJ4XqfKjnWU+PXnrqa1Fv6HPzHZhGar69hYzf3IHxtofd8Rl5p
HcmQrGR6EzPq/BjGr3Egwd4DoWkMKh1Tfn5W8MyItXYAZf2tc7PGe7N0yiDZgWEIEWYce9joW8rk
PsukbXy4BF+Q4fp2g7/eqbLXq5bSnK3njAt8QCnz4vMGyG1XX9YZWa9hDTDzTE06xm5NSQPb/rof
AczTJNCuDwac6kSkEtxbhiCGcKchAA0KLEG5BrzM6jtPCNYmZSSAw61tIjGuCiV4g1UlKVAWszTG
Ek9uv1i/hjOcQo1wzN5yz7CkFIrYbuvfDAw540YCZEH5jo9w7VFdroucsAbb7GRMp0J8ZYglPn+J
I9mfSfknPQ24PMAAW3OGwFhKsj7dPHgyrwr51QwYTXinrzcS3fcRRt5LvOZL39Ik7cOpcd4sD6nR
u/5ZrjXNara39V2LLdyDtvKeeKTsrVHYUKOkHLErqYCG+D6Ju0T73A/zxHVL+fPPVPv/sy+wy7Sv
hRvsXBLJnV52OSsDapzOny60lgZeyVbkOkRdduGyGDp7nxOFOamJNgjFD5wFkB8fp9pX/5w43j2m
pmXOgPFKc9QIvHjVOKlkLI/9VnzDAt6J2lrY77b+q/AXL9dxr7Y3hOJ7JdCLfI7Ms1yS6c3KwpYc
hflf252nWj4sZgs8qmrmLMMMjDjOJytyeWyduGRRxemnMaQIb1Qk9UBhByQ4R/Mfjb7saUZ3FBRD
/wELASwXds7iYU+0CJ9Ov6qH5/dFURPl61dUqc61G5p1x8L87NULQsSYDNbZVdqH7jEGZJqViCjz
fqjtHv956uxuOAB2Nv0xHZqWgMDPngHs7S0LGEDaT3a1ppKiID6YnEjEyx5c+5mKvKgSsK8U7Zcp
k5TQgzITT86rsOmQI+KL2g5+KCJvq1kW640S2lxrHTslDMfr3jSwZnjsNk2HaZ2DlsBDtQLWd6As
RZjTCXyEcHu+Kq6J5G+NWMJdCwnZ4Wo9cgkQHNLJQGOC4joG0SA6vH6zq61D8dz13aqYf5qGL3DY
w3+dn5U3qmLvbXXqUh50Au8R7goIU0MPG/agjRr5yFCnD4y6ewUGUHFEaXykXNawSgMWMappv1iv
n2epCTX57BLROZTsSkzvnmg7VunOITlC4Q/PcaFLaNxyNyFrhL7nag9jm0GXg6rfBfkXD0wqRLVd
prAHFqV4D6osmydgb0Qcguv3Z9pd46yo5bkvsqWbRp/oVVr4pz+4ZaEkhi6n9rupHs9/MSlxdWua
fif5QPRdtoAnw7zQ3IbsUkRoxkrscuHoqgLFhi9mRwbhL3qX19VkxrNMCIFWFHD3ZDxcnRqVg0L9
2l6cL/sR+beGIYBP9gvUG3VqHPgt8/8uDEJS0zUpvJQ+lszbykwQP2dAlvkteYDbQSyKf+xs/HEo
6QqE4j70KiCsENSfHKAhKLfJ9zxZED+MH3HsuSxeeMEGy/Ns0xEl3hT16G5Lv9Tt1Lo9JUXUKN6V
xAJZIGBnXnRnaGgc7IyAll6zYiidp84hVr38njEILhwyZCaz0GwBZ8zVq15UzwODlF3LOy+/VcGU
mkV7Yp8u5/Bqa87fzlbPpTFHx+msicqA1RUdKSPUZIQx0reRkUVlyQl7SUUxmNEQCmTm+fLa+bIP
HpfImhWo+ssq2L8YzuQoHjYOkEeWqs1qYBizMShipTY6sufMM0ol81FXW2Bgv3Ykp5zRM+fwPzq/
q7HoPXhtkIXvZgEkZjVxrP1/T3bAxSusOlZv4NuOp1InWx56CmfugbVNtJEGPqCNwkBnGVbCfqMc
eS3NcdxN5Rw5fjBIuLnbDyJpJEjYocbOkJqBOCNaT51XjnVCklms72/pYTtue23iN32Skq0iD6XP
ccZnw2Oc8uc0MjtP12QN+VCAV0npXZoGO3huScxoFkJph3VbNNy8q20Cl0Fls04QySk+U1YTBKXv
gmUZlHun/fE0fs517tEBQmKr8S9RagYCasEYkh93LtLh8Pt1EasG75YJNITvaiteUMcr8Z/UCtjv
+4yy6fOCIOQau4YXDqfeqtwylS2qxI4wWrkrQVoEr8nfMZDt5vtb/qE9333PwXGCMWs4Mf5UUHaL
+lrZQ7Qkh/T6tUp6nR7OHWvqpI9YC4/wPsE36Ioc7lGYHqp0UZa2mTnYN6cgi+2M0Re2EKfrJXEn
qRH4TXGPHxWdTIbuFki1JatvU8b+YCBTyGHFukL1htistgAqiWDDa+RNXnxP9hQ+Yw7cQ547Q8Om
Tpt/PQ0AJ/keod8xBDWuCWTkyPQRG1I8jArwONr+g/50Qk3yBzRR5zARCFNpNUh62eWEEaLq05fN
5TMdxxF5oTmqQvOSFZwDzx+mONoZsMQ5VXUA3THJqyV89ayrYSTW9lhWje9Ax/CRsDgK8sfaCL3T
VTPfps6nvjqvYq5Uf6mJa+fgReq2pCh5iuLmS5TcPOSMiVxYjDeAqvSqVXdwvUPbuTtvX6czsjSa
zYqfzBilu9zoK/0Oq6nNh5Hj5HjDC3/K639yt+TERhZj+icQ9KdtKqFaeMCmeyf6H7A+RLUkTyxu
zlJmhUutKrMejA/0EiKQWGYC/C2d93gnU0r5wDyANUXy2k++40cE4EJ7I1TYnKt8znB7RJndCFmI
k5247HQG5uoW8lirOqLxFguZEb/cz/7TC9gVfVg8gYgtJQZalqMXwOpHOAnAG/xMkRsk3gM2g36X
Yel/kAZm+h45nUUxKMiszRDtGPfiEg8mJElbrj1idROqV7oFZkp1gTzJu3OgpW98u48DHTdL1XOo
ZP4iNdSpkYxXn9P2DsYD9EHLPnu9NyUktWhe8lm7DIu215SG8SXQl8+FsR5YmYIUbcc8POXr07Va
V6rcUd8J4AVwD6MXNhXjCwL8rPPCMHoI79iwGTRtZgVfad/6BntyIze08MMfsAqeA34Lmn/3BOfL
G8RLM+Mdg2egPcf5Hsz20V5wTdLfnIsQILYxCIOrpMMjgODmS8HvHGFTciYYF3x40N+Ct9g0fPQN
Wh/y+iDttGkrmugqc9gXTme4b2ebFMm5DFwcGbkAmfUyH1QqEIhT6WNjtn/1SxUoxIn4ldwvLOWg
yp0lVSV60C0NiHddJ8RBJFEZNAEfjR8Wce+COdNH676MIqRSkgeayHHsh6lTJwf7raCRpk0frpDC
qIvAzFoA5+iG5T76NK8nDkf0+vYj1drXqBU4eLBdy7CuAXD45sndFuLRscm4U/Uj4jc0jdKsF8L6
3IVaj/N89ZTIggbHXC9aWn6V8qOOZizGAYXgLoa9YqL+23rEdlfP0NCiV6NcFJFoFxX8Q8QgXIgg
CYZ+n6W3fzshkWr63X+oGo0pGQeJi/sZ6qf6aYcwkKS2xWyJRFYkNarht0HbAk4M4YgD+OD6l5VE
hWlc2ri3f8pyEodXNVJXV8j3HBWA5k3yMPw3wl7RBD9Np4d/IFRZwFm4PBLaVOQdLsXbphEg+2+h
ayqzK1TkbezJg92SspjSJ6vt+YfQIw6LIn8Q3DCuHZI++muOY0Un8VA087iPjrral5LDjgl7WME4
xAr1gnIik+SLtegip4FPjOSDFNj57iIkrHEncBrqb+IR/QAxPukWIVx+VCaEYwj8mSMEH3UAYONg
mHZLrbHwqJ+quEDEpPjzKBCsbjEfVj0YPP1Ct9D3972v0LMLi6YPBRzSvT6G6FU9ozUbisYn43mc
+S8k7tqA19drnafieDyJ1JH0SLRgVKdsdGu98Lyfg51cB0STN5CB0TVtO3T3yeZY76EavLXpvvYM
UOge2Fc2ZSbk+Q1l8uq6dF/v3AmCFqTOY3fOXkve0nLFxDwxARQL5IajpoTnXM90OjpftJGkNoYL
kATJjt8mLvubmddLQnthvQ/AQAtq3qS9gIfFKRRwU2zxuHeDmRL8p1aIzeDymp+l93W5l5tqySWO
tqz0R/RQpuyZiQAE3NLiUtySc3O/loqbyr3VqXY2QPP+7ws4ihKMbXCOQE4cAfjcPqPHeD5C6zo6
ehACpNMxW/Oy2jEYzgd2dV6G9XnamRCpeYJR8uSnejmlZHhTBCyphExY0ZuLY2sspmpW1xgqdLQq
LxxL57Nlr2C9aAX0+y3nM1jdo/xrYQBWyghvfhQK4jasqW18J9T7vbW++LPYWFXaD9KZbETKujfL
wrvnOZTR5uZ3j7mNb0YDI+GYiGsYhonxZvWRQ4Fe3YQJcZ6kEX9K08tFDyvKvIz80IvhAmzxE5mJ
2WzZ8Igw4bduJ4258RgmtXEadE82reZ0uq2Ax/rXoHAweFw33buCBiabKNhztXHHWdqQqd8VkVTd
lymogYTug+NZzqhWno9pIbzkf7S9YI6FvFa5CfXyUijmBO08OU33vmd+CbveVpfiJJvmOJujbLpy
jhsUqqk6OTCDR00+vxdQ2xfNKswKNEt+VLN46QqXxYZs+KQY4tU1QN+rKnUaDFT8GnvvX2bwOiWM
TwhC+TX8PhFkFifkMHP+zE6BvhMvn123J7vmLOkJcqEFngbPqOyzyrOgmmIY9Vd0He8PVRfUMHaS
9+9cVP0i0QMtuhvJPZgCgImkvXuKBiXCB1J837PJFybsgia3hrbOUsAQDZN0jX8kjJsIyvLY9VR+
vdRItvRzMj3g8XyjedTTe1bFNHOvVxyI3X3v6/xOQxCKN0cjsZVPA8Jo3VKD1u233CuN+WSYjiAU
RyeUUSieYqDU4DZsz6XwhlHas1B7leq2A1uv64iPQPaHAP4MVWPLch86bun13nIIRKPBZ/3cUDP3
MTBffWotjZDUN7gj0Gwgui0Y2DEdLaTx8HPuaMTaPKlhu+rwS3huHhxlNKa/BODtlEwrmyMq8t+E
R0/zdnhMbamYQLIq0yi2srAukc77hSfXQb93Nod45fng792qKpQbVtfsYN4i86uBwlM65boRQB2Z
1YS5dmn7U+ND1TdZgNyqDf7h2EOnRjfPddsuuD3sRPQ2zI5fiyB9qo6uHOOhdQmfoWh6tdMGZlY7
vnEIpi2gRRPTdLhBoKc5bI+//rstLsriEbD/qOMKX0L8JBv17goRKiHNurBm068khqdwse79R+Um
3MCah6hNlYPJyn73MzjevF0habGaBmtWPyCFYk3LOMKbRCn0usNuNvwEkeEh7TC5ER6vBARVQN0J
MmReNI+vFgbgIizPSTVglFJ3Vfly+pSiZEdBAnS+rGyRBXsvk3hOeWlFj+HISuKkNenPQ6DPIHlW
lKyN3xpFmpdNsChFMsxj86qZpEQ1F0//iu+X1WZOzFNrs8k/0+gesGO94rukR+pRl5qv/RweXmxs
KZ2pKpAzT/cQwzaNhVGhxZKPcG4HTv4V0aFoN4ofFBvNkpQGXHzbSDqCeO6E/V03a+b9q+/bcI3J
ncY4I51sLjhEZI151MjsdO/eswKEvf7szcj3YaP9L/LHhzgJebNM44esYerRcNmYv6t+rQtG+X/X
DZBiP4/FooQL87swDaPAByZvxxURIjmZZ4xw3RwIE/d+7WnD1yziS2IEmdUEXsNbIQToC4ljCJij
uupP4YsV8nAFVU050Fd62/8hIxG7BCVcDfrukRoQmV8UKK/0BTb48SzLEdntM41wBbDVxKM/6xib
CHhFSr2lipG01BjlKPJ0PmippZUCcpkER6CDhxB+qACF3WL0V4TZ9WxtTcS0OicT3bCfYM2jryVf
qJtQyDeXKEwP9A1+IWTw8Hhc094lj2xkHDlgSfQKuTHthKE4AIQDm8PPQxDztfrQL9PKfJ9vUQhi
pmldUCiBdl2y6HsPsNtotp9K/4Xlu9w7246863KZSSjJoZY5hqaIUkVZvRfktn/PPFQSpXdUp3Rs
5wt3ARZlEuKMwqHM9TtVbe4lBO71vJwTK8dT4GL9hY2CUjg4CMIG+qmbSo/SI4Au/tVie/1Tsx+7
fFggoguuri1e4so+yUSWKwcfWA8Bi4yxtGHW4CTFQ94uGH1xo3S2VJD35AMpzw2f43Z6p+6iYJG4
NOKjHNBf4h1RWLuR96DF0almrqlYDZDpI2qAgcpA0bOKWLQ7y9yn4jMVXwFuJksgujT7HJRikIaU
VwckyChXIvkPxrtnGkzo6eLJGea6Zo1GMFAnepiun25Sa0RXxtm6XXbHXlSJDNKCXCoepxcsoURA
C24UP1bqUwZObPgBRET0X0AK48PdG3exVtcwQ/2pV0zGeQVh1TkpJa9vBlroaaWpW097L1vKznKM
m30cD28oIEnjD5TJ0P7zcMCPKQpuJ5VUookFN+6l8OF7VBwY3hgQpOTf8oNyuLHx4zL7La+bqQlv
rwF6ajoBHxQCptWg0An1tHKGwGhAiqzOWOz0Pl8GmBF7OQmmKepgD/jVLAIIXxegWQrPZiN5QeiE
6evfjyusvu2AaqB7wOeJlwB8oKrYr4bMtWMbKOtCIvisCwtSR8uxyCZjOYDmycPRsFeOTBFSXyxK
A4PYGHbq4FcyFI1jSk/WK/YhhL6yZ3NUn/n2qkKFYukQ3EagqDDU3dsrn23GZvgK/MDo6wXk9Uul
0JVsZPxOgtrRteUOaYw+n7dpL59SVvIq7kG8EFyz+NTtFX9911sQGyYKEwDSIhRi7YeiO05fRwPf
/bTyjq5oJeMb+IHoLzyFKGXkWI3K8CoBruCMrfCDxUItr0zA1sWsdur6jrWPNIcGxb/KwBKddsnk
rgXoyOhUZ5E3Q2JtW2+V4y0URBxUcurp0XN3XUE75TuBodUxJEtAjmEnwpIHZCMbdOGiWK1XCZmG
Aql/7ztJ2c+MOaVRPMysYZNj/r14icvr63BMhW68OVSlIAYQ23hgrEEsQ7ZaHd17i1d0QDoF3V87
YfWk9S6FGy8rOZ2pAWuZBQLnoZpkle2Y10dHJIDVm7RvrqajSbr+VTo+UaRMXonJKMMhq6n3Expi
3ZL0TudyxG4YGlefUuU6azzjBd73AgP7ezmUqaudsx0CvsyIDq9uP8RRbse+jtvMS8USIs1ljaxh
mILZ+f1fVDFx7qnM6EsN1oZzKCmsnVw60sAxvsw/lK3KzcMPu5SGwRcjR1cmQ+kmiwUY6KlvsCjL
xT5jjC7nufxYEv1b2lzmCnMxIxCV8CfstjJ1k7TushKjBX8tI2F3lUQHIuaQL3p27DWijL1Khnzr
Jkh2J6gl2B2uIzqwyKkDkFe0nVkTbQmCIkrh2iygm9kboY16OMwZI2NxiQfRJ60FXjvBFhJM7udZ
uyod7ev6nrRVco88K5AxqtHiZ4lhK+Bwq+PjwhkwBuhSjIJZVG2Hr7xvCxROho2LkaZnYZYG0H9h
/V2rnD2rv7dEpVf3nLRUaDX7rnR6Rs2gFWKdapxusiqNt0jQJrV5d3wB8zjRT9HSXxONQTIDlNT3
6Z2dPus/KPi8PZI6bWkfV5MPGFtlua8zBoQ1w8Z0xOaKA1hHa2GdFGgZWPfRNcBiqLp78/MovcFg
qduAZbElfS8u6Aq9WOkPc9zd7z8F7DeSLmarcK8oK4YtsYuZT+3s9xVRjNv9Liomc/K+I1ypTh+d
8PCxUdwe46V1I7Yi2caQscBMAd+KbXawaBw0z1ikxOcpi3K7qnQf2idRTMoKiVUPKcuIjyc5DEAx
mzHH4NG+caS/dV5j10r8YiiqKafirBBgnTws8Td3epO2dw384ZWvVG0Oeghxh8rU5MkTCrtWYF8v
c/1zq8cyxO9AmrZ/rCVWuvyAB6mBbpOlFtPjEFV0EB3jwVtzfyUH+JxiD3ldFoF7uAx5oHz9XqOu
eY3rhsXS2kfE6MyCKYmgiKYS1DuaFajUPyCYRN2jOG3nABcXg9RUxqTUW8yh9YH6G7IiYZfV5Jo+
jlxAlew1B0zcxW0cJiPkh5QPDlg4S7tsQE/wHnCTv/BX5RpVLNw0j0QvzYnyPa1WUunm1x7Wb+Gd
iVLK5Byc0zGUEBkaYteNHC3M7wFvztbtTmaeZeD/E31aCb/YMivYOWxg7JucxydFAOO800+E3sbl
Zj9uKBJzbexbyXc5lohSgueBnWsPvGi5sdomfaPFqlDnsVxyOf2+WmSfIFf2Awf8dBa6YdfgScDQ
DH7sbiPnaY67mhv7qKvehgodv8UzdcNvOBjEHARnXl3MmU2SD3O+rDyY9YHEA6gCW0Mu3gfb4s3r
YZk2JRPIHLwAc9lQWUzxh7oGF0hy5+2RUl/UvxScNFpmrnntWTEtpSQUAdKZR+ZhV3ve1LpNx/gC
0Si4uHadc0i/gA0VJlD6ZVZr3e9jSInDSx7f7Q1AvgS9XNGlKWkrsmcFuPUm3D1FU3cSoGYa+jK9
AR3mG9RooBs2eTc2p5dIMXMmfgwo3zck4NCOGBf+tgbu7A+kq6uVcUguSqjy0U1+d986X+VsVtQq
E9VCRA0ftDPxk8wb0xLxSaKjd+jP0mStYR+5bG0VXIo4BamDaTWPDlL1vgGI/nedF9KodylV8Vjj
xO3ZEwxUn5Or3h17cz1eU1eroCd9fsoVlvqlPXZ4yi2qZnXQCARPW/2gsjwxxR/ATGpiR0gmaWGj
GxCvXFdWCkVh+YNVapfm3DT0EfjWtKnzEfUMgApZ3WUkDOhjXu+B8X5sU1Kasg6s9UQWGXGq2G0t
vNZc2xchC390MfzujtCQdXRX51oBVvb62X+aAd2G+Y1tSWA38tsTpXtrk459Tb1dDVTCfXlDMyhh
ZO0emmSkCZ8ivXHvNPP4Epy8TWNbuoHy2gqJhS/wsqz2cj2r1Sgzfe0tvZUd1lCPc1M6ye9QLJSl
BygUDcZ8X7F7CZMub1+jl1dkmXkRjJ1jkd8D8JhsSAnbY9jttbog2sTadk2Eoe1M1Y00zG7yU8z9
c5+jfGs/QPtUHHiVHL0kOSdIvQMmwQhFRvScunLvkRM78/RGGJVoUnqi4E1srYcHO+8DiF44uO39
XGBjUiWsI/GP4/XfJSLh9TW2oFy5IG3K+qK48kGxNCJnQeCExNqMgg/drZegaWAdoeVw/L19nooU
BpFGhpz5UfWd2DDEWMpgB8wttLg5mBNx6PFzEJTjiey7qvSbkmdv8FHXiztpIfwmsfOmDUyoF3HD
58U8BFTHM2ux9eyXyMei0ki79wh4kYOT5XNIVFkDjFtT3kEbaINwrl0FBo8TwA69iHaANoNHWEE8
ZTQ4igv/MsJrKGdYNFoFmn5OJlhfryHULg7Rzk1ZbVViSZcsnqTpkmIazfny0tmNvtWvitL7vdHF
m1/Z5YPPzj9CJZOSEQ5vYkbVIf6KL0e4DBnxH9tHuQaj4B8XoyVU5H0uNmaVsvmr5NASE9NRpvze
wg7nXDvTCeK6Od+MNVA3R1ys8i9hz611QUhEPkHsbrpv1MiYI45qZcRwj3ximL8fg0Wc10sW0hSu
SFWYC1Kv5mM4uvZUzrv+A0QXIA8OBGKfnac93729qh6ILm03Oy4dG+VZyvETDh++/0r97be4t/gC
fgrYbjTsk/dErwL5WL3SQ/CS3bF863TiOnBsquzuKLpppJgOxBwTZSBuKTP5hU3Yo1wI7tKprWtz
PnPAw4yVKVztTJZErghC4zulGGwe0VGTv5zZWJiVmGOWi4lZ/DW2uxrCyVgJ+25tQfGELBQAxXDt
kGUbPE+zudnJ755rvHQyYn/FbhC9ePvxX9H/iTX3WyZ0H2NXLz+je4J4RUbBDzERwtIUWrmrzVkd
XkN4rMDLVSnPF3QbnU1k42caCLw+DnYAuHAF7dolNGfzjKxW1MUR1XlWXAgyorW+xe7/Fx1ag69y
kAun/wOflhspC+fxrR78LpNxdhec3Nr21c+969Y/EGWIjFnxKOkP8F/PX9nqTUo0998wsOH9hnbi
OjceaZXWc3zCsnL7FWvOrXh+elbSZD0E/RaNupsLMYO08V5dhJrwMpdODa3Zy120TjMK1b0GQ+qy
yKN1NBYZGLyqvR6vu5JfdqQG0I4qj4EwFggFAI/2wxS3rzy0Z+6JIrjyrPtP3ULAtqKCXigZrOpX
Xa2SR3jq4LkuV9Stqi3OoIzJaCs4WvW12G6fcI++LZdN4dL0Xn3IACBwBxOaIDTh2T5R8qxhDJIw
syCXRfatXxd0f8euwj9YcyqxlbaJc0j0qqt+M5yIVnF5ax7jpJPWI1fKLJz5nT7vuLs7jbfOtF8U
69fMGMSdg/6v01gmLnuxIptYHP4JnDufo3BnjB6KVkjH8BRAAolflWOgaiA33FEtvFU+Z/f7NK9i
4mmwfHgh+hGeBll1M7fQP5vUrQFKTs7lMkGQC+ACbTNSJ2qKA7/iIChHfdLR4qvDjLTimWsnuQO0
2K2XaF7fFNQLOYvbw2sn5/G3yPNb1wbxlhNB/k4OREyUS3E47hehPMAsqQ9hctVcsA5ttjBJK8IO
TrIlraUuq/CxChX7URPFCpnNK5+jxQFkQfoVtLt3JPmugjWKNuR5CiDt5CqhkAav5+DckMvDbuZk
EIyQirobXaTjTX0zh1tE+2hofUP4fcBypsD2rjt8LE4bjIOC370BpQ+vGdmjPC8vHiP4mqXdFeXS
AV0d9wmule/Q8Rww1UkidVZEX70QUd8SQaW0tcFT/idVmg9HAPQWktAmkZNtmogGcmaBG7v1+XwY
mHUgVC3N0pxa/p/mdUDr9l8KQZfpRhfsg//ICxQsUpN8P1F8OFvo3HTAubFhS6+1SgKuf/s55BbB
AiPyRhdduz74u060g/jrC2pJZcBYt9uAd25gU1YnOKu6V58cFj6UkYUbrMdFXr10pIBBLwwcSXWi
Jy3+iR5ksbnysD99ZNPr/tRD5I3ECiRnaZCTNhEN+zmgjMn9R4wBdHRffHqKiBTfp4K0yMYW9J5N
vhSNaVCn5Av3Q/kwGpOI6oVrT2JHVhb2y7zi+ACvEpyxYq29kDnN6e7waUK8KoD5+V66FnzlLwBc
DqlKVJNDbAs6U1qQT4tFYmxsm24nXV5wBpnngc5TatlRb8GkvwmkkTHB8laDT/i3Vit8c2EpOMz7
8E+NDJtTto2leQHMyIaujxDHpT8OQ9mw3eEyP65/QZg9Pl0/o5J8WfHLyLtvivXOoDApMv8ainuY
WW8mcNPu0L/E/q9KeDocykjmDWMLYCNllFzZVEOCvVZO+W2aNqxJCZEuEty5ndKjkb4fzkB+C6eE
QP/8a3dXsYekoJIjZgBWi6rewvc1EUZSpUUYi2uGpJ6VbPf+fBoQnZcmc5sWsAuwAsqMEbYgbkJr
Bu9kKHGs5JwDRyij9C8bsEWMCAHUOjutNSgK/ModSlGAaszQ2SsMojh7nnYlpvL3sX33eP35O8/4
LHDIXp4oeRjKtj5GNLthP5sAlJs44lRsP5VHwJVLXjUAGfobsMA6ywmIvH3pvtyg1st+xiv0+YWr
ujeuvsWwBVFxqTG27HF3JMzVieUpSmqoyQC7Q5KARhKSF2gByPUlpqR9e/Esaqsx3hHwp8pLeOuw
+xQKX/VnKnS7SteyYzu1GT3zWicwMeMq/sCgjy7nTE8BYfZyCoQziG4oqCWH5pX5vxmikhhLvF/9
VLzOtUsa2h9kaYHX6Kp3DwzspVjvenTdNdqEAneHbAbi5/BoxvG3ecleOoT+iM5fZlE29qvgJJH8
KL6AXC5gRv1v9Cg20ovFXOJf2yaPRHjfOx4ioK5LzXTst313XbFfDyFbjCM4t/SqQO9U/jFvDKQY
bM9FN4pcyfIkvamfqvq66GsyWaikSO9ADYqIo9W+SjwREVuZEAY9kMlElnbcuABlrXUTerbdzHZw
KgeumaDNBU6Kr1ca5q5CzBo1F6rgD/uvkb6l94xnQ24WPYhW9XewcEPANCh6MMLwl4VF8+I8TK0v
Jh79q2+4Ppt+bED3anv0a7AusGJybloyoB6cXIGE1H6mDgbiGS/sGS9Uze90tj++7I2XaUgM4X92
kMrwJ6iwchLgG9J57Uvp9CjpDrYYWlUdC48NjBn/Sg/XCB+N/cSgh3nTlBNBpUcBZpoy/h9ksM5Q
P3mlvs2U4MD6LR17WCz6jrNqCg+nqXaNwYCPhoHgYkRJeUMDkuMPmRytzhMnHGEIsga5rw8kp1v6
zcpNGy9pJVbG5SJo+tKL+4v+fwcqPSpxuz0GEOfvuYLXy+LkIC+dftz8WcI15Y3Ge+X1c6HwMrQu
dW1fDLctla5fBreEdYzU5ruNKvjx1oUlPlz3k+mTwsLMHg28O92Ys/bJ5Pdu1yO6hvQ1Dyykn2sn
DwiCE2trwo9mDlyGx71DijN5jfRIjxgTa/qhlDmYWXjgOJwDVlkKZEXZfnUuy60HN7kYZGtarjXn
izrCBAhsJayiVqf6ebP8fX0dbJ7JCC/3brJJZ3OmAhmfJahH7ZwGpLT9ak7eAMj8l6cZN6VWHSuQ
Kf0FSxKbv04rcYJdu+k9pDZO0kXyKZgRBI58jIwByVadhkAF51QrQGwKG/jMi1Xd43bhN1T6Wxdx
54+jHlj4OiE9ALss3oI0oCi/cjPoOZkHNt8wArG6Y0ZgV4wzH/LUwbPOHcsU6s9AnOTfYKWQ9xtp
H3Y8QFRS7dUwr5lZNlQe4jooZsqb60IFlgLdAj0IemPqqkY/r5DrrUkA7+/WfY48OZc5n+W36shg
d2MZNra3CtzP4EOBvzUzIi1tWU5gPU/gTAaVZmNreKYXS/OTGB8qSYHCQLaMj+KC4qRmdYVnRsA8
z1Ssg4n52Qp92+tLimdd/ZJNoBoG3fWy59Xm8rB20Ucs74dQbaw1bs2mUQcJsKnB3wcMIlExzNXd
fTJo6rY83fwcl28WuNqWknsopPqxKTytPKja+CacwRUxqrbwI95iImKiejOaSBuZberKvNyCpobg
f0+yYi4aPfU8P19fL7FmEx16po20liQa/40Hlw4LSaDAsbJbkNIYvRCeLVSJDaN/uZZin0a0ep4e
Ksttd3O9xYzjfkm6a79peKqR1nk/xOawVF+af8cH82VEhNDN0Yr6OFaxsUZW0zbIqPC1viyTQkpg
5ABO/j/Pw0kVL7uJ2uCyz2+1lzZeUXfMEkaZ+eAGngWeb/038c9veDC8sR8xOA2Uc9dVG45MTBbD
xGLhrClvc3+t4T37G8lABJ0su4z2DjfZlRBIQk4ogqbb4yB+RM/g5w2ePrMVOiqeRP67rOiQ+1Hc
ulzhihE+ryxzkUPFCmoRRumfXws5Nss7ONgES27hEtZfr6W+gKxfjweiASXkFkTONJUJLICMKRbQ
1Ly+W0fBcPeHWWIMR2KrQ/I2GvhfasM6xCGPpCjU8yrdYUmnPAG45YBnNyAb9Mtp0wYDkDaswG0E
kr9dx5QiyElA5pHyMD4bENourruBq90oCOMWyHyDW/H3zQJxQ6/VkL2wdRiItNssmzmOu2C0zycu
KZBAbQ4Bd1Mr5tRXEMICwTvG4pWQq3TbhZlLH1AO1eSTMIv5jVX8k37eq8vLIFA1CQg+6wKvH1ok
dphXLZdQepEW97ea6fkGO0tlBPwoLWOrOy4eLb0ey3xLOhhPc/CEbj7ju5wYkoFwDtzpgnRlEA2C
Ihr+odFkxr0/AlrtRCutkEPBga3flsQKLOsl+/QjwqQNOI/UMZLPHiwAb/jM6xWCKvA3wQqHU8Y9
qWrbIL1aBgbY6AzUNB611VqEqLutpeOdhG7VmiJSjzgZKniXFOpMvHTUVgwDYDp0A+34nmSoC4//
NhWP8eMWDxD3qoXH2IpZUhOnmS/cA2Vga6ZF/2kUDF7Bu5+rTJFApSh3oHjY57+7G5S6nqfbY3Bk
LRyo9N3krN0aoYFDnjs2+phCS5H4XGcPeVIvSe/3XMe6hE5M1z3cK07d8yYP+gfvP8u9ROk+YooV
s3mCdIPgJTBA7jYuJ7287xX77wZIwHszx3OIAH6/ZSPGDTNMxkL8TECl/aKyofzVooXOt6Aj/REE
9sHTSTySmRVVOhmn9h2sCX4vF5OYZGLiOyV8qZoQKh57XoQ6/fjinC8nWy974VUkdLoLnT+m4cOn
jUhN38JtLoUaxJ4tNPszyp9b+kESKzJS3lsB48sG98f7PzTHF0g1qrUzrKg1hscYZGUh9JhI1DwA
rTVPZRl0i3xSBCAAE1gFPjjfAm666WPbyLOua2w4p+VnHit5Z9uZPh/sL4CAhQnSzYWx/3413yhE
IJDyrzdgvJ6SaukwmanDb6uepJOyMtmpJwIcvqatEYDZEbukZ2MO4NpPVWUt5q2OReY3kNxFd4BL
58zIsNl8+cBMCJjSwDtyVFwCJcCSFHdghDzBtvK45/6cFit0nM4h0VgJ2oju9jgrw2CgOWOGAPed
pdCOUJdgUzpzy96z4EtE98SwVDojbUP59J/jrX4IZuKji+3zjwYczvHzc8OqXC/+9qiXA/uOWAyV
050hlzTIK+Tloo+jJboipC0cPy6eieGhN2+m/JDaM+WVNgVCTZ9iURwaM6ZLvVMnLQ3ZuF8qwnpJ
Z99DrMWEVIQB6B8XpHdYHULKNtV0JfFYeJarspisQOC7ZTdkuzXEtQIAOQuYYUIINQ77e7gp36u9
aFh+VF1cR2MPep/UxE4lhGw6qrewULzLKb8CVIsKvPKxcvhjsf5M+A/HZ0soWm8u1i5r5FUn+LU4
ekYSR75+7tkk1TOLB6P/Z7C4aMnMfeOiD0HjQTeSO6gwlpRxyXKISAX43j3JDwACHcQVI9uTW/FD
uAw+xTnSK7zQWrASnmhQ4No7bAxTLknApGHpTuAdBe4loCTv7Mgc3exWz4GDBldlLSkF9lzLWJKp
L62NR/8kQy42/xRrYnAlhyL4XiSpGnO4UpyOBjyA2BJ/ZT6LDX7JyK5UQbs9ZdBANNIhvPxX4WUL
tKBWVZsrW9K1dnoD6ULeHcy3QjYCsSPp0lSRS/xC2zEJhCdaU7FEDhls+Q9h08TDUA5js/hE2l4M
dM4946AaKpjTceKVBnWfLB2JTW3StN+zh1uWzlVfln5ioJ5ScgId16dYAEmSwSu9QTF3pTMgbVEr
OALZUkEgs9DH8xSWF2gLDbtswhioaRX3/SKRS0ycGhfx1OHkvqs9kasQ+EhBU2Pp6JOmGJE1sT2w
tFotFArtnoEHS0ugV5A4kTudfUjicMYxIrkz/6P88SaLPVm5Zi6Dp84QEkhkYuhVB5XX0m9I3UEd
2hQskmsFYuHVilHs7Bv1FfWT+5BRCxxAGowfkVyaEkGMZdtnKFeXH+3OND4ifH9X+UluNCpbVjmh
jZwH9DgQLxLSE5xQ+L0Cgvm0/Pw8Vy+BFEl1AQ4ypco/CcdnptGTK2Uc/iNwPdI1AnCZW9EjZSOD
b0/fNGeeTaLOANkMGLhvAnPYkKoJc8g0LjYbHjh9kV/u5Q7gf9vv1M0arvT0UBo7QrmUanJOYUww
N80AIQ9CAHvFP7P3XrxRU1vFmVDOa4eEuuHEgO5fCz5zVVlZbQwRLLH8Su0IGje9i7BGbvnQ4OZx
rvNjYzCz1CoJjdQ1Hw7sBfYjo69WxWxchd1RYf7z5VTN2M+GraM6niKR4fYhX9nQxK55cbI7h0st
7HnU9t2N4gAj5AukdvZCYed66tTNiricsoSveu/RJfLng8kGUHmhO2c82jIdjc3IylBcebxG/X4A
6DNBdkbFHI6AR0aJueLjaoWxgP0U3tfQFLI9ueIi4MTpYm524QGbbIh07y2GMCp0ofb64ThQL+N3
7kcFAaMA6djvAV2juwAQKhMEGhnxc4FujPa4aby7tucRZWe5G51hmxCj1jBgCeV0OSBrYJRmcASV
cPegAMC+emDhTm3suLJ3xI6G8dFB7MJxUb/xyqGJNmqlPw3ZXvth3TZqEtd4pkWbI95mmp2/CQ01
FgCwg3QgKtmXO36mblJ2gLoxjPQGV0NlEkwJTYZ+/oKNKXhj/f1lM/sqLisczjqlgybf6bNNkMi9
khvgFTtFRajPnbZfunElhKerrSwPkCCPcu0J+YEDEu12x4xNQu4E+YirK95oe4IUaEiaSVEO0klS
0Twz2ZlBbujq8Mewp67tONZpUyYOkA7Vl0FJ7ylYAMNxn7qBJbcIcBlys2hscLkp+zqNRGBm5F4m
6HD4CU6FRXB874stZ3bmKvz9wDKNK4LpRLmuUIoQZOyLfs8d5q+gu7uKxLINsDikV6ayGogtIS2l
KOSWefq0UwoRkmfyWQy/3Y0AleYk2Cxh+jznyORFOqU2xSjCWvMtLdOacO5RRw4odRDh9wukuSwX
qrF4BICSZT8CT1AhzbMxq+EE/UHSMLiBeyJehy0C8xhg8daFqzN6wckO5CCMPwo0Hfyxejb8A83N
EgH3VxINvUfot5m3RgGbDEwutY+j+idCZ/CaUTyVciJP6u/p15O31dyy8v8GJ1W3eWqjgaj1hQrP
HRW/VxiBUtWOieJPV1knm3if99cxI7noJN1Hc//Uh9XFgnLQKF/CPzRWzJYElGt3VF/XiSUM1HU6
XYbFrHWO8XEJ5fQNWQGqlQVo7XeTPdvqKjleuHbwAkX+e7BLOREFbFED4MAxBBGNgTXtZEjVhIpG
LY5gnPiF4rOst6+jQ4BYr3z6zhN8lIb2XM1vlU78FW5WSWZYPTcclG48Iqppq5WRUPl7S3aK7XWk
aGpKRCYbTIP2hk+8P+CaegzlHcDc6N4e8YLYuPfmEkuM5KNbVWyVYUrZp9OVSpapQakEjtuDS7QP
p7JPtNdae8mVLo7KdNhAbsMopCRl9oTeWZeXdURpwFqTS65K7LNtXothB/T1IzN65ORyGgS+I06B
en5fQMXYo6OImfbioIQF5ITmM/KtnsaYwIo/RXihkCOqnR1mMYnWmjz3ARh/yIC5Pfh/y2qfSszu
fwgZw5ZdB41tZeJJPkJq+ruHjxcgnWEA/GIs5IdQNGINp5g1OhE85RBJZ4jVn7hpnrrUXcWTLRAb
scV9XKjNwN8dxGGhifi9byeKx0ihxkArYCUwI8pK99dsGDkk983il5B16vBr4cIia5nJRW66KEwL
pXsb5GanABqfCP/LHozOcBr0mapCzk4ciXF7Enr+MzcVPjNXyNJhDOy91P9mjFyT5xwKCLWCPyrH
lV0XiivyHztrjt8HEC/aMtNEin726eedhI1QFa88haqijhU2f9PP+zWMX3jlAzCBfcVW/ZpfseT2
sqRvovpo9gxc7S1H9aVq05Thoi23EPn3AMOeRUsy/20+D/FDVB+E1ZeMAr+CIv4E5ulkPK625zFa
OUYsN5dwLVe+qVS29bvTznVSaKRJK60XFaBn15RmHcnd3LqQqxX0nWoZ2jAPARzod2caTG64mt3k
I1Hm7+ebWM/humAgGcaXpRP+DTOk/e1GxjxQOWp30SeL2NUN93IGVwv1r+y/+B8NgENQERFO4fSj
s4EqR57ywMyZ7y0zfv506u4UL4pvI+cbZuyzs8FhRnvC2ctzc1m4OIB1Q657Cxe6g8QdN+MzOzIW
cvALO89/TzKZ8lzBGFm3YnZvKhWO2DaqnE9vI6JV8Bg8iMkr5ZCmY8Fyj/rvrIZwF/6Cq+Mr7bNz
oVUK+Ogcu4Zh24Z8Ke4WwBYuqfkq9BSWORnpZWzbGpbEzrAuzjy5fJ8tNGEX9wkg15epYu013YWC
AqY10UOeEWQzn2UUbVFzRBr1Et8OdGJkAu5BSOLPRqyBSaDZzvCALrYFTyGtEQhX67yuogEbNaPE
JSjcmXgjgtfEsxGgOVJ+I/Cs5G0yFC5maMAwqIcbErdNLaeRXG7L1oH/YA8MnCcAhRU309+UGTsd
kU31zJYAI8WStIXLBf2NmmEl/Ym3Mj9p3P5FK367hjOX/QHposunieuhaYv1aCAwx2E3FL3LD9VW
VAqQMGoIX77dM45f4Pn/GHzPqI6lvMkzTpW3U3ArYxpLWPzCwlY6wFS2yxJ/cW0xSSYMREjAM9qf
KVrS+0FvixCP6C/J6SXkIr+OR9HXEklGStO0GDBuG2MA+lZdV7Ld+6P6KJHiwU0LRCzVxMKQ5415
HxfR84fInO/4UqBrg8FjKEVHSITfOpD17ZpASecKz8zuTtslHDZrggVHI2rhUpyiOko6k5+gWzzb
Ysrh1KK8fPHeyuW4o0OmsHJVRIhfgGdO6lU7A+lamSdK+GiXZMI7AAlhVlA3lrrBlUmYJzZ+Hjir
PVPbjc8wPNcPHxFPuLZpr0uB6dHZktxfphr+QaCFP9KV8kIN2qTh/5Kzb9WKes/g5A5gQyHN5yCf
ifAXvwzBQBOOSnklxwQmdUX4+hVYy5Gv5CshA2J0c2Vt2cwDzbI4BUCTdhMEiJ3zTBaJosn3EWqP
lzFp5exBEK59Qgj6l4Duvn0l7EHQ7/lnlDHtoCvRxnuq6HH96zW5JEYzEwj7UglnCYIvGb2lE4vD
PxpjRDV4aSq9NApQGgUdJNPkmh7PbFtJWEJTmTJxoybccmUNGzMd0AF1tJIGnd/KyhaTgMUyLBK6
NVxRZG3vrshFEce0NFdKj+fkcKQbogUQWDLacoW2LQPEsN679lpHpkaOMY/s+k4emX0ZkIvcIzG/
ENvudjkVriXE7KV8EcvnzZbqv+H/Nyc07sBZn79QYHr/KpdyvwaXEb/n+quOkqGvwCr0CPcmsD8L
BEuhM/JrVxgkg0+oNEMWR76irdHXjhEJhVCf3QIou3Ved47SYaFzC+0zLCQEoDDBBXNIhmwEtgxJ
fPmJRw2cG8uvXyJxmx47QIXRN0sw4cV6s+h5z6mh+DNMYKF0ODjJb5majCOxc/x8m6VIbMTowgAJ
gXGvo4TqxY+buNkaYC+c3Q5GQ6ETt9wEzUf+s8Ec2jbx7Y+RA9OYx1YXAtyyAIFz0WnKenN147sC
OGeNz0BmBdIKxCxR5uCFmnXz6hrWlucOdjCUlj0QWEIq3qiek4e+ZW/DbLqKuZMcJdHtxzA2E2ak
nK44xqsbmMjcZySGqYABfRNkuB6fubfGn6r/3Vlku0Zy4c6RyNvEEdSobAEQajvYvZGvSQtlNiXy
y9psGRq/sDULtLBwtayAy34QPYsep+pGqPmr548vztPSibdcUwHPJcCQPscprYUFp61hWH9SyBgF
YhQ6fGfppkZDlDUyUS8BdONsp02+jAF9gx+nlayAkBLwW1Td7C6JxsYyQ0JMO9jMUy80q6J8p+Rl
oR7lUwK40RdpBAG5f9ArR/TC64gYlm/Lrz1EyIV7Gpzz/o4ZcgYSlTlNMc3MxSM8uxsMJRIr6Sdt
vkGCp1LbhCj4xvXf4g2id3Os3RmV8+lMOgIMQvEhqyA8rrioDq10PboFdiNvwfyYeC9mAHon/rJM
k2fArpdc3pjrXzqvk5jRyF5gw87MHEvpU11KqVpiM9NTXvqh7SqUK1AH4sjlv0WbbHhYb5BlVZpr
NA7/06a4lGq1qerou7nSZO+QjAIVfm8ZZ2VfOX+qQg8i72HM8M+hA/5mCzELSF4AeWcwsw7Z+bMp
I7mitiWmRRVKXtfJAmjlEBJtnW1IkNi7XrCofOrm+HVqsEFrQ5RDV6fxSaYS3giTQBbeeqjKjqer
IgBy2wMfbzhFueS9RdO2AxyJsyO0jLaj5lx64gKRne67hepc/lZIkxq8uuqepMiP5kzs71/vVlxb
Sg1Y4U+SMNL852znmDl8YRc3er0NitgNa6PqUaTWUijea62J08ANSo1klqAnheF9ByG4rz22vi/b
cU38QTM4rd9SeTODrQwhaOJ1EKMivTYPkUArzGz62HPJQQe1q23EHQO/aZkh/w46Pm2bHRabKXHZ
lH0chF6IYjbLcdmi1ti8QrHMbkL89srysLXaF2eEOKaDj6e6+amSbVCznLuxlEAaQfxzX3Xd/NNi
BRNssrc2rf4LfBl0rDAABdzbYcK41K8qAZTLz8sYkjXrIXi4DcWE9W+9DMsxe2ojHVVLMluNNM9O
E8xT8GAWe6dJqeWWSFApFfDBFQXSPj64KL5dSuVvgKNW63VwAg9ceUsh+21n17/slqvmkABqBRif
4r4Uhjs6A2eYANkDM/jg/asEWxKlZqljcXK/Q6W/twPBVIbDfGhvvvLHW+umn8TZJ+9ix2B1FrIU
QiVcW55S+yJ2/3a75zkG6xCxrLyYgR4Q9VsWZ1+5gFoYo1OvnwKYFHHB2HT2q0Z7gQ8WeR5cq9DF
gW0myL7CCY4VoMRA5ial87kRu6nGgErurTw4kcfL39em9bDSUuJ6p7PnZsAYPEiQRwqdL634VOPg
GM01G4gpZLl2IGXSmyMMB/Yb0PYwWh21zztiydSn0QVfj/zqWo8ny5HkfgS3UrAu+I4u4FXqYOij
mUnMSOTmFHQNRNs1jOd9YJqOjXHqZyAGxFROIL955J+6T6wTT042x/iiNYn01i6PpxjbsZut9yox
XJL2hekREscNLJMNFTTLNQLLaSJhBD1Nd22dgsObUZkkZ0KTZ9jU9eXLJaXGfuGj9eRq7MIJDEKZ
DwMgy8y0Jlb8kxrtwZtOzqcCCnTn9u+O/7vCHMyrGlhAcHXFOpfuzjCf8YXioxuNqXslEzO/wvFY
B9n0siPOZPrwEdAloCE8ne7dI0shfiWQ6fp9a5OUlN+chrXqe58memWEryysmB8HkhPugR/WI2SC
xEBb9GidohNPS7YnIdobOTygQtLoLQ4nQ8h3agPQqE57HN/EYoguAoilBQNS1uQMBj2HgW0gogAZ
FuQhUIfpwM39jeTjVi7xEo8yWD5erwz24cKS5053KpqE7UPU/WbPp8OAsd0MxzvCbzwTKBFnKFPG
r1xDt+pJoFCdHnlqdtJ13l9hRMegOJkU6gHLuHR3fBDw3CsYUnUk+D0uZ2toBK6q21TO8e/2L6sp
gv33uVL9w6EOyyV3ceKZdrLSzZ7c3fOpWlr5QQpJaIqmQ1aMDyG0+thZejz/T2qt9kbGDHqyZDSY
lJ2rKQf4NE6M86o3j31H7HZVe8hmC4ZhoIbbUX+HQ4hQQEF9vJ7KetTsw3NyEwq9rri9iuXQ0Z4I
6p6aSWGOxV4eWesLiYHHwX/rHw5XG2MU2Eu78BAJbkanDBPVs2EToxUAFfmmSXDe7tn2K6PTmCjO
JAuWccBM9B0W1GvBDd4kB5GLkbDzV3M9LlTgv7cRN2Da5ULrRfN1k2TkjGuVNAawI8o8zncwaSNs
bzO6zn5bBMopKHEzhQ/imq45IxhGs+Q351X5wv88MAtPd3Pq1lEEFp7c1Qz6LI0hyRZa1w8y5RiR
mo5Ey6ujZ6CA7ZZ5O6zhtkgL6dYL5QxlgVK9Kat8YNUKboaXcn6ghNIzNdgnfp5pvI9OzH1/HWmz
ZsnLQa0CWqYsT+3AAtbkMic55hqjAtBthb6QHAK4qBpMwVlNsOliWsv3CDhLybMSneGaE34dz0rV
hWH5F1z2Ox8dSCz7L56RXLm8/G+vrSGtbpExS/KL1coUjaYiruXbBadFB0n6jxdgbicv/HLIvx5z
dSbGD719ivyHr2I3LyP5r5D2PQOQjLg96sYDnFc+ZioQSo02JYq897EKL3kSiasNj3bD+u/guxG9
i+LL14HEuTuVXIyA8Y2rx7JW59Z5nthamvVcoHCdDoNZTVzBYz8DJxvB8wCizuXFzxFrKNoDj9Cu
5f1BMlWAYRtDqA4v/iEqwpukut22C996C+E9AprQDtarKtTQAyYEd+dynApjFlh9YkhCrHJGC8Nk
bBKyvMzcpCMTKGkYJZTXVuSjoCpCdnFRJnXkaQWoh5wdXY2Jm0Uk0uyfHguxr0n5VGaOyqoolsq4
nFnHi19Sp8ghK2dTIWASIYxPMhpAWptEM9ockCjxzfQGJO8rny9igJmCaBwLzxbzxvsD+iVM90A1
oOGm76yoehm6jFArGF33aNgBb34U0adGyqILx/KQHVk8KhhPm2nAiSDFaOiR82WuFZwSFtt9zZsR
6ttHKSpqasF6Jq3LrQbqvcN4fctxtnAHCCGQPlFAVk5buaKzAnNJhn42TGx8ce3m2AUv68sDfnuY
NWwtCsjsDkuSCq6wWIoXoe7q+ppU62J7+qnncwW5Zn14C7IHu6K7h9gygnCdkwblvPJnOFMs8hlG
sBMVWPhRDAS6qSzQo83AgKeP+vQO6I2smXLEB65wabikRWMQ9R6wRVjGtULr1sNrYx/Pd1j1hA1b
Xb5Uerl1np2P33GUZJAnKIJ7joYuX9C02fP9F8AvVIWAnT9P/GfJGxZbVGxc1Fh1j3jjuEtvDbt2
1JVG2IBTPCF3GG/zh08MCAqldWvjhI2+sVgupyWF7hvPy7safNt5ZkXibAeziuhjGFuzWJtLN+2g
QhnahrRC4zkwA5qnamplt+kXylkO5aF4v8OD4AJSTWAnfq6XBmxugwk4UhGzlF2bmsjUd5DIQmmr
l9glrXgZQNFNsJGbU0ec4219ta8Fvh/bIDDYyV3fTLBs0ra/RcMAezxq240lKruMwdIP8abJ6fOU
9pRRQ682m2qnNWleD3yI63FRqeAwNLEXbODFvcmL4vE7Mp04ww6R/3S0hAgODbHtaondpuD2QaZt
BvV8N2uBLBdVqS9+b/icA/Hfg0B6ZEue9vujnzVDlPsQDLIRivjlQ9Vi65CVoHJwOCQI4vy8936w
AovxfBGYySCUihCd4nPTUJx0xvRMROE0F7T94XH/JY835bum/RICXpbjLUvTxitX1tfmA7Ttp+x2
SRn0pklp9ihImuJclZfNp3jctCzB+/XCFDvNBHHVkd2OxFEo97iaHGbZpHGvWv9VMIpnpABufpPx
XPGNWY8S0oG63+MwqcdC/VxZaK8FlTw4JBeAiurWKWP9w9fJh8xtPYrQayydgZKo5w3CW3QKZyT4
2gWbymu7yeNwqI7k+qHrQqGiXyIFsbyHkDuSHfhUdGO8ttzmPc31EWapBJcecGnLtWcDntoQvkhc
Yuoj/lj1mQmH2MOUv05bsVUQNE8YJ2koRyy6rsPMMALdDc0K+QCneQvLbYj68QihPPIrsR4lVrXo
GruwUHq4gWoOZ2GF1LBF55Xsl2XKl0JvF+y43FJEScZ5uS6K+TmQHZ+boN6wG8Oz4QJTvsb47mo4
l2X68gukf+tJ6JwOoXbeSzFFmstoF1Gr0eXl4G5MKwYHhXkyzcsgpA9GHgvFSeWV8QYzMPVM93b7
wGUBpl3EahoZUFBOIaV4wSWREGEeu5KvcuNVRq34IiY3SC+np7TPyEBo9IOPEEznR0HGjL5PB5sp
vuHgfmUybZBJ/blRo+GnLRs1c6KLBQhE5LQ2vFdk98Z8lRbA1ns2PU6SRnL3kVLVW8PCA7aEEqJO
QhQ32NyqaEZSr/qvo4Tk0qr3sIwPJnqOYr9ebt8xHhif0zXpfth3/rishgW6qjK2JLhfjW2okL2n
MJ0iiUsuMHV2IOJjT9f0J0j0b2JghrCXs1mloLf8PcHE7DbwHRGO/AsXrdVKO93CZ/oMvbV/pXNK
RN/+7H4VeT03q6jyDBCheuJ8h5CSWoD8bQ7te5bXzmA3ualJmHrgRvummCIRMAv6FELjxYSzDYQ1
D7uyFbrSCCZKLepmT479RidDE2muS8JVTBqebtvhVHLruhpZN2aE792mXscCU9LJVG8dstgUlGgB
OpB3smLr39jxTZUQN9G5y1jAdnTeeT8plcCCJT8XcbHF2HA5D0scr9xRS8fW8bnFFjQ/EEnrqpGE
jzpbCASd7m8s8vTg8T58CCFmDpZsxY1WAqDe9d110K/1qwcC1dYXVVsWl8QQnz4bd3Amz0BY5xz+
tP1HOtW3ZHRIG7pII0DAjAHYZ+cGkSlNrm+CBecHbGIEId6sdbV0bCeMXkWngvCi2VUbVybHFv6h
u/6QQnfiktJTn4oeBiIe9nxrVndcQnrIqsMKQYzT6L3AxXro1+XGSYKLTAA/7nfLBPMn9W4KbA7+
RXS6r6GGOUu77HM1AuyYNXuD2BpumMc02swDruJr5H6cJyDvVrnL+qlrnvNAW5d2FVJrLIXcuNVd
63qXMPU+seWFFgROzCAUjGcnBGlS3kzQiPcUBFk2JqDxudX9nXzXMOYsA9pR6G6e/Z/KYXk9syvf
0MYQJ4uPOPLyoiIOgErObIvPjYClS8gdpRqm6Vr1ZKQM0v4ZCtC+ndLtvhc/jNErw67N7LYJN11y
GcCHgy0xI6vEQspbSvtA9snH3EuhQszOf7JUb4G2fw5MFoiWjZ3QFC0tRPRGXhjMngx7kMkk9PaX
DmDwVLbWzgIcziDD9ce7n6c3yvYwRkCwnRwLNZ6+wZ8ntg5M+vdA3LJQTRQjTnjX0/inOcC2SzlP
Sx0aHdJxwVPj7HfRxDU45tMw2ZVUQHXDDEbdN4F1E9aLwjg+uLpVpGV0fLeruO/Z+PhkJs0RvQ4k
RNcI6Ion5zGmLcUfJiyRXyC/Aoax1xOg7kGBxtB0LVhIIf0RTHmna8unju5n5ezmWbkXwXeuiWS+
NYltf+3MdSpxO5BeER5STkNSP4+hjzyfZx+sAWJHvHDtEJrUOJVvZolsVIbXeSRNiP2UjVNJzgYa
OKSSL5XUPURKpuTUOpSuAx40SAMcgHWCDneKfFXm3xUnbfu3+oDJQE/a/96kLTwev3wPhiUORsIF
Jbq0+F8CISm9dqSd40Ct/kkmm4ORRE7ERCMqEOs8d2F78KtVJVx7GYEAB999ZyONrwt45GJPMVfy
stX+kzW35UvKNJ9EY12YfaJMgmONj1hUMSEHvyo84ucTb2c1r5/ph6WMCJcbfpcNQr6v4pjl4Dam
uEqV5ar1gNGUrOsEz2vToWj/y1nxkK+IXPWa0TMN25QieigW1SZzLIBn5YwKe5sBB9TSkHDUBNR7
nIgqil+qOqNe2WuBWHwj99inXfB/5G8BSQX7e2MzNK7ctaAodhb4m8Wh1TnAThqWXgriuyAuQqJy
liVJpcAXaFadfyIvDxSoOIPbVmVKUuY3cZP9zgs1BNQhvF4lCL02N8PscvVnMhNFfVBkrdyGfbmz
L5vj2FSBIA0jEwsfobzX9MaPUmEFEKQ9ZAgSQFYeyq5fGiGvyQpVfErR0KRhpW4B/biE3PO4Fs6j
Vt+0m0CJW7FzzAe394X6pukCEtS1jxQ7tmv0cJuHJ1WLxkORidmYMESC0dda5GKUsDogEyXl7LYz
RE9iXiBDGpUbHjQLReTkImHmRQdqzUtez0w6OZ9VoOoDQCH8REV0xNS9PuChOvSGWJ7G0w5JamSE
6p1WvrGhNOL1HI7nZKxD5RrXyhTWip0ivMzJFrtKxTglndDzXHIyPXOh+xOet1hQ6cmhmFlTLg9h
X/BP4aasf7ZXzersC39HuiT11pl4JDYnpLPu/LQdkFjR9rggfZ2GFNTPGxz0jyX32Bkhv2BV9qRB
flr7qGcluYrpF9U4uMG0K8hG2w1PuR5CHhsui1DbB82MQiUG0oBuiSrM6za7TEZMXXnpK8nEitoJ
QS0uz8yzOCb8U3iv4fEVxzUpFOrZv4DtnJ9eT36Ht3sTSDp0MGAZQauCFBRkDpAeCGLINQS1/cBk
4r5y+EWNa+Ers2tR9dFbXXABp5dGwYW06ft36Z96iYVFJx4DlwyYYrtPua9tkbS4Ig4YVbAcEZgc
S1Zx/5YOmcmRSUxxmP3LkMLATh+Xk5KnIRZRkubwqohzHhwNtP1DOxiacDrABakLWRzUuZHMcl+Q
Y77K3sivIbo33BxSuqhzZJdwut7Q4tGxOJKHKQKhJ314/9UluphAyHDKmfUXUm99K7CVPWeXVCqu
P9WajJ/5N0wlpW34XSuTLRFkFseP8ztroIkydi9dXGd7XF6QfV2a472kK7EEjEZBq+urhr80GbdL
MUFDAeO3xpcRjq5CYH3qpQ68d66wtC2Y03JcgfynXR6zzvFdZy5nzyqeKJZKAEb/qsB85F2Grpls
vCNY1jIUbwEg8Y+mtiGgNMTNNYY9UPysyI71mDzKjTT0WyVaDQ5ZwvQMAUDPR9vpYF3waDVbrDRQ
sgKdgRxW7KujF9/7fGBK8Untz6Knexu029NqS/Zda02ZA6qWVOk7jjhbFpYYl6RI/0LN6Gej4tOo
bts6o57XagR60ojrQxjI9OQ6Rn90TTgctOAfcSNZNW5A6cbToP2Dj6u5J3az51f/WKdPoOX/tYBD
Fsld7BXbRyYniuG4tUiJXHl+RYyi2nAYJZljJVh7YhMmVSlOl2mJHoCBuD2VIetT1dqQ0D1l1zx/
HPcmpXXYKjUFCvYfmsK4ZbtP06ThF+iiYKU7XdiBPm0ylF3KxUa5nCtV+6di8pt2ukdtf0MU1/w1
RJ4WVQ7M189UgkwD3cNkQ8+YNkCIiR7gUf/naROXBlUE5Gn7ecoEb3s3oQ5l9AfpTSYsAxXfueDQ
tqy7KSDXzNLJv13nuvVz7/rwo9+bWBkQk7k/fg/xMDaCrcONfDkNmWp6PoXDEV6cN3dDmoJhAubN
k9xqumbkFQXCUPl1eqXrS/MCdC8jlyVikM7Lql3nlXGM5xZmT+0ltNLnuh3jVFXBJCeNFPcDN860
cUiAJR4KHxprUIihaDmISvkO3mjI36T4v1YqWpiluZAYj+CyR3bUe5NB1XXGvvMc62R5ammUgGgl
3bDnuT7DxVgRID/g1SRyIXVkHJW9w6kkmuwvc/em4Wynj9jIWCODrPb7vgwt1B84oxAaWiFnv1Yn
8YFQHN3c2C47GrfgLamGl4jmHh0UMgRDx7YqEJH81Q58iDQWDM6t6Y9fsSiJ+ld2jmQteAEhA3I8
ST/uLlBpzHsFB7otW95yT3EnfckMra1DaIi4x/BnEZzaGzJOCMTtO6lh3d6vgz6HoZM5mMyHTn2e
AarKFuSCTc7eIr8BdBkFAUeg2lyBf/a9+uZtKgc1UBdaCIjE2o4XNXwfPsi4cKb9Sm5Pakn6A39y
hJXyWhl/tVdbe9d5Y79Oxp8XccbpvoV38TU1HFbgh9M1YfOKxcWIh/NYSoHS/SOg9XUTkdrVa9h5
H0/myVv/ZNYt17HNHa2pRSnP6NWvWDY8qAT4X9YbrShqFoxMiySy6uO0JYoSoZDfsXADvGy550vk
uvpIW7qt8qI59lpaENFhq/tG8Hu1IT5RmPY54vJ1Se45dHpSPn5C5DsbpP+hYvJ5zX7NbCqeAM/e
+fZBEK1k8P1aGj2yMHRqdRDUgB2c6VNcEakcZTnzRr6zBbz4cIfgat2CzeR78/7/HCMYBaJZULbN
Gco2Hs+M1d839i/3TomPpyX8lE9G+ARZ2aDWdYjbDr3Fm1Lxlp4+cHlSr/RDB6+K8ZAHJ6Q2Y0oU
agpvYc+5yce7ZLFstuITfBlyFnfhdB5RLlyTUp3/GQipA3kQIsD595DmWwTjc42czq8kEsgVA0dQ
tR9LPTr3c24X8nRIuGYqUptaaMOdi4MGPs2VorqFEGZf7Bhjk/DegAQ75H3K5112f/Z/ZuUjXlz6
bJMn3Md8eyJY4+4BjHP6Pff5DQQ6Jn2B/gDmzIKEubGHJRYgC2vApsov+9PRjx4x1wgrPtGRYDZL
8KRGk4DKSXFjxQGNNwAdMuV6n4gA6TRw93Zpx8EKqsyBESZiwwGu88muI3/T+WgUG1vuZC4GmGCB
4w0t4NwYgEVa1n7x0r+ZJpGGihPlq9kihjfffens/jxFpIRRbtDNclyixYsih3m3juTnpPeQ7bzF
KDjVN12/gKK1VE+Daa6tEiXSYDp6WP+1ukHAQXelXi6sPezowxZ6WKIvcq5P0qeAm8GjufvkIOOf
Matqt74QF5tolzfO/Le4sVARR1s3XicVBDV+JhfiVYVg25X5FfS/86jQzIjWjC+rVtQFn68YiwOm
5e8A2GPfTx4HA//x0craysCXuWK0cxff7QFJfxkQJhr2Xxmp/GtP+9O7pZS2ckjaC9+YlSDmfxcL
+2CEDYNUewJaQRXdolwPFv+AOlWriEineTAqvqj7YIQh1+OlfTpbrCDaZY+5q2caBs9p50TnPqOY
McLfYtkVTaSkzZ10jyVyi2ETjnjgyyHIylm1335ozlMxJZ+ApRw+9ns1aNFZbe5EvB+lGe+xS8Kh
uFYxygkHAnY/+k4U8NNPZXZfEG5C31xoxU/Y8gSh1jRoQ0fpBc7Uurc+x8dnMnRuj+O7CGfbSloZ
q8i6QUVpB7atoWBDUVJC034IO0EEXJH+fCdzS4zWjnXjR/edrNOyeM3iF/YbF7Pxk4BKxTWq3f8F
5aU2UlBc7Pf3qVgVACJJurGDTEaZzYLSzExHQ4dTmmYxgHG6ZZ8uz1q6dGelOAHXFHIMJl8HTjdU
9IAcKLrp8vRnR6l8IvibOgvRs37RA9M7D7rzgnDahdW2JtgiYh+ij6Uupc6gxWmYPspCxSBEKAdY
yocbTqcQ4fcCUUIbQorBMdVH+Xc/ug1Y4zCzB3K+XcMNBmtzkryVSgcls01GV+MC/SfKZiWO+IMY
jtIDjWg36fctqzfMOVeu7apyqMQdU6kWD355CXbuwga5yW5KFHkv6WFr02tTdtIgab4nwhxvtvJK
cpmmPCYtwmWT9qrIASSsSxLej18MUAxzAYnpDMsMcVI0cJyBPCbiqC//+sTBTnSrcHqmMYZNxEQM
K8Pk2Do93fIkv6UsFlEETtu0UwrqLPX4isEAmj7vqo4QsPQ3Pi80Mj5S09FmZ6bavbewDbcQFWuG
t56bqTpoej5GX4z/bjqFW0ybf7lw8cTXNL3Eyf8fNnr8aET9SWDLAiFafpsDYjW8mUAvuJmvbY53
aXPjbbXpGsvmEmB29UaZNhuPMEv17KZHUDZuoeTvUOVFJrRG+IMLcubEIKebrRbwOIVOlNddTV+N
WurfdGGDwWaMmp9Sh5+gbgps9FzYiEEfoW++vHcRrAPL2SYQzXfvzRBRZoAm4qcecM+ZNHoqFscC
Ok6GBex7lYnZKTOaRsuvAEOv/1lS3VxVHld3FZEsTsAgligzMv13CWoNVOCf+K37E3Gw/yp11YU8
fCjJleOVuiqClRPLvtnW8EwlIDSbP2cXCqeEH+Mk6qp6jE0o3gY6oFdtQuPx1bn14/GD6pixyy9b
Y6vHBMUr+rxd3Bfwj3rhDCLJecUIWzvLfRZcb8DTAJiPaKvFaJ0jwyYbSxp1ccxVSg6FC9uQxqbW
HwPIqH5Gn1FA51Me9+rwjryhkqwLZrAXbigNCgaWJM0eb6vcxTnD7SAoql3KDgKWQ4egb3kQOdFs
Rzfijh3NpbPt4ZY5ZlE2Awz2bND2nzyHTiKth7yJExvm0419sdYyxU40ap0FQxJYbzcISgHWSMbf
5lrDJq+PGUbnhlkGXuid8BSmBwiLN+PBDNCIPAJEm5HQ6pc/nfVunaXeCV2AGqwVjxBcLP3uzoyE
+LKWHQw9SakQvF2x5+Foh10AVbGn60Cuga+DOrvxUJzf1tFnzYlmzvpM0TUTwbntCoVquXsnaqZe
62/ULCe6jcvcechNTgcED4dP+o34ADFUpZsZ6Tnir2ZYOEu9tVa3kPizMN7HcT0d1k/ohxe0DiCd
ncz8LHH10DwXfirkI22Mfuf+b6UoufqIFrDZs/33/eMbWF3hmP1cvlYJXtQD6hGJhWzIcREWeqb4
+gkE3lER3wQSm/fe/Sxjt46M5lq0Pj/gdmLR4G6oDIxjc09PkuoQvWAHE7PO1Xsfz3CobdVL8HSs
6dk6Aw/JXO2SWAiW1nbSL8vx/cpy171xmZvkWsCAEDurxEN8xDhqNIYZTD4ADYH5jIgeUHcgnGu6
jFj9An0d+p+gcTexcvi6rZPdRykPbapM8e3MiTo7cfwuPuHrNQkmMl+P0uy72oyH0lgOd7VhEqeM
z6IZQWf+sqef+0sm3XnL7flz4bggvuS+nm51b6WZW19ZKv3CBaaOMVS4FmYmLpyDnoWPhwCENkjM
EFRuWXUhz7UiJeCgbKkB3B9NRn/mmAFB/kHvrob9CpEk8SRDpJK9nQY0Pr32HaxxhHvgu23uFoYp
Zs+J5jprBw1py/u+cu5ZLKoUE56n1prtA8SeubCRPjleH2LaPHqCdGe4GxFWLJkxbLyb1MsvUgnQ
iOjENKUj6JT4UmcKhqipdrzFw4rGkBwqTDsnkP0FQCmPJbO3HMGlXY01rZvJvW5p5QsCitsPEO/g
ISOGVJ2hlqYVQb+X37YEGdLckSYh+gBQ5Tj/56/7C9ZqE//v9n3kLff3CQ1vcf0gumjjnWqsrP9T
v3WK7QVNMN1S89NZv7WuejEnbHhOK/DMWeq8nret8ic9rxIM35Z3VXs1yQcllah9djbhY617VEZx
P06YPBfCQF/3IjltOoRotdth+gV3N3/Qk7nmg9ntGRPOflc2sqOLMmFqgYGsl9N8ZUF2tXfvoFpH
fRXDrqdN/4PpBB3SLgyU2nlp3Fr66A7SPam8IJi8AvrBlRR56U9pmvbd8tEje25sp99R/WXrLlYb
xHShRj13d7SRwChm612eIVpaDrNX4xOMrUPGolbrtydKcgXBRfFOHDxD1s+1gBVfiUBnVJqz1gGW
Y4ugnYVrVw4KSHxD+t9CDw6KyNgbQIns13PP8FZOdNSYFfZKfh9NiMTx/Mt1DPyEb8htWZcIB1UL
zeSUYdSaBeqaAgLm0gDBzII2edDlagEm+rz9kjIKOmUBD90ZO3lE5okcKcvpTRfgeRFClrg7nGVl
EFshxpa+2cr/nGrbCn6K0JcgrJQ3pDhvmvJeWEE1AWWtsfDu2CMO15lk5StLm2J0d/EBU+0T5lDm
PxpLH7kizs42W5dpgkzLVJD7J/deG2CxQnBLRuXvVY+/EaEEca8DWarmGuQoat0f4ELQY7b4mot4
wV3EjX2mgP7wbg43MjmRaM24QGzso6LrQFkvyy24ERwNfHWe4Xb9vTs1vT6JQQZRgzAhLtgDTfWq
OcOHpor9pgItrHTYwXFgBiSq2EuIfDNPQyJWgdU5nIeW88BrzxejUMt1m/CWDvHT81MmdC+vvoEK
/M7qCh5XGtyT18BI11MHL/D3QOq6daWixdVVCq5V/UkHNgwti9VIWymVUloNDQ+5P+/DhClmuRb3
qnVscT4OrQtBAp9dQ+3uW8CP8ehanISV23ddszJ+IJ9egyES92QoXescjr4T2ABtY1viq9+U2l9g
6+gUfHOMJ984F0d2ZE5++Iv+9Wlf2HmJKVIAlOjrK9RdRjHhIltbrdnspSIUSny6KxIsDy4xEaUm
CmH98i3viQJ2eZr2egUolSomNZNMO3C5zrbNqxFOSYiNpLsfE6RL/nZ5LB5rzlcvvZnrdZTU8z3d
K3SgIJHrmoIjKCWeMbpV0NaUxeOFUZWZgiADSgGyPs6AhY4hxlnWhc+eUAY0ahzogWmUX7MF2ZI0
gJnXPcv+GgN2pCb7ozE3l1HQI2R4q1bdUIxabZCnwYuPHUFoGWuAhdSpl8BRhngGGmvvIbwPAUg0
D13g04bhXgowCNN73xGMI5prG8NkIhrwfaF2PuuR88hZtnN47z8TKtVeUjMwBJQdrdHZ1lJrbfmp
8eDJEYihNOxn0Z2BkCKaG+Qd0I7b6MQ+0QeS9yt7h2+9i7/fqGK5xDh1GQhFt80CZtcCbalSNsZF
ma2RyUQEKoojcF1JvKjSeU/Tuu+fwcvvvQba2PGTgFadDAxCW9YTfMSB+4vNCfyIJdFMMefnyTSo
ugZwsf7syvNZl1OeFFWk0gjfh4m41wOmv8FHpMTyv+EEBkQBm/eugp+ovTzRwbIadzIjuPwynn2Z
UCZj14MiFpJ/+YFDsOJprGRBT/boshUMqDBY0inhQqktx1agNGxB+pDPQ/yfHtHMTmzF8Og8cytW
adJgbs+ZOpn1jgQnHzXBrYszyYZOrebvxTVQybZ1Rh5M9/9KCvRFTDnLe2jYS8wdydME/8p4W6xU
HR0oCrqdNv9C/8jqqMxxGbRUiMvmSCjJeLsGqiXAcFmDgcEyNkrJLzGxLXnkXcKn3qyOoD4FTV4v
mmRN9WxXZn2Uf4y7KFB6iWgfQd4joaaa6LtH/IdoT38rVBqbfRIGaTmx2ZVRKa85Ro/c+QhiAZIO
Ovs7G52yhIl0wu1t6MDs5liSof34o322Sj2wmR0rAOfE6BqIAB1rjRS3F2iIttr5NtYOB7Sg8ii4
HzJGZnfRFYShbHMF6fCdmMBJuMSVksBTYx6CCRL4AuOtFMlv2d1S74pNqmLOu4mEEry1IITYgvJj
1Ca+xSaD2BCxszYbvrqQbSrG5qv76n/FZI+xMoXeL8pfE9e2ZIdpTReHITmXKPkFtrddmhXhsMx8
IeXZRL0t+84Bo7dLnitpEydQo7yVNy2r4PsaNFoxfIGt9V4/aqfyx+HYyy6HvdsDbXOySEfTxif2
6NsVOLjF4Fsj6CIHj8PvccSaqMCYULHfKX53yGh8Oe2vOoYFeEH7jlzR79ahZgnTpI/2uXc8ALTi
9ISL/I1ksSLVmUKAtuyDKsjvTldzOMkI4NJtr5QD49hOfCebaBABZlcFmFS/T25WjKJF0s94clAb
nRzNf/V7fK0D2Qf3MLnL/fhXZdoaTiXk02CzVpV3WEi2KyysiQpuVITJiXU7SuMkBRgiHbY/AddW
8Po3d9vvAgapYPJoOZLXiHgGFdaeKinkrMN2tvAofXHkpYz9yrgMdHSHh/YSJhNyt4uvqlR2gtQv
3xXsAkzZVAuEHZEm8RlsKsl80ZfpFSW8mAn2DkIcOKPYF5x+2dqUgaPS7rAXiG2E5q/xjw5SOsYR
CTA3OTvlfjWJe09ZbMpGwIXbiC25Ub+s3xpcp0phDj731lr0wwpzpM74MKKhqZlJC7jZERI6QkGw
dUrGG/s+u8L85uHiu/QNdBNkAkFElbsQantKrHK7sF6X6ypPXW/rYPCnFhjpWxJCQARiFRbr+F2I
KsYbJ1Suox4xw/YJLUniLDftK6kFz1st2j+VY9Paz3/JYiEJ8tL95lR/rbQzsJpZeswldLQAP2yR
U3iKUlaicA/SFCXOx1BlT8zB3XgCDYUXiCmCbxOYjxWPpXa+oTTYWoxc3o1P78RJZOvHi2z3AJEy
zJFiG3LhmKgk8Vqq81wkgWsFWBftMDTsrf/hAJoi2Liq2SMM/yDTO1ZOSIDlfhC/cQ3DIzTMw7dS
kXLN5YKcDOhyeXe0H/l+1eX4qVjudECV7lYgnXDT0yazwoUwaSOPR73VQgikAo84NP+nz0OFTKoQ
wp7QpZZDLWd20cCCOneOs35dyQsRWZFVo/ppvHxzmOKRY/HetnjnB8j0yKj2T7zbL7VyqCZbtyMG
CtpMQgVqx4RhnHGEohVxU+f5F4Trr6VdNXBrCTDka/92Gc/KYqyW8smQ3qsLNfc5uNhomrp8jF4l
5LsnszlbcDI3bKNPrAdbyLbxkm/QNa2nThuMGTJ6XR+rAGAEJxcokEhRPyJTleEACaNI+PX1nQQU
9Y2hBkjD/OHPfqcySiCkuFyhBNDnVDMrbeVwwR05RLg9sMaYzHMLAGJ0iaXwaFWzgjCM/qp4QV8G
f/9Z1JZG+WxE6XUBkc47B8+1KEjz32StIneT57JcmnUWsMNj+H6Z/nb/8GoB4Cqp6viOkJFJfqwu
Xr3F/Z+m4TIbqbHjy9ebvpLWv0kxI5SktSsIbj3AixhvPr6CLp6REr7lJmvS9LmU6Zh3Sx2xlJta
nA2cw8DgodkPasJ+U8aokqooXMPLjhK+0rM1Nmgq+uONg18czd4QTxDDwWTm/KiE8k389gwxVB5p
6smZuoLPfmTyqJ2+wnBy/k8YCuLtvInjX/+OzuEBrVjsqX/G6TlbZc/sC0dFgYoluPHLOBZxb1Q0
fA9PKhqyMBBMZeg1Fno5Jb2DUHNglr64Mk+X9io0ZopJHdZ4+iGTivz4WYi949jpE+cOwK4QBQrx
zOIqk7syRTF3Fn+S6DCY9yPT4ItBIiOIZ3Tp7nxt5M4apPNIxGGrsN9vef/BXn5PN1L19xrJ3pp3
yzVtFbf8+CLzcjuUgzIXtYXiogLyTjQBsjPQtz33eYgxjCQyaAxbNEwqXpQGrlYKc5IhRd1DAf9s
HpF4QKihzoxZBIWEeMbw9SNNu+s5zKEHmycqsaB4ScQqKgpxUW2z/LXiwSJFb67bZEOBEL5mbQy5
qOtbRadJ/Co7h3YRQrv7XTvg+nwjdTrhaokUklp70FUWMxwxp0N8ghEYPvuHo8VgTD925iaFTP7C
jPbEcqE9gAHuyZZZU9nlf/qoK85sz8J8z1BfHjMCo8NQiKnlgn9ZHRM0yV7JZlSxu0sVTrdWjZu5
haoNsWW/n5aDmfRd0GqfcE2CuqY1ldA+jZMYHIPQMoMbxouznxea3CLZpHBO0anXyHdKve+1auut
kGq3BLZUA4YnB/ZxKNlOrhrLnrXT4OYzmJL4ZST+rFz3waTP80wyJBsYfMZ0c+O8i9N/G5ugLmes
fG6UjEN2KTMQYG5MzAacnbzlMq1a+ezBHkXlc7b/ZsuGrX4bvHgf4hityp3jhpWd4vCKSarlbOci
GFiYm4RJjDKQgD3O6YXtaSzt2++S/FEEdT4OL7vzLS/b12yddqmOTWrC1pWmGxTNxWqKthLedNHK
apdFxVuCZuyJNemB6DlPChAjBx/Dxe7oLUlh4lrTR04eUsAlZm9w+Zbn38SOO6XRqruS7GFcE5C9
pPBcVqthCEy3J1dlW4ALaU4TuIlNlJxA+eXSt6QAhxbn5RROBgf4hwPyDQKLtSM1YSsYJyNHgPDm
4eKBejo2DhQ/cgjEmW3uu7wn/WgjjRFduVvywzdWT7HBOJjEVI98Yga0KKe9V4ZizpwMzhIv9dkR
4iVltx6IsK3tO3RpazPnK8ktuYFXrkOHcd0FichCepvBQHsBWCXMuNGlGtV2JHVqvFKDGE2ydlVm
CpFT3kcEIovkTDH4j+2BQ2/kkM7+Lc4ydz/AE3sy7K1ZILCwhbNkQDuY2Jqv53Nt4e9z7JZAufjM
3D5mIXY1suXEO5aypkKqWoP6kWCDk1sluBCiWSO5VJVNPYkpXA5xXeKInGg3icU6jwq02aHvP5T5
bfIH9uw0pg30lWuWlQ7fDHgLqG+BZVeUGRC7PWLwuCnvBLEfK8airFGdIaCOIE4dAM6dJTn7Dznt
giKmhkNBow0AkM3bPY2465756G/dO2AechHA8uovvIbpD/igg4P0gV5qh+puis7C/s2UiFBzy4co
Jso0RLP+WRM7k38myNOcAD6iUBxg5/eDVs/NWa6g2Pz9hBRAaRZbV8Q7W/yKa2TjH6j18Loc235D
5IAz6kZavIo4I2RO0rTWGTjB8Eu072kGkp6elMDFmBs6RQyl8Np1F9RgUBJ0W3ZoNhFvYYPhQpKt
Vt1uVSRISUZ38z0wLMWYi84fmYR8MjqECTr4yMJeMuPAIDZbSD3dYp2xZEe2x8DMGyqE0srkU2Xp
3PTxadqmr2yEghQhszS29dZ7/VZpj5yzBHOmmGJgZXe3P3YtELvog/uuL66trwvSi4oCtBYkDuUv
F9RKLTPZlNSLcJuK6hZmsyzT9jxWnT3CrxkiHBr6OPvPZSfP8EmUYqUL6NTkrzTdfJYOs+0RKAiv
fGzKvPtz5xDRqSqCmAcOhjQSuv7yxBZMDe4VT4FC3+s3L0NyqFLLWmOymFepmUOaz71OC/0ZLbdf
v5qLjPiceMwrFOaGoUBStjVKBqUQAnxsKkYbItZPvl6WNmGHBa3rbeuYHkxh/GQ7f3QF41AWx36B
TWqdN2D0JhdEDBZpK3QHDeI/DA3wm1TJWuybOd5GHUYSOKkfRcQvUGw+pUHSDwB/EpnlDbHLsj5j
kLMvbStgmsd41ROamUxkVKfEzKHERC2nnCrDi7goLfDV0NzDOopyXS7VQur/os0Hx5dOhwNQNGIm
p/1lBdGAN8dTRCAqu+o5qRbdPEhLEiiamqIVrIPbMcDuwebdY8bsoncAFyTS5bOvoyKI4hvzzeW7
VOkYOMXxUMUxP4QbPYw5x+tpTowsDlVZU20qn5Xh+GDWxLz/YnTmelhlBrXKXFaVCov+n0giJ3BF
opP8laA9p3o4uf479QK4iAcGRXLCx1/CgOQBSX7OwzjEVCyaMYJeJgOBMGyLv31dZyGT/JfcN6HR
bzORN0tn4MKXwHThKOxWZzbePl6mXiJKfq8jB/KtklZk1FpcYxRylNncPVYJ8F9ymhCz+t8TAx7h
7nZCIy7lO7P4bBKY1W5ZiDvAxvG4ALh1OY8WLSX0kvOq35I6QK8dQf0C+R4N9mGwudr657AmtXB+
sj7e8yBYh76mT81gDdYGNMZYhBJBbbv9pp/EoVUJjAm/WCUCKSwf2Gu8uy2rsrknbMKLRVlbv+jo
c35NDcmuqVN6wY6t/Lz2W/Xe3o5jI9DZh0w/pAF/P0+7uWjTxOOPIzbQ4B58J3io4kKppOk8TNGi
6duQ3uy4FlCFVCPQqyj0UF+gzLaiHeFdux6y1dCeKSmC2Q9Re2D5DNSHFPoMpd1goYmHW12hHd+k
Ga5EFA0l5KXamSedmfv4+U9eclLgXn6ptnvh5bHJZeeN6T15bf+8El21cyob7OmGOAU7Ke/TE/f1
EnapKLv4cjzWfer1Z6OMzHoDtxPXgYwyyMxjpXTjKmpMxdGrASxzC5KKcgkYfiFToQliBjr7PqAM
sETlj+cd8Yeb1Gj1tJqduBNqIuQ6sioUqF/mZ8dHttQjlzMKY3ea9Fd+CT/WBD9GTwrDPjwccXhn
H7D4NFSSccvuTUHPwnzo85xqZ1y0o+BnBe0VSvbwKelw/ps8Jaf5P590s9BDPtfFtC+I9n2hTDxT
b61A0UxLGE060JSsermZ7YfLtkQgz0x9FwpLJM6JWB5DhH1Z/rDXd3JYGMkOzk9u00IfwA60x8Ya
eFu9ko45W2Gmy/hgdz4KaabSMuaUFqdwbfaccjqC90956hCLeLMu+YxIPUWCDbYH1lrq9yFewPum
Og7cI17lVN8uqvPLvJqFEz5x7lFoVc8AUauPBrNf3REscqI1HM2+Mhf5aPHQDwO7NHiXu7GDPNeO
duSpZOrL0yhCUJq52mtB0mMxHOu41foM/dAkXF9ypbIOhoMpYtk7/YoMlByIJ6tzGPMXjvaQ9yUs
qw5p1HGjbUeElh2hyP0e3Z1+jN71zMl3LyODSenAhfiuIAhKokbYYVHnuN9jrjyRip1ir8BT2tMk
6WffxwMr+KCgXfhxP6zOmF4Dza5BiJY6UfPFwowxi6chjB8RSuDALqxVRm97qjM97Krc/TKnq80+
GPCekb+ZwX7wloaHJE9q2KIuYySkiJ0bAp7iIqcwavPFmwmSCyVg0TjG9hC92AOOYnBzCNvb/1L3
mWh75cNI4vgAAdJGAuO6oQuJNrWaj6KoQpzCTScwhznqAYcD/YJyfiD00kDZCg2qEY0v08wbHccU
0kogbLJpD6fpMr6Sd2ERl4HP8jzMYZ53XkLakkn7+t/3gSkFiquXIGvEm2DuWYWN6lm/IdgtN8y9
Oe7D1qfGi3tDIB9ML/NLwCFJs1YAstVDmDOuCvTRX77OOdCPOj2Mi5OEFhD41F1Z0mxolTNk5d7H
ZqMgsQwUGOb0D/Y+caLmIKfZReJaojmZsJlKu154pqQsUPg087te0DOXxDltKfkUgV0ZRgUtNPcH
gW2Vr//yy0cqllWFvH/F6fza9EdzZgwDOdVFKgocCokKQOlwqiwTDsnAz0V97BJu4zEZkv0FjtEw
LpB5ICjj2oXTtMf6CqN3oIxhFuFLcmclvo/qztU8w4sI68I2qT6SfMapgCZEI5I53az9kZHaDJ4F
nquL7JLTxqjlTWtXfqqZLLHBast5Jr3eBWHPKJL+vtM8i+3om72Xj5JT+abwDAwgdYNGCut4eiv7
FZ0F7KUtZR1VDYTais3WRdNmuxl4XuHOgY0nVyDjpyo7ZX4G3agt6e2w5N97ES7vh8/+UYgTljou
n6QZTjJWgPc1hehhJlmqFX9XGWi5KKjLx0BzsmUtMCyoK2t1/dh0ZsuHytMTOqKPaWzsncCoSbCg
4FcDUCF3Uzdts4qLpB7qF/x9TvfwOT+e9xzuEFAjNE95RHskpeG8HdXM6WT9oPtK+k6K9pPI++yM
cbsGddoDt9lnJOdfkM4u0ymCRJ5cAg2ZQodP1DzDvMzhr3/iKFPQXmUFdoXU24mk+8TY+HdGIeFf
aShRHYLdnUF9B5ePscZT1/mBp+CFNwBxEBz+eMdsLPgNZUK0wy6NA4pcftC4H2JHO01SFkHzpcAr
rZbD1snvtVeScv7touafYcpf9bwg7idJtqQWJcmwkdeb5aLXXJfJZjSGW577fM3PgtIi8nbs6GM8
p3GolL39teprdHAwXHp33JLPNCZm+T3Rd2fMWRryUy/D1z8JNONY8/GJ6vJMfs4J+AOnO7SKBPPs
HbSr80nbgQqsSvnv9gY7+83yyX8zSfEATabVT2QWHXAskudbScARvEYJBfB8FfMXdzPF25Ly0frj
pd/A7p3oO/8M+V81oIGh/c2JUxOk2CkIXV3m2hC6+obDKHXdeIOqMNaXdGbaI4Xq62mo6+sK8Gxm
8DdB7L/ewFs3LPV/lOQUp4w39tumzUpUvn0K62FFtCUYXpjtPMOjxRrwyhVaAJ7CLSj4f2LQEqjk
cK5sQUT68nSpTCuiFQRZPX4zSVDgZWmG+bGL7LLneNwtfsrtJGApffRrkrLXmy6fIy4gVLuv50JD
sxdyHDzJZ3Ckodb+2YC0TZqzqVSqgwEUwy7Plm0PMbpVS6jNR1VnJ5wzzOsFb5c8lt4U4YHSpe+F
FGbB/cBooxjzxl7r636f1D27AFK+ncLseVg4gEssptFQdfIFSW8sZeBCGwFUIofJyiEiyRxuAbsT
1P3U/sAF6q2oim7KQATFnLsAtH79Zuv9We0vJcUWfXKR5EP2lffq/x0/wjEBherb3erROi+jKdk/
jWntwlcMyHtxD7Kz/2cxQR2Z6t2e7Dm+LC2ZfLuw3Fbo9HzqxZ/Ap/0qWFia3E9Ht/uk6Hc0UsKU
WoRg0MJCxIO724lW+s2IYXD7QxTcjT9n7/hfOytIGcAUXHdsssUtj3E0WF98rY852QbG85YR3U5Q
Z+RsBkU9AmaV6voIMubvZEQJvilaqf23CFzGEVnyq/vL/CsfTG7GIRA5VAOdlOgtfd0o9ciszDYF
Cmk1r9Ro2eH7zxbnosKC5p2QaJhtvLCxXBYe7Z+QluJc0H2c3CEdpzqT/T3+au+rjoBgmVn7oSTU
RyiV55wRS+6UeoaMafs5zABQvNIusmkkt8e1FQOb1CBe4o9CHha8TQNMbT6yP+KwucPreO8M5arF
5ZIecGDnA6gUoSJzz9OifvmFHQHs4uj1jykf7wOFTySiUowyXmXDdHyp6Ve3pjY8S/t3fN+ymbU/
sjoLPUax1CCwvd8H1cJ6xb2KHFiZk89gN4c483tMhCzEtt0PlzHeopgNMU1qC2WXKVjDK4PcvXG+
z7h29TkyYH6xyJhbtlu0AUUoyHakph4XTzofvdcHJ/1PyJ6p+H0theftEplc5i6k5DCtQ6XCPy76
KLFnuUvR7azZ7sMbXL1ekn6ohFVyq/lvniB9/nVGe1kK68PYdVzEeT3YMu7RrhRMXMgbQfGE/PUa
S1E2FvZZIKAmkMqjqmGAwccfA46ypik+Zbi+TBstbqokMs1nsiqJCQnAeyV9KMGEgS74ObWm1D6+
AQd4zPqD8l6pI2FleTA24xX9kW1H0FonwCKYrAROppe2eKaRRl+8Z7YN63jhBQAebGR9t6UavgzB
lbSJlabFxqe6j1y4TDPDoUx5CbkU1DBbYdAGR0mNCz7Nnfa9BaxlJTx8LdtBD2cirO72uOJrpIlF
MPETC+CkBn7iPzM9sB2RReCWNYuHRunxX/FGFNEhEvEgNp2xxBO59dzpRzsxugXa1mXgw7DMzagl
z2BVqceRLjq9fZjbU7UJCUcAw6XuHUmj++V/L5c1mis0yUbMXWlbyRbAvWN/062HQkYcHjfFu/T2
OGulUBf4ZB0pfj0QfydWLGkUZLwB0RYPMAshmNseSJ4IhdZG1E74lFNzxr9bVGQDp5pLv5FeSIvv
whjWlD9bTas/3q63N4kkYm3e+bPWJS4fFDdSYpNBEnut6qc3kdK8M6DK2sfe//u2FAWxyESQePYF
BH8SJAeow2WLz5fFwJSid4gFt0Ve2E5wGsjv/1NeTT5U22I3aWHsf912COWluzY6LZhGpgYcx8EW
UVMWvLohQSBpoA886h8fn3hFdjF0s0JusoDAvWs+cPID99QLQyJS5axBCIDlkIgwwRmTWSGNjBLS
X+c1IBFtDOqP4xr+kMUwGE832T+twX8RlKm2gamx1EeQmJlMPOauYaHua7/jl6lEnGVNDTBcIM5H
5HDffH1HLwdU84zNQz7aE7PkT+w0zHHRB3uVxEkuUvzeCy2i4iqwsjJ+tFGY8U0kkwgFOWsAvhcJ
VP4txvyRJSzYK1XxvwgSbNPdGBSKMxrBkHtgFDuDyNJZWq0B1Ym3ldXpww5lmzxjqdJV9RLPpVqf
/YeWyTNyRqNSKAzxLS44G1nYv9cSTh0RD1QjijeHojx5sEo01Npw9j+jlmMDsL2PX5v0qnuBjtYf
Adck3xkj0Vq60HeaeTQ9XxlSRXpT6XTcKW7cDrnAdKuFmeHT93NYmihdas704bSN/rH/s8Jce5rV
MA6ZKuEIsWGNoOSkSRcrnR3BSxxL/+Hio+hIQVijOA7FM1tDuZHAl/wztjgojUmHVQ5dlGKlpl76
qjBvx4oC6+xtPqoIEvhZpZdPxJoVI73eXoF2xoJpnYMWwyCyEHNN/94xnZJ6pqaKoTR7s76c8xPa
zHsmkOL4ZFMxtcOKcc5ScW5ZewEa6AlDP0eZ9W3u/bnw/lS8H0zt0QOZ9pRAMXjaTM/qCpt2nddf
wUh9lmKMBYRNO31lQCClxT76hIO2+Lb8uTKUXfdL41NMe8pDWKruTzhhzzLLo2Mdr94ZM2l8xLwh
1WAamxTvUp7/zH6uPAfRPBWQptXP525bHMxhJgOuACrsojJtBwwmNrr1ww0SrAZ7/I3RzEgBu9IH
+QsbY63CVLFrnFZ6/5Oo5PIWWYJTVj14Up2sqbgwqPyLVfBXfNsCQKkxgK4MK24sR+FXLS/7XmCY
qtvXMVeBSQGdg0idlK5YDR2y41xvJSk7dc0mjtTCpV3DKUVHuwN12WC7q0vxBeugdBnKHThzTAMj
WfZ7+4y3NIWdOOAhdUhkZOCYez/OgZtcYSO5QUPvlOwlIF1VLvLuvpsi2gypA7c/P+Kftme8Tv7U
hW7nH92fLk7Tl0tFipbqhK81g7hOydoOIemGyd681Qn3hNuD/WRymvabMtJuam5+MfxJM+F+RAle
QdBaT1NXNt6Lq76+coz9JiygRedPV3QLDuuybLhUnEbk+3lk6EzC1Lz3zJhcfsgcy4oEP42QhP0g
3h3N+fQmtfmWz4lfAD+iGHnPT3vR2RIh8lynBEr9G0gkZoKozj6MoSfFcvwBdCncptdm3sBUWyao
pj/VpWc6dAgUh15/hvPTIXyPdMGV4GP1HQysVPhkuWhFcyszZH30Skw8dmeqmCmoKQhaMU0LZR07
o7oN42j3EEC8CFQEqwMWJ72Go6ZwSOoCGfe1INSM3ADkUpKHBCKHbnRJH5Q4WITbpAbmZSVHt0ZK
lWPB0JWWdMDjEgM7J255OO9LUnOc6sKll7wWLCq1DgZgk6J0/4HBtyXAGdpdo+UHij3efjKTwXtf
aMWKzjcyFLpNbVBUkWT1O7WIkZHXcbUHzMad+qcL4doWPY3O5Kp3m87PFxVf4tjJ2gscdJOXqDuf
pdCWMeTMILXkhMoV2ujAz5FuK0pK98Ld1PeyZKTA8Sv4riM0AJG2C39B7WunSASpDeM2CCLgPQns
qPPtWTNP47R9jDVOj6JfFWlDOJIlQN4+vF1cXwVEJD4Yyg4PoNeWjUr/UgY+s7P5BovRVvQHVUWz
Bug/WF40C4DHma4fx68B1GErRCcvhEEkc45UTbIbFf/s1ZbmGi5rgInAGPozdl5xmTWsSBwcn36O
iSJgWFQN7ezDJ0tAIe1YKNMwoadrhOU57al/8jioXtIUFzjAxdtq4BZrsyKDIK6L8w2uFGcF4K7E
gpXNbMIyN0zQDwZapa8VZQqASp0fOf4E+HneKKoLG/GIoa+JMq38tRCLW2yOKl8cfUXU8n8I/OjQ
iyJOZcCp3VxO4iZFZNwUgXaeoXuAAS94/ycmVmlRff8qdDPuDBU3piTEJm2TnQVzrMF+4l+LnAMw
6U2guzS2+5cgL0LRz4XKyf8u2iXOOEZpIY3UE/nrZjtoYOu86tmR0V5ctkGePqaC0/u+69PBV0Ep
OI7ZZY9Kcpq3EjKSG+SoB8XG6teZcM54zywhnWN4bV0g9x6QY6xKUFxlnOGGEBB6fy3JbQ3iubsT
e12G154ykDnkwH95IDsyeVQhQ5HhTQB8b1T+jsVkB1Q4PmSOkHbrey3ywuzwRPSKnZlPbb6EVRZ0
6rhuhSFe/yqr6N76cf+MN/Sv1Av6zna3wgo1ecIkgIzhL+5WXDfw6x/ivOSwKKIwpTLp+Ww1ck3A
/FvCGfJgTTlWEqzZsBbe0hbWlnJNI1Erf5OpTREiVkbmpl4WV4tWW639l0xc8goVIF4OHkP7kD9E
HzWph90gFd9gMYxh9LJFZC42naeID+rcGJexflMEUtWgB1V+qRohUivokTPfvHuwFJE+JuZEtlMs
IE+MoPhcONOH2QE2mIPteNTAReLN0qUCX6UxvoHff88aKKsJYG+bsjAUoggN620yjE8dyYPV1biS
KSWPauB336mW58ivHRXxwAwem+DVe0mT5EpzEOO9KzrhgWAhgJSJExDhckcPHIO6FJlbX5rYAIzj
4lsR6YwXCOm4q1qDzynKai0v16lYddKFHQEVgMJPZr6/JlrGIEYtc7AM9eANwhJJDquGYifGoVce
744NeVkI5uHVKH1MTEdMhKHtP3UJGBaszEbKydT6ZsBcw4DilBNQHHJEvbzbN+lXNEeZBIuhik5D
kY1//vP/RRj0GiVuzbhj8j36i2OW/H5tYme8/sZ76yX/1bTGf2roh1ih1tILhKZvBouTs76bSrlB
Y+JPPT+Hy4H92R4HoGOQDqY9Xexjp5RLPfWBfxsoa4bnzrhtIwPf3JcSGOv5TGgMJxbtxlenuQAO
Og3kvOfWiWy/Z9xJ8Vw0CfrRaTKWfdIQDk6yex81M6+r4+oZU3b7zvWnTR2B9xS6SirKdmOgwVKy
P/NScuvvy7uRlBkBH8X1wCFVMGGmYwZoljF5R7HgrdIWi7qynpd/rzwnzm3+OWdMNWaStYIiSRGb
RAm6i00fQrxQXZcvsWzVM66f6cgym2s0FqUShhcPQVTSas8k3KfbQ0PgqoqPB88R94yLwVL7L09m
izOpLDVvNaZ7CLufj5FkIYnngFJxbE4h3hzYNIK/7opc7XFmnImK/o7zFkPkiHcGg4OcRCq3zhdw
x0PdpjYLu60pHZJF4acZIE+r207hnOYSIwC1eg5GfJ0kuGB1FweOX9ZzamUNyzKD5+KfpghindTL
eT+bVy2WZYT8/XuXx+x02ZQGmzwa3riZADBIRYlyurV+xoSjKVbmRwJsSYQgps9Z3yp+yhjB+KIl
sE6iR1UlprfxIfxw+NW0L1cFu3MCz1munymDcbB5QGcJNAEgMeWwZx6nE1zaI8KVmXSsL5kzNolr
iFQSf1wkJ4u3ibCacYnuBvcpUNyUWWMGlUQJdn+IDIlOPqKUUqPYZEJ7qjm/e0D9RQ8M2GoB9QuE
X1tOi52Sk21Put3mwsGbWgpmBgdIHbG8BA2BTq5zOv24EnGlvAwdivQeHeRUVBM0BzzZ5WSw5k/r
QpHuFJ98+R16IXg7TDq8gYikIpPt+OJE8R9LOO9GDhBgEvoIEjYpsyVqXLLi9vU525ouMIWRer6f
sF9Ek+2LTxOx15YroVsVL5Gv/khoxHdu/X+aRPQBh/zX0ZLJ6HFs02zzhNjJIwZ2TpMxRiWzxIFs
4S6OeUSpFeC5KG/z4SrzvB9G5Jt/EnZd6dqEGOYuDvwxZ8ASnPQfkhvNWh0Hp+p7k+nvZTAMjRxJ
gkRVOk3vlRFebIi3D4sNOh+ZCl/uebii/Vomjf2rbJh9CU0ItYikYYVwfafjGc465prA2aqVds6o
vwhF64MHU4u/U5rnP8QP/ClpIR90HvgeHnDs/WL2GOkz+7EhpxuMbLt3fVui7iZbur3xMcDuTYOu
v7iaF85UPM2vmjJ9/qI91Fcbs/UvEo4Qh1y5eEAr7GDRkaaRtZY/vWWtHoRzQAdsnMGlHU9z2qAY
nihCezE/kOsT5CWfY1SiJqbO97n3oo32ToK8StrtdhFhKKwnX8zuGFhmoHRh10zVzdd0jRY4Y6d6
vH0mupX2N7UAiz+GID9p3MzWQHS6nsuWPuSODUbKLCBeEdTP/hxKjoPLbsu3Z0WDHZaZwXeH2KZI
t6li68aWNpuSMJjRMpO4JsQjivuJwr2A6ybu+ilgivydZWedKZpER0OahlHdieSRQDWmJIISRrJ2
8QO3Iw0pGvlGu9MGhCmXw/qfEyPXd78SIQj/f7uowYfekQHDSW1E1TXClzQWrUvYXfhWSEXEEKSU
IHdb2gFeSyg8WpIcusZRYaGoaxDhko3B9Iyt32rdzZOgyatcY8mrDX7s/tQtrGf/1zmNLYuDHvMe
JoJU18fEiBXQwpHsgKFYOchgcJoNvz99S3AYCyBEMU3TLUWjwMjyO2YzaK0dUmHr/f16NqaYM+QQ
hlRd/WGk3MO8xaZEbgtux7j7jfV6sB45q2rDedOujN40WFx5jtSCmORXNmm9gxjo9o2vcGJCG9XO
mraXIabXcNguRU0p+M+uc6sVpj6gQf383P2NLSpzkW9jmQCUwpd2dzT1fPrCoL1mN859VlEZxSIW
0r2bu8TDdO55ljaBvYTsdkMkbJfm/MeV4CspXsK6b9p/F+uxYzKGl9ES16htrssPYssh8BYKDS81
al7dMcPQUtJtR3RU+gmcjsorZMLkp1Fbpvblr6KycSBkEBbluqFKv47YVSDR5SABn9onuRAm6dlJ
nxUc6ZRuzPq2ek+3x3kQPE+gK5FMTsxj6vyykEF2a0IN7VYTrqfZIek/ELvVCdSADjIso8HQaa3V
hLX6Zmui4D1WazMc9DTKBZS6MIPEhrtII3jh5J7kb9QmlFkwcCKP5SZDgpKeVmbxv1YnipKR4yJn
7VteW9X2APN21NHoBluyeYLaOnfawXJy3XRE+9AaYdTxXAcVTlm8/G/KVrdLXjzblgFDi8Q6igfy
GO9lBdC93mwJ5jUoJbZ/9pE/wOPzUvBlufQMdhQEMvL+0/1cDhy5deiJ1JTLbQBac/akAyrNnTJl
gqHR79rFUIcqeqK2B8QN5dLstyEN9MddkXFUMdTjdDri6qOH2b9DZZzLBBbGpIc+Liho9E6W5h5s
Sj4nCv/SzuqwCyI+BwuPReWuVsyGMZ2qR8u4ORiFeq1SBmgh6fcpSJnl5S70OxwYWSgb4ViUd83+
X1swv5pEwOOGRVgwUgJgPtOw9eMel5kH5Xfq9AjGpvEfivYeRPtAYjhFoSUHgPop8+phMZ6FZDs7
wPIVElyzARfx98voqycCjLvJ46upKvO4MK+vGQDEFI5g8e4hxG2dy8q6TCvwwLxTA9dUhKPZdjgS
FzXy/EbNf3qgO5OTj751hGqOsmcYZoCh+KPrCsbIslhHV13txCxsg9jT4mVDNtClZ9HY5Rsuzv7z
a/ePt5CStzOtn9gFs/OywxQzxCLguZYyIKjigD34uk6i+5wGLSk2FLYNOhPnCuOHMBdeulJh0d1+
5mM3DLEpWfbm1tendqt7xQ1CGuui8Mdl5qB/yszBjLUqeWcIAll0vJFy9aEZV+RfQkFeubgq/o4q
8bn5zA6t2k1k5e2ESlmgR7g8KGRFNjpA8jq9lZHomEp1XfWUCc1rmkTOKFp2VsYxSGN47mT8pnYm
85cYKpCt++Lu7n2w/QC160J0fLlcMDDMDQF+35cbnc1+M7oms+3prDHLpNwnRYjBav3nCOfSRQDg
Cnbex/S31USDVTmf+WA/Ie/2ztRrA04SZFVXIpoA2oCo4YNEss3rwexBUz9EfXTnrqp2f700nvsy
IDr7ZopLBs3L4+Lkd1rZ+OvgoNQI1K+X1vc2rwaQK8m/kyUbosoyDRWO28J5DCGAlbQNTnf7mMGW
SUrs1yV0pZ9EKzHVIpRP29RmptJLDXEcMV5Jj+VrVwFsG8mmdwF3qMc2y2RKB4qOq1h1+mSv3G/1
Wgj3vCAmMyLpAhlhpOpq4GuE/aOyFRIEhagSqxrFsJ3/dAMN8SKS30QXockZrj4YnV+TLKoUlsxM
Vc0pqGXWx/OTIjrK30gz8od3e5jF9I7V8aY8SDiPHx6U0vqxuWYFuSPasemnR26QMP8+ia5+EVQd
gzqv1/iteIWefXfv00hUiPGDrHJtUkYt1oxMAaVDqxez9XOq7xE3g0eIn7QRz2esjAetPO+1q+T8
Q9sCSMQDVmmGd3XrSyFCLO07Fc9Wu/K3/RCc3ydAwiwS+PHg8oT9Kh8pNAvt06OWfg+spRbMpt2p
fAv2QzJrkvjgv0BTmNYHAFkWO8OXsON3UNX/TeqXEjsyFnJgKcfpddp9J/0F2ushCSaW3rNH4Tvk
UeaVPE9T7ejToIazV7Q6d6sFRBgfXfMnFGI26rr0W3CSLIQq2+vjhQ3vZOtOeDZMRMbhPqM7XPIW
KsVfwn/bMf4HokrdHPanDE5yjqYDjuHykbtXljFQrosHL7N8WgZqJUY1C/MYPn2VuFVyErOUmu8p
wczT+/uGwuwOS1WScl4/OdU1xqksQXwybB3Bhkk7Q1qcnesK0SqGlvRoEaUcDZlGdM1B9YAMsDCe
12lX7PE7AxGSl7ltXrAyo1Ww98WOwgkdpPbr4mzBgYZWmuB4dYp7SM/v48K7w30Z1Wv8jeUbfE/z
EwudTIlXCMeTQ/tv3MnwpNlI1Px86GPoEwkpu0jqiixmfVvwni6bG06FdqAiPUEHCL8S/byjruGj
VpRZyb2OkbrgSGZDamilXENXA1+khRHPJn/q4Eb42Upw7rDHEJjiWM9E+xNLcL6pgM3Y1AJUS8Cf
AftYlEbewYWP8iOabog32ElfQSOysMUxnzZ0i0JoWrWWe5InII3o5fiIf5z3/gxdV6pEqb1/wHWx
t51YpMKw/j91M1DJD5dVA+cg6Rv7ntjywl9QWWp2HywUiVUu2L2lY07zQW9Btv0rwCgiS1vEXS2p
dmg7R9e8yMIs9l8AgrRwVMjfH9Z45IaklmoX2Mw2+vauBgXJUlL+sw56vZWrS0c2JTBYdH4TCItG
JB70GreCViH0hEiixRFR6PIInZMGpZBbAweP2jU8xL/79MBru3l9tFNvmXZSP1NOPGpPSRAZXu2+
Vf3t4E1WW4i6Bz/afpCL4FRuDvZiiKQLymgW9xau7Aj7C+N/fY2s64mDDgp+VMJUlGuo6hMt5yfz
w+b52VaggUOsnfg1XIQHdA36Gh7OqtB1iW0RhPXPh/c+LxHZg6fT+Dv01UnVEfk4itA/wyPvLwCE
0mMnyEUZxS3JW2AHRB/s1wHFnuQwSrDxBvJGeIWO6GWIk9eTct/76Rt09Uiyrgj9uSOSYxDngna5
U532RLdMqGDoM8hl1UeGU1NrosayCwg3Boa6LYmvy5sbBeheS+TdFKeGBzdeG8+gpSnNrIR+we0q
h9NKB/VohKLypMLyMcUFRH0fpePaYGBHtb0BUnygpy2LHsmlcs1ZEqvmAUwVDv4aYDruXhqvHYeX
K1flt28IbYmdiscR1mepZliVtgkMKmRC2l+KOSP/wtdRIZC96Sq2UkFLCHdYE8rtTihL6gSYEFoa
nzFDgolFCOO0U1DY7xyt/GNtPyEKMexDgh4Tdxkme0S8dXzKmLYWuptnBNM+kOVvyz/lcs2hkDOy
CvqDxYS+RcFx/Cz0lA7v1s/FSBYld3RGDnwel+zN1dtCp8i4VhTEMKOgTjM73wn5k5lgJfKX/5Cb
9XLZjOx6ToiaKTb7Yf4Ff1Yv7JdeQFp3M+7n48aU1BcUi2ynD9MxIW4weRmuHpOKi/L5vaSJDtj5
C+DLqFaW+TYfiwaLDcP7vrwpskjgkxLXiZzYebN3HoDWjbucP5CCdwQzEYgaLCL2mowVCP86mA9R
O4b8fCxVSYISnwvHjI/MjqIc1pJ3lhfHK+LdJNY0TSD7Enpz5s6ASW6tJXuvps7boEqTN1JcO7zV
DCWr3t+Pe/IJVRml87cWrWh6HkOddF6/gM5iBKDIFzMCUfPTi7RKo+m6VJ6VPM3xQm2eKBJkyUGd
xJgOgokUOGvY2FDTmakPIBxMMaYL9RWSr4r5hU1IqsODB5ohtD7NkwfP2UY1BmNWyB4hNfW/rSTO
haBS7vM3mnBgpi/whL1vbq/L/sxSzTS+yLpdqngVpBI0m9HW9GfQWqrdYREtc+tE2NlO5bmpr6Bs
cloWhu30me23KpzQFRZPkY6xpZLQFohTw3Qf7ZbKlpbtIcTDhmus2G6qeQ+mnifaKL8aSSQrMDC8
a41kCvehte+OCYTsVM91YO1v3nSIZGehrbVGCbV91EYH6L6Xc34lXKAiQAV+bSOlAmLx2F2xJ6Kj
HXXRdLVeH636E+dnuhV/3Sx/aVfX+OHNvNUaluRKIGiZnlRt/nE3lc+unJbgvpQO3jLpIaXDMZag
Mz7fPTFthdJiFK0l7SpCyOpHm/3ze5hRq3rNWviCFQ4ypQ4hvlO+lxhe2E4HrgrcwMwpHp8Q+tRy
LPKEwy+GikAIi3RUqB3BwljRLU1uaTAyEjP+FM3u6Tyub5tmWrxqFP5dwSo1FOw3GbqHMz3sQRKM
TE8OX/HkmIvYm7njMkYpnckUutUasssVlPPkFFr9ZCuVsIy46K0rLENSZ7wNfKoxfDjdbn3lrvMp
x8csAnUm5sXltTTEnqUpJsU3Vp7msNYXdKZZy4AcOvoGiq5THNYCoW0kcGIj3cCpTjK3i+WolqHa
JA+wGO8CxEQgGajfGw+FVo6kxOr+WwWq4T1eiStuJq6lzmofrxqojCTIY/Vvgbvx94NU6kRRmMhe
4kbu8CnlSW0KMjv+4SPWiAUhKtZpAh2pGBmP4ucHSW8IyI3cXtEms5hAo5KEaB9Etz3Xyl3sxyuH
BUo6kXIUMmRZsxiCiDH9qwPzpBUF6B+Bs+vxCQYZoiMhQZ2N72kc6vvmxAt9xyjT6CJLPN4+KOKT
DcJtz2o/wYxc6Ta4qBLGdnVr8+liVrHDQu8edrM9yO8oXWTmkIUWWRHUHqBJ3T60qQJPnC7L18Mi
mig576ZJWbIcXcvBP4xX/ZiV9fxEUiltNuLvOIWT9TfWD2d8rdXNuh6oG4XDQrE3I6sbNvgMi17B
gZ/9aIhZdM1FqpQYmL8OBoxHoC3pUKO/dq80yPwLnDUo85H+TDucsNXG74iZz9ggae1FRau/fT9i
HpS9eRBw4rYvAoQr137y31xjKoRo/b6gNhBvQaOx8J98CfKM91SYk5cpoMxFrgtJc+UZGhAQ5m3h
addEr0SDhOAQqelqa5dCrxXZDzVMr0exbjc1O57znBKrhnho9Gdl4q4XhfLwx8OlJ+CYG+30Hwr3
Pe0eVWe6ikbIj6xMiUWmWtrm8A7u1r3SWoOxSERsL13fKkaVwZKk/kTbCahSvozl574jGeLr8EdA
E/CW5XM7BMg7k97Ss3+efqzNnFFvTub6x9na7EqZe0vIpLYSWfZyBqIl/kcEajfDZpOL3qlR/bWa
QBRaPJiumzNFfG0NRMkXdauK0MqN82ICL+RR/JDEyYCkNvjgwlh6ubDjKMDW3vRNpUUI0t5QRIii
ZOYFu6D/mhnwQfY1IiPhsAo9POoREEIc8OqGzVz2NuNPHwVPLvbt+iGTEG9NOzlrxbLaDSroEdG+
KEh9XULXKHsd+gKmOtYSddtmwP3wL/lB6kqd+tggB1ACNS/4kKhhWrEKohdT0t0MW6OaLl1eLkWT
HxY3l2rs5pO6DCh4BAiTbOsjAaem4vvfBaJiUcd3GRYTJrzSByRoG2Igfrb82UakTVHORFU8Lazk
DtOvLALF34nvDnwurU7WKUzSpAq9jbF+KBTcKV5ZYrF0plyfOyQ7vJqWAFXxW6mZNvD53eJ6yC0i
xgzFUuq7wFCFclNDG9zsaAQznO5qX4RQLDA2pPe41+cxO055cGmutAoLmlIfCiWrEeTqRllvK70N
lG1YtuHR7q0JCTd/1GKlxhxdlzP/b4ymBoacOCLPR14DXkR6npdBuCDcG65sxSEMH9D0r7O4k2RE
3KLnLSD7jSftqKSjaOjyhsEPrOicWPznWK44TJAGENNFu8SJ8D2WC+cHZ3o1f0FGiMdyXlbkzAFu
HtG64v9UzjBSduqXvAcNoazLenwfMN7Upk5ZhQqZ7T1azafATglogFj/mY3xLJPBysknBB1MSP97
uf9Tarx3EjMRIgX+oKsHtOAUSzZ+GT4QXN6h8ZX0t7j1Vw+snDN/vAu13xuHY5S+VWpRSv3OxXQC
/QP7CIKTUKifDFzqvZZ5EP+j0Fs7vGQctEj53XITyuumHWXYkJhhB/+bbHUSn+ll5g5B/uKTXZSo
xmyeuie33q5OoIu5Y3VpLew4i/neuLczrfy4lOjC8p+XevXEDEKCa0JQc4lBqEwm6xJ5cQXLKyu0
5de0KeIiaBnj/HAnR2pvUNpXaseHXVm88CyzTChR16vqlyxeo2f9lZv82UdExoRTwpYbe0lWdTl8
sjQNLGi/U0xq1IXynBj8gyn4ANYO+WfBzoBMEXZpvlf0X5U09MXBIUtuA5DoUVnkdmhMf6YNnyjf
CkEGvFplVALMyvuktIkaQBRkdUteQqNWLi+iR/1v/RuxBDXax8MoXqahky0g5+nMaNwLOng6ySMP
2w3p3RiIk8oIt8BX/Ea2WUoVwSuZCZnSXhrz6D5d+pp+D5+P2LmMsPK5SRiVTtzNIaZEo7DMPZWO
vNIFQhxk0TJTT5WbMYl8jCIroFs2ETEZNl8fRGwm2vjyI/jIH8Fj0D+sB5WpVOXn41uqP+xdIpe6
EeiJudBi7IZeVmVch9CIt4VnqyN7Yvv1dIo83Mq8JokrnSSeQzE1/iZI5QbHElUKFuXucTmBF7Zn
KzyXiPp5SSqwhontn7dQfvya/SwyZCKQzpWDqcZYd+F4l8hSQ6nGKmOMBcPQ3P5Kjtq6L6Ftg8VQ
WmyAhfUoYrGfjSm2eEdyU1RcT52X2ylG0y788v0nrGxTaGagG563GVSeww2bezDJShDXUk2zGV6U
YSAk10C2KAZxemT3yK4bfo6/6aeYVIrxGzDVuCQE1MomnznehDpbaOFVViZ1Na2VAMPi5s1Ykl04
8GTgIm9Fou4B/SfVBBOJfXLCO9nfosQWwc6w8ORshqm1++GxVSFFXJL0OMRDMwtpXnHfOgxAPF2I
1oeCcQ7fw6k33+h9GpPRT6eZGjGU4kPmHWh1etNzKWT5UGfXqkR/zok9eq3Tzc+r2Zdfr3A0Y6Nl
OHl+iZFRMF6veguKKUqDFV8aSi7TRYdonEaEVJSE8zJWVK9xR1ATNLdXuBybDqvI2xNY1mt+t4ca
dxKR6nD80aUSCHhs29pdtGGyhI9V5AGB8nHDP08xLJ5VDj/l1AAiHiFmL5SGoIJ/BhmQoDQaZin8
EI1BrB23Qd5uPzxSqdxAzZd3mJvQzcD0T2e4aCLGq/RTCEupN8ijasfXWsrGDilUFKHWC3/Z9WEz
WH4jDqXr5L8IvM9yCwRXExuwv7KUcchwsLO3CRrWvUtd2JyTKDsrnYToaM1bRjDaGTvtYFnb8z06
MxsbGeRHV49f9WH6YIl/EMtoBWREHQa7glgDTp6oQUt7TDW+zaeTRSIOrQTmSE3hY8YxmTvkd61q
LIPXBFTXG6QjNGU1c+PkbCh4mgqQu6fdVnlsJDuaRxKHrRgLa08/StLo72KGBpU5lFlCQAup3mPT
OT1fWO3s/khJ4SCUfNzQcmzABLFrkGh6mRtzNmCELLAv/W3J01RJJya8pY2h4+vKArrbCZ9BYxN1
xKaelh4hWHUs5DkS7pfFsw/sOZ4qNAnbRIeFeXRY1GAB+hopuuaNwsTN3+4Qik6ykUEBxVvRnekX
sPGDPGMmFb1ySGy0/ILi74nTQfEe8MOUGu3e3lEOMAvovIaR4e9ttEL6b4tE2Z4faYib81mqZ8Oo
4gUgGtPI75ZeNpw4LFcvzfa43CnZ/aWIBUULpjANKLpEf/u/fDIJloFE+mxFBm+tft3WIN/OiXst
vGEbAxVKcEEkOpkAsYWZSpcUYDXOqKgGIf9iTLs5eXyF6IK+2hBNcfyMzVgvYvlm4CxpQ1KgSxJ9
4IwMHcmJQO9g/IUNsh0pSBiC9iG+IwYFa2H++xKWE72Z6ByiLgx4wPy0V2Z84yMxZqiOtuMLb3bT
Mwd6EW5G22nZAcGT9frpP26Vh0DiRl9JIHyqyray/mWl2lyYD4oqR6gKBD99BbbntWce7LL2J3qW
tpWNhc4Qkq7MblPh634QTpxf74aCKXpbR2MQoprBk1qKlu88YE5ZltkUXbUhypawgVfzOThwWMyk
DAjk1g0yLcDXzjWdwZJKep4wpvfAzI+0ELDcpbp9Re+pB8467kfeIyuYHp37Bsjw1qiajhbAJ835
NJ5DUWhepW5jCgGohrnght4gerd4zzVZgSxpVrHcfBSUUKJuTBVG8uDEqhvFSjTwtwtwuJ2vMwCI
c7yEqf/ysuyWcM66pzuf2Mt8FXqFOnYMxTbDZzX7eisRcb+GkFU+XkwInB7gyYXm1a7zldFeDBBp
R/NayrLR4i4gECZcl9rz/Ls8oM49E3R9+d2jpIYqsLfYtpaWgKMYkjksNEUEtEQ2HobvvzdamFIz
JSj8cPo8+tUKyYgfHUWk3CYwKoSBz1lPIWAwGQANKSGppp+T56x7AO4jOcSjoodmxZL9448yb4G+
TSjTpDHCY6PvDHRF2YkxIYLOGibmTfI45UFpF+r5vhX4tDxSCGDBj2w2AmLvqKVBfdEwLGfDBWKz
QYWL00ZNFNv1e7iaTwYj6JSU7JlZDxEYZ0L+jfHrf3knD0LvXXZ+zuXhloTg9uSCXF8SJBh3b2lo
gaAcf662XSmKawDyV5ikqXXuwNpaYX1jzaZKhprWv/NPk9vq+7klvBPGSW+XNmuc7n5oXc0xg9N8
77foO/t0pwCY/2KgNKcGEOh5hkTJwk3k6vsAvpho54UQPF0lQZakxAeLtCq2NHGz6RxELFgxwNkb
vEI8ZWz7/rymjuLS6uq3VGkZI3uVi5tHhRliWSmbfG+sNycgPESKTV8Pn96jGl5nJZizRk91tQ1M
PybNZvx31M3Aemws5EmUEjMisqY2WTlVKIdVK7XNccfgk9Y5tmyfdB0qdgqFVD1oGw7TSg3WWAGx
Noe15CAjW+Bm90dfVlZ8U/0v35zLkhREip2gw0lFoeYX5PIaYTla4zufTQO81XkBFSrJPwPpxHPp
uZgFGMND6GZxSjc6zetx1pHlprSZdFyIUbE0+txRTTtdy0yzUfUdumlbedDioSE5JRNPTmGTqug9
4XoLaDJF7VCUrIbQvwFGGNqvboE0AIOgczOKVr1GkdIHxfZu/P4NWFVNSqW0RImjqIO/r6IE2quk
5bl9s0au2GYgOxjb9fGzFrAh0bo26Qg1I7oGE/RAp9ThVwa34VdtqX/57ZCz86KG3zstPyeuL5Vg
/01p607mbbb0eU7oG1VtlC9bjzfJOCQBsBQEo3eOzOCcT60rFDOMHAHpc3E7e1cNwg3D9ky94Lhn
SY4kUxYL/SJOFyyMaXhUlA0BNtoJPzrkzy82lyUbuL4sTTbLsYYetniONK/vG/eCghGzqHtDYrfQ
jLsRIVAygawD1FIjf9CA741KOQvQtQUy8JTMGRVgO+gGVqoIs2sr4Sn7qZgoAklT4UaefHRSZVXP
kpchE6CVeZ/lpao0BamFdTGRCK6sae7DVy7KKNcSknBV5UXI4LdQcPbzOvGRm6+Uh8XgYx4RpHkB
GY1+OAMe9lx61Zmwb7K8prdspir+/q4vYvoUFfcQqAOzxs/qZD3TtTf19TjimrDz7i9eBzglVqMv
qMZEY7CJfSscdS3ZHIgxx3bbK+XeC7t1EhlOuNTD3QGHUO5nx+wYxwXhLQNH+Pj+poB98UXWBzk+
EB1JU1lbVXZQKxUp9dVnFdDMAz4zoTognJkDtks7q6+O42NCQle87zI91b39hlMU0fbekrKiPHUo
b3sa4jyWwAlqsFFXlNS/iJfWySi+mFl9wg+l3gTm/fKmimCuCE3a8A6+HNHsQs3FKWlzD3UNcEFr
cXeOVLeL76rlsj3APzyTffVgYmXrAVRY0PzsQInez/dU/jTmmRMnnl1TtctlZlZQpawpUp95jam/
58EPY2rZYRQ1XWkznLtVmp3TlKDWq1X0oxD8pXhnGkXUzlsti/jieP16N4AlLlp4BuLDbTTYQ/gS
5/QUJZ49MiEodjRiuB0wk6LyTtbhmXSEZBTf2x6icSknpuoD/9LBx2O3v/y1OOBgi97OSzOJeoTS
YbWcFAKIUI5CesBdVgEUHongBywJFAE3EOD99xhGTd68c5on6qpLjC/m6rVx6GXoIixrT70UO1+M
/pKu7auIxZixUo9nxd9P0OXf/3aEbvxZBFN4DBmFZxw5IvgOLHk1KopJVTmcaGTTs3ttnuynnliE
Q8wF+hmGWwrTJxfjLrC2fEit6anMMgHuSgK4I0FE15ZVvjAIVOjgeiCuFyQfUraosmmliYx1K4OX
U3cV42RCtHVhh4OIfNVbqMSMeYtcALHtLtd21HrKQI/YWMhZP9MreF1KbFkiMwgGBZ+7LiTqUvBK
snz0FAGXxe+NPZrh696o9m1FTt/ZkqWQGwcb9zFBA4XBYuNY/UtnvIligDzJSR6SHNABA0xj75gX
IvEsSOvvZR2E1kxNbdqtL5hUP15OiUT6kfYvSCb0LVnEwpdKm+Xk20enJHVUtNdv0N5MgQichKBT
LPKNhCqrCO3nk6ubckk/eNP9E9wZrvnAh/kT1Uesskp4L3RY/Jgsi4o9YF5cymXMz7RLL622BTJ3
oWuNkM5QRUqq9V7GlYQLscjPZv/YJwQAvE7U10En3s3rtawwJe0BsZ8+fL6ADZM5DT4Yse1EH2ZA
fwJC6THxMUJzLzD11CwaqdgVcuMnLq5Z+UJ8I2lbJasCCAiCLbHVmeOHFVUfaeu8/xSX5/tM4xCD
HP1ePyFF2VKDjMWvD7Z+yuKC1pGrtWmP9LJjlqz10CTbTOqnx3n+i5JdpegXmNM1mh7MtcFEtl+E
9mY+3qGGwRhPTwosDV+zWH4dHmFtZ5KdM1IebMGfYPGLoFazjpxzm6hwT2FBi8T06tWbKqi06hJn
k2WeIHKixZT1LmkuP6UBgWgAn1KrbWmyRItH/KSkA3uo5F7+R2ghI/C18RbAcdCzWed1utEGihU5
HG8DZzejnvuqL2hrBWFV7OB1TXRfW+2IefCu70w2GTATqY/SPE1RrXYhrOLo1Vt7If7wXGBrVvRc
i9+tM0IfzYcZL2vJp0CXjfMTptCTEWEKCSU2p7sbffOxa/6cZ86zjFbsf+rH4b59PAXoxS7b9RHD
QdJ6/ca07LohicqM2zVyqBsjNvqKzUDZOL3ArxNztCbUBc4HOtioE3vXe02wVZ1pkfhftmkmAKKI
EHa/guHWXFoNKysq4e2REp9g+M5zim1ZuX+ynLs+t9OM7zJRxptBnLGPyEkRFHCfj2bS2PmSVDVc
8xaevpRbDa1DBTt9Y+wlvcJGv2kRrmGKikBvlI7SWgibX1FSxasZzVoqZYW+4sK5Bt4tjTCpH/SJ
OwuL54QRpK12PDkBHgubG6EiSY6Oq1bSer9PUF1S1qbmA0lc3vk4AVb6gq9Kay+wCJauFtbuAuDM
6X74fquZYRqGIy5SZbbJXWvW1yfojTdtizkw7Iyw4iyTFR53n6uV9GM4kcANJkf2PwDoF2MycUpu
RN5W8znZH9LxPl0vuUf19sooVKEYMgoLo/kDqv3IniV+RkkdA3y92m+6PXb7WxR2/VwqRwfAOdfT
2D1ITdQqjv6Iu/KotPCXHV3Zgr+XnlSiTdtY+S1RXUb4YmlijgLp0HGqUoYZv1ykKSt3gjXvWgVw
oviFDXqb3/EKgqh/AVI5HaXIAjskxQzx4m6oRcO6v0DV9SsD7nHr/XTp58RU/g0D4//8vOb+6Wxf
bQGAmABW/Jv5IJVYb9m2t9ThcYRKRhegDo+BS5vpR5Q0bTHwMswMAiVNr2yZ+Lq3ffPnwP/lBRDC
H0J6W03P6dmVKqq7nLzRDkG0gyl8LvKN1b7mjN8sqb6g/rwgDefDyKT/TdBF7tfB2Wc5ZOyZd6yD
hlhZ2ovcQ+Pwjrl/Y7H5Re7yiKv4IlM8ry+CuJ4p5YlE1tcIbct10bmw+g4DGqJQrL15zE/aQCG3
m3rTVo0YnwJz2d/JZWBEJfxJiihnQCp8O+fvTcEVmR1X2GqI611Q1Kdsh+CPVNs2xvx+2l/9CAlT
oafbHjY4FMQQUtmy/2u8Y+vbPmsih4/aJy/zw05+E+1x7vmXmXDcNZF1N/RL+NVzjm3C+ED8A0id
Qnzi2RS5no1AIDY2uZjLT53k3PApPwQ+Ki+f5OZDgqTtnPS55VW9GVErYtWf6pvofMz/XgFD/ywz
4oTCayr/t0cNh4fafTvktqoW4AWNGCy8yJrWb1z3bZ+GuIL8pCabGzr6D0n0x58weGVxH2/N3xtP
MaF/t7rnfC8B8gHahNFsR8l2fRX6Z5I8U/2u2wEZW4mwT3qr0zpYJnIOGBN1nB4jch2GQ5jZI1P8
ZxskPsaTAjXJBmnJa0b/xZtV6SUc2kKNNykdK+siZrNxiqm7Mjy9P5aGRSFl52glsb8y+sitDK0z
FvrlYvAeEf0MnmXqzAN3skdlcgsdE6MnAZ0WJ0dS7WTTDvJp1NoNf3QpBs76FJRiz4VDsbwI8Ekw
8t2yo3nz29M6cbAfUaoPr34lV+YMBd3jpjv8vaCR6bKvjhTCdvHXv+tD/8/YNeCoNgBtsfmcv5bE
lCCuGKXcWW60eXARkllh/BfwnsRg9O1QglqgUlt7c2Q9r83ZwBMMMcBxwiHqH5HdQ/+1U0+2I24r
3QSmxM2JNjYH4kqU/ypz18AHSnhNCSR5juU3COyIU3wQTTzJpWml3LfoVgAiYRDUI2+jSK7rPvOM
qTR7g4a5Dzq1r5Onz+fy/xfk76B9+3YYlMwOkwsyBseQdI9SfdpS64Ch7nuLadWxDYd5/6KYEBKj
8yb0a25h680DcjW86od4T7vm3uW9CUl4sDlybC/mXnWv8u3BXFoynyGDURcNd8TpxpMgbcc4xcfI
wlrNvFRkTuIKbqv5xBkv9DQoWC3/ffEFSPzPSX/3VH+EmfEcOKwdWaPj/D8pPHp7qELtvQBBHvg1
Qli14Hs1WlwEYi1YJRM/SY7VeRYGrIjHqMr5LIZvntDr8cRG5FDo4Tz+5q/BmNps/ngofl15k3Sd
e4dHU1BX48nANP8ZSs3I1JHt6AcfWITGLcaKhW7UQmAOEMMv5BTEzAZ1/S6c6vFa5vZMmQ6oqB/f
ftwWX3jnOVzaGBk69HzBlxrls+H8ploDrs/a9Jqvc+5BmBipXjA1ibAkyD4OuCGVq6E+yqsmQvBc
3wgqtSeSZJ84SgJjggPQDbA95MNVFmByK45VWbiHiMQ1L/e6Mrj18s+mmWXyOMvNXsTMQeGNUhuh
CF0jWqkuAP+MKTwFPwg4Z7ZbAp9ybkrjgB13qwO7KuvMQaY6qYCsiEGpouc3ZAWxsnS6CbFVqs/i
8U7ChXShajbSTTKyyMTeenRk/0fR34Bo53BzQF9++QxnprTMuY3vrRftI+kLAUkL6n9ZxfiQ9Jtu
00CqOJVvwQ0beXPeHY6Rfd1edb1qYkVrkg4rdBxPuObTwDN3P9oeJ99Qenu1wcxU8etGBat9GpBB
6CX5wa5UugKEVBzr/fWkpE1Mi1AstOxzT+dYlEL1VICMSNFQ8aNerv5bflTd77eeyk6+9ZY9nE3m
H7/eeifzdgvW4GQWBtoeMCgl/6iDFwNRjLniM0Ty6VdZMUYOIxsrQYUTLeerxhcuX4Uzg0DLUegJ
f3zfox64/xOdmctpIAR1rWcoFsMmyRPQ8cfpjrlnfFldxRDAQOSKM34Z5Ywtc/AT/WG8WmLb0JcK
rZAaYwGRij0xTRF5k5eceDxWhFptK7FDUXYGm8oNB2jFdSz17IO6vvYA3ekl8tF5sK84D8srweYZ
F4PoaIe1RHFKBT6bXuoOGvecqHPpCGUhZmsLXjpiR5IjDFMfuB+7XxuHpFUUFoOeWO8MPLvH3soe
M08GSQjLjs9vE5PmDfZgM6vIPYfph86t88kY9DD3WfBPE7JN1pxS5/9nQrRtWKe23EFGrcvcWrWN
xFoyuknGnlYsDzTRrlLuYIjFHmQui8Qd7NPOcVhRWwV6L61I9mVROmKL++ylG8SXTjub7VTV+dKE
DzdW0Tsv+VQaTgvN9ntQ1dj/Er1qyl/q3H+Egq9oCYNT4QO62JOIsdGwri3VfYkKkhTgQJ1euIat
YkwdRVEo3K/9eCjDAZfLSVxPXylAXfpo6y5LgGlIOr7+qLoSNQNokjd5OLYvdFwU9NYtJWocQoyF
/bB+dCUafBB5doohHDIFepmJjbBBiXYmQNWhgEgnoXZDSu/HZ2bKAC8OzR5tXO5yoCBgco2hEPLy
1L5f33bE1jz1Hj8P/3pGwHS5jXjXCqmSEQ3/hWAlwNOSKH7HUffz/K/re9qEmi5YnpfLZEWm9GXt
xfMDtgdEHcGSMJRVY3ZRq2OPEaOCPVYU7khXsH4+dEMDteQQmLKcmEgBHgiCj3tRT3T/fNib038j
Tebv5rpUwRj/VB+X3QuNNlJhIHIGcPvjIFgGM5dHvCqIivZzzk/ebYLFAeM/y67jvtaRBoKkEbdm
ksRSDaSGFImSV0xEzzTIoi4IVONomFt5qM4M6fI98O111HDdfQe+AdO+iQKk9eby2LGaAv9k2HRJ
DWYZSKKiKaBBQf+eagqB6nLkZCWI0InQACYVI1XWV2FfSPsgm1v+7l+priDobSoEAIR8r4qHyytG
SRgq3pCz99hBDKw8Hd/F30sB99Y+S1e/mE3ln8IM6RBPsazi/A8FQzv0udS0gxCip3/+rT9IaKxw
p7uDk1HBDMWjSF6zVGOsPN7j76kxKgUfrxCMJ/4sinXr+gtz0x+0ayXU8DuriLuQTzHjvhrPuR6B
Zoo/IJ7/qWY8y06fdRi/CaOGSL1CLh1eeYa98fnwSUuyJYheSVxCPEybMcIy+4xOFSAMbF+impkM
TGp3gRu94vY6z7KhBuxmr5EK3YvTfn/id9G+v1HZ1bAznTbsD9Ov2Gs0hBjPEXoO4H85O4KUllLd
/kmjueWoE9YsanY6OI4dcgbtadRNm5ZVs0wlRlGEUD0tuLJVPQOk6kDyn6Ec97Tcmr23WydPxEYE
xhwrkEcBuyYvnfXvTAXlDILvX5iBhlmkx7Sg00ENhGbLrcQRoYajQpH0Av9D7FQdq3nHfeBOtYCk
py1HwF4uYQiI8tgSgFAnC+k98/03d0KQKFs3u0LAyDlnX5KmZYvNQTLq9Q77ysS1/iNp0hBiFGoU
Abmw2d3YaYqueB8wRvL5VzvIf9U9bkPSV12/9fVSdCPByz2Co/lr2pr5SquHNZ82DMFCgt5epLxw
j47YcGPuX9LxmoEw8EfxnO/oNNBQFPsSqkrtvh/maElb7D4N9NrOx50TNpi/GuV6taPrKXpRV4eX
JbOs1UEQ9gm+mc5jszWHaQFNBvzL71s+8Th8OfLHggP/LFyWVs5A42T3q7sOtAdaZfwnKyiLAC3x
5DDiclji9PCw3ekfDVCI27UJXym2VTDbB4t09ynIoxK6LwUDg79/8fz4RbWJ0gQ7zmncs/onhXip
F8cbCAK6jKr2R8X0rg683TrJch1ydo5Aq9LdlZw3RraV7oXBCUhueSuw/3E2xKqduLBOrrq8pjGy
N/7HhEnhzWwAPLCjuHhPYb2xKKUtfg0I7fSSzqthoKG9IQFW7OtMeRHzwr9Secmg6xwM3N+coRaK
U0r43Ull2o/jHzGHTjK4/ftHNqnK4JMaZFV3LNVcdln1ghWnEKIavV8WUL8xRk0rMfEYkCJwkwQn
Te1KES3ucJNmtdlNPRYNGDktjBsJuP7+QMH1vWhd89/iMYeZnfl8g0cPUm7bgr4QsAuNC1rKcmTK
xnXehXOURTMqetrFKf56K3VXUT92siU+mfW8jVjKYU3CIRBdbnZJ2J/SffA4mO6eG3HrUQt1Lf+y
PQf/GW8SCJL/QWyItF9uI82bB9voAlI9MhEX5BAjjY7M//7lD7OOlgWFF2mA7I8V6jGxOe/vQApw
2ZqQ7BsdKmT5NhG6TkQZZp2ZNJ5N8XcHzGPvj2aWRA53kCq4BhwWga6tGRvdgso2PIyTspyHKzuV
SeYf86ddAazwtJkQkIUvCW0XpXV1qBD6j02XoKP9Uty4n1aO/5l6YERf+DRax86Mg3u+8CskJJgF
9gCloxzBbypgGZGZdxmH+kQb8sBFvvwTp5E8ADQ4kGP/kRxRG9dQS2GUEIdTh5H2v4gN4ahXRDtb
z4nVcc575zDlDaCcebViNEGlXLytzg98fIAlcadscJ8f2biesV0jZtjSgtelS5SKGjsPpNBHxQLp
+M/Cacmx6+CS04RNYb3YgqDN+gp2gWfdB9HuhGKE7/lSaaqIS2wv9pNby+JfbB00k5ox0OVo6UUg
LNpl1rnb9MS5FMY1WDCN+ahSuXQcdMmdomO88a2NV4hqFuO5wuPAbEUG6wLsBF/yGJmZa5ROpBB1
JGbTjg7ZIdFMckCKkpwy82vmjDIpWUqIuiOprqUo7OrexeGSnAoG/ZDcEnljdVMttXLumN6WzSjI
pFPFTgEv7gvpLv40BoF+yoLWs0aAeXtsBCNOxesucCT7ODK7waab+y2bvXkW/xSJk+uTN7XFX6qA
JoGe3CITY46YwgKIKMeTV23WmAFQsMnavMtVFxx/V8yx7k61WvEFAbxiQE1Pp+51mbSpQQE1lEYv
TWkC6sQ17jLTvS1FxJjU9NmhLApoKUEX/1IaNYo0ddldWZQyyKd0xL4H3sbKCwOH5caRmAMZGZ21
3tCWzkLmx/NGJvTagwiMRgCkf5H3HE4ie6Guw366uKCO5r0xd+V1jbigW+GowImWGB+h3HaPq3qm
NX98VuoZqgP+OVFs1fkG5EPmjCcf3/nbmQN6z0p1PSNTEGRN8MsD6X6rX7w8R98FtEcCz8u6eYM+
oagAH8NErVra9OZSFFwoqMnla8ANwB+6yM2oEUrDj5rl4Gz6oNM+hB9tlAZ1iYG6+dp4TEGy7Oak
TBAtHTg7CHLzLXYhhvYqmdTeYUHLKY9y7KuC709AyNso3X/0oSwrRw+Tr63MzlpMh84LrB14WgL5
4PDbkN9uFNZTm+5Jab0OEnE+9mn8gWtEqxsTdxiygk0alF8DDjWzg1ZHYwiA08XLizNwXkzJHn9o
Ty9lJ6Pe/nehVNMF5l/jERuG4UuVJB2Z5G84Eog4TkPCFxestHSlDtU3gW0U1+NlRQXeTht1GLFW
F6v8PMFowHZpOXGfsSX6QQhxRG3UhJIlVSyBGKe2A9ukPtatrJbj+yu35tnDW1P3OS7qGediS7za
RB07b4TQ+fGRHpAPLSqelHlFUPJmRIYhcQpgjOdLFKc2PayBoKtGYqy3dn1fSRVGNdxvgQEJzqxP
neNI69nm1saw64Z7+SgxRh9iW04sbbcMkFgYHOLTvT8ZU/ZerhuqaRG7Vr9hEKtroCEBYspfvh9e
zUU695vCovZQWZIPHCF6jyeCZv4Q2bH1LaLH2onJUenTfnC587jOPDNozjpyHQQJVedNZkNz8kYX
7E/peABcLVgAsAdCBkwIQmV2ujv2qxtxANhpKHztrviVLZVux8iB1TeTviutgC4yWXXcRFSC2ALI
xr0R5qpCtLL8mDjazGjWL4cGVSCnbKka8+LgbPAcAEIPnK84RljwinPaBKyoA9vRbWVGrCXrXOgN
fSD00M/Md7dsXIiYlGaXW5iznuDTGRADQUqGpCtaiyoZDXO3Ljk9Wc3LGuY5DxtnPE/qPyqDTlAc
pDWQI5Yy6/MwD3DPGfiMK/8z6L9b06rQhYIfuEfeGAtEmP0/y3DH197KniKlmagP6ZOslgi7PC81
Wiz/lCN/XGQq9ILw/zfWBKgm45gQYZ0uwST7hT/9aUzs6LiiAhas8ujIo+/h6NntIbAcvxxqsT6O
KX/X/mfmnG3wjkVg7vR5u6ol9Z6wezmSJoKEe+L6VPiLryUzYFl99gD/dZwSvYOYKMEaf51Vhyfn
taKcMmsSA42RzNwAaUxhUkZrp6wy8Lwqdz/A06d0+e62MKIjATIb8ITJyzueeAprOgi6eVVOqG6D
Gr/DD4iStJhmfbYTldPCAf7O0AQ8FC+Ms5coR+bYKWUItxxGlsu0giEGGqf8K8CMoHK28XLwpMTK
yvjZUZr5xX4e9s+W9b7kwqy/O0oA6wK+qE2DIlUhgQqLzu2+fCgN7KWyW10l/1TrYeNaVj74T5sm
JChxvPsfS4rPt6sFOCQqN368JBFfLY37umciKsnyaM7A7pEiiuXcbiFxPL9cQcTEZb/vDO4Gfs4k
d3kySWPWyu4mXSx3EEzev+hVgPKqe6nKPBM7pSkhWUNEN7SrGMnx/oh+tXJ7Awh9Oshgy+KvUcPW
nZASSM9FlTNt1Cj5W5IAYCis8Dl7Lx+mTLk0HLiKEHyVeo3/RIz78HC+VqQfMGHBqPQjTBhGoIFU
PzwRj7jJaLisIOa6t6cOG0hpMJXh1P+4YShPlgsTrONVwM72muvUSB/B+W/TWp+6XcO00jTSAdPy
rk7LIFmTb24TwkGrZ3zaOf3QmMxZvYg/fDCiVG4k+OrG6WiUDG7+IDVVKrt7J4vMk6C7TeJsC5ho
q7i90Ukn1Ae1LsZToPYVtM1OwlmxrvgeFeAnwwTOJs6GYQ5WKQeJ0bklFT+nSt/ZWMPQRkL+i5M/
y+BtVDF5QPFshirn0o1nMw9DU6NDKBfb5vuqHEI/DqnJFyPny3XdRUK7JwtzPHGCvnbKA0A5zUol
0ZGttxVww4xuBOhTENZH2pp+qwU9C6mHEHvgnl6X3SWg0zw0rIcRrVpjXTU2vOCKEhTDU4QJr9O9
ht+tFHuGLeQrYWPp2eBl21xEhU+os4Yx1mzLnQjwS2h64WIvMA2IMSt4ZS5OgHsxeVxtKs1i3Nvh
N60QujAd+k3v+88JMO50O3E1w3Na+C4mLJBn/03OXqOwI3sGhIdWpMHQieY2bn83wycv1fp945/2
hfDkN1jVsdu6zo8Cac0W//BWLHb3ItJd5B1GMO3cZy7UKQd+sh22ljRc8V/2A93jdksj1/tmD76s
RMn1AMFFXmvcz7QV7At0COo1HrfZ74IlT3+RoNzKpfxRvW3O168jjA27g4RLZcWD2uRYcXKKL5tb
/2/XIkHdHKk8sUciiSi2+3oF5jldutQFWvyNxN73dI4RZVX7S86rghaAw2fUbb3w3+xTM0jF6Qzu
apVpNqDA2fZCwWTWeCzhC0hsbhUfGX3bqTP/m2OAVqSHZDoM3drnB2+X5Ttaf156d61FyGE9FCI1
upftne/NJCEoF8hFAIWAaBSq6p/dYK6qt3dtQgugJFbVgkWYTDLRckLxzS8jwbgKnJGoPeXZs3f0
0R0juhWnGqFoCm7JxuDXzuxjMCEn+la8N3nL7MKMkJ7BDYFZbnMPZF0lukumyMB1Kq/1YB5mltJL
3uTWLFiWQWISa+Ka6iy3DrOx0ZoW9aRzWP7Nrk5a3XfdbEELBqrpG3s72EV1yrzlNDEOpwkNbzPQ
Ap0JEcAFBAI/Ow+6ARcvESg9tUaQiN3zMw7pMJ2N2pInEYPfP5BPAXV8QmR5NxzKqPYXIeimuHYe
fhsojjWqT6RJVqDisVG41H73EHGSzBPm2Dz3ZiWoQAuhzZcgotRvCDPFN683rKFt7Oax1otjIV7F
tHGpiKgWLC51uUZuzUny0Yr8NX3KCZ8DXulK+Lwmpxi6ildEhSzW8RNwiC570RwxGW9SyyiIYgH+
o08+EE4M5Oqc9HCR3wkj86ARgKdV35BWAm8H5gD7VJu+2BKpdu06VQcaQDdKzMDs0EcXm8CEZMjP
T2V4dzd3reoJwKFQASnmlCsh19qCk/EeoqrB9e/UNtRqdA2Rjc1NwAMrQKlqyXYCqTA7iAQvNg9j
z+KTDclXpkOr91k0ysE/N3t6zvSNA6EvZrlrBMy/8gN7l4GBkwmEm4BKjoKyr/T7UhGIiIvY/VEr
7q2y04u8XDqXpEqj+c7uto7372dpIKwERBgDWN+Cb8RTbXezY3SnV4UbuWWowQ7g8RvihpMg2pNf
PTZacDJqhfA6OTJVZPSKZ93EbmoRarYXbCd282kbeGnU2LT8cjmQK/uR9enQur1ZWpIN0goyiIJq
dEQfNPqAINHCLMr0++iptNAb0OYoWt4clhB1TMB7jdS8v9YBZ5Lz+RKCcumHsFnVCM5DO34jMkWz
r/+cWrNc3YEURAMMOkP79Ea+ya1iMUWiVx1NXXJrLE5hWFgJFPvrFhJ7r5IeVy4D8iRa0NKPfvhO
js9qejBzOJjPbb3UtigLTikHEB+ZPCAG3rzsfeoSiNyz97f4moeP620ys8Ybgj0RcGLqcwWdJuhY
5Kzkn+s927yOQpYu+hSD/K2zNWvmadT8KRAV7FUpipqReGl+ooRYsbtpV1VvNMFKkh+d09C6KBof
BCiTacOI+cc/WE42EOcGxywcpNzQaCeje/FeqjzjSM5LpVzQY+CQNc11I9du4YQG7P8OgWWKfKfZ
zwpL8Veu56pCxdRoqtH1MjSs1lQ3tXj6zSFvUu/t6o8J7ezakGVmbOlWRzUX407t329q+PPIdmr5
UGFhgIhDUX3gBB305XaiYycDr9snPB8HDq241Mzu4A2nAkv5fHaPDcS3QsmOrNEbsdbtZTjXANDw
mpbATb3yQyJdzKoX9Z2h1w1qa0mk1AYrJrAUzifYRo+T1ALV7walVZC1G73EB7DgqHSVMpQzZukK
SHG/OXNBqrD+yOuNsqj+bMEN5kuYYiXHSIwKLw3KUldIylUHxIo4nkxVCtXbrpuGrmzgB0Oe+RAr
SYkDkD5CzlC+4TxYrOVr21gAfAHj4+MYkb89X94OJLLiPIjYC9mcZvFiYBxjnzpS3jW1nVYdKSeX
RwWYwRSXgjjfka4+6/2zvcId7ORBse1APEQAN9QGT/fNOlXGCMjcBHR7d049kOq/0MiDXe6zAYJv
SytyNt2WxEpcxqIdHHEldy32jGTssG8hJ/aA6UN1+OgXY9GEdp6b4PqyN+YRlWO+NL5weaUK3cZY
0H5CxZ2+iAS2W9iYDelrhLeItFVVtro7LYQ7TwhfvP6Wb85iRKXSfvY3oFUVi/XZw9NqWLBEZ4SP
4vj/44iLb+qoOlO+md4YUAjdfLyQ7hxjvjifvcaMLuNSikeXjbEnnvBxw3W7ywSok+lPBVLeuYi+
44f+rFdp4mehS9qYw2FnNyMfHI6t9f3ADvTbcVw4G71fU4MCXmBUxNs4lQDMqj/sRJH6A8a5xJCR
nhKQKW0QI2XAtm7wFAb1zRSw+fsD2cM+We+zAXFMePP02eAjgEBZCuSyED9Ak+x4vysfLB1KD/AB
9l8LXGwcCelHf4djeJida2KVds7O/GPl03QwEO/H9y3A5hHR/QZ9gTPYMLgFFYw33JEDrCe1dR7N
46FqVc+GWh/hghhnnlyDEsz7ThcHwL2CM8M4pVqR5HQ0ZnfIK6GOKW6cxEZH4a6E8QuOMyZf9U84
d2HT4vDWsj2pJn4rQN/kVtnxmExoJDm158TI9yzPEBMramX4FlE6yL8RTleHpaIWz3Knki5+SvKg
aEKVXXQcPARAjaacMLxpekxeVroMXhvVH+Toh/HcWA07Qo7WFbzXzbDQ2MOSrB+8Hq83O9w0VO2l
qkPivL7Jf/vpKic0EV09rNOHtYqYzU6c+OvWX9f6gR724WiVDjBkaVCZIOLBeG3x5l9NV9Aqha+8
Zky8jlYTuMRYbXKdNVECFUcKA7LAgWML760wQbKpNCT4BJeJl92N4XDwy6eWwyWpLA98SKNdlIBD
EGOBlyESq9kzK5x/Syqwj4duLfFYmXSraoPaa4euHAQ0Ela2S1LzInn0LlJPZwXcLIkyKrRCkmVW
NCQ9UT7r2PIBdatu1oWchDoy/U9PNOnB6dxJmiWa+gY2UNcQbKXokBo3uKmIwI4PunPu0MQrpwjZ
Ni6/QPGAkbTV6a7NsmUz2rqoliXF1z1M/RWY8ju9Z6xKCKQBXNngtzLQf5jGKVNLglfMruhnemR0
KHD7Er1Ug+ksZzFLmvGTpXxzRsq3T+6+/buTQh01G8OwiTtQv/J+aboJjPJETwnWESlUzfjYMklI
skGOa46G5p/u/Rc9UMqDVU2GXM+ShmZa4pmJr9lH6zKxiFkxmUXAZImhywi/ZKkdvLuKw3HUQQbo
j/x0e3KVujyu+s8vqPIAWV9Ls/Ptg9OA466s7mAeROiKYUCgkA8Q4udiSj4GjAw9lLH4tB69Lg9i
xcVmjT5fFA3v5f7Uai+qgeFyiVe2rvzYvcUvIMqbe+diNw5avGWtmCZ+r8z7Fn9xnN9jZX6p5F3b
nasDZMqveRGgml94odC+LsudYnmnjegiPb+XhCGSK35wxvTITMTfGDvmzg+X11iBIv3C2ACADAAY
GLNp2rZ+/AZsfzmDop1pZRoEm5N8a0szX4uNcGSDinhUwl6IyqTwKsrVVGAKZ61joa6hBD0XRzMT
h/xdTKL59CWvHBDlO8S5Xv2muscH94pZrTdCou40+LBe0dDtK17kAyZZGS+xY3nuu9H4Nbb9Y1fv
u4kVni2Vdhh471FuVSLGoDDjMRN8D9ea/v9wH3A0ek0yrwNGVUL9LmwV1fztKX4zBvU13BbTT3de
hYAjj85d0E/d90mP1OM4rK7Gtm1UTenw9pafkTvvuiw/M/9fINUgfnzWK0MWD+qmp1bwC0Aibc56
xIAjtuH1WnAbdvb9S7AaZPhHxDPl9R1MgaptDD+cJFkGRF5OVfqz2osE+u9x1jy14cNZ0rcf5oLQ
7CaNJBpEnbz/9ujwyNyYZK4mZZWere0XDSVroDLOcPYZp2GkpYdFjiyBn6vk3XvmzmTkvtbtmhhX
IFr7WIPs/v0sBXWFs/mCo+iaEwjl9wB6eQqF5k7XwT7O10daoxVM6OPBDnDoR7qHPY4BTWJhmpeh
RtI9g13bIYHxMonAVyiFjEdr4opFks3mLJcF92XN5aaPaXE4SXWqen7DlTvczhdrLbTVSbTMIyKw
hD8ZfbbIQ14ounigUu6nypV2Hvzv5sxchDkHPVY8zCZwI0eCcSwnqqmYx4PJ/wmYCYqHQJtgQUGo
SmRgHd205T8TVC8N+Vp8IvY9xSn0mC8YvwregTbbSKmAenDFWQWU7p6qWsuZu295bNOAEX/vcP+v
pZVgaUwOS5Fev9nbesp9mr70FUUaBwDQIuOp61tSksOalFLg9kgruHnzHrT6x6shrS7EUzDq9RIS
BFxK6LON8yBwv2W2rS6L8niq9Gjs7Rn8Hr5nasUNjAEOGvE6G0sWHrCgVEdiq0PdK7s09DF7R/z5
FkJuFOV+Q2MTuUPVYTtthMMp7QoMCPI5otfSUDDuqlEsRgottwmks2WSg5XsUKMkS36/MkUSzVDh
kRmsgWv5wh/6wvCZohNofqr1kHwItDjfmVqXKcKg/EXHh2f6NDvAvHC4/daP6y1a1w4HnRAYYsd8
YB6vRmhqdbwwvWKwRjasAU9vPPB3ICk7rxZeDNsnGQekXsC7N3cpy0qXvUQUHC4kC2geoYPqeTWi
2UqjnEj715jk+YT7fdoDS5cHlXWi9ls3Y8mqP66Rr2ewOAubuq/PkQp4MxVPjcd7r9aCEAUgbiE0
SgHkj22D4wocN3amBhhh7OU5BRb4FhGmCuFo9CpdOksKIdKE+Uu2lOI+kEddvxK8EskD2wDO6AN4
poYd0uOZzg0UTeWtcGsZHPqoNTQfwfkKzAdtmn8Vv9UURsnGRKNzF6c5qisy19ngwYPrdlIElBkR
mQqVi3SBCCE+237c5HOUFAJmXJcGLzK5fU7BECHVuZK+ZHuMFUdlJNbnFpR9hY6jwUI5vsA61/3/
is6AwZ2o1oQ3j51RKijYxeungWAATnl3uQd57GiQRRu4NFfknFCUaek4R/73VjyTEJ9jjFXGJy1L
+QlePCfiQl5oFbQg33CleWrcHhiTryQ+TnFZzS7piAEBf1xxQyMb0xQ7aN1ibSl3Eqn5L0gSxrfs
Z77tb8MJn1dfhiysVVqR5t6H1+KcrC6opYT/GIKeDqs4MQa5FHjANhswYuwe6NYTuXdiSxFy9UDT
cqO+2FBuPI6bS7uVe5c0AkwY7u+7Io95/JUpPGNMs+YsupQjDFqjQ8wNKsJkdxfBoBuYCUsFEZlp
yKDz1JsodGN+zWI/ACPzdAZaLfRkji+qhPEVVnZG9fclHudvJrh2dprN/cCdw9SD5aNpBRp/Xd/D
2KGGL6dQw7JNLbWC1M3xtDd8omGYKQA///FqB5VB/xDJ8SWQjFQiU2lz3MNQdLlOf2bdXB49HKyA
jAwUFTsqZQzJOAwtSOJ9XGEgu01VpwKZ2pX5gz4uOlpFwg1JtPV6/I3NIuXIytXJMgxX4Q0QZsVS
CxoOvFlDvWMgrMd6QSEcec3PknJMMIEYQ4/o9P/qczEVqXjJtkrYblpA0GGeyLMBETS8mGhOGvFw
YuHK3ZFvXJ9snjMrI4uEpRP5v++fUAuz0yFvskVTW0PYzXA0w5wSfO12dJ1rLu5LGZKyxPRihU6C
60t1PChEktKfp0WEoVuMZZBSSFES+t6lwdrEwcfWoZ5JFRj1nl0Nk69DpiIRnS80vLZuu8JCeBZ0
JixanVrl4tSk7/uQeuTKoJKUv4CcbdtC7lh1PlIMPSBubSopGyl4QKjabXbgVxKnUPqk0a6YS7wq
V9cw94WbRPk3+L+ozkq1vZmp6ZRaRHR3dhdZCCKIL2/f2XoicOobkm+LvprQEwet7U0hujDHtfZE
MWtzLRXmsORnxdePv+Hq9+DfJ5U0sl1Ay+lxbbPq490WthoVyONMbaQkpxMCsDj7740BjXmnRN2n
7hg3aB0OaoaTux6ziV3wKWCnvpf1U2x7FV8mxeCzH4NC+wKhhy34o+0GDQqX3EEpIIOrmCKaDHXn
5T18I0Zp5socrlGXVP0MHSxUoVBy54VE96q4UKyouskzQHJk6K4RM09GcoYTl6W0Vif13/mUw6lW
Cq0awbNFHSZI3d2nF00ekBSoxK2RSkdRL4OdZGdFzEz6SrVrBbeUX2cjc599cSS8kmYD6m/omX1h
5Ol83PU1e98XbzpIPymnSe4q3OLgmrkJQLlniHsiDqIT47pOUa2WDpPtZHVPNwzqjgHv7pzfXAfZ
n0Nj0/5PZmuhhAMuWwV4Uc1Ji4ceh9QuxT41nCSSHmOIayYOH/u1J0UGXTv5Hz3G6672ZzdoUXfr
JkhdpvS7PJkrkm8wtY9idXhwTE71swrblcPoKwnxCgmFQ2o3PsVdpwYeg2IluESzpyJUDtUBdjRF
PpCRzvBL7MvFzPk9mW5rZKx3/IiZNlRVQgBVhF/yKvrcTEUDKxtmlE4z5xOSl/PoCDWhy6lPGRvP
MUkbfp9IkI5Uxl3NopAosVUhWac6roIizk5iulfaj5LdWdUUaXyJu+/t/pb90KNaXDBP2LXNX0ZS
w/DlFPPZLMHfwGwmR2bfDoWNwgfddwg4D+V4IVHHaNW9ATcV/QWqXHLX2UggjIgnQ80ge1/TNOcT
fiW9B3Z6su0N+tKnQlv6E8xSgoAx8fpTUsJBX6tRYHo3txrE9h3WAK4FAbYc1N+mdQ8SLcDEs5+N
Z0eWaloHUWzJ2QhJKNsRX2Aw92B7c7UGMaB8knED5mCt+zY+w/mW+iTbTW304CEPa7fk9/dFyWfW
RiKHlrV3r/mgJmSZBIaJ9CDFL7+XHSvzH91VXcB28Vu+9FEsWYYLOlUyZ6ySqQyMXgwK7RVVXpZG
lP/0lmya9R1T1OR96TzvMfIFzbnPpy70sbAkpP89gJ7csvPm+BtqjyFehJ8iqqxZvVdGjPbD6CNX
c9iE9jjadNOHCB1/o5fAm3aj11AasVbnKQEmXq58MBDK7C8uhpyYEh7g77C5mxUXHKIRn9z83kHO
lGDTcn3QNFDqwnSzFn49/XYBd9eLatwY+rH56Ca0ZjmzPUPSK8+qZ7PwI5wHwDUKJ3DREmjMVIZy
XajRtPcwbA7yQFV9AZ26o+nMWXo0uNH7AQyapuwCYZNAYcANPxeDpq8ENgKlFGgGu8/uxw+Z75Nf
zn7JzVigEhRTO5XOEH6bts+0jJU4sYab1U0Q4u53krM6dd14HPFwmCkEEYO71OH56EoND4tO9VSz
qBSPrJto4TSuBdMubNHjX3qlTy32Z3V4wsifhJ81kvdxZBdV+a2k609dStTYPU8tPyFfXrNPQMzf
z0MW9ZHqgDZFmYtCy69qDO0v/wYWO4MfKU9SWI2GPzM341vn0SqU5UUbuDl9v0Kxsed4bCXK9xZG
MbB/VSksdklv2cHH/8ROKPqgH/uhNp0XOZ4N4QmWfUAU+Tf/E/e7H4is1RsIz/8t59DhmyXbIWeL
EIXcSA/rRenLEsePGmvImJAKPlHi+Y0uI8Rv3/Hif/niPlN3zcKXCJhOY+JkYyc+QADuXpRQ3oHk
/usVYSqGRIvJ7q26W36kzTJY0Q1lAF3vY2sigOsWIkGLSNEdsqCfCoLP293RU+w6ytPZ9kO/9jCH
BLvTyC4Qc3CyyO5/waKY4z6Du9ZTPSaDGwe+4zaNWOMb1PNJtcbTTdQpLfwesIXMHrPT7kt+jPWx
aTj2nlyfz5saBHARNRBWJHC++FmUkVknfXVq/cjj60LxG4WfbRh68cwVvTNWb92JMfgvE7gfJFlV
1K8s4QaJCBc/dtRW+s758UGAVaMTFLxyfIVzI85u8OO6dpr/oPLAwccGkhD0eAQPQj/yffifL/gp
i6u4AA84PuPzV/y2MfT4Ziyhsbfx4UmI8sQkuDA22BVe6s4MSDwlKG9rwPJr3+1wOxZoiM+9B1MY
a/BSyUwDFmzskEEV86ousNVahME9JqCahf4FMLv30GvdzWjcT5aW2HuyJfQHNC9iKQgVmDqYQIJe
wSKcUtjV+bBF1yZcjBm+nVAt3K4ZHIhNTOHzoGYgTob5fKwq6xRX352mSJx/GZ6KkuXke81yzT+q
aHkt8PWcdq6L4F8kOsZwVrvCJU2x85HRMR9/8vdLIExztzJfjphLCZNjHCQqGwstiNpy4kfdST5Q
vbsp6NpIJjOVQQv7NlBKjJADpGkVaRGTpuln89MqoSf0+u9Z7QlD2U4ulYSlP6wtFmwz2X2hO/P8
O+9vJSqmyPQKOkiG+FdjEJ5icwO9sV8RqMp+ApiJfmLotWucv5jxa3sT9OXDqDmu6+iv4sqosZ99
J/bKLdWOPv+NclWDqIB8v1bU0MWAjS+AvGF7CI68e9rpUQb2sKMTM/Uh3JmwB/V0oyq9BoSV4ADv
VjnlKjezzbeaJuIM5FqgjokSYaArzPgBkn6+mkoGViDgiAZvIICw3JCKmEM8iyaS+19MQPuhsIK/
Ls3rsKKO1QtkzbVXjKKHsr+SR2eWsxxVUxXwdRtDlEgw6gVXV/GnTxS6WpmPVd1rFZYA4joETxrW
djog/38McjaXy4xquS/SU24jJRL4bpECDRhlmubLQfBRARtcd0cuchkNm9IuBQ5opQQrl5VtMhA0
RlZ+4VGYWI6uuWLeyPMhnm15SNVDOhDgWMyBmyErbozab9wxgUwwptwZJd1sumRhPX401ejgnd0K
QsjVhVXEm/AMnqDAiNRnr/Llg8J5VGurATnhUScYaQ0oYmZD+v+igYBAG80xO5oUcMy8rZNyRO0R
RLW7t+keNrYKf2+m1VVG8DcbVBNViGsxXjhuEBEZqbB57hbGPWRkyQxsD1sS9ri2XvIXMJRCgRKK
CXjtugLa0QckthYpb+GefZlm6gYnwZLL8LzmGH1o1WczFQ1XLJSr9lPudEKQ3qUeVjEXTl9gXD7r
5NSqTVC8aYmeC6i7sETv+/Dpvl+6k6AyG9Ga41Xkq5XGT/sXlU3gE1ssZ+xOu7dsmc4xeBjyjVo2
H3V/T35b7Xtm5/Nx5xmnT7I7OV7OsWbDByqok1uQyaE3dBaFE2Ku44xwLFy/AacH8S6cVMFMuHod
y4g0yyyg559aJ/BXMPonhMxouyTqWZKEAJEHymveMcnjNO2Zec3WUkuaQuOOeJp/Vr4V45DMEtg6
0y2jNayYooRAr4IuGNqfWV/F8DHnKZrFCVDO/tHpEto/njsMD5UoFrWwN+8icoZPwT9fiWtD5OpM
ILD7dOTfgwUPca0uANszvBbanOt1uIlJ2b8dvJC/62C1ia9se1iH7S7vTfEhcnTq3CViZbReQFMf
EckqfrD4bzRuJyryQNn29WGcubc9zDGZvQuBTfbW0YlGKqs5bgQwO7rS9Y3hJlKlbXpSdgFzD9AG
owPAHxapwXUVdYoVfySOBp4RyirdQ/NqC2jsdSKRyFRhXjrkA4a5bjHA71bY4plTAWbKboUt+bvC
CKbhLVh8PvjvRC2/0gIcFFRbnLObBs1olp+MtXcw6VAO/Cybj5MfrYsOmy0GCygMu36jA6//2hyG
Pg4VVRX81O/UFtKZSz0euiwxCUoW8Fa3HZ/lAfSvPFpWfkgkfNj/cnbdOwOoNIC9wYnnnJQ+fbLu
snzGp41In2qfEeHs5seeONDWBKEgOSvo9MPebTh1sxt4vbin+qtQFPI4zwfLGP94K24Kwh+p9uBP
itkSrqbNlmOQQJSLF4cwNFEgrEaetJUsYh2Qt6cmGaF7HSR5f6sN1OZ0SuT5518XAWW391JQfe8I
gnLF4N+mR43XGpFHTDswiwUi4yEGE7Lnmr+5AAlsv1q3LtPJcN9iVbV9S4SG3YEFzS1vpTCH75i1
a37AW6SifMMq+4Y0Z8aRS8YmGRoSjH/RWzuwnFb4wc4rvRY+FDFZq8xc/EKPs624yWVTs/qgQ8pd
ErrjJxU0+y/fRjFCkHG1a73FQCGwGQXz49VN9Faz3BMrzdHOIJJkfXmhq4lWWUvOym5ogWNPuHTJ
rFschhzm2o/OqS/LbwclklAPdhGtfyxpsevXOgxJqxrEOniS3WVSqFMt/p2bc9SS1AiO+bQmXQVy
2XxuvYU76+6zqeG7RACmK1h4dkkLQpCRC6VcbWhEmZ4dk+UrLzF5ZHxyLT58Vq4StUqiJcz9LHSx
OOAlLtCGEKcvJXdKnP3EiUri9N84v3neBu67FQiY2fBvjXtKD5S/ZgudaxFRpjGPIfsQnU+LWJ5V
5r6HSiwg51a3goN5AorEtcvwTVEaO0X8/XmF/f1oRRZDZpYFjRJ8cAFiiVNiDPjW8gSZ2+ZPyZF1
qq224pdPSU6ajqe7biE1l9kqxAy2JJLkUIYNfMkPSmrnx+uylVRsC0MbLNN7lUcHmO59SB8YmfU6
p8YR9Am5/nTaqqpb121CtU6fUvnp05VOhCEzCXDv2WItLByaMDHg/E89oRs7nCzLq9L4laDvgkTr
BAAxoFDL1flwXzWFD6iDuYIZvGVKcozQH6j5Q8jSu9Axh5sFoQx5MM8vrUVVSO/pyUj77zPe67eG
JAXLEaagCTq1/BtB/w3ECXBrtcoVn75QTSo2XIe6fvlawULC3EA6d8PkDvdrA/T1COZrMvHrvoUP
vsWMLzvyLCMi4G8Liq9eAd+tXrqaNOg/TgJiWwPG9UCmmv/Ii+746Omh5dvx/FFIHH2tRBd67iDH
ssXCeRV0G76CH4kB+RlNaAgdEUWZFV5+m6ByNyideqbwH9bqINErxIw9kAlRwJE7ykY1nPurafiV
7WHE0W6Me0TcLeWTgXwu5Ie+zgfYSuMsf4OB3sv/zyoHMqAkOOdDKtgez4aepWaKHgropDIwJQdy
JGPegQ9RiMsgci1BKnGpjvHRVOdRn5U5EAP4BaidPR0F/F56+cjnxfDVlotqPoJtiuHzjnVH2Hxl
S2ikwVZP+4/z+zq2cSNTtuhwfCs7BIE0iMMUa8B7FCfOdB2/dLiNYLHd8TLeEm7qNDRRGitTmqAi
gsUDNtvpl+TBBcpsmloDG3TkzKlkNR73C1u2z/N57FG8KC9gVtfM+pbiRvrt75dmQ9OMFAUFVWJv
LF7osb4izPWHHzlJGqoDfdbXkhvWMjQuP1Iu8FfpSR3S4EnIb9YHZq55W/JCpThT60fyFCFqjP4J
IJ8kM0BxZLkuiGiJt/X0ZyssupF/pV+Dhcj/h4+keHt9bdGq/S9MFSKImwOTISIGioTRi0yGcAzx
lcL4dWhpctfhzgSU+5sY4X3L92MbqUgEbKZoRiA9THZw19D88TXCC3AwNdD7RYWac1PadoS3buOg
+ME9KI1Kcwl87DpUugYXOoEmWPmMPZQ2NkzTnZaIwhiA2ZNP6qRVuO4tnJOk2pdbtZqijQ0FMzw4
g5t78iTaBcJK61Em+AqHqltcy5H9QAt6C3usPtUcAr2sLOnr0oc5KA5/D6MocEBJeggddT9H5rT4
NZmUGok8/2xT48cQTjNcLgv12O28mPB58JTptmLPsrNuIT0/gHp7plQ5/KHlWA4iJQS8aWL9gTJz
dwHnTJccjbebgGDrNwMn8LjY9m1dJ/JcD6vtI3el1+ie0xLWhj6Starotg2+91oWpHch0irtOLOP
ZsKzBd+wI4pQwPGRYZdB1pPMCaLwfvfVi5hWY4Qwb7IylffAXbslHCSW3PF9kmZQAVuhSRsHmUsO
4lOY/Dax+hSpE4VNhbJrTpindRfPlmALgMJjfDz7Oc59wWL7qgL8a1XXS6Af7B8r5ue0eJtBBN1a
8G5FVB+yhQ+PyKNSwd85z+4rNCMnXSBj3QZFW/N3h2oh3QunIpN+3HI8K94Hwg+izqDFAByWGH6k
YP74m8Y1ApMsTeUUzYBduWAetrHKsidzTQ4nURBbsn6p0f6WYjhX5abI1QCEF2m4yo4P0CPGNpsc
C7yCQUxi7S5K3gvBY64Db4dIi4DOEL7x9ky9tD9RA/EJzVuATarRB/gO6lSpTqXCY7LeJJM80q+x
ev/NCr7D1IkrGZ7dPWKMQ6VFJ9LX7LQCHvn06uymwGX4p5xYGZpHNu+sFZQzNcrFjROEnTqmBDTv
gQdgMNHh2UPbU4+asNbg9zC1d7zQQHETxUOksDR+WDMVkj4vis/DNzZJXDEm+0/0VufAOLDe1m5w
5/peDPnebqKKkE57Mxu6oLzO6GR7SpWFqYSLrysZMgbPLMCgx4owNzubsEFYX7OdHQ8jOhjfSQ84
AP1OeicgkZdrEqTefmfAWnV0ITeQrWIClLDuVZAYP9idf45Lnzll3xdP0qklPXS8Kpa1rBn+qlbH
6edKHgPN56Sv2V3g4daiYnYZ4++CcWorrDHUPuDk4TPvDuU5Q2Ej9kVvhnmWT/YynAscyxO3Hus/
oAekUJMGXyBISfWEekrqrYe3qmL2GpOMWH8YEBmQJo9WiaJ0+oaZoPgqq3AhEBoMi2GEdJqVlwA5
ixfQeboZtXNUbdvNgcnjpkS9ojgwihZZDjCCqdCIqu8EtNwzgLM41cTt/by+Tjh/GDniLdVKeIUs
ChzSmJyb4Ats5fHXgedXA3BWTvKQt2reOyS9ySXJi4Z5Ob82c23075f1F+2xMIRluXUcQW2IdF+q
9lumGXpl+QDPgTgrd2XRTUo9nlJt1D+1tObB3oU6MjBXoc8yHtctkKn87C2+3GMjXJWBUviyB2gQ
ugniKa0kJwf45tjWNiX6V38ORvPK8fX377Z6TO5guOAN3hdbUHQmZlfR/20SEpz4UcT5T9XnHHvC
2fa1UWxQ7XJlrLf3HGVwbBqm7wLW4OIQnQfKcyj7/9SQiIL/uQB7ZuUX0SFtH25jyQ3Ht4LGBuWT
1u3UdsnQ/Kt7ka03BBFaBYZZLD3x2NSHUNKMYA0MP8UabJwD0nx4qFNzQOaFH0hXTkgnOfdNPdf9
NhSNKx3X6A3wOCs/82Z4uUhTq8GhtFuudbwmkAICOljoQeIQ1iBvcdgf4K1PO0uBS5Y/xadyoQ5e
lBcOCMnXaUFdba+2fzqmybn49cHgN6QDEfgX3ABjomVTaKg8KPdb+qxjIPo6/auByasrAuU1Myyr
G72tUyekUM+0+gv6/4EfcZ8qXas7BUONt3c72nYiEBU2j8UMGNlEVYK/DYA6kmcmWxnPhLGABAN8
0VetWlE+BQ9AAIprevrnh3YdeP4wio8cgfoyaB3/HL7E4Cliu2qtm3NA7X+Rh10pRUekOYFKmtX0
Y25icha/GsR/W16rEi9rfcmyc27mbA+AZCTtEsMKxgmyfE3pG5Fv5Ma5f+cLlFJbckSGyHWtLgmv
2SZ7QEsAhg3XrBsKOMNUfUuJU2tXOb5fL7t5g++ezGqsNcsd7V7ISWKWegs66z6Bypkzvfbyam8o
3CJRRUhiorEcQVvxAsOBaVBSHzJsT074LGu7LH+uvfbU48seMVC5TAiZV0YlqKAb8Qig8BTaqLwL
iQ1JNGXm7hmIKFg+Br9VRim57N3zYDFrRVTB2jct1IybuxHlYsk95fsBxNs5dkGrIloexSINleUe
vzA71k1J4GXwvjPH9ZyBvmQUJ4BD/hmmnhjd58WFmlMjghLZpyJchw+5PwszPWqBHh03yhPXSL1g
oYRaFFEUeuB9IZARm3HyANOkghQq+HgZUvEMkOA2UF/lJgC7rnrCTN9j37g19aczn2UlsZYt/vWB
EcDqyMY/5fa3pugakg/IuguMW5DONqbKXFeM6/0BI9YCjndSByf9N1HeHaTlzqcLwGa8dUCs/QKo
SEM0MXMdf/a9Zse2gqME4TtEwavS/K/QhdgnLBa3VglQTFYn9HLjJERKgKE+xnH5rGa5uQQv2mmL
9I67A2TrXmePsfVSwUin9k/z47XQIao03zx0gPzoVRHRDoKb0Xk6MYJa1BDCTBdN18j0JIORiDVg
qruzRFOzCpur7aFGs0CkxW0KpguazUeW8AQeHvMkmKPtHB763UzWEnA3VQPt6QULEHCIMT5vdN7a
M0/AFfJyIEZyAak9QL7qwsRYmqjMvQi4peO54Ts/xX6E6i1v3BHP1lK4HXtPKiMXoS6Sfg8+bv4z
WncB6QvKSXmmdrtOoRYkaQ2qJP8ZobafsGFpNYg97cVAFSJIgyPqpGR2k4zvAJ4IH1tPTKYDJ6TD
iYIIJQW8XTISh3bpfWRBBMunHtuylso9m7+oWRtHrJNJXTYWQ+aAaqH2CMC93azKRjN0eLrII0XD
maxJ0SmG8ohhyFznUOi/797SC2pAzZajy0M7UBrsQVtfwNDHQFjdRuKpIqmalO5DKV+J5FuB+xnG
gGkI9CdWOUCe4+hqew+HzCUv1DKOr/yZQRhky+efDj1E5UoPGeH0Zl9wTyGemyUyKImHD24KF2JW
n5UoBd3uAzm+lfO1wZOEhzF/GdBhyduPioRKGkjrBeFybcoWkzbaFxdhTgVwFd94IHXMoAgS0dCh
5zrxrMwBo3A8X7i6XdBrKHtZEeHBJlAQl5P7rvhXyKiy2lU2va40qZEG3L7i1/oa1EnaVi2+Pzd3
coqEa6EWZpjM/JXSGlYd+Bh3eTn4Es2+VQGQbX3bFFw8pOha+RQNcfG6FzZ1qi4s64jUPf7bkm02
w1PKR0GmBnIZ9H0nkcQTJGs6NMVHwhwQDl4Ui7dVtYQRVYB3jZDqM1lp/4Dn83XCKP9rcwkAZaFV
uDfy/bUG/HiuUm/z07m/DnJyh3Q2K9/QrTnd2llZXblqudC8T5ZMZDDUZ/8hwBUzjq0W+8RUVy7G
7EDV5BfnNZri6uQN1JPn8vg3JWkx9tjjTHtpqE0IN9NpPyXO5FFTWl7+wc/o/EoPjjepdFUh0kJe
tAcQI0pNDmcvgjGPi+UVkleUTf7l0zPRN78PVtjbe7oYEAX8ZX+KcXp453M8pMY/xETXZz7MuE4A
LhXBpHPiGQ1vTDyV/E3KKpKG/3PexYgaL8akxgB51RYTsWG6QIDgVt64D+ikRHKndwc+U4NE1Tbe
LUrs2ag30xFkByzQD6+CO/DOspei5Y9p0HgWJ/YagnYevUNmqzmwx+LZtBBhF91GPds+Jxcl85Q5
qRxdVtHbayqallTWvFsPK/+YUqCgBProuOQOKY0TeGxSz5feJvpx8BbGl4O4MCXwyDpW7M/YG2Sx
BJPfG9IeaiZKvFAOua0M9fPAipJEPXMOPsC5Bce09rxDFvo3lnQJ1u1Wcw9btXcPv/PNUaLXbpsB
q8esj+y+B7KoQ25G7rXeJW+2EnmDa2LaRj+0vP5c6GnEM0NfDWyPKAsALHGDVQimuRtnCQKr1Gpm
Y3NXWWnWkqgJuoVLUmP8EAlpj/BXDtC1xU/Hg++0DA4RnzR2zBzVEUn/TXpJ4zrF9Cg+XosF0JkH
MktqWpSXGIbbgi0+wn6Ieag9URAyggsayIVY6Mrw+tyzBYLnTa0euc9L/TPl3PXSxDH+Vp/Yz1fs
gHvg5B+aO04CKMKsvLdP8uxGP9Aq3EITSMjoIyIcbNkPEYAedaO2BmBeEwBc+ELDBr/8czA8v2pz
xkW+vYXlpvZotwG8ZN4XmG1RuPAo66Ze1jHpAMxSWC6ikYUKuskHqr3azsj5Y+EhvfO8e3U/j3zz
X5EKegTiR6m5x9lFqdMyk/L7qOfFcYUzO07EZvR1rPImySKHQMKdIX/JfthBGw7uBgrpgr0rk+Gk
aTT8wiTgGzNSu3h1jXZyF9Siq4aoaBNMZOrK7I3ugH79q3tS2O+qAjp3D0ApKBGU5Z8vkeUYgwBH
0tHry8GDul6XVmRFv+Ihcr2fTU6rTN0qvoiwK6xIaSRNoHRwFZtPHahnv2+rdFF0SuTWzyUbLUhX
2CSvBvVFu6l9oPs+hRkX6bVY1Q6ZSEP5qNr3XeGuMhqfrXw+b6GSq5wq12cPqaDQVT9C6lwdT9AC
pOmNPYku5IFU2pnqqiWFDAqllhWWbp/kLqGS/PD1KLBOsRC8ghVyzl5KAoNOSSGOls55AV52uCOg
VMiMspG+MfJvZ/1zBFdXuNY9HgMkC2IhE5fVtIN//5Osbp8XzgYPVzQ827IEPEvC27tH1hfDQnI1
1VxzwWuzQRm+kefXPnPR/0WT+JwTy20JDCa3p3Orund+geLuGMDPj6akvFLI6nrxG5cnHEN8k5z5
6UIu0NvfM9ODEfuYjrcODWYNziqsadr5AJcZR4cXXU+MG1huiZtfBnCjHLei+Rbs0Yh6ZeeTKwGZ
747bwQDOfYD0otRgradngxrNTjOJzQZrxParTHzqKhmPRtnUC329kqSCgbn6X7SVnR66jWTudr9B
HJ/7WONfk6Sd3VB2Ixb8cRbNY3JLTk65TDvG1o8BM2uabguxioXroZB8sWVJMCrFA7bs4yMlhSR/
9CRA6ST0wiwQOR8/X9Laq1RPIWg9qm18+bcBY5i0u2qSnMXeGTArZOrGpkICizIOVIq6pJpeZqZA
y0fdGBhZGujOIA5iPbt3BwkBaw/SaIpvFOgXyVmEd72vXZRhn1mLY1HN/1CclyOW8HbauxMf4Uev
N7nnFrQRXvPyBUaoC1B30o8NNgwes5tv9rQV6gzlCQJYKL4WdP6UPhCrM92jUqjj7DHlypB/YuKt
HIEzXuw0WiaN13Ny+XZh+6O7IqSsC+0/szWhmBELGqqzozqYEcA04yxQZuNl2UdfK6LXughS83rV
vPZcUcPMkR0JRgWTy61nTglbhZCyj34Shgsv4Y/aRXwPnpBvRL2357nWOkA1VKD+bpxiQgkdSOEU
v4d4MMvmfSv/TgHs/5330wVBAF8Mtf8mBYn5vVcYAOtThvU/t1SVdHUKWgsPIfsJjPs0iMe24zgl
QarQYCv5AMEW+RJ90pHSjWR4462o1YnMJj6TJX3U4S47rHs2PIUnz9+opnfodmFOT/UoSHd9QGqh
itP3tZ/lkr4YpD4ejdCHK5P65IRDsPuVmFntWKaEVx1Yoqeb7XJG6AzrFZ7euXdIXVRkDn4v97bS
cAdrN4pFDv7xzpEBzntFJ4WFtY75MEL0kNTrSDOc5rkhAMqNieg+2cKnZo6XdOpHNcGpzvza+QbS
QHSPcmMeTWhw+zyizmUo4Twx6xf5HF7z34cXppjq6N1PhsncGIA/phz3BgIN7nDukMNaZheUbeiA
A9uIyDnPtspWMev/Kap4mkiZMdBI+9dRRm7rbqm3W4x8r2XBlQPViI8NNOBhk00+fgeH3doNxw3q
YLizy9UyXBv2IY5Qt+RfuLj8HBkC/ibjUG7CsKoj47dIQs+aCdE+RjQbwYYdBH90f6JX0o8nOAjw
/bwBTZ19Dd4o/cM8grU0EIvbzNb+6ytGRvbRvpK/nOoLxetD9BP0mrRo7p7F7NeyC20gVU7vyrTy
HvsB77w0MAU696RmkiZOnXs7PCIx4HhfYNALs4H39k6SSERvURU3IdNJ6OYdnwcAhHo0MEVbrIT7
gkwQ1rpf8zrW/u0J8VlvkCFVW9U/A6Oc4A5L3izcnjp/IVATpVeyMrsTlk1v3zPpVDrzhOUjpIrZ
1f//DxXgbhIfgJM/rEGana1h3MJZgPMe8sOwuXLeGC8Bs8Z8VVeOHOrdY24x0GBky4Zmo/rTAuwl
Imrz36TO5KCHEqMrH5eTtItwbpVgYwKZrhCX02z3G8kfKgDfFG6a2ZZnQGqwNEFy4jjuW+rTRGTq
o0A8JlGfGXfw3BvO0XR/IzxFS2INzi3KJWb2NVunc/yZOE489ix9PtdNgROpBOVGXL+W9RGdtIf1
de/nKxzYvduH+vAGo5/SGpocqTFpKGxqwkDT6MkCPcuegG2mz/OW277vdpSrqfL8DUuBGI3XXi43
YP8E49jw7aPE675rYraUgOZ4axXsP0YVCJr8aMlh0phue/7unuM01HivrybXUjZQaxrsfiqr6dYe
2Imn3MSJPPwjTel4W2Ind+xc4YHpwA74C+q3CGVbiq1dzeE4u57KFnRuRm3DJdauKk8Jsda+3Fe/
kiAeX7DgzNWMYSujDjrUoRmAPiIA29RSwJeIP5/EGuhmy5W+/OmnAz0h1GXluuNdco2m0FlJ82Ea
d6rOcoxeRt4u2U3hjhudF1J1oQm6RABjWZjbTW6coQYwbKLha3H+yQ9JzilPT/wokTTFYHxXbudA
oBqjJ9LuB2dKDzBo1VY+w/rYZokmVUopECisiZAZiZycmAElMo2BK/uWT72sMCAc/L2vYRqto9fl
f3ukawNcaUF5KzusH2THM22LdRiJUFTSmusCDMWLqpWqm+GECdR/dKFdNa6QE7B0CSUMYSgLiAWw
tPNF5Sce7kQ8IpMbk8RjgOd4He79KvgBM4zZ2bJv9ONknJHbYkimvk1l9qZeK672Nwb5Jf3nHItB
hU7yPbJGgF8DypCCu7dQlmELvuNf/YHXL8fn8Z1yqd5J2nlLUB5nowiyMQnjzYs2xj6MghiU6DtU
fYTuibX3bcZATdaZDhomULyGSTXnBw6i/gqe94yKOhsXtWRPyhqClv+FbK5qaVZEpGAlrfCCWOyE
LiJAmHF9v/UuG7jHwW1vpohpTHh0mdBNnXYAngPn437F6BHX9htShaiYBxupf6pvWpoubmTYRqKY
wMKCrlq/3c78cipmLPEATmx6bZe8uSTG11CH89lCMyh68u9I6Jt/JRX2/QvSmG0JEgxMf6BPG4fW
VGwu7AJgIFEguAgPCdeSVXlN+Ei6gAcNAi30JczPjc+b8B/zoG00Rns+VW8rogl8ukTaHvfsTpf/
AfwaplfCQIT7l1uu5LkunyQvpaKuWOVYTjujPcBM0228tAt9XLelvGwPzUkP2kZqhXm+xI5It73P
Twz2xGj+DmmJ4jfLE300m5g3sCWQwTS1oKfGuto9cN2zel71lLDho+Y/7wT7f3aLbtFcNu0r21yS
wxpa2XsbYog7SEtWh8zj1CECUFIKncr3mPUhCEDPgDtOIxrtKteh9SXc4UneUVEruQF7jdNk37hi
o2y1jYAEbiFbli7KMhVBW0dmFVM290gnIA1BSMA+Th/tEyVTsl8jWkANICP061XXnjGGzyD/tnHm
P3iDR+BPLtgNdTFt5W05KwZt9LRu2WQw+s78P3cmv9O0R+1Ii4knVjdB8s3KPRm8+HB+pM4QmDIj
dkCKDp5XKTHKkha9hssad6Q7JtSAjNMrlWHv1AGRHqU3sv+83giGbvAgxZGObIA3rg0kRmx79zLS
TQqHVOHqj+WpiiqAZT1Zu0nzn5RGpFIOoP/rlLXh+tzZ7QuRM46iXkjpmELQ0ZAZSnbphw2UfEFz
0jQKEtfNCsoK4E45D3RYPLoYJvU2FZFTe479tKjje3STxWuyca2NSSM43G6QErDdrnQR5hcWcjxn
KN3l2KWHrK1WuKWRNz+r1qKAo3r76k2XKOg5U12gqbeZGAYzEcTqNHDip4rp9W1NfynuO06M007F
hJmUdc9EYr8lqrqXfcXNo2HZw56ZV7Xoi4ZT62xb7M5pStE43AGgUo5yQxq1S3LQQbpPG+/aDgkA
QRw6+aGgoy3e37iX2EKpr7L2X0UVqqB++x300bSmuNdSpGisHGivkJJXvu8ySbwq0Xu5mKWLYeWg
XUdQlLrUAs6QMg/1oMpuLsEKCDVzRixSfiJK92PZVYitpZtnWwm3EWT9Rpl4PEWbwa0Wo9uI6Q/5
sPf9LGSNJA7LvQjLYtUJcUf3hpy6hWywaUBDZL1ZIGmFEMGuiyc+uq3CoD7kO83mtmbqIoonXlpe
z4hSEIBkxBi//8YDG3B0XoHX8sCH/SqJjJ/Xx/vgDA+twL+3/TGMP+IKnu3VCsI4TdtoxV0QI3Y6
6Rqto92UANxB7736vWWXz0zpbgtW8MLi7YPJeWKtLcS0xzZSb5REI12MA1z8TLLNNotLO08qN2EG
OEmDkD9cV+R7jnRq1AF7zcGB7R0749LnJXQY1SpvfCdpvuoxuhsGCYTjdAxKOe1uBX2k5nLA5HBc
bL+vOXGyu8NjHlDkZrg0xtslFS16XKuZ1igwveWEWN8KvMCDSAV7wpJ9hicbHutCS+qcVDrxPw14
taheZoO/VQpcpHe2V6gdGjDM36+2RoNHyg5rJq4ZnF7KDNtaZkze5Z/cZhJB8i3GQcG/1165Ow2y
n34LEHF7kPav1zCKS2K51O3ZRXIaurEYhwYnavqrkHYlY1rHIcbZ0U4y5DhUokWi18OAS9ZVDDz4
FIqSBT36nFu3MdVqq3+OrI0wWPWeJQg0zGZ5HkY+A+40Y8ilH7nuGJ2b2hDj75DSNjvyIP8JIgKC
XjhW8QeUZpLA6e5lAj/7WH7UUDVCeRh+vJgcz28dOSzS4fErZZPi5p7BnOBgvy3MxZfTyc780e7M
iC2UEp8tfkCRsDSo8SdYIZp5qHB8ZkkoJaGwTmN8VsmRw86i/Xhvsmn2/RQwPr1SibECOx95ekss
UlanaB2b5Q4FZwAOG3mBrgYdU6KIrc2Rn6fjmxK3tGlQmU+zf+IkmIv1mvlPdS5FBo8ihh/SQ3y2
gfLI9w38Ow6ggHRSGO4iMCWYqCNponMdOUyoXFkw8ZhyvAC9Z4grUL6jB0ndLE/cVQsucP2SRJ8e
OkqFSKwPa8Z7R4ZDwCF4SgW7UuPWucc93I+6CW8vmUsD7DqsmI1qD/gwBmJiuWWZEZUEebT36DLM
+Lx35GMD031TNB+0Fy6WSTqwYscnuyLd7aVNIyBUEoWRtSGut+MrrQ3YBi5JRy9hxxo0qe0fcGHn
IHWxh+/I0WYI9UUwaehkItoLYmpZ0psLJu54ljR0Po1cLQ8l+rH0wsz9CpcCCNofa7FZBRTyKDnu
m/xsVCPJI+Out/YMq3bEiuD5n76+/1dax5hz6KZyJm6Lqel9wH3u6Yq7CEiNO12C/fH56MmrGUnd
1j+fDtrw40qBY+AJyWUMqzyZXcnlHtpTH78kszQ+dTXobe1VNj7Y7zJU1Xh7s6zsAOCwBWyLwSPL
Hi1fpz4jrlOP+ynk3TX09fn1S+jGnQVVtbZ8LJ7m4DQ30xjPv6w1wcP7QabeqOrJIzDXndY842jQ
Ufpccqqm0tsAxn4BDcBRPcjWW8kjcJrHQ2dTOkmE9RJNLz7YvkT+LkvpqGmJHfjjI2zEwE96mQwE
5ViEs7vGFeHY/PoxaWSw3VKncHDyGzyxcaWBKwDfbVTx9Qi/9UFJMBQ4tmF8rq6GcKw+iLGyyG75
zlh+ckoaSVkOU70t5Fwz6cUps2vvLijLNrX1iu9Jd0s2bDaA4ZwWs2H8SVdCInW8EY5605tgMb1T
FXtRo0wahWBhd7Mtm3A+f1WP4v0Id/r4WeTLOXZKCu0Mr0hlP7tXxlLhJ87sKQBH1auNDwiRYiWr
Jy5VgtTrob+bFhJ2jxJTFTMB2pPQjZPZBCbIyXwrDLllXB27dWDM7ycJtiUeHKQtm3iTOM9ASObG
CzrJ6a941KbiTeSs222+myyOGtpNoKA2pSr51lXYDI9oexHx6eFbdzPB2Id2uYkDJjaPc+4IFSe1
wlviDiUxfyYa+j8/9L5DfEjDgDsrVEZSAmExU+oQ2cqzFpp38OWV+oPe/axfdZ5KTcGI1VtZlbLN
/yFpO834qqv1jusoe1mDcLc7bYg/zwPoni4wyCtltOERNmigHB8fPsiC/4UguS5r0PtHRXEElEjk
Wgbe2wJpjXKCBFCwAVD2r8WQ9A0iV/EJOcbETKOqoLFeAfK/TYKD+70pmSdfB5qQdZz5lL+LUX8A
q1UQM78zMbYYm8RqJ1HgoFMK/A45bDo40gtajMnuSvvITK6N3QqXsKwipkF/C7gJNY5YDsZtoOPo
0n8QygTvbyrm3254cQNpyPkDfRoMFgGuuwcGm1eKTDOk5vtkB5TWQBfNWJtiBKGZPujX3IuHs0EC
PbHihfmb3TJsXq/VmjT03ZRFnlaF3Dqdf79U8RE8fRkuFNrRIb3dC6KjT1j1QjJO32N3FUP4R/sc
JnkDkjnPwVkyrocQUk32RXNGvd5FJpjgbRC5GzlIJN3fjFT/sqPVfUFQHVp/zqJAl5XEMUo0gC0x
1anv7gdIt1B7aQm/o5UHtxNvOW5lAhhg9sGICvg6RBgT2OT81sPNWJF/JUX3qcr0tiidlNPgJ7eC
eIb0nLZuLPztcscv/aC7VAkS7v97sm+NNcYTxsKivDY0MU5ja4xbWh20BzCZ5EZKTSWryHVcEerl
0yQzZysKmelm31RIygxlQETga84SI7YoiY/wW8RJDqMaeUpzH6YWKLDPukOF3ijr5NfnAJKM17cE
A4R8z5Ywz8PLO4St9RNow6U/6fvNWG1TLfii/waWYoLqpZCEpKh9ujlC15/C/bz+0NT+XLJUamrq
BTlHB0b+7Se6zxgHUlTlb3WdEkTxZAlMQMGr+ytX/BwnOXZ4z2Kw4fZVZ2X9okSwRAwxdhRljJoR
3hZ9r3tILQZpQzetfkoZuTnMIvyx0QHLbIBDU7g4puaA7qKuOzskFJJeBCcajyBW/eaEOW1jhrhM
iU40ZCLZLczwHWYZdmWjY7epxrQ86pRxDjA5lypIO4R2v1nE/Wyf95cPwZSD9eo3MKmudRkxf2XN
FwtZDVHI5TxxsRzOWnuh/eOWMIFyHT4dPT32DWgDeJlLVjUJCrlCeuWRnUjczfILwdh+sGhmxUhS
yf2m+Pvc2rD5HGZjIRYfQUxn8dqRQr2YHo6ysgIo1MvktkgI/3BfbFGKL0JGBWqI2yqvx8adHDbe
Dh6cQLMfw2Ta+05FuYSX8Z6GffJQi/0CxXahcWKBsibhh9q3Kx/Dzgz8NbGChMQoVVgvDU9pAzT/
Cd5H7FdisCPgIgMph2vfY6C8o+9KT0gRXs3NDlhVsdpQ0DW69Za/KLF2odrmFJ3DxbOBQKQPk8Ok
xSQ/3JIPy26PduEjJUmHetkA9BkWItNPwY1s8ZoOit7Hsb4ugpArO11Rnz+99dAEgaTJGWXPIkLb
C0+8UcJaizFU3oi2gPlS76jxb82TVcNp/OoOKsqPwboQz9JQ9DAORS3hZrJj9QqxkRw1cl88wa65
nNGpTLsHM7rrH8D1AkwDN5qmrDp9J8wfeT0eeAJzvhQb8tWBSecM4bHrnF9pewMV7k0YpZ+Gjwq2
hM8m1jdn5fEen+YtiCjegldJlyAyag0cseD/a8QlKGfG4+w8d6Wx/AZ18ID8LJ0CWnXGJiPz6wSa
oD9v9DAqBYz+xtlLCEUXCgpLQ1yioZWRP/lGnNNYQ98hJdFjicKAWC2X1VIb+px+4pgwR8DGGuM+
jP4Hpfk7KOz+H0vV7D33TbydBaMMuF0YR00js/0y/vdEyu4bDF+qmnmM0zpc2g/1fE+Q/7ZRU+0Q
63FqkSbVJVnQRKsVyuGw2pPlQmZLWQLcxWZsRi1Jy5i6aBmImCJmqeOh1WHbAd9P7FRwTpTSmjMS
G7xuvlU1KlF7/IX/zzI5m+LK6xIEaARSxmzDhGhyF0XpOi0eG7z6rLFxJNgvlNjLPXx77/fwFaxp
zwBGUmjTFYY+j13TZt58r6gcb/kZbU+Ztb2iYcqYP66erDqJQUN+jg+iUgqI/N1PI0w8Pw9ojKY0
zyH2T95ZJ2c59I8DLKvnJ349hMH11l+ACNdya3Bq3G16HhPrFFaVO9pWcYsupxnUxJgYvWcI6YZP
iAejgHzydTV2eWhfSU2njmVJTLy3278LxKqE5SAz+OgiugtyR1XmrxpqeL5VLmpUwoyoX+WMfpLq
PYGB1x4zLBQYpD4PENwtA5P+nbEeIMdp5ONZQ7mVnSus/Pg/0Qaer4tgZXKIw/X10rR//cp++V2l
PW8yCh4tmySULZGxCBwuUzArEpLf7aDY5RZ2HQtDSCZTgu9+tTHTTWwxqMFZMAIBOeJUwO0fyup5
W+3aARUYU0EhKLe57dmSX45yRcP0i8x3WyzZVpQlMx+6mtbCXxhXbVkboDvMD0Nc+1QcWpjWfmtC
8jfEwk6VUkIAl3FvHciCg2MDcfNrOePJBmvs9lKzS6h12idBtpbtHU9zIayu3DKFBvHQ1mDqcc9a
8CSTHAkbIW075D7qC9lgxTJ1mWuMYURJ6IgjbysMT2o+Ldt4q001s96Brvndg3Mcl9XZRrLpJFqQ
SnIbT3MC+VBCkf3+BjXAVVVNxSCy6lRSD7s4yZWD/kv20o2Pj0R+Lti59ulnMgZ9kLJQF13/y8C1
qISxDsOjX8JeNkfiwNKYwymUUV7NVGMGeSJAJ047u8p34b0QZrdLKxnuVnntfZvleyiovnLTg6PQ
9XchwBTk4flDJyCmFOz5LrFxvFGZUvQKnL32unb/NsTMzJOdOBvRDBFxwbTr7MU0fAbKbVSIuxgn
IDhA6gMCXiZMOHwTXnk6DQYw3gZK8f708hTFDs23RK5ZNJa+ttRuYHs9BCjMwLngzsR+lGc36dk3
bA3Ew73aHE8QyJzuSoMshoQnlaBttbn5RmH1w1biF6r5CzXW4zxsV4vdkZy563/+I6E7nHBMIVIs
KVeLDOwVN5NXLtW5AbwhZXMTMFkdEi8Ryx6hGmfx+28sgHliDTFz9ave4qfldQqQKXws17k/R7zf
HcNX/rrBcvAfO3d5bMdTJUxulSxrk059YU0/XbfDl2em8A4pHGukJp8/eyXgCGPmS1JlJ/Y4HeV7
ZCBfTsxvyBP6hyDtukxpgLpHemrVpKLl1pUgJOLekglS3SmnA0CxGyrPGEpPaZkcqBfxgqIXpKa4
43Hi3L8HAzl9mr/p5NvTNd73DNlZE0sehwLNXF6HSHhF5rr5qO7kHaZgqefvZ11C4QClasanlDe2
QPO4ZpZ7lsKhmxw1iMeGamnju/cdqFejIoKGvPHkRLpbg4w/yLZXIfiDAGxOJlwwnDxOo1PymWLJ
6i5XHEz9qKFnWAw1kIV6M4FBPvrB9iD7EGxSnzECSh4fUDUVGSExKJELugxxft1NuxXkOerD1l9z
3xVSpMzZqZ4W4tuBMT8NjVChJswnvJhsyltxCKYwtQgGJmFRGi6xW/plb9ZDHaF+nPpJmlxkIuZM
s6WRwh1OES2R9a3InhoxCYv89rR4GX7jH1ZE9favauvmqxwOmu6nt8GbxLCCZoKEYQLqVzmSDolf
3bC+IP8H3ebPs17vOP9EDWTv7RvYjhOEVov98yLdZv4YmAbouOOjA8DwIEsCTlNO2DA/+/d5Z1K7
umiewaV6BvlcQusqQkSRNyzO62TnsiulI3UptkHSkTQp/jhGT/LidEEwsufH0dYaRKwRFVD1q58C
MICrYIwJksbzjqcBuii/k8/PkR+p8KVvOgPN2YVU1EcAbMPM6JyxY706+uZgOaf8Nnch6Fm1LhfH
ZkpU4TYPgwR6PD6PBNmatm6yUf5+CZlWj1wHvrxRzh6HTEHQKRDLIMjojykLGCyk+QdjpIpNiDV+
vPBV3DSsfhWwa78lMvXONE0v58ngdLjjO5TFdRfoWRZds/m1AHEfUuKtNtxW33agFC3guTeI05ii
06cwgmo4XPxAS8eyt50hi9tNkJUWP7Se9aoPJF71UtYNTBsc3LmgrqcMVWSEWV1OoRFWiAgKd6H9
PhRXLfXl39RuqprsI/vHPK/vaptmy0Gz95xmlLI1CZ1tU+ISqkr3qh4JodcbzGwuW+O7TExXM/+p
jSZMZMFvGRQwOGXzyaCRzdPiBbK9H6mmR6iBIiwMdjuxlSqnUkVk4rEl6GPFwFs5OH0FFken6PjN
J7d15l2uUt+RjrZkT0H3MZkXJQLHKIIonxH1XDZiwVDw06QoJF8HnXiNxldBKWMUTmQKLJjwtrUd
ZGtAUY7cceQsJxKrBdcNOt5EVqMzFuLFG/3O3CvS43fcMHnXg7/NYhJjTLo0NgMDzr5qj38KUO1q
0+eb/FrYes0DHOUrMkdKIJWJD+JbvUWGUBw5b8mUQ/vUMWVmSpjujgFrOSMPuctccVPYXWhDijCO
WNKJHm8LsiogBRpFo/6zo6IM665y7ovCq9Ibcg4Jqs9BBf6+dcICzQTFVNbmKtOM51JVOkXtwRMD
SKMEKjAV5ZuRJ8PvsH1tvWNCsaYE+yewlv25h23b02Lm1LK0rsvGjpQOV62eBeO3y2J43qKN6Cop
ALGxx3aVWrap+ov8IeyMpLvfzX9A0+IpRgl+BNuXIwKtPkM3j8NA3L9OebyrDMQOCC4nXo8C5XCE
M4mWojQYtN4ESTaVeMhs8rE4ZXlYzSc/86EwJW9ijtsqMYS4aHLRH+6R+LcsM+nERugp5rknkx/D
nTFRkpAZRZARisZzqud0vG2HoEFHZYHL3ZxonEETQEEwGEaieqi53GoLMcRpm0lxhVmAgEYQaFp7
PPW1cgYc+pMS2senSTIQdwPQSBeQUvZn68T1LkNJx7V/45auxdI/2tMnQy/8sGoEAxGbRNQznUAK
ya9QANjeQ8nO++5NT4ZNUZC0KG4UHG80gX+ATibzV/cq7P7ZLBTtOGJFpZLVa2cC7BEuv/eL9v5Z
uCuCAq6UQwjG494e6LjytYsMXhS+WWThdO5XJrpnFYMbZO9Wq/Sj5yd0ROeJuEthM3DOBAONh2Tv
7FvRNGKDaHkseI4T4GKescOj3LXL6AEnA6JTbHjT2x0yweMWcm3r5u/7pz9gZTqpeoecevFdXka1
sA9X3QDgcY1FbRg8fomn3c+FvSiG2bSWBl9gG9lB1S6vatvb9ApGm4n3/a+DL0D7Ny4jvx7I773k
fJpaVPqaBdSXy2KdHtfaO1VtOLFk5L8xANywzy9KFCBjAcySulVCGgvVNMAlBVZzlhzov5CkheQT
Svi1iC/9arQRJMpjDeJKSAgeUQQgXr9UKGCUmIafoWWYbA0t/f3RyKIg9VPT/Ti2xWCBwm17Lf6v
efM4okU2+6TCaybX1YnKgjdM3zBqtwSSl2FLy9xkEg49z5v8OzDpEUOQVAwcqFppcSbpwdgKRkgs
C5ZVOvg1erBpomRJX0CWNrQBbaYVJO2AZ79zyWOrQHi8WmaSJYfoojkoRNKL6WcwZMmt7yzZ44IL
CATKzQZ1xNnKJiYutOOkAgjlAAmcaVjr3CoOJfoezmbMHxlccW5CQC5JAj68HCOW5fULJFlhw1p0
gN9Gnt+cMxRqVrTTzdIbXlKY3xa28gPRHoOGoy/cGvpnOrD4/xf8mRkT6IW77LnNXWvqBVW6VCc6
6NrcePOsQpPZfXDf2UD7Sxpat0qrbKuaWLWXCnQ/Im5YNF7Z7sDHwPxoCxsNAqYviqvOynsjzmOp
gfX292LlH8FdYM/3eXdKNNvD1ktt9mxNt0UDXG8KyMO92nSlfz37SkfyF03sf6Rf+a5McmVMFyS/
8JoVzDkA/z5ESHBZcO7ba9Ed8XvRURzPDzOtIHAegQQvF4WiHf9yTE3EE2Bm9qUqLE/tXg09E1Nh
9V2r8Vfl6CmlcwyDl6xw+lOViyv3jVF7pp6rwmzg69G5feUh19Z2NhS/PjBltmm7XwSX2aoyIn2G
zF+2IXBYHhOvwWyf1sNmBXzGT58UGFGMbEVoYYCOIxQtFDssO78ZAHiMp4EXOYygjtS9964t0MkU
ksgBZoPrNj9NbNhuknxhqkAzif10CKA+yzFPplGDKhN2Mduqf+EKdVbpTG6TmzLBy+uV6+5DKh1s
1Q4IzyehveJXFWpU39hxAJN1R82fHEFjbNhReCFVHgxSQaiM1Gh7boI7xEWAYCqU8dfFKqPu46aq
DPNUeBXtuEncjIz6lRmFI3R+bRGmdqCkrZIcFYcPTHQXWbPi7PdmkroujoXzX0AQ2wth04uStzlf
nSCMcEurgr9mVekKqYZYHg/wGbCrg5MOWZQGci9r7212mShKQb/jR+2/aYBrerH4snCEB0fSk7fn
kj13xjX8zw+fNbehJ/UAb68WCPUOLJLquPUcnTwJF0UAcATuRETpA/wtj/zfm7t8yd9OC/xP3t5Z
gX5gePj9UA8R8HRGKdLs7y5J1TUAqRXM9/BjIQAgEAPh1JPoBYzDVYLxoKssPYBHf+tzxr+Nnlq+
ojBcxNba1/5f5acObRsqZpD/MbE2L8AeVYufuy0/fZxT2MylNRe4tYfgv7v76oSEASN2znxx2JWo
9WDSUrGJ/skYNJV96JjJ528PhGvj5sB5j65m7SfOTE68UXUsIwmr2tMzwGl/r7GBZdx3hnjaCM6z
bIiz+xeVZYpyLirArenOrUPQRai02z8uloZ8+0UMmsdEdwIMouWj+KA0bxQWMVhAyj6LX4mp1QJf
MCLr/b9W+JqFB6bsXyiBxqLNkLLpw1pu8zV1899jamaAN6SecerUsIop7QUufX+9F97pl+MbtDtz
InvDF2rDJKm9HVJF+1gAx25+ZrbueO0hOe0PWxjMLBrjfDJGHRZgfdLPZd2cbNROvBnqy7UdCoJD
UVb0VqUz3HpHXQC4Opz3l369UaK/zI+dOSx+13cJ8ivCkBSLrjJ5GYI9EZNysg2+lmn/ddcToTH8
QwUGNOAFm1wBn2Fn+Sz3UkcD3W4HQnBEzuWiUC6ZZ8cFum8v9vtmVvhTDq0cBMQ6TXSnxzORoSai
U5giEyXzD0M1WJ2OxfIYH9em3M6gXzL4ARTnUT9YwKVJeXrsLIGhUGrlq/PN2d0pyEr1aDlLj7r0
CwETz4Q+q0/VU6MfmWQUSKXol/UGhIi9DHs4UzTN8N8XTGGhueZA8ZipKa6mP1fSKWAf6jrba3CJ
MpeTA86tH8zEpPans8N9LfIQ6jMX10r/lC2OCKb3VQB14ldfgTM8GtMO49nZIiK0FpXcX64Ej2BD
ZM1L0NUskKWvK84mcSOyOqdwvdZnPgBXSJUg7RWFRhrjX3rHUfW7D5x7rgveXatcwb5Vii3L3hsw
cCP4gl9ymN/qgT917Sefu+JDEn3jR+CrQchPOFnhsDPMoz7s9zBVFahNV8xJ/ZJyF/ezktbDtz/w
8YsE9cot4hoV7ChW6sUrv+rVxTG8hTkmSDKtVSsjW31FGJ1UBfbq6MPmaHtMYob7+cUyJESqikDo
HruJyHlzHMiwGXEc5ZvKdU3hdYPP0UzgzwcRoPt7PJBxM6UCbIWT7/tJVJ6E1DV8Sg+l/73UUgus
2q1XFh+KYhkJ7iH2FO2LTyZ50FmtgM/cx1rEkV8+Ap99/semN2XfdYf1bb8ObzX288jgxZdJDcu+
8IvRky4QxMK77gYKu+ZLQ4vO2IQ/QBa96v/I2ZWBmprZ9Es+1vBFJuwUZfNp2qY9+/qSizRl8NSm
ooXh6UduUTFgEKYiZKBXqaNkpGfOj8vxSiczZjfpn7T3dFggGqx4v0s2pLz1CIMIO8I7FKOtqybp
FG4zFh1wWkLI2AzZ47GuspT7OQbRHWsAjrEj0FaTpeGahF/XiyAlUitixCIQGnwC5fpqoJLiU3JP
jWC3cUPFrXvsy4+cKDfM+k9sHkRpq18tGYuALZXx7K8n4eN6/O/B4cisff2K1fJVewYJdzkuhR1W
Q1EwgdUhca2uMaY5FDsswpmxKD5y1rsmlqAFWz+bDnz/gIKVUlOdNUGuEr0ZPTeLgXgtvmPboRtK
R+vSm2GxBXP0hsAVjU3wEKQjJL/y3tuqIDe3JaJO5W/SyzjJP/VMp9aKX4g2nosEtRVZV+n1cQCT
XBh8hYtOnOyrhH4hnxgCdw1+CwQx7kS/ModAIKneLj3W/aCCiAYRJqipcQcr+ThrOaKzLx7d1UyC
qcgJ/5RdPWSIF4lhPuVBvUyLvbGuSe44qJQ+5LuxBPpD4aC0rLEU80Jqt5w5VKfHGGbXNRwKUilc
8MY5oZQUuZMHncValBCT7zC3wPSiBTTSe6DtcTmTbYcu6re2I0jYbkezMLpChojfBA/KILjXV4cO
cxeOlw8YOvv5os9kBSkRmokIrElk22+Yt/w5mwJyMV7Uf1N3zxmLW7Nt4sSNbieEbHr37+aCDBs7
fAxvHuGXF1BGt0HNwtalWJqcoLaLR/pNxPh/braiqCmD+FTXAdkMihDQrQ2G7t3+dZrExeId2fep
DlSgYV3o/k62SRRZp7HsTFrZBR5Umfe75SZOsPDHlbmu3FwLii51cyUED1NhIeaHRkUeEafpQPsJ
dubtI3iBxIh3CMBLL3TO76u1ORB0GKohs8O9SLP1fT4u0jkctlnsbI5U2S49WqafYV4Mr87pZb8o
vMNsApPK+0pThxkeevs1EN8cQmt1UvSuYvmsZpqvWlciFytwjKRvs6eMIwJBQlycZno6OAZzz8Y+
95Yb3eCrQMQBxwS777l2QeCApzyKR+oSzQELt3/L+74o4daIRnhZd8Kgp4a17dG+YWL+hkdUl+3I
z0DusWfwDQ5Ie4cGtbxhcuFC3QKifh4jrS7eeIezBCocdzN94zlutpc35esxCtbd5sES5P1WyPgm
nAd/A8BefgVnNlgIQ9V23jZnfKE21IabtCUMTvw47aiuRs9tjnGOcCXJ0uvhqTUZn/I7Q+ijP0CL
lcq+P8hq1xoyaRTiR7yPrDXlnTaFkfcubpFBbPckkDQmAwpakSdQX+sFinV0937D/RoZhEYpFjbh
HGX+RZ1qfC9bdMfAKLEm1zNZ28SVjQOP3Yvi43xfO0i5yRJgqLw9/zweAdUIHLX+4AuKI1KC2GXs
ggxREunsO4zwdQcG0RMqlmO9Gu9qlwXzcJqaAGZeeERzVOT51mBPY1REaAzDX2gJcGjMPUernH3J
6gg0y6O9fzJkPoCGuae/eErujTdFVKrkGbOl/DrqgWCzjpyx4cnwQtmruj2FFD5Ft3LEHbSG/hOm
9Y6q82f5iPQVHJijJtR5G6O1NZn53nJOE+NgElMdKBbEmhIuQM2z1TQadf4k1FwBzoQJbjtQnkSt
e0eiaYGPPIWC1X2Spxc93UqYnLVS8p/yI11w/1mNUIX89eXo+wnlhVhXHj8bJiTjOt7+2hsUMJqN
nRGPAdgtwk4h+lpA673gaBAd1pJguhTjkxHXwg/5Szls+lxRT7k9jQ53MM1hS+jPQFqnKyRsrxWb
wzfGxMvPHoh3RNN1fe3GDLXdEO6g98DHaDNT0LO13tsarXYi+YCwMeoJFjfk1hozgTQze4btsplo
lDvy91+K03RQyZL+PfW81V78zIlZ/4xpJbH8yxRjpCHLq4uoyZ0S3ErDWbKxd4r5/lAh/gmakLmg
/L5eJPiZ0o5ptBb8UG8HWX7j7jgS3YobVyiVMzO5TYl4qlruyn3AV2KdvPORtruQcw/mi0eXGVW8
KTXUat2uIQlQFcq/scRR+Pbrg6mlNZMZX1ZalPlG8Xh+ew9D8hYoY2CQtyPICd+HwRB5aVmgfCYy
flQXoOiYvg7g+o5lSwe26odlHBTu/ANv2SJlHMmzG1fj44tTzrTKfBjFSLsOt+/Lxqi7kTaHTJx9
3YMgy8N2Imdb/3B6cE1LemSKczxisWfnh93Jj+tTYfLBvawpgiyr12R8dkn7qTi2KzHf1QHhPEoT
/8HodjewWAVY4WkP8hni3LVAHPd7Znml1xmmCTsKzFdCm4gGlVyYHd4YZGNiNxXg9CdvqHztXRJL
cPC/CTzxLUqWw9XmY57JbehjAZ6Jg1BURxye9Sx+IhEsfeirARwAwLG7EEQ73JO6ICua0B3BdigU
sr9Hbc2uMjbRd9EAjXCqrGGU5k1TLzHNWROkWG+oHTUjMIq11oWjDwhrB99aqnupFXEYkqlRB8DN
XDxUfM798YnyS9B+kbawoCcVcmZSbkmkRJTmj84eDVRcngPNQ1h8UcH2ewYl6ROyMIUBJojNxfDU
e+x5ie3vDJWhryVWqXieVJHtIsB74xnBPpAAgvt/hilKalt9PcPMc+u3cR3aW9krYfQFZMtZbrdI
ydimcrxgYwEd/emz5J6DE0BOrU383eokBw4+g/MzSTb9JMrcaD+akuIHA/Cl9MXM4b5/10lYzxJQ
fya0Oy4AnfbJ5bNbUFBpdZcEOw6zs+gX4JDQxXWZVuwzqw2PDscv7PgPLN3W9mLZ51hjp0WjwoIZ
kAp70qlYuNBCES1dgUg+EORzR/GSRVKKcNOus9p//Va0/NfDcmENVVP4odTvbT9sSc6tjSulkCaM
/aydOPIspX8orRf//yflzgrBJdXQp7vJdL7YF+laDpjT89f+gVQUgud0JBt42aKTpbHGNfBUdpl6
qknmn3KQ84pYB3kKt/1KKmSzjC979zDQjq8rMVPkJ9wlycH48iBjFIOmCzzANavcNsrtqsFXxkrX
3NQbkT1kLoPhWa/MkzjPk1nujt5IkTpHZX4Iok5acCdyvNdg5C5B334vSdVIFVAT52Om0u5mGelK
tsDgACVSX1oVgh45539pBSuAXHg6obExAr3j4gvg/70WTuQ8Y4/4onjikfHBIuPpg3nAciE2E//E
OxlpFtTP+6C2RJxIDq+75eNIKnRDo2/ec0xt+xTvHuH64RPJ4mI9BTL9Q5IwHEv+3aTA+aOn29Ab
ZqTjNqmnYD6umOLOPL20UH7Buw8I2arTxPWXOb3tzyeMKH1o6cGhk6TxFW93gLGPUXjuYfx0LSiC
Mo/JnkJVpkyT0rAUDUOLoAFADX/WwYo7j6aajQTTFXWrNdo7Ay+y9CstDeoPLtFO1QeAEdJdkgHM
ezbm2WoT0Wumly41cCEdqBkpyAOXKFiQ7LllWvlSH1KIbsFBr69l0j1iHa879dsdjN4fuzgY6u5K
clwBMLoRdcS9Kdi8Ktv7AhfdrgLo7JEyK2r7oQSVx+osr26eMHNkXZAI/VORNB/RbIpeXIpBZIax
7b4GpOOpdesg7oRPkE6nXWWwGVYmseyKeaUZIh2gOxw8bgN9FDdzEFqBUDvGCvNwKnt6w5Es8W3h
fkLkeX10fzbYu+GV2teGnyHWEomrBzSB4NDP8p+//50uULGVMHEYKaxqKvMqokkPmUx+4NiDpxS1
jSf9olFETtlnKhWRM7N4FL7f7b39qbqv3Eiq/lfMGkxtjZMzWKILgZKiaCe1xlDNbiRpXYx/VMdB
ROJmOv498HTQ9m7j4dR1eCMzIf33sCYXiAreVXxWSM1Ac0t5JoesebTmbZcF0vVxGrNhLKp5eZ6T
z6CBGqSOmJ6h7J3w9w0XAEJaLJSyuQO41MLixk/WO91e7SlUdLlVoS4gmlDozpo72k7TKDuJMfOt
5GFrU8Gd0VvnKi0fav6uoEbCjcSZiTCKFCItQKUmJn3nnypf+iWfaq6u2jk3yxdki8thGMWmrVPY
yEmPRyf/qgQOw42WabenxtdUzt3Jpq2p4WykMLW+KGJAgslHatiu/PXPIFcNzljBXt9tBH7xTt4w
A1y3GTxeEU1Q1piZuSv+jdnSr5HYVw2WH7g6cba3EQuVKwEgbkCkRlDOvYfDF3MsDC33GhDw7+Ij
uAP1emcY2Lnflj4ry9new2AOB6juqgskPDTJ5EWumQFLVfkuPtqjHfYGfmr5fWlqOKruENN2iJsm
A+yYPR8a+u5ZxCmxgL2XB4qaCt/c1lYZdB+fStDGgYGinqArDLTBTgSEaSucviMhO7DeVqeNDpiG
/5n+QQyrwNxgg/MriLnHar37TOUui1V+P76zW3ZVHt2dqYhZCuSVJQe53PqzNIZd3xc5QR8LKvl1
ilfD78XVBgwTO42JQZXF7TMGlsKz4PdOj9LwA3GscyXUhxU+WBWatof2eUVWQrmzllgD3S6RGlfm
YtrTw0WhXssl91riMfrNQI07nNQDbM1HtTsTAidj8/IuXqknBTOar6gzi4reEX/1xVwIBkKrrbFw
qma6OWm8WTW+W9AslCWDGD80aZaeG/rI1uZPAYrK0y8N/QSPRy/Ws82dFpdVjG4zKvnegcvXwuiP
advjZP/mheBHPU1sIVOW2Rg0u71YZbYVK3LoKHFREZ2ihU8RbTfP78+bLtZHlB9PQn4yZHrEJeR4
auCze3Aol3tQ6g07GqZbTUeAvjexhKulyCpSkPscR/9WTEDFSoxFsYDVc2fp3eTqFKbiQf4KBHCW
tieoe+YbepyX0cb9/Rb88WZVUDWTd4vJlN792A75wTP7flIGBUp4WA8D5DE93lhvVfbP9V0/QlG2
KF6NXxSWHb6m0C4FfJouqurRF3gwQd68dICTebzedChYfcOaPe/MdokDFjm3Tu8AyezxRIp6syOp
lmHm4crUSznbNOlYXNHe96KORuEQAKG0MDO+VAXfz6QgrcenZbXah6OByUlzetlndRR/mAkKhEox
7s4XEYCLjrsadLAP7iNo8bjKH16k/ZXKprgHSdIOauFJiPohDBZrZaRyGo8HwyfMPbH40Rv7JY5k
3SD0shWW4eGdWtdYpKgc6XhQOQZ2e+LhqLD6N6OLRAwWnFy2ShCIDmdQlKZVHwvQCtTYys73AZq+
KVGIJYWsFxUv9zxbaMX/YrcSUPeIEDFSjPA7fB9cGNxlHdN6YpmAPVilJz+gk2JAIJeDKMEqJ71O
jHpIHCgeq0maUaRA0K9AJAfrJMjEm/HbKm4g1ii/xsxy+YQC1LBtFPetECTIaW+VZzwPD7kV9QFy
ReptU788NYT9RF1VNHUBs85NwfEeRfwRVFCGBbpHVjO6ZzVXv94iQzzsDI7gXQYLOQVfQX0//NQP
jP3lXLOxxPLDWspOEK5xjUBxhkO/7YJxMYqr6iNIrTdLUpCsXE4qXA1oGrUF4cCLJQZvExc/0vcI
7lqoSUIy/1P5RAlm7IJ0ExuFOjWw9f9lPvuAoXGF4Bz5swmvpJe35EFNsOD/Iyc/XjfECtBitP9a
cvqdQ2+vHekGEuZZg9R7G+4Vuc0anECiiEAwPZbuhd4U3C+oxUsNoE6YT4KddHGhrcmBQPcNI8Ow
C+6/pa1+31q+qS3gTlRDGYT+kAZry9s+xiFkEYhYJIlOvibVAtr6tYFq4TJoln2AC+W6wP3Mp704
RjRM2z49Nj85x9EmtFzPvjHJQIRigP3oiuM3J0u69xeUJbTxaDpuVB1QIkdpR8YodyLj3PC6S1gY
ZO4eqXcCGubV1JKMIhz6PCujzBROWLJ/m/TUReFvz469CakGxVealMhiBrKttjizQme9ZOnRaR38
+deaqpiMgTkzDBFE0K+PwZP4HJgI4rYgIgObI+JajVzFLT/TI5GzFM3ax6AjycfK3KKWshFNh9iD
C78P1QAmo6frdI0rCXpdGufaKRGni83YarrW3C6XOQFnrCKQHte/KtUUd0At4mQTY/SAaMwmkFaf
jO3buD548bkftjZn+0nTDkaRwt8JPTh7nHMGA2RtHitgepJweei++OxILh1KUHz7WI7oYn7d+ZaP
dNQg3ZV03aVH83LQp6jzHtgmH9fSKbN7e9293wOuRd3A2rYGK17wf/kizFQ9WCFF5SM0wTGhbAoo
RLJ6zk0WsI+NAltVQLFNVQcIUfQeBYMOCmKFRt4hp3PUrPfTvBGZbL0Fk+4Pj4nXLBhP6FuUjSAu
d5F+6PBdcbNv5m8TG6AckMVB09pjQZQHMDySsE1HG7tWDfpsozI+FhU55W5Dpsg3s04esFLfF2sE
8aMlglLP4Pl4teUVygLTHSqoN+BPIclY0hjo40zvOebME7smK4k3LOmqQnMUoG/wGilDUblqePjv
Oneh5KSFJuVoKwyrAv0/3X083kw7b60/MiLb/gnEZlbNbB+TmPyYW65IPieoDAETyqsUWX5h8Spb
lbCIzA9fj5rcWOSCRyR1Wqsh2gkS11z/B+RJVaLBKgTyj0jPvVAOQrLMl6zIpE0PqoSFAVk6sduG
hbqpbK3eol+ct1aj2bUHJSS3dEWE2R0r+/ivuYgkvwQJAQAuLsVSsnDNdBetWzEV6b/KKDFaTKPT
W5XWOLt+tmGZlb94O48jjU5owJwbwY5HdtIogg4vIJ17aqjaGtGvyULmFSdsYewv8pW1GBk8PmV8
pHU/earA5yLsklobuUrwZ2j2+JPg+vUt3TPSiD82KlrewL0NYsFbL8bOLqe62LAyZuEPVGLF2Aow
VutHCx+ZrI1UDfAHFC05RCF2gsISB9dmavJEGS6+VCqkEV+Io+8+cZFrCy0Mt42WQnPEOLT1DVcB
3GX90RdSiXeMLD+iAujIJzT+pOsEA3St1YmBaOltc/sNh9i2iqLxQGrPhvoKcLsDv0FrgUikCdFx
gTNHKUnGh3HIDVXproOq0R8jfHldfjW57LbQY0YKaXEuTSC4b5c+u5R8nC1ieQkQ4iuS9F6oSZul
kVkeokklG76p3+njYXnECu6R6HBgLPLgrCFR5GY8Rg4SdmIZGtTdkoQOkzDu3bRPVz18cyFjDgy+
PRMiPLDc0YS8qJ5rkf05mUmj+xRKXeQi16stfuMF43VPegMLrzzxj+RqMd4lytPGq/2Ui66EbZ5r
ZiQSfh0upp9Yh4EgJrOAz6wU/3EkNcgsJKLp+thuLwWH+XxaExTVRRhb0T1QrMf/3otd9K047p2P
jL5nYt93Vht8cvYp64jMr6KWXhDLRHj1J4UXo3xH4LU2+lmgb2bMXbJfwk9MaQ8Y6FSSTORbVhYu
5yvPoZKqb602JBXI+A3hzBe5GSndiq3ySnUJkByGIGR5SNB59nhh7kK7Jm49GHRwboJV9hphirbh
kAQwbltjt/EhbH7+tyR8+iiXksNp0fon7tySbmGT7BhvGe+pH/6fqQjuS2dK3mGpIJ/dLpU0erTF
grIiM9QK4U3d5sAkQWNxv1puXXpiqtbH2Y105WuTROjTr4/3ks3gqNvMVaJwsbulc6QDbivtonAk
/uOnT9HQXfFDLVoJqKJGh1fKTWNTOp99QBGcFy9Q4DmXRg/Aj5Vglf8jCiMxN/u1JrpxxOLUI/GR
BWzZmTm9+bmg0SPoCQa78LhpSRO+iGWRF9/PA7aOmP6tth7rt8d7lCvS08Z1+TxdZ762WONOQ/Na
VcjcPRv8tup6hJ8cWjk32uvzfKeCX/4dhv+h3ZCZKLP1GgWwruWwB2/lnrQt+jwciPaAjTK6WuGD
r81e0auIaXv2lzfalUyBq7yXmbSa26q2MGczKdEDcEp0dSNOnWrJP/TLXVD2r2teQTAyaWxwBdxf
Pf74ZcT9GOvo13hQR3UPrYGMKjxdcjp6gXNU9GFEqIB6dalVizRtNZ//PDQPsNFhPY0oOyHUPuSO
Dlf2H7R5UlLC/EOffvWBkfTCMTRh0LWA5ac52Xd+IhG5iCQHsqY+YJmXTW8rdHHRZ3wcIhMP5M7E
A1XQzeZ+C9UgNXTj1yHVtR/jdhaPV9/K8T91wvWne04boN8w1rFYgGVsq856upP3AYPjeizyybYj
pWVNhFXR9xlfkvXlOISqh2ZGk/9xc3H54M+yopQKcHaSdsHNOYTIxfgJib/rgDsEPOZxLfNyVZ41
iwISkAT3nG/hjGlxEmJu1sqnzfCOOx4iXftNdS3qMRDWRIJceI6jmMOvpV8P0w7BCb60FKCo1QCR
AkaxegZuTduKyYx/i9DDpJf0GhtLP5MHLBlHYFJeshHXl8Y5vRkax2H0RG+UuEWmxNsnqVilQE1z
NF9prju84Cz/udddkUlPtkGAmb8LdYh2vKJ3xGEf/KAg9X9YSITzyGnwUhwD+N27dl2HMAZsXYpx
/m3PlhI0rwpcu002U1jt0kjpp2mjNDvqFCaEtcdSE9Cq3imT5CTge1mBKd84s6MYW2hX5l0UurX/
4CuEhuNXtekhXsdPsLu5YAklqtVONSVL43aBsuso33hSZnyZGHMzRPOgwQO4DrR62bsEp43S9pNV
p0PdY+gewfOosfsNmjRZk4Ff1nuO6JnLtyb60zuq7crEqjLknai8ApieJ3gsp2bzg1cQcHnnIzmj
ymv8rXwFrqGA4RYaj8vdCLGKjY+ry9mOVpvg6F5XP0boy03oNlQEAi0UZYS5Cx04j1pDmOoP1FZ5
qptv/gbcoviRwrMqjD1zXmR0CVHp5E1uoKOnTKb9Jf7uGhJmi/K3S6ykm05zG9DgJ4EGo/jazXtf
3UoZBMrSCt8h/uBuguaI5YmRMfhDHf2xixojdiENsppi3j/JdGIV6ftv9lWwoAAstnMwZhk/Ywxl
UaEel1IkhOyrd8Qklo5JlLFgOA6Wr0lYKy8B7v5WjsbLJBTcH1hyTfKl1yljPEwpy6kdFsjkjbib
J7DPQYtdAbwTXdeKnJqlko4L9DJ1dbXIw4KBHVx7DeDtQRSQBpvDhJNs67Kg1S74XY/Eud/f6YHr
Dyrb13XuPA1rZK4S2jcYVSFpZE/E5o9mmgR87HLCtMibHDD/dVIhXnJA4gwJZL4EfgY+T33hHUre
Y/ziOUK2rzorMCu+4la++ZtYzjrqZYG6gew3Bb2tUM4Y6t0x38L4A4wppy2zI9sQaI+4H5nzkTrA
RWtENnjBOeGgC2PMtDEI/YpKNZiYWteE3JjpS2FjDTWIa5ep++3y/MuQB1QM/u9z2iZsesQxYyC8
ioIItveJd+R9bTSBS0bf5gedCAziSXjZGzr7DIKXiP6kfruz0LCaNf/2b7w2vZltVaUkxPmno/yw
WcgAwZ8WsY2DxBn1JJb0tlWuVj+yv4/xv5V+VOvpaNV106fRKCStXLpg9jNCkJSu8A2HdwU43k0J
DHx4TVEEZKoyyJ/tdoQI9zYhUx0ZGIinh1cMJbq/LRSwy+xxJyCVCT/xg4wsJOIw1Vo9ZzDvIn/e
uIVLXCpQGunmeisXl/VVaKxCM3YC4ZLRvUdG3ogpcO7OCtdwKP/BARbcwdbeNuTFwS6/whb/c2xW
JAUc2TSi0hctzHfVhLJvN5psFYHwM5CDCbqGzu2a4mOgs6rB8l6anOEnHmd9oDgPjiHuW1poHddG
ttYKT/4hRd9eWGA1UFyZiJ3ByNbjVYez6QE1uFpB7i3id1fBfJOJkbJsBAAPBCnLfDl9aWWpELZP
sbevpm6JuAf2AFbdscnYXqb2OQcrEn3tqW7a3C+eyGPoUrbUSvbqjCvQ1LivpQlPeZJdrrnfejXv
GK8ZSC3iZr5NZvZWVN+F+roBSxyeZLejAVcZyh638a8RJSevb3uBJamHNkAERxvLUZo724NKm99e
RNL1DV9Wk9ayPymYFvAO4hya3DLJLPOKqDffzzCIrnwuIzCx1jmjl9HAXfqOe5W17Ck/KJiKIbUm
tTzHaigmlNR44ErZl1ZT1Trup1d+gwmz6drTTt3Ykj543tKQUvnkFNNbgl7f5ftQafK7weYiR+Dd
nUWb9ehADTaWjD2rGx4gmuug/37xeyjrFDEMlnDBVJpw/Qt3HQK4KT7jffhexFuaJ0LjiQo3HdT4
0fN2b0t18jFcQoMeg7Q2tKpOywmeg0oPXGsAn0parigN6OrZYnFP2G73FkzuY+qP68AdiVFIv5oF
0DRYr+8cWrLxhWDgMDxsFz7QFnlH3kr299LyBvtFAYzAWSLnapHSiF7nkxW1QKywmPEuYSIwRQWK
EZ7aXM+3HdQAEo+peZ+Ue5RD29rqvjakxz4A02lmrYqcxzbqFXHLOHXmww6lI+un0MvxRjZpcQgF
RypmIRlW6ZXIhY6w/cqbMels0gOiPdLKbHwNCoBT+c+ZWuglLAwuf0jg573cHgJUebkpf8n1R0Mb
siKL7YO4IqNQLo3SFIUE5oUDwBG2MTpGFoJqZjRwlXEimHUa85z6GlBmenTWBwKecFk/xG2Jv8o4
Q013dzrXRywDSpqYLPRwkjJ6ZRcoc8SCE3wsEOPYW0DC4twMz8Ru9oVeaGf+Cben+HAmEWTBg3b6
Xo8rzaAKeM9fFfQrw8SJ8XDXGHj9vVJBp3OzIUF0ptm66/ONnfZv/ZYCqaB5LJMvAcSmecjC05YI
9xNhDi5rZY8+WXX/Jhi89ddmlWOGWlggh7QXthIUBVa25yFJ+WkKK7mbsC5M9bUIe3HjCz46r/EH
DHxwWNmCnf0xDHQ+e3V+IB6dBWGC127UjRC4S7iV3G3LLnjniu3cz+PZnED8/P7xdcbYQ6+PHFfg
GN8ohGUPGjN/4PF6g4jQar5tnukrhFshkBmLetmpeItrEGOtTKJKgs8ktQKeWIXZCxeHNhU9MEZF
uU6pePx95ZtoXd0k0EK9ySp39VRv/PC1Oo/XF8juGIgaQiCmbb29WycH1zrAyzKSKpqJ4YQ4G+m2
8DmX6G7fAprHDtkUw7CRl8jiJ/yuWz69/NltjPnqhyHAd74YTL8BnNL4P8EKwQnNwr8qoGLYzL8W
G+uknqbS8Mve0BPKlcKZVqhCGBF2KY2HyElORWItxS/jEUSEphjXUrNYCgyA2dMteImoLEpsL/ni
XhdrgwYtLwr9dhpIkIcoGxzVTxMIvmtmpHdC0aZUqkgB2UBdVBS6X9MXHB3XhLtZRurMpAdWah9N
lZzBjJgSlPUYAJGZ+EE+8ckkUkuDusXgcGdvutysBACZKx/IHaJplkfCVPZVLkCu0jpatyDKSYuv
MzBRiNs5J4Tz9Ix8UGhJUC8mRcIsmljIh6OY0gFkuprJ9jnO0uwYHtgLuUWkEj7BPl8+pgHeQqwm
+wq96bs0onGUW7pwFX0WIONqB8e3IuolDCVHS6zJf5Qe7X0n52DapffuDQc0G9okz/FHS07Yj1he
NE9AACNVXBJ1jRqSlwRGJ/fPP9mUVKykjI7GdbacMFpEjYiSZJa/ZsK7JrEiT92xKX/09JSBTTDL
TfpcTRPJTW9p6/QbpMq2gFQYQww8JGLC+ytfqNDNn7Fw+6z6IkFkf1QxVfBA5xQ5LVVwR2H5hk8W
gCgfk9Kw7KQP/f2wlS3nPBVGB2qJpv+2XSp9OslJliggwjvKSJm4ekVd9T1JntsecxF5TCychVY2
JzRnzca3rcB8iWsiPZE6+X5W3JaeOSCmjtnF7wYsVl/NYge/0z4aqnkKaALqz516WdprEVENnpct
2NbEdFgkN1B94tXz6KL0RjT3/d1fDmMjSRuzLYiKxnk1yIfkL8idio+4rvVEdu8v2rEQbByJlBIo
uHJIfGqPkE8qKRlkFxFOs2pcTqHNOaoomD5W2wBJg84gzzmr115vm5DOqVxNJ2JsdWpQuba/dPju
zCKyS7WuCKbUhDZFe2aE81Ue5K4eTlhvRq85/id3zCdW2Vyk/EVbMiw+Pk+ZDZd56L+wqqT1ViRq
YEXxGRGsXcGQ9RaZ7OTr+by66hu0uAqra23ZoZjm6xqW0p8fWG/KSt3qrVJzZE1l8B0P3FzrXX+N
V7O8JkscI7zsWEx/MVxa2fOI+vnnJn1UdX2ZcEf9fCJfS8YDYDBmaStiPBe4b2RlOQKq9wRxNA98
vluqAZVPuv8JhmoC3cghezL6RGThZJSp3C0uFLE8vxeQTufejW9Pv9Ub9zJAlqIxTptYHZbRN6Qi
jC8EuM9+zV1xXH30lpOBVy0exccN5Hp56TrHI72d/12FzeSaDvtzH1yXek6UisdLcpebjme0HZFe
46w+74MyXJB6y58Pya0qyVrayV6+XO3ObmrwpSE0vpMGothvROJ34WTrZvULAFiExwzPFNjj8afe
lAt7mQY8b0eqK/pxqWLu9U6gGlUh061/bxqO7ijbMPMQ5h4LDonQuG2qRXAqcV15y2lhdBIk8Vk/
ySZ/kN8OpWbUBE5H/Go/MpVBEP3fsoQuSVVI86TpA2JhpqCYsjFFgsoUa3OjIcfzqrIloGC7butV
wvLxBqY6j7BfM/HL3NAxCMqV/6Az4KyyfxNwQkgCkMTcElyZtgxaTga5rqxgkHXp1Puxg3wqjsBa
vA0ri3LdfJvG6ssp2QqPQ6+xg7kdXHC7d7KXTa2P7Id6whKDouDqIVDTQe+0HAtuRMTg6h69J19s
P0hrwnUFhgRxgVoFJpyewzgEduYN4ipSEo7IdbIzefdK/j2PZir9wKXIKV0ln4N9Zu+gcisMIIbx
bFCjsA3cYAUdcywJcY+2zYUBtbw4+uvo8sUKfsUhsPIU5W7tQkHlhBqtOyTVzJkaYPO4fA6Elcfr
2/8IzyrnnkC8Sy1CHl9wQIx0bld5X7j3Nyw3cAa/W7UO9q2muI4zkqYGytjW4DlZ23vuUBhsB9D0
5Cy3jSOOPb4zrhTg2ZvcgSXN1gW2OR/yyS8BTRAJ08+hr2rSwB6SvZK0k09iLSNpPKCkP6kUZuaH
P+v+E/zs/QGYB6OyJQ9ZiLtqpt7gX8/euwJSrf+w/nheZkam/rWcfZS4NQujaoLH/T+LIoW1XrrR
dYwLQOUWs/qZDJsfKIdCBd0A6jXllCUKdGVqKWvkUwPYI7QLuY7Z/IkLFYd4SFcM9byY0LZK564I
3bHW/F96mx1n6ojXdqmnOKZWFTjXTZi+qAGiKo7wtImmZfSvlsa94ENjPb4bpvaGt/qJ3gs81yLZ
L1yJ08XkA4GYCamJ17YeZs6EeRkEY/vEez9E758s/KjxL0MS43SgWpZ4t8zm/uhi8ggmPvb6gV5z
PoVhMjQGt9CfW/uDkw4WAfgIv+EdXlqnr8mKAgQ0LveKeqcm0lCFXdeyOJQ4a+U5L1MS3/U1IQTG
yv5nGlRuvupHJRr13+GgAkYawmlz66cgXFtbGfA/zWyR6ZaKt+JoL78QUlmOCYsPJLk6FYVthwDb
qehg8FrKcjwTBuhJ6e/9siWO5Ygis5YmIq453/cWWHBtz8f+FiGdkRIMxD41zdAyivRV7FDK7ExE
KSfWPWY/ixsAlBXJ0yBqfCcsGFCyp2JYEmHuNi7Ax0h3rlO7G7PkhxcXnhIdepdVJpA1T/9udiwR
LkWGvmHf457vxnweTY1Xf6h3+fVSRskDJ44h3DObDayuNjIqMAAh9C8O44d9f3tFqW57+WNjDNPy
JJgYacwzBeZi2I+kroNsvpdHiry0eTqq2OayAVKu8hBtV3KwXjDAhNHnf5GdupFs35Mufd/Ypshf
3McT1G72Go7gMmlVvQqeW4hUAeO9XIQu2UyA2lDZcEscNmisNAFTXqoeBc0+lD2t6TWCyBOiVTqs
neppvTi+Qogbg+r4xuobUodGzEJgkYWjz0bwA+8PyW8GcdDCR79hVGqmOZVa0ZFXDnoU37NqaFEW
6IZLEIzjROvDYVr7YrtXAlWNz338nbh0zVTVOWGZnbO67qxe4aorcg29fCnKTTi+z1rqI+tn7eu6
SX/cL7MoNOof2gqNOEBxA9D06MNxtdj/NCdcSmZilvaapD/ooEYXMpQXTiXRLlwK3QFmw4Fi0gmR
G1uduFI4ztCWo1rwgFiWqh8nG/U5WIPGy3MnQhikookENXzPICevBw6tnxzqDzH7GP8lH9BNXrcc
eT+vHSDUa0yxm83e/oCTQ7qVHFNiHLjyM/TeCWPL3GuqCZHBb+pRD/FDmGOt9XzFnzQkf6iXH7ip
l+md6mqKm+sldVP55OpiKCYnriAa8ssPkRjn4xinE27kjKN5nw5JnXq6/7Dn5+4v+7LSQBtZ8mFk
slfPNqWC1H4oWJJPgM4PRYiJwwI+7LfghL2FMV9jF/KSVvgdYpcUEnAoiL7gz1BTGaf+AhMZLvcR
aP2omRqtp1dCVvIKYpPH7/2sKWqcJQ0rs3Cn6hEfmuSUidMxna8TOU8tUSkhha5W4WVJeJmT+bXF
AdrwJYMzGH2gzdg2ikDHj87QYliWYzJUirdRJLHdPIWUbEArOmZIvV+HTdPmV9gRYOQAltQqAiYS
nBrA294rDXf/4MbN8PtcaLHMNG02LmH55RUVlL95EyYhb0GgVeqGISnndG24NVaJasOAZh+Bgy6l
EwINFtMC2KOpb2uX98xP1QfBxxbAeHaZ97o9WWbe0vjFcke38aEnDfaxkU3al4OFKG2MuGl7DHlx
evnvUU71WVwhRgblh6pD2sijMFgGJnst7gw27rZyRuKyf8hYHqoQ/OgeZ6NmOCQj854BQSax675H
QUpmzWqhnDKliuXTBJSMW+3TUr16LkBKUVEhSsqEoz125ApVkwhDr54YuvGIjuIHSrX2M9CEsqyW
0z0Ik9sOIXDwFc+HEVwFHBJkzQ8FVwc8cD++8PpNWkV/E+4ayU8ri0Vo33MMdku4zFYPqQs1jXzB
Dxh4CzRZMQRBPUS4B96ZyrmQm1VUT4TNqscqJxyFfCmObN0EWVoehAQJ3VlfCS5Xs3q79PWZuZE0
JiTwpiJlSRWdpaSIv1zeMZ54q32FReWv31n54q9ojRtIK/4JNV8UiVbKZm/3/amBaYoPm9TZigIc
F4yZzTucDeWsfE1e2QSclAhBfRWS/XGGrDNB65MO4sE8nr3/vrQvr09zxR0b3igB/Ch86XSHjdtq
cd1ZpYRNfQaCZJPGZ7yOKKZLFeDUY6UPIaKkCnuAkdQErs2mZFkY3b9QHieCNXl/aFkTgwa2NkdC
u5dHMpqNKSZFxd4PQ7rsp3Cw3rCbuex8emniaHG0n1cyvR5WqcnOcFqtOpv6TtMjoQxBBwJ23+AL
B8jihqU8cA91pO9JucXb0d51bsKwXbzkwkPZRUhZRuSVVuPZD4aUh+/kFOquon7D4Vp0gaRPFAh8
GKO31M74ft/r+Po08eD7OMref9uJcvqRRoRuzl4ice0g1+EMjhOcMEcnU890i41PJdVSDFH7gXKP
U38LqSeF2JNz2y6xPu8XACqbsa5ha2FgSiRI4bGG7jgk1arwksMTd90FE59QhfrfXQPaRxq/S2FE
d4JAYlMem5LZjKBPQFnouEBspvGb16GrBS4ykbCKRavMTf3ahcFQ5APvfOl+aQ6QPYusKIQ63pqL
Dx/3zsgU9LER2serQpw/UpyVSKbKPMKYieaLXWbSXpR186ybAxe2VBLz3YvlW1MlEFr9Pe6rnJN6
D+tGprRT/gRusLdRsS8iIjuxzbX2AG0MnJn+TsOVm/2P+9yhkixb6tehO77s+dI9mnMwP9UMI0Js
T7koodv53tllB1b+IdGeFjjXaAKFV2/7YdfvmecKmCyVntG5ph5u7bSIIki8V1qlLwtNN51WXogl
qisAzTzhuieRPb6BcO1uSjnKAbr9FhhAYYC3Vn+6G3mr/43tU0Bk/2n5VHmlSzYXW8v46qhBWBQ5
RJ23X4xw/aqBsrsnUmTfxb3wpH8mvDW/EJVYOcKdTCqYu4+H+VBslngDR3Q8HspcrcYfxPVUiWIq
6UicRPFueSsnBztonISHpX9Lx5FcF3bWZhdVW8eYUm+LUcSpEXTjngykaEvux1J+E1XYuxK1fuKj
SM8rtFDMJvMOymRYQH7z5+9nff0tyBE5a/fQmyNhkCsuiSzCWN12axOtHyg5VhQRbrBvjdrgmy0d
X7MOyMLPvC2sYk+LzgZ3oCrQivhEPbziOtBrVko7+2By11wnseBWX9IPbX0CDtP6pYe/KGA9+MCJ
FzEkGcawpzMvgwbsHV2uTaxltZqvUdA0k5bc45kfGweHL3ttwdiqWCJvw9UeAaKmDp6qV8cejMwz
7eEPGTxgQdxWLbpndi7shvVW1WSk8jDHJ6u9+JxXlyVkt2ZpOvGERhCrz4i3Uk40bg0BVPDLOCDU
cdafVuROK7C19Ljrea5NWvO0z+n0eEYEmUOe2w51QWtPsErhficInBk00ouUqBFThHdl+nTy1CDX
2650yCl2yDwypUed81vZDaZoJxKcAvMkjJ5RyT57PiZdAZ2AIspPg5vZ4bsHOYiCjYTHydC12DW8
jLLGvkmaBDRiOHhjFuDouQDosalxzWqdgfHRAJDBVNGU/2QpJp4FNnkDMnWQkSavqCTK3sWaDTHb
RCt+MhPzn2bBj8FA2XXfHVmJx1q/iwypt0gDIWEMyAi8m3tAOhlKEmSZEecXz2hIE34+Okq1ODZW
WWtAVJFBrFzg1aCDGI7a8mk7BZf60Gkp9FK3xDVqtw3GnbzYLIYQ+wyz0J4b6f1u0EVMbXvqBlT9
XH0LO5Wm05DkFjvfEcRKZw6sPbOznRtzLbmMN8Z8ZdRMjo+DgaWrVcsCo/Q0oxq2pgy/c2t2D64z
/STJ6KboUFlBwVDdNjukEJl6OcrYGU5Op518kMMK1ElWSyadkXwWU+JCMqBU4aCLkJQzvNWXBF89
gP8o3ldf9akMzELsXRmdYEPz1z5DeAQ3JU5XGi1p5EZsvS/jSIP+ThaHBOJMWkc/xgwNsia9lIbb
zzvZsorlrA5MY/d127fsA1myBCGo4o9qpdOEEniqcexMRz1ZRP6dRQfKgIO5oFUZAIBh7cRfGoxq
ee/pq64HG7jbF4Cr2HT/g+Cu7yuTOleMOBuED9NnAbqVD55LqYv6uYwKBMudg+c4bGz24LFehzMV
kqTwkCH3zhrfKGm42+vfVMO2q3v7bSBkRIP7cIF3Ve6k+I0WseAuMGaw8JDINKYs+CyoWHEyeNCi
402MEoegNuUPEO1VLo+PmWJSQF1byrFFoApQPdlVFFW3Pdm0UNaAJFeBKl4xH6LdrvhBIKtVtwwm
QzXdxx2/ff/f9MjNS0RwYHGkZQJYmfGfwdUT3+DhraI8K+NYDHr0DR+7y8AEmYjmnwA1os6O1Znv
KEArQRiPzZu97JLQO2epQ1GTrzdr9a0LIPb0Mn5RV4NnrKSMq4XQoUU7K0YaxauEltLTZrLqQApE
oM8NwCdcuBiTvJjfBVkwgZnJry0FF5qZ71yl202DszJxpV1sWRO38jPqOqDhxarJ9n+BxoXE+7k7
+kj0GXGQ9Pgu2x4F0weJKHXYIJl3bGONu9OZCj/edSkeapC3TroYT3djwxlh05I5vZyCvzbJXxUr
y4ZVphk+vryLT4FA/DTT4GqXEue3dY9+Kcrxs7TWuGu0Ifkorz/af6rPrymnPFhkpuzgYpWsQO7A
B6lkT0xPpKCiyodUe8XKM/Iw7SOlOhnckA6Fpm5hYOorbHLKU2PBrfBaqAKWQbx2vlJJlo5W3NSJ
Va0Ftfh9qINCominBwSW+tUOlVKYnEArPtW90kHCXxBMkBflkGo2CZkyINDKYxVuwhn4m//L4e5V
1dQE9RwIypyhgkAazPkmS4AW4sWYUPYxF0y7MvSlpndZLEjZhhuOKTWSmD1K3x+u+70IATD9Fx9K
imluDV8tNjn7SjIW9xJsxznwYRzAwiGBYBay1UvZglPUSq/h/ikPnWadQTie1/HPlny2t6vwhADL
ZV9/hNR2S87FS0KMY+bHe7gLwLVoR0WaCXm/lVjOxmsJ5JD1ST7BpJRgAxIQUfwY1lBUX010IUhi
XMxeF0lHu6zdFP9HiXO5jTUyUEuXqqzpIG6CIJh58lopDz9XIF0ymlHXdgVEoo6ZRVN+QBgJk9qY
oODqCtLurJbuoZub+vFsr5wyoQn/G3EhABz6YuP1udZePASVgrbY2G/p06Jvem0YHXyzD65adr8G
amRlQdLwngNI1emr1x4ykrycnzZl6g6MIGoDSoZcc3CZphvrLVk4nHa7SKxe4jF4GpD0nEhk0ZgL
IWF2KqRSZnpzpyD310+9kXS/PzdzgaDt4YYAG9rQVE+5kyPMqFWKosIp9sd2M4d9rj2So+EKKmgW
Tjk8nTRdJgM5SdeRh7mQbxuexCDyYeWjrW3QdMx8l39DI5fd9732c/7jvxA5cJOXL6ejM+2FWU8n
o3SgjbK0ytf2ZpgWQTWytUx6GRCZLhpgOw24cdYam5jdN5SDkukkmVSUbRUKbzzjthP/s/sxucBT
vkVnAOya3f/uV4UusG9hErX8/oujBnJsfZ4u7C+r55hWnYydOvwLTdgvyMmqwA4VY+bq3ToJp4O6
oJf6SBWO+Dqa9rq4B2F8R7epet4MKh7xBXCnM68VxMSAyWk6Sybcza9bAkFtIBNRDd2d7umEo3Hx
fw2XZjhP7u4OwFAWoo/lJYnSA2QUZolFRH8j4xdStt9SPGxt/rz18Rp6ZJD9n33rV53dDhuSmnct
7aYlSyjtU/eZHwzyVZ7oSBJjyU2pQV13/rege4+1+NGRoosh8AmVPIGyhuA+ztIytKOpnK4YD4Em
xjPlbAG+qqQJZ+ODYaqMhM3DXOGABcbD7/5Q/dmepfnhjFIw36MjATPxvVGrjyteGmocV93JCKJC
Hy2q07gvJbdLt7VQPNzYToGMFlrbpAMrfoKgP+2mmlounl1wslRiPgZ3bjsgJr94LCkUQgfLkxmj
AueG8WXpMx5OiYoeG3+vUGNifr5hAFppWwJr3wXNbJWK5d1KzLScqdoS+TKTovDB/OiMcCXONc/d
zaC4t7Fnx4bNgFlWwq+1fpqdpXHDqpIigC7TYH7S7rY3Xl6Jbil9gatduzoQYC5GeX5mGAqZnmwr
TiAH1rtb3qbeR9xKYj7h1iQd5E0IoCKPaozp5dx38dsIOhfnWWOjIG1UCu1S1gBu1/VXk/8pgr03
E5p+c/zAY+Ce1X+J35PRyEoNl1lWzhpt5i+bToI1BLnhhOzGkYGQHTp3/TtybtLBAIPkD04cPnnd
dKBaWUdfqdmZa0HqwZpeFVBqEjxKxrUk6RdRsAMmaHulhAJExPyMWK01L7sc1iTrPBzNd2UvrEQ/
O+5JqHs5POloG39qN9c2/UqGA7AgeSZJTUtSxcDBzxlzZyKkx5azffiy75RHWNfqOIEgQvbf6FBF
IMq08mIEcNHPZCOnuuJeN2MAr4ay2Yji5ozlDWQ7X48Qxj4z3lxq0hMGw0wdZ5P8ae13cmD9SaAL
8v6UEPSLnxSDgS9E6hH9hZ6crU986gW1sSv4lzMAe7g56GDSwVT5owEo7ARduvvRttikIsPsq4FD
AZl7OBoUhBXpEnxnTU5vWJUiMelrC831vguKSwfVH1T8fHpXXKxLBA8X/NTBtXb9kBIKczUmf5ts
2aFoOtpp0pGZRDo9QHV7ZUcHbpqQ3QxAgpdec767igStSNvLm+JgqfL4hmqZraqrXxG6d/vs09pS
Qu5Zw7p8Ats4p6YCGkOVxx6HceKJdzCoML/jSmiZkMDNO6nirQYFWEg53+6IfRhuNs6c2uunn7iZ
1SEk5brkB3Ugo265/10pFTQ7QKMiBhG3ktsvFCCObalD9ZSVZK+ZCfoVUxfkAnQObNIqB2lfiodn
TfHENvUcISyJBnN1MwfWrmAAs+7yRCbuQvdDh48leONrNu+AsryOAgA1a+UfvmecwnsqJ22qm6jh
qzLGnUTNEGIXCgCwjHK+DHINi9CEG46jWWpcjD2lsgFf1qKdMavhUHTr8GV7p9f78jtZ2rJlnMDv
BBr6/7tqI1FJ4/DGyYA/hu7ZpG6wCbb9s+B4abrNwcj1Fhc6vEI9ReVATtpB1mNOy3xg7Vt7LFCL
f0oH/g3Xh4Cy3U6kV+uDwxLuXaS1oVqumk+V0yEw2ksb4vogl5bvChuMInYAGmb9wE0HAZ4Xbxd9
mo4unOMHqSvDYSiIPOvEACt+pMOTr9p9UNdjGCZ1pCZapVcCpEri93Jiji+QfNH8jFjmAKfgos+Q
tFLOe4M7eThOkdnrUvr6iojZXGQ62vVlzNkXacMwx9K1E2u0Onhw/y9fRfvbBdVQy7zLmqHpB66u
YzecSrQVbW9kPJSWp240H+7TBCXPc2q/76OKyWbRSWRT1Iw9Qb/lqZcpqYWxZvT5jP/sazntUTFA
ZQYy9qfRoK44Hwr/u1CGtQAVST0OBYtXc4fuDq1E/L3QhV/2ZStG3kbolyjjCDcSekDAcQHcHiPf
due1bnoLApmAEMs6JrwG+g6qHQOI/m7hgceeOojXzORVfJ7jA8bcwFiKhIbbieRD+7cbX4vEfvUN
ocLAVLvgRNHLq9n3d2yeZ/EipPrtcILn2Na7zvwmZY12MbXUzodZRxnzIsW6M2WiiXkcBvgI7gpE
douOGbfcZqxrGNS/VR6hjNu7PV4ouCP0x3YJn5O1+zz8TOEhkXc8XLxs4vFPFOX4cWBrU8wU4WHq
GByUSKE6KCnmVhbhBXqTmuNVf43SMhHXYl55F+wlrM+EyeBwatLPITHshj3ujE3X0kksTFyn6WC9
lCD1Eno2odrbt3kKr3EbXoBFiSWlQPqrNX+nnR+9R8pueR4YWWwdmZr1rUjkMI5isgWrl7MVEuPM
wvZIEKYgfK3TKULbW9+GfLLKL2V8KD6bd2+NGgo/Vq4eBECNVpYNvNJr8ty116ZkhTagXAfV5wPl
otYfHHflgtLah84VEeikjFYZzSSMziGQabIykSSebKzHgjC5qCJRaPogCu3fiVNZxbrPAOea0HpP
QRkLdYmcCyOjpfzGoTnTVOyattudY8nFS1468BDfZCnhHDE8V8FCEKvFxHXRHlXq2SL4P+BZkzx3
aZzFNOvonHFplDP/NRVYazHiZU0wSHtbxr9WlKwJhSLzQmpBp4Jz+qC5McnRTe9+AyPlSlfLCSdb
RsjezZWxiQpEfWz70MSEmCN1VZ4OH60fUocPnpROF/JqjULbz9zUwoVpWmY+bNJhlyYivHUKUZ7+
pOpvdcoNm9h+/NYF+pq98UI+1tpugRUGZAh6ki6G7aEmoKc0qJ1zWok3jRP7wpFbKiNiVTlwiv9l
iH4zBvviedXh24UaGVAcWUHpZXa1OVKsZXOErHpUfHL3fCyukCdAAZ+eNdFWbXuoZJODTnSF/8Wr
ypTN0Ib7cVtz3JTLwDzd881MHn1jxtbzHLSmn1iW7UW1C24JB1fufOLUMQxb8FPcBNKPH28hgXxB
jo5hhMebOQmIGvc/fcopq5SnuBAd3FYZdM2FL52kLKHCWs+S5fz8ATqmC/aBFHhCjMbHB3zQ7n3H
LsQ4Ox272qDrMX9AnnHpI/cni6C/V4S0NzgKBbQ/Uhnm694LOfG+OBFTXQupsCe7hAzH5Xd4CfAG
yovVLTp/OjhX8Z4UbGecyb8d2MxDTRUyZDNnW/O0JckJhoLTpj/576xlNVbRiEPz4/UNJQTORmCa
KOKfGG4bx4ZyA1LcaRN7KyzphG1z7wV3VhH5ECH7TLcPRLiZtxrH02aNOP7zlHAMyY2u3dDEAL0g
nMyNNY9pxyLhfVicwKznYLoBm6qDKOY3OYOhFYCtaEEdiuOnFJzPjgSQmqAJ+xPkcytLYW/KEWvV
1KJzwqrb5lf6i9b6EbZIDUENoztfmmeBR4Ngdx6S95PqNtGSnT+qKo5XHLhODLboUljfE2T12EPS
VbaViHQ7Wi0hKN9O8tOAyNGQD8/h4pqWPoqmyNVM4oFbr054jVyZf0SNfqJ9Zv25y6vpo4jjNjTQ
Jzd71OvYqv+VwA1RdA00qWyYOxt2MjCLrU+obEUJw83FgX6mCEEtAh4F76NYC4hKMUO2TOw1SwIa
NfUsxav5xUu3zKJq5M8C13LaEQZzJfiI84uMVmlWVrJxmGnK5XtBYCmlIu4bHr9kJAbh+6w3gB0u
YhE8p8/FLCo+FSLbyBdkYUVzuQsvQ1RJ27Lqcj7pWoIDfrao5MQEwGgNXfCjIJRbzJeAtPAUznkT
QXEn5qw1HIs2/R75fK+mtabwIUYyM/sg3IJRy+EMLlEx9vDUmOgR/1Vx8hXHQJ4LlK2PAB2csAx1
vsUOfFiOt6M/jbCF55krg4bg4xReL3Zk28FOJ8z+D11e1KT20/rLhsd1cXuFudQDARTIcXWhhpG2
VIyFgNJLRheImQqoz+y311qml1jNIPDutK8qlVc8RIYmOflXtSeZSEOC0tlQJp+s/gGfxUDCNF7z
v/7Dk5sg41KdPIYmjJ0zzpn337wGvjw4vknaqJKSmvKUuVS9tgaqsv+lWq5tgznYDsLi5kWU9Xql
I4jFeJ7EB6Tf/D1YfV8FXa+6Rtc1kCugUAuVsjFL1fb44JBMqLh7KLNuq6ifi0IDyws5fADp0TyO
cK0pyaM49lNgpDT24dUauA3VYteHiNV0eg620bFYhCCEz3bMhFaQDHX6uRdwqOOKnEfeFFktZA43
OxXJ387LgnJqgWQ6OSi6ntnFzI/NkGVDdtCee4H2dchCuGazJHYr+w37ZUUWtLcDpnornt8jf0J4
NE4dsd5Kqg4eGCB5bjc/3XpsDezJgTllshq1nv9qnpbNYsaARQH6agUH2OLpf5UF53vWGbtqVSzE
mT7V7J0rHj6c2dZGRSSUPmPfCCnO0Xmc9bUWQs9iYor9es/TG4nQGR9Y/dV77+OnwvDxCNfosn6Z
P8e4XdJfT6Z3cHN/JAqd5H9vq5yxTO/mtafVIOP2Ntov1ZXlELb9YoSu+0xrxzRLebI3O1JCCOMy
bcR9TYe2gTd5MyQlhPGgxcbtU0IMTqTshNA/phQ1iwCj6EqroSR2TKhiuk83WVlLoZxfGIr1/7BN
9vMClUov1DEx4VXTcNzuefIqq3W8D5AFUOk6ljt9Mgkvq5tT/Do5Sdn+OUfTX1yz/rBNc4IcqrMn
9w8zSfpG3mkFmmaT1BhRvpkodzGGDkkvlTRocLU6+rEYzr7joLCoDfNxyacbzt5qUwKytpagGuT0
WYbsJT8Kc3cJyhu+EeqW2T2UkeSg9FMEzz4IhTj/Wg94u8veXp9W1/R8qbcez53kT7OJFkCaqAMI
X19gx3+NKbEO7JCmcjL5uiagZAcn7Kcgv/HNR2S1x6OEIsL7An/feYTtXrswOir9gCdui9ff9kDS
p1kSBU//ORlE5RHjfLf18TwJv5h1VQvcYh2UZwzgZtMPb7NU+Oyc+4jPgH2VP4zKp6MjRhyBGpWp
Kfl9nEN7eVIJIXZ3syTPXVT7Oa3JKL+1QRzLv/oXheT7JnVzJyA9S3EwDCcLsu/E6alS8Jnc7VVd
pz20tl6xj98Y6yaKQ64amJs26u1EH0Eccq5EbMTwvDKUveT3wVBTXWdSWgx0FWgQCBnnlC5FQ++A
2kCrG0eadP5ygFIwTRkarUJmAo4aYVw4s6pQC2YXZ6siKk5y8Pb+lvsMfYiRn5gP0jMuYUT1TVyv
I7U5ZzwiCzhIZ7pCPBGs1sJjphAc9thjixF6XnDLdlx7tX6G/UDURxrlL3U1Ep0oJss8+kD7yKCs
Yb26F1KwW+JFaxFf53YNzGiCmp3exzKDkPN21/rLWD4LwjGAW2uOSluv1WDPatF10Ih3WGUSRUPx
MKK2QjmHWkkGP6pc6xeliHG22UKPCGfmxhkxThyehItrDMsZqLNMR17nnjRntr/WUtTmvpKGuZlN
zq9IewX7qcmK5W+HkgqEDoFPTQSnTPWo1Cna03yaMSTht17LnOwkf4xyXPRnPPibwgVKGT8ibCd5
aUB6GtOheoRjfc3ke/MXuE0sb4/G5XNXvVyk5x+JkQ1veBRHJzcYPOntl39eVW4hFTecUWGjDxIC
Ifd94SBxgtHf951Q/iALJ5acXHyUGWLbF2aUDxaHNcfcanurxVHtqJcWMzrVnjCgDhNuywxg5O+d
8NfksHP6dKQ/yTpRXqqy+ISgCogvfSKlKdy/1d18mF8Hty+p3n8JIIcRz6JU4HpOSQUUHoE6lrVV
Zg+6QxpWb2Y1/vSUPyKK84FBt+2rWlNQaVdZwiV6c5z07WxYWWBodwuaYi9K1lVqH4c8WMxZ5HWx
Va9UC6gv53XhGE+p/mOyNEf+qZCaU6tVwk2dppI2hsnqnJF2JeO81+M1drJlwyRHVBRw05ZlYIfS
UL/v8yDlpqW2RwchrMl7BQb8xx+qbFUE8zoMbrRz+8oebHh4YAaLeT5dpeY/uJJ1g9AkpqoUOio1
zctNpAlLeSRJ0vKX0pKFSNjo4aqMuMPAM+SQQLgzSqzb2/J4CbI2KEmdp7tU6HVa3pWzyx2N/C38
V90S0qmIrorS3P0i63LdTf0Mw7ZljOeeGsGcJ+3+vZK2JdiXomUvl/1O0eC2lN90WcCeQYyphkik
G//L1DgQtYsulFIJ5Q4Sc+tto1bBYcH28duFIGKGekxjMFbBh61Ubir9JA50HPOVjeYvPdTTxOIh
Dm08rTwbT6J2kRj5iWzLGLfz/GjXtQLr+cnzcDICZCNTbeMu05vWihd66/R2HDxhSWrQ7PUuUzER
dvKh7g0hhnAgIDa1njuQa8Qq3KfY2bavso9NwYXSpFt0szbIrqKATALp9v9ewgiZPPsc7mrYdgL9
ouVvhJm78O51Vu6DCJSdb010+0FltEs9HAOzA3zJMcg8OOW3n1gyrFC7JU4QFePxhi4QSZIcRCE5
I3PyvpKb6K9WTt8g1Ixkpc2TAvnxkUVcD/m3yywT7UbDfuJApKiE/fz22zz3AQlnYC2XECwZZuJi
+DaA8s1QZUX3HP0sY1GxgZFHjXDyD6Cne2mfngN0IXaVJo7oP635Bt0Hv446tCVDvyIsLcVrNKcA
XDkcALS/ZLAuCf4/r8P5Dqm9gvNPjajlg5Gp02wOLAMl92qSkckv22na1omcRim6NJDuP6WEDUvZ
FoHv3HD8ftMAT5faOSKYOiMLJKRdaxRj/h2BMQOlgtjMvUOnI8WjxLYdiUjpjHOwSBX7gJ97AWV2
1LuUeZKlRmknjlJ7C2OHYsqu4Z1qh+9DGjj0d8rJ2qQj5VBwAp/v/t4CfLEGJw+Xnxeh7nVsm6Fs
iFqt9S4r+ArDxGZS6li5NeuoPfmvpAnBz+BanN2Vo4ZqJJnlc/irKz6mriCsYyldBrggv5bpuZE5
ivNKE30Q6o2/F9jn5DSKiwMZ5qSrEkXbJiVF1nwf08HyOkfx2AKRkm7rx+gQIgH+loWJKxhPSJIZ
Tu6uLuL7bbD7oqvPXA/k/1w31JnmXt8n4rGbOfHR5AWekmFZfPazQa8jsB/md9/OXngOtl+VkWmA
5PNBpTMyFieG/HBlhtmK1Vq4gipY3bvLXSjXibergBNTNOfYDfUaFyAQk9tmaIrq51ghFwB0Cc8f
HbopGxNXvRv9cic/DLT6byaCccDWuPLwO6Jk59tVZt2u+ateJuW/YatN/hWgASsyzvdrdg0p/gzl
z/am9IIxYXQFkGQLSNRq3a8noJo3WDzS6gMxjX5JrY+hD+W2nzSNpvNBe//ublEBINPH+w77U+8/
2hE7q71EqbVvdgRbTY4sawnvnGy84vSTQ24XA9cvq+s3nPwdXTzxvIHDxbKgkyuQG5egicUYS4KY
OQeP1sVXWnp1frpr/krDMmgngVCSKByUSm3vIfnUw3f5XvuVfEi7wsq60KEMsg4pako+feGjT6CK
RS9ZLJySsGDlgzjjna+ERi66GmrwEibM6hdWgOOcrgTwV8Y1JvrEWCHRIpxbdDgNZdsf5mWzCh/6
IM2jsLW9t3sl18PiORZyVW8IsakOWhh4X3fceJvaIVGBF8iSPn3daB+MLRehchtFj4d+C+qvaKP3
2K7xOk21AGOpH+zZW2G2ousB1J0xBxF/BMRCwfkmxKp2avN8SspG1PRv5QkYOAEIbFUOfWRn34Sf
4tOz2bGv2ZkeXHgYde8ww6eMpaAyqbQxjOi41jnfEFzda4zDqfaot2kramnHwdsMriwpO0yjpgEW
3ckAYVJKUgrWuNpXcLwxx8Wt5ZNrFjyIHAt0DgXoV8g+ZgpjlYDj+V2s6o8AqvDZYgW4kkolPxSr
Q7/MdhVwZLqgfkQM93vfmdTs7F29gz8GH3bCp63c1bhn4MORkGtrtsmnPpYlyY2kOZGct9F/cfv1
qvDR1AVUYa+PpQTWH4mmrmwswM/CPKBjrEgHFSMjnHiLIR7B3yANpLKXjz+quiQMgpPNbt5FcUzx
wHOwM2da1zEZuBdBU75JLNnnj9cdI9T+ZZjT76sUoFVXh9b6XIqzFSRv1kmRbmIfqB865f62rC8a
y3yJo0UK5YVwcREVgmrQGqY9VPhsLMo+dJptPvfaHSMBlT8YUYrom/YeUiv+bm6KBkPR7AOeMZC3
OzhhVits0g/Z1y4OpbG/86AeWHO+iU0F9lAUC+dku9k0TbAkfFlsIxJ7zgIwNH/E11JKDl6n+vU3
42MsG8HMl5Vt5whNOrbbglGyttEKiATVKRaUo37pzi4o3CduoM92ifzthcKkTtYHU1QmtlUePdTs
MX6rhEq//rhTKViyXX+860kd+yCi2lBhtVKSuf0PiAR0XhQYt3BsgEkp7DUSb0qscqxskNnu794B
DfTXSO0MBm+bVAiDJ7NkHeZx1C67opLs67PZ2T0aJ0l4Gyyr6AEh7W3+LJCiZb24kSvL7hr8LHZS
9Sh6KebZYVW4Sxql35c3l8iBaPUm/UzzEe6AATM0elLZkm/UDIuawzUEk4T5t7fCbEJjc4VxdD7Q
TJwjsKBO4BCKKTYIpV8ewI0GkHSkclUhWS4/bExVluZldneT+bJqHFAtg5RgHRLtXQyLb1S+4GYF
mnWl17uWU2uDqTFipz6aU8vlK2QBX7Q2lzYpkAnm6QipO2/WRJR/YXUaCYUdHlZ7v9YEM5IjUNfl
UaapJU5N1mlHkuKNn+IOfW0URkpomM/riLx4cAXw1CLub2RPpNTJWz+Jl6cZRkODov/ENpZv5mv5
ChuP4V9q6KvyX6wMusfeSlLHYdWRPNhbnEwfUZuAXUKT1oUYE7Z4InGSW5sgAiuIHBmV0FUdfsCg
lwohRp8b2I5I3glcoNKZoPXRr47WXbQCof7re8m7YhYNFiDh0sLyYCZOV5/mTepv3YM2KIc/8A0N
30OefZql6TlN14MgH74NCJmw17JIvtANiFGbpiYapVjfYGcL2nfk0dnCQWBDO4S55Zp3X/gqD5hN
ZtXewiN/qEQdlRaT/0ZAhWwtlZGqzHXJ/9LDuh5Rcsxa3yX8zedtx79CAekFrFn5l2auumAVuhXb
oXDfUx3dPqDYnxUjjGT97lQk3zR6iYS26ugj2NcBQw6g9UgzoEjg/sLXtU5CTAhgw8DTmUCelu4b
0vrnIGOmRJmoDCn1imVnDfbJ/2m2bELmj/G6kpaxeYHvRiBioZ6U6mXrmwNJEqXQNUkb0t5+Gk9d
bld0DcN0khQtFwGt2ruX1f1ggXN2ODS39j41JA1RQHf+piUOQX3yaAKqFxsfLpV8j5038LWiKwUb
PIKUMgIlLtrpzhtBFslVKd40nh2oPrL/zZY/6Usydnm7/Dh8AVfhnsQSxJHy+yap5AVxUcMdq6vO
I/QVlKGLeqAoeGrTyVu7NT5zW86rH633ynNl2A5DLJJva4C0RyOA5Q59fdDFVomh6K2WtjdbKkvK
EzfqRrZT2MX+BnailEZ4NJbII4VCe394WLh0Y8pdFBmpvvfrcSL1cRB6pKo5Thh9oS8FIjweU0VO
hLYvD5MlpDIqXkFtJ8JJEW+VWd4II5U+7tfNEnVJXI5cNtN1pgZnCJc8lpzs23HqNFoxpk2xiz4o
A5IB+rkE3Aioey06L9inW09x7zrluTAbcrz5LYyPgVQ4HcTcXlg+r85Pl+8JYk5+qWfnvkmpL17U
8588GhHwwGJiF6MqahfN1y9iLz71gjym5lwLj0Z8fDSu+aLj6zNMh6E3UKfOzVfUD0HKeJnrG6nD
TbNHToRrTjp272ZPLlWUdrRfX3XsyL/D6souRVm/o/WXLVuWInE+n0Hisu+L0YnfjclGLplr7BS+
CQ/vCKcvAsdP5tz8cwQwyrwvgWuJw3vgnAPmnBiUC6zpHADZZYyl1pOdaHSOq51uL/RduU0QlFo8
TyGZuN41CEmm2lNvebhyk6b8CwkQu7bVmwP/t9l13ZhTvlkBWS7IiMiA4wzijdyp1Vizymr1+Tba
5d6dNngNN+XDH98TUWi9pQdJDgXvdEoaT3Fq2yAGBNVD0vLVflXPBKB1JvteQDl4UccONNHY8Nbo
sDwnS42jozsxXOO4zCTB5/7tUI4cCbjuNndowbjnhJbwpV3dQJ9V59Z5J3UG1qHoS16Gm4PBlT+K
wVSLwEACa70ZRbVso70XDmZdSN9jTifUAzjLzKtqScxAtp4utsmWLRVp+4Kxt4RMX4EE1O0QMwcL
zp2bp4rdSM8UEXUI6XVd6ZBe8dMFTrjIA1DIMHb0bL8r9VAxdzypqOeprOZ9PiRd1RJbcIjgnX6Z
7suWnNk6lJLCG0hsg0fzRPiUiDfMixcUMYxfjoywTf/Vy+ihYDOKIiiT+lqnOelpC0p17m6KXxXV
ndS0V/bkihav7xceq78TmC6HB2p0GNqk1FdiPKWZFhONew3Gzsq/6c4kMkqUnns3uv1FEV3+iwYC
ljHSkQMqJyAQxbKNPg7+jpfMvf2JIyP8DwAa4HOBrheAXE7yj79kPhUVRCqHWnFCbi+gm/mUer10
ua03cqTmhM4Y+VKV0jUm234w6OfasHGrRlHQksqwB+aweMbAPwDMPmd7XIA943G4ZtUU1osQsSiY
rQOAjZCy/xnzLpskJkgzjKA8jPCk1SuQUN/ZeaMZSNZ/YiR87zuR4oj/J4TPoj3cyo3V3t6iomfk
U4KWTSdCNhf+HubusfM7OPK+mnD5n7LV781TGidkVjDA2RsZr8eNtEnBNMYgZmkHjqOgHb7jYAU0
2PF8KLFJj3onDHF6eaTvkTDjTY/aGxy1rwZzE7RlVIMOk0KQ3rFgHgfp1iXfpxu3+zXr8C+n8wci
dz8g64EzwHofckjpmJHZPpRMitLQug/OaO1w7yVEVoYb6erW67X/Y0XDwg1UfuPWYS9WI7lRXtla
lympkQkYHgZyXqJ7n36h0RPbzpGOkK9FaAX93Sw964jhOCcr/twNVvKKa7kFozZbejD9nuRiC8rx
x67oknfs6QOMrVjjg+24cBAILeSthRx+GIm4WnWOKz+GSUF0EFHez5AjaPAZxLsW+83zsgB3tRc1
1zW8swOa9oDJ0Fxkor5qhNTT4n3DitfUSprPTNdvuVUhg5RizGY3Iiwl5NwXXrwHY+icF2Kr1lxf
4ExQc81udsI2IXb/8wVh5iRwJ8+ZB7gJxF+f4cN9KhMIAQhyjy4UOtiNm307otJ6d3+fEWO3Drz2
Epb204EcGh0363xqVoGmIY7+uWJTKdrYAEsxxoxtsdnEOZgLPNCfvmDIIEwbAQxuPz5cYYaoIg2O
S4Rh6fYQa2lK4I7gNpS3gLSY+nuWBQyO8dGoL2bvAnffcED+KNCNn9kZsUloCwNYU19hoBXRuO6i
8TNREB4CErO8c1yIVbEj6jxg/G9cYruafUV513Vr2z7W26/31W7QHoavnhMaDze0EswxQkMf6WfI
KUgxokvT0Mcos7hTbc94LI8xol5GfhiHRFo9bTkqAnvn4p0yu1elHTd2Pmn1uPAjSpu6lPngDExN
ZryNHYTN+vmY/UGTVQLgpdrJbGBtblt3BMBQvh09fPQqYbfTeFs823fwgwrMbmJN/EyNi9NxGhtC
iy5nj4w+IDt56hh+PpxZOCuS6ADGCVIC4TH6MIFAO26iYCI90meXM8I1APChe8yc6H6iMeyJ29t9
sJUZKJbXQkqNskifJH4UL96ulhUox/cYHI6GXNQzjkKyz0Yvvzx2qSonaupAZd9yorHmeCwHyuFw
Zc4ex8yqOnlMQCb71Xlz1OOjQ070q1vnb5qOqYPCP+yjBpMJqq8Q0ot4BmEpPbGzosQoqri9iFGZ
evpjZTY5J8z+z0d+K8Rppzun5Kz/rE6y84zWctaxbmkIh2IAXmLZDU8RD/fccAuD8lvIi9dNc36T
etV2hFBsqWuwAI4/cAEGt7yIGUz55qLRD5Bbs+rBC3sgLS59jcaNVbJGEoreBj6cczZVbn+ku0i7
5cbZOeKRWvu4M5vvNUK59wQnTzGd4qrjgJh719XJ6dUXOaEWDJkIP1J+VCPQM9T66yZrjyAHNKpy
nXaIYYHayIw82yZMhN3M0ySIS3CpHdkTlKpQ49VgPpJTQomtox26k/4kxkTu2yJjU/h5mqcKZGYm
iX857no6IhMYUFCkPYjrzzjOYlE0aS1x+m6pX4Ta9sPBXv0vjMAxcP5T/NgUYtWrVjqQqr+ua+XZ
KMZwCn3kQR0sSpo7d2eUUcSTEZJ4efv4nmEeLJiK9by3XWdaNTJst5hdXrHDlSQGLAof9J2qTB1e
ajmXv+njj2i7cVjm/qrQOhL1ON5NQiJAhQ/sR+7Z4f31OhxGC4sIKGk0iJvoTn4+OsUpTsQTnuJn
bvG8bOI2n2o79jHS3Cn8yQeCJmJcm22PQuas64WeRE1JsCDVJN1Co5eIsWuNsKq6d493/7Gjm/nd
CXu3wadNJ7xEn6lds1P2FcBePzCh6LW2YhW87LXpqrDfTbOqxSp+GQISQaasJ/5CHSFIOQL40Q4E
OG3cvxoOxo+UH9WlkIKN7S5HT6SDJKCAj5KgTOHHUD5kH7Q0a6kUy+vL4UyJPetmUGeYvs+4n7lg
+HttrOvoe+pVz1c6wlSp3Nh8wE9zLBeSIvmbOfZ9TZ0L5NZWcWqnLmt8Q/JqeZDcvUi/QNMXAr38
GKtRq3jmAicE8BWAeZ6cW/XoFDjHM3eMKow/VCQ3byD+u3xN4udqd3DhaKcXxMf6PHZ1CndRJaax
E5oGXkwP4yfGjY3pV5ruDQQkw67CbRAic7msjeIsRRwKBphilUevZI6nE96xk0L60MckB93sBO5H
3GRNk0PDk3orVDw5Aww3a9VIz6pLDkR02Blfk343QG0+08DwT1ci+QrenUBz3e1svBUYP6RboPDL
n7p5riW9KzlQOraq++RBEY/K0wFBE+WCR8v8hSbY779XbmaNH1cRSTV3ZyXQ2mrXABeQgeHvCGgn
PRMD7W3kjmC5bR2KtOt7Uv5o3BcYGQutkmmviD1W+3V/lEZ0PsBOWPnUnwD4e3gSF8fWiwvaVOCv
MUYDAKChyI1CxR+/IltVHCZN5gFlrWhynVmxhZvAymXPLa5T/V67G6VA5foUF23vkn9AMuqWlwiS
NKabzPvxaZZyhf2II7HTCCwZM3IiYmMf/sb08EC7Y5kxKY3Hw6VOxJrzal2KpmloNLjlMTNtDLa0
mMQ8e5ZritEB7YHls5kBqbpsXEmSHQF4WxZf68mykGikvXqq/K2hgKjg4PNsP1nOj7/FLxpxj1bI
Z8s0rFBLmo4Wi8Asei8ggqmuyOY9aVTsgsmTMkyWSnC1D0l5UHitgSxwn06Q9XuLA19H2tCxDcgP
5i1jngORV9MrF2Y+6xNaPJm/NmtZMls7S8H8AoVrhBNGkuArzsLUJCMRbWwCqfT333eR1o/RoFbm
8LodIzQb5/Zfn5iqSlA9MEOmSeJg44nDs1c45M/xiGM5au5hfIuYLTpuAROG0guSozuF47Rm1YJr
Mu4w8kxGdBUG5xJfeyoqo5wksXH+wPtT0gsQ+9xLbbvCQ5I+9aA3CxXDvz00K9tTMtqbXk5WODRZ
7niJT/Teeb/wvmWXQY8WF+mC3VwY1qMqhtcVRTOGFo/yxI6FlRMF/i2Gcc+/rK45oSfBa3sDYNXH
Jp2C5v6SrjoPjLFoVpHtgoN3uh+Sp4P5H3jNaAga8uipgwXdCScs3YiK7T9V3MMN6jIE1hdnfkUb
SahCyQ3UCOzYlAjZxf04W5UKtxLLi1GRirpzg/5urbrop2quN9Cdi597R2Pt0QN1/NzeIZ1ymAz3
KhIVLN8jAEyE/rRJx6dEBhNcMZ0GHlR4slnP93Ygb+4BtkVfGeYGcLCTSeLiIQH+1dV/w3D+wyIW
hPbGRD9AZfvvAINP14Tvr5ru7kn6IluSaLr0Z4IcUGexTFZogCI9BXA1TLwKTLeRMnxEvAsJNyAx
V5p6QqPNqCoYKHp5euNnBdvnZnZQ16TsOf32k8XRhvRlowx6Rg7mTBuGwdeuzdBX5eUzDDVWSLiY
VOPGxv3hxtdGHNdL5LCgzJ7d4FilJS2XnWo81rktqendzr4nhxOkHHmqlx60L+1vvSZcVzf7jD7Y
UgTy6SObIvW/PcN8xVZSqyXvM9uGKQcKENFe/KQWABH7Sld0fDOVa19ik2QX1CEmSM4JHUjMqvSc
zjWB5QbJg9nViK7q3VNoS1tDCV9iUStxF3TusOkGZbhJwJSQ+gugGU4NNPzYDH8o2haILgMcw6FI
DoGoBSbThu6KcVTbOk5AyTDjx0ZTfrUS9y00cU9j/mLOgtKzzpEFC4nMxKUuxeZnunLNTC5jM+/b
vNJ3gKVTWitB02alaYYgPneoqHPTeLGGYp9v7NYbAA2pxVZtr7b8b7yro4NGuMiw5h8j58fTXXLi
dGpUWHMo8o5+wb6UOlAM88ww4N54A9DEHEJl8TU0/DrpkBS9zOSJJ/oayX050Ji8V9rrrplHglTT
3inZUBr7vfIppJFzlkM5AUeVR0LZM97TsooBYojT2Yg/VYTAX8pbYcno5GHwuz485051kKL0zp6z
UzBqaDntk+8ucGrqcgQ1+AKVC5IzMErgWcXqdT4xuTeJ7lGC8bGKjvpmh9HI0rZNF/lJ1hOXJI7p
1M9VqYw8W0GpBsSPqRL6o6tAM98jBSYdq+p3PdY+cTNPLkHp15x+U3o9sTwVrFmEVcJAdESVEyqv
zItHL2AtTs3F3Rzxubwj6LNgIRCiAcXcBlncPzOtg30hjVvov0aq/sAWcSF5sqZvvE8TX2fuXszD
g5MlGcwNEHPH6X90WnjHubVdf0lguDAvRqCnayLjGAbX9ccS91DwSuC8I9j6aBCm3bEJFENu/3S7
nJEPDGR3t8a4uqf3/GVTQmCMxlqJZz/FCT4UFdAhGl55j2UvDwYgnwLR1MBAofTKcc1vWxKLDF6J
kWZDIIbBeGTbLN8XHV3YRceLQRguIUGTgETptCAaW+zbw3ZFJnYfBxvyXcCJl5MHHpINFBeGSAC5
bPu6k+aqaxtNDmLBpqX7jqpXFufHRxnzW9cRt+D+wlFzhVJda6iqKINlY2fRgq4QvW2Nsnu9uxwC
ChQ9JX3YCb7piABIKCBTULOJt3t+bCHy6K9v9XtD59QSGivP7o/3mOnAxEALYqT+RAog46zC1JY8
ulyH67vAXdJplNhUotSMBWu1rECMywx+a0m0OT/GHfeVJCOFeSzECOSqh5co/nPm472iPN/j84D0
Thn4w/TqlOyfOSFV5x0jUPx0MhjZ8QxK5H4Sr1Dn1VsVuLFx14PykdHghKAV8W50SKsKQrMI/xlu
sm9J7DGj7tyYPUn8UqWThAMfSbPD1Yb4hRydSqKANxPzPhXl3RYVA+T56pay4HEeKxTA6L5TRgKv
s3g3vCGlnwNGyY+wFk7+7gmF81Vr3LIMU+X21vc1X4WKlxk/bPz8+S2ZKULzu07YpSyi4ZwqVChK
CJKQRQ8cYyJNwrpi377HuWwZFD4GSjO125+LJKhRy0AF+qsDIeCsZYflfecQB6wE3sEC8BmFQtJ7
YA5q4C2442ZsvtNkjInkz9josSg32r0M1v5fR8g7huuG777PaYbJTyPFDClxPyFUHmqIXVMdWMMZ
BaAxWUQPz6u2Ytj0Cf36p6WRncm7rGXd5i7zHtERAgkIX2fWoJpCOdd8+h7CqPg/WlGlDbDB7k72
qcjvFpG51Z0tpZEtDB0yB+FQVvQglxjanpVLxMrmSKHGxjjOixbG71Qd5YBqr57RaszeBc/7vZoZ
Q+rDK5CRKp+wElti5qL+HswLzq5pN64N2+n8+xqd/e2yBDReyLev9J98S/HrpEvK8jF1aziFq0dC
fanPpzTHmZ657qDvJk4oRWWwFFEeASdRY+EtYgMozkol5dH/qmYWa4Y19zO6WN6lVzL4qg5vhEvu
n3grOA16k4Kqazmh3IMySrU6H1H4jOQLYl49hNmbodYHj2Ta7QNhC0U4KL9SoMQL9CpwfGXQgf3w
3l824/oPXmxW1iV2WrL2XaF77Sdr6MmGRHrF0xAD78JldqvV2o+2D869dD20zMihblbaL4dU2jew
Ix69hHTUioi3pxiDICdsSgA6EpTXjh+pzpVVzenJUbQqXFeCDyjS8TfJIQWvmOaDguL6vA1HUxlW
w6JE88/1Ate2YCgJIAG0Je0or0Pd3REVx87EMe3NkqQYIDru3DJLH01y24isYXp0RscJ3pvZhHem
Z/RB57kjuaD5PCYXWfi3j+FgAZmwKu3vO5HFAOyRWmBvCCDsDPyKn04iUWzqgyvyRTijigQDZIvb
ezH13NnENpU3t/96EAvNyXQDvvShpevV5wiOyQLr9/R8gj1YV7Dh2N1aO6XfuYK3qithW21mv8rL
sdSinDCxY35VeF7yihq/hbdFhQWHSqovHlz3lrBLGSd0ce3f68fTgSE6a56OqspGcfdVVoUHWQ95
IVxXj/EuHyeFHIgmjIAOaK+vstEaMAd8dGaOFQSq8LAZ0/kk9xZex+bWvdsLJJarkjlG2dhkNYAy
b1wuZS+joytB4HEu66GFZ1nH4xXQ6TvvdrA9a8pgVF2xcXTX9LdntS8n1KIyoHYxu32EqXNtkFoG
UMckyJRiwuaHD4XhtSSVQS32Ie7L/w7x0P1Pge1MXda0mjVrDvNu1az6USA2N/3LFPT80vg6ZR9L
8ify4RzIcYVVV4FXZOQwzKQHSKpMvizDqwfridmyCBzhpk6j0MFtQUEBjwmMoT5/D+hY7jypR9cp
6JoKKBa/qnBtDSyDbZiO254MOLWyhG8kKn7sYSVmOVzX7LkYhDmqrrJf2xoy8m0njSs0UikAECjf
YWIHgvdE+ud9aNIwXYEd7ddlQCxSMypmbMuTDe+hz0PWzLPEoHJtqKvrIZL9fNo7z8bKCwKLkude
MbLizPRP4uErg6Gs+Jp2PoAXPBLXllg6efpdBbHANOsj14nQw/1mew2WawBt574XrFFR/ADeJ8gV
SCPYGLxj4RIuzQhU43qWaFN/wyoJKvK3p1KX6J7ljqD8R6hA+PND4Uw410VJAKfOWf9DN4w9fthj
uwHGrFVPs4cbN9elMF6SXITBbHnXT+6xXQNJEJF1s1bVU2yjdiNb5ZWMbWg4j/xRoDzPqLY6dWjd
oCkHiM4UkaTVvT+vaw4yAs7j6HDzcFD4/vqmTXANf+JTxTKUAHTqBnLxRvHaSn1KQpHOUIdp4JxV
urCUBHBCMFiCTGaf+CEhTb3wfc5tfgE+p4BFMspCR6UPORgnezV0TVBQuZcZb/sYr/sKMzqcz3G0
b0Ehb48Zn5XSgub6VaFnREtnVN63xISBrBRVsQAIGYHtQ75AxnhacV9QvGR4aGXsD8DrdBOnXQ4C
k0dq1uIojqZrdaiWaNAfkAzDJ4igfaiF6Qr7FjAgf7qOgan4LguJqSyGomordU1yrsGuPpnI8y7o
yKIFOji9N3bAmOBEdb9ASbqvTyb6wIKJmobg8cfEBBdSEL3cqwIu66pP2jFAEwvVkplO15tcJxLa
Q6qIMlU/VNnsiruHDuTHt5qojC/LcSzH52rLFGq1PBr7WyCMJK22fzcJzoI3paLZM5PrKFdN9efu
SxEdnC7J07TsAZtdtFcmXzsGQeGTxJCH1BDpvGCxCcej4+F4So6IDP2SlFPu5IwkoPZlCo2kv7Xj
3xH+8Gcnt3VE2Q4VqCp1BLEKpYgrcn/3AnFzKrcqf6ZPJc04o0Gs/sTGi+s0SXydrE+qduncn8I7
8Y7OPFsmBS0BBaxZcKwxYIhLG4hm9LT8Dsq1jhUgOIa1uNCNLXVZmIpw6Ur/DkdhJpuQX4rHjmmg
INR6m5FgpCzeETUPtPuC8fK1WUSZ35Jm8x6458Y48VQA/bYJ6Ps879mAlIkHg4XJhiSFoym1drP+
rK6hd0zGtYQ4dLhLgumtf6tQipzBLHuR/xrfwJDeyphKAR1og1srz1j4DrDpbKacSjI0w9qVELRL
YD5UxZa76KE01WEzeKLLffVBTF/Eu8FhYnZ1c5XBOvCqvKrznN9IQqCzQIiffsye9dciKQIpuHek
LzWpP9v/Ke/KBdm5AsUZDNG+wQ7x1FpnZuALwAREvffkSBaQd33LDh07ZMANwDfUQDGctG6zKQZV
bx6x+XgakbqLe7GI++1slvneUIfu4fEIEp+sMumIORt3e/CLxW7o1mSvvI/HMtt+0ZBBsG49cEE+
KaAIRnNJkVpN+ZR3n6qnUgoCr4NlO2hHt5f8JPZauLi6vCXgc19UKu90mlAdm7fNA2UP50wt3Ba4
cPbcLyq4HRssffjfZ1G05Vj1kg3TEoE1PdPJpcMNbL4ARYkTYYSRDvsU6sQK5jUK8uL7f7qCZ+xP
G5eGMudYp0g+66ugnhNUW5fNUdzzLdC4ijlx12nXDxzpelxI/S9JAVjNk03oKdIEP+sO4hZCSbyb
ijmvjH6I7pTtTTqL138ygLQKmcjfFgXj17+uCc7Tnr5c4tr4aM1R/lTZr+d6ENh5A21XCKiwvwdn
tjax99GXWj7/oJSMOrmeTSYZmKxIo8T5xdeiuujhmj8NNTk87mjd5/hc/sMwSmW3pKyL4TjfxLEp
f1kh9rqhTFwxRjqHBWEYNqOym7kEJS5go5JjQ688LiiJn2sqIQimog7lMpKPgyhGuS1IKvKhBuLT
YScC7heL9clHPfNOX+zMmIus0KpATRpNqLkvKFpQ89VKgPZU4MvpTi4Mahej+EaWMDGqEYpqS8mH
Q1D9EGHozZDI64GYppAqR+naS+LKaUOl6fi1ZutNSX1T5tCUPHrp+CQgmi5WGDg6rzJaA+vxXdQ6
fewhDaamFd8RhbanK8N1OFiBjpfXx8mcnPjkJE/zW5rlT7Ldb+i24pVMGkEUYIN2C+rtmxs/T0K7
9W0aFqNsr6gpJT6vb3PsEb/we2fouYx35UXieS87hrTNAz7/Wdun40qnV+CyMd7feeM2+lWJYwmT
QAYiEuSBxvR0IMivVKyi0M2UD6bPYA88ksiKsWfd8Ua0vIoaEQOv9qHz3ZP6a0bXfDCcYaFGuI7P
7zOUdWdYg4eRrzvEa1Z4h5ZNqFrJa+JT0bwLrYZFajKgiV1oNt8YvhlczkrSoqHKJn7Vk/vcU8QF
Ku2QjO5xDnHU8sRwQ89Schr31VZLycJ6M3f/fxypUZFBUaeCIHzZYZKAdnMzCx8u2e0xYDfQRh1Y
L+lfb8bPowv+xKObh2B5CXdqwhaLkjgtyr7Q3jUNUf9F4W1TvopJhc/ciazEpUsTsY8D2+g6w0Ms
KJ3ZcwPoTWOT4FbnHYNCXWmBVTCohqNmEBNIKDPIEIZsiUOQ0JzV/2xxzpqMPHP0trqYlctOwqw1
UlNLXJMAPTumLcc7gYgtSYDY4vmw0uiWMzb1ZMcvtdDOjwWQWtAGRFYTnY6oE3BwLwkZDJcDbHof
tknnOGFuWdoHdkaEMhn0hvPXiy0WGj/c8cvaWC7CFzxSQ8vpN1Yyk+cGgwjgXrIH3k1tUNUBas/y
xXKwiHgKqbgUGxxZ6Zdnnhhsmd2e4BHdYc3xX6oPFiyHQp3nEe4PZXiDBFHTp4ELEw6krKGaTHHf
NgXT6jED5Y7UBRifqBVaPr5Sb1v8CvIxPG0ppONed+3ichnAy5w9lw2W2VULmS0rqDZRv8B7X+9d
Jm5Ot4rx0o9XVjIt089/sCJYmYU0Lu1qhKE/oDVmSy5f/ohXhajycxklOoxJAOl+ruNmCL0xZDmD
w9CYxgaExB1ETDr214CNrG87FDZspkPPJUczNH/tw0NLqScbcvQDH6N9lkWdNfhQe78F9BExBSWS
usq1ni0zpxRIdwXvA86LXAF5tZ1yxjC3VD3uRXzjGhkuFGEcZLMSW8SgubRMeva70+hZ+e1dR7kg
XYTDa794FBWyJh8f+3m0T/DLUOUmsxs8xH7ZvlneCne+jLJPJqYbem06bPWT4C8+0kiAqbBmX7j/
XI3sNi4iDfrX59EsmGsGIQ3KPCeK2Cd2GULYuZxIT9NqCn7vVD00O6/zQiZJ9uZm3OXhKpvep/UG
lkr+s43z+DlTH1P9RB4+LnntVtB4aG5kTJfiUY4WV0epkoYzwLig44ctwJCCji6wmMm0yGXfAov1
GRJ0Tvqmz2Pc/LWWnwKy26XSvmqANyfl22fvdDFsvww/NNpDWQbKw6VZBTBMtemnN3k44Eh0MMhH
ICqCLa+iaAXcxI1JAMyqaEj1iIu4btpSqMz+D0tb9KbVx9JOPix5MiiW25Mx4KoizSZ3hZft9D8y
xZKNCE2IYNWJCfZQFZ/mRtxzHhYEoG8o8nX8IsPXryHzIEQP7+AWsb+i38KzZ3o0dgICiq9Io9zW
ZlT50CPv91mdW10F60s6S4lc6JmISZU9JmbFX8wsWTvvQVUl1orH93rRTwuz5obzlM1Xd22yEb8n
cfgBwB9T9hDaTRqEUsdHdKp6UXVASku7EuQVHYYqrMR0PM82aXW7PY2pFX80WrEPAeDw4KaFIe0c
kgCJ7ZmDAJ/+/aw8pvyLy8MDN6tbwXgvnBZGagaB7XxBb+EyXkZPALHJCKN6fJkrh0l66oGXJkMG
DLrtSyHI1Sz7D5Z1LeFicXECkDziLlY+W+cs0a6LwyldDp09EpJT/EemMFNYT3BKkzVnIG8ogZXO
hYXZM6WLpjP92Mu3aZQpRhT0ktCLS72nEfvuWOozWi2WYrZE9WwOF8MJlsim451yt7ZDsiPGw3jA
uFJG2ldlmPCDSQJph2a1lihmhig7YCjR833HWLqwRK34IsdpIHKYiVlN4wiV+4ctNSHjhdndK0tC
ataUUF4TI9NDU/O9cuSlLu2AcC/xuojOodu8t6LVgKwBVKIHe6nwDWlNWhZXmL/0Idcqiy4e9Xn4
JiiAeOnhF9OBrrQ34Fbd0Zlx0W1we58oamlTDETug1PGIJiDkpo+PcYS9yRl5AaCnuQW0kvoq/lg
JUKbgsKCcCsGW0FHUfUNBU6Xah59ghAznSIioi6lpFdicuqGw3GOFKX38mBP/6I1k1SbQXzJF2Pl
7OUlIJxj2GyDKTJt+j9I0z+MbVSzHVPA0FP0pdcegnJl+QWFhhOSZAHRErxZCaehn8NCCMynzS8/
ZrEym/GW/pGWLL5YSGJJrLeOgzupwfZyH8iv6C8twAo5OB75QW8YnrNIq22LKEHYB6h3w9k8LCRk
m/DjbUWDR1vwLXDiSr1wtaT1xop3F0NaghO7Gfe6swv/17NylNpxLfO9CuzHpsqogzToRT0GqBEX
+Tx/WL5GQYa2oCKDuQoUJMsYmmqPLznP09cJD0FW+UMZo6jT8UN2JI1zw1XlUHMgsybc3iseABfD
5EEVv74/ZyxL2xyeuzUJVNNeGN1UWvnjNS/L7LDaFja8RusQxtA6JSasEZZxlCuw8IaZSUmHjjsu
nGfvShRa2ju9bfVdPuoL1vuhHVPRbhFbzqxGdFiKiHLEb/gLOE0kGKoP2s4iFGo0g8MynETyToMv
TTYgL6VofPCBfqE+B6EdGNpklboR5rM2S4dHwR13VoKxVlPqQuYYWYfSbk96rUOHapSVMleQKdLQ
Hw8+RL6Tg8XUoylDxe76Lb8JgAWwss5v4Y6tbzuluytfIl28ixrfL6K7zIVTuWj80CBNbE6+/vjN
dTx1Fx8Ujc5dOn74UIBTRIsXkPmxIaye1ECNpZFgimVGBnYuAEYBqtHotbQ1pgIcD7l692F50GT4
lhzzhHbs1pSikYBG/QXfDEFmWqqmT/GBK8ge3o5jvh1kSLOedoKaaMO8909C4rDsWMaRP3vkNFdp
N2wp37bKflvy9m/JNdU2e496D5YhR94TupZzokFYBCI88F6QZlQkzxezaSzJ8AQN/BYTp1ZxD/9Z
QD0TwIeiA/w4MW7xgDOwxIxS9NvAhTx+Ny42hU/nAdELv44hdWKPdL6/FNLMs66USl3mbtW+F8BQ
ntRJvjRBOaWVJxhi0BMo9+csCm7EI/qflOihgfxotn8PMGaa8lM2C/n2YrBZiu+bY/iivAuTizBk
gCPa2/9N5HJq2W9bPv+Tf0/SIrFRK4LBzBQKZ9AeEHtwxVlYy03OPQSgWTlQfzeXkwIV84eG5B7A
EaGeQrUNNVNV6jyAlwyhulHebv+nKfXvu8B24slXU5kK6EmOLor81Q3bC+i3lIMuy9OtbpRH44PC
CjvRhKD33Na5yW0EA7jTziK6KsRzJkH0GilDCMGgDS2/kBE7go2KQnJdHzTpnYpJw0LgG2TmV/+G
0+ZYNbxFSYwatatyJL37T6uxepXKGpMmmZwTwR/RCJu0FOxBT1VVQSb1hjI90ID7zrmEbrntVlss
i69XGP2H9JhDOIwER+QWOJ2eM1Z4f2fZRfjaW83GZ22aCRdNXkbquerzoCSfZ5EK6XaTnck5Dkst
b+WUYM64vRcM00Te3HMF1nLjX6AtaG45lmdDtilsZnzJuGIXF9IR1e9FffPzS3jrRXt/mMiJUyH9
lzOG3NPnAtp/MGrr3uX2CsT+HEQYfiaGC1xf6S1Th154MLiQ111LDu5JvaPtqD1Xwk2h8TIXjVMb
WSqvPjsHBrxXcKlZHx4Flbp6VjoxVaLvYCVcA7CRs1kxiSfcODoeIHXnW55ixD3yFPFTwtjSnIc+
aKBwSk7HUzYllhtCahOSLvEGSN1GM0Trqh3FuTEF+T7e7Vq0xptLadjZERzMsXC+8murcwolpagX
+oiJhZIuu9z2UPpMEm+es40Xq2tjx8C2o5LSaApGnXdGAai/vNU24vgVV3mIixu/DPDJDvW66kMJ
2ta1UENT+mCSSt3A+19eDYDojAXrBxUJFbjDgH+plYTgE7nUp6SzHAa33bcDY3cGk029U5BKzODc
HFRDDQpg9LAMUp68paJQM5ftOs/JhTvTT9knnEImAZb9CAbnEMISHntZSzWcCdERw5iI6xxDMVnv
PfPKlpwQB9Q6SQGHOPFpNsKrQ7SieECTU2PGJZsXM+8Vt2rfAKQ1/mkCDx9S5vTJTVFpsjTMpCkv
v6dzN7dAOju9gAmgurC0GJTUBeG5a8/8CTtyT8BOQrRMnmVFiFYCPz5m2x8eyEWwKxDB+gXh049m
nP/CV0jJ64v1AKfGbRYKSSL+/FnphC0nFUvWspdbLHXsnWG5xJIBmSCuD/e8hF5R4pEu0s/0XFZn
W67jn4q+NoGeAkXmJ2vgVGlyM/4JJps0uPd8tdddHqBu/Jgfk13wuMEnVJZmR/9sBRYr4Zyowh1k
TXtg3YzI+0cqRmsWBuDdy5khKOSun7Cg69BlsxlKWpbMmorvD8L3J1aFMLI0DMEJGZ/g1elhJUMf
b98OD9CN4NMBi2yLLV0aQf8/4dEl8yzdRptwaw95x7EaCMtx698Z/bBnpUkYNlnPkiADhLC9BU06
MPSrBwDq+hZv6IXQJGan4so8icuLLibf1s72T1w/5LtGKH//sgk6No/qAsehHEQPbhvdlt01UqvV
a1W3FUXNPa87QXOmnVPyiGCEEHMjBIeNg4PoIOirN3wc09btHgOrWc13bMM4JlHhl75rGRn3G87b
BzvBjmdWyQg+ip4htc4Su2WNjd3CsHKLFUh6Xpvrq9fbssVMaVuALwGwh8CokCS0Lgxnvl9SLuJs
h13YZv5pJm6sCstyxi+u/g5NQRQJVY4jYY7H1gIEBgPR6pdI1ZH+NPOWLhU9XgbPSPOblZjYbg2j
F0oJHtuDvg1avNMj52EGf5NPKXZzepQ9QUgInavWq4qAsfo7GFGuGMlr1FWLc46FLILclztF5r2l
KezjY1qeCWHMucMtPT3sKe57vHLMsX/yjBDfdOeQQcOM31O3go7bgDEHDDabIDz5W2N1QRBKeQzt
VumWbrPwNffuQy7NqK8YisLeMI1JKV1lwhZVetnRSwB070YC47ISgYaDr8Q5p603x15OhOA7VNms
B4dx4Vw6ymbq5+I+/ttOqepjmWcRcgFixt7XTWE9cql9XqsjEI3HzJmRlWyjUrutOn6C8+Rp9a4Z
7ym2mHrktn+7ah2cU8/2EoFcP0c0AfCkaVMfAHwv6UtdogeNd7TF8frMphDXt7IFvMKW8rvBzeZp
OCzVe3C0q7poj/f5EUqg3ZE4TOU/T/n31nN+VVt4ke/91gZJOFPYwlXN1wkNYA0DvbweJ3g64MhD
CNjaeBJfszCT+CFHjh0lT4bBja6sJFHKuZfFyfbOlD/4luOC9+H5q/NUX5GFZ0n9tEecrXfxyVOY
16NMwEcA+EntNJOjCwmpwZv5RYX9A2REifPEtD0nuNjXg4hdwmHwcaasq/i1L6eb9kKScMt+Nfc6
KyVRY8QrhpNDNN0f++an2gq1pAQDiSUcHHoYLvIO+VL+gJPbf0h65J3s03DVdpzrKwJg7zr/H9Jj
46J1+sY79WYOgpyOA8gGAHrQ6EYpUdoIus+HHQW+3Gjop96GNywzzY3WfvuSR330WZs/vfJ2vUEF
w6gHua3Bra+ZJgGzcdJ2Y/nea1Bl9lKi9Bp6buXtHbyiR7JTR0fy6rhU9ALbFmJlCKPnUjTRihEV
Y7+rrxxmXihrc2RUDYYp5GmT9sLnBvJwHmpQM7FmzxvIvltPeZMIq1h+uquuhGE6iMRxSvgDcnhs
i9TI7UuVDESmyHzNt6a2ThJy08rOcDlx4cjWcLpeKzgEOLJ8g9y3ysz+wZoVj8GF/qjT9LLbzAn9
3T62kR9+k/TmaLUIZ87kidUgom/TrsQWY+5Ncn3l7/7BSo0/KxcZ5HFyrQnbHF6rDXBtuq1XXsId
zGsavio1Y+BFuQxARTSEzbQpjDCHG70VmVnH3VZOK+1SWr0jxdhMdBTt62P6FvPoR+WZVP5hmneX
ZevnBYcEgiRH743kLUgCNe2RNs5IqEPULoDpy74ukob+kBbT6Y2uq0mdZE0Oo5GMP93RNeZD2ITk
SkQaWwb+fj0K4HgrM/3b4rGSDQ9ETjY+zCkKPNtifVoOjfrJ23nQglm1ZVW20iJOEiTtQnov2b9Q
Jn7DeBTeP6M9jfNQf6JmbA9K0WqgGO/8woZotQXOdDvACgc1eAFOmNRfMPxLSW41WlF8of6BUWfa
TK8diSTK6yS+olNS6GRtuKmemDbL+RiQw+mB53Fto7Yn1VMTN/yHE1SOxtx/kAQv9mMIvhFF5CvM
l1nJmX4IBra2BVJx9wPOVPSeAEg/VHA3aybo7l5GvrPf0x2uwfRizHJEK4zigzM9mJI5U2r3WH+l
C/5D2jgYJDpSBLUdA94ir3ytmekka5sDXtJU1NwFc6UKKm8pRuZT1czTovct74nOJH9zgHCvkYW1
0RdbU5IgaBSyFmcGj6QT0LaIOeEWUt64WjBMDZQSXiv7sg2O9F2j55kIrer3dle+IZpxeGXC20AY
/CA8gz2ifLAJurWmFgz5Fvdh9TG7fSGjmRpRU2haLce/N7AVDSI+x04HohO7J2puFTtuSj6LeHXn
G58B/EPzJA9jcCR4ykFxcJVRJf171sh/w99NLx+midtehFQETCD29D7Bsjfiq4pjB809HS950Lo8
cexxzgE94hmZoZzCfom/sTxSGOhCz8Abz6vXiH0Xk/Yj5hS8Jyd9hrL6Xf4yuAB9lBWDKZjyBqfb
Vp0GwW3YR8eGfeFU9BtPkN3pI60IIfclSvZ1imiLC5ojeWGTEH6NAkzRAgahJLnA+GSXgq0Juy/B
TCU5y/SRYXLVTfPrzQf6GFqw7vW8eO85d3YVx94CygT/Eh8JKf6CI7co2mwsW2pqB5OZFklCN1u1
XiPxj3dFXMhSNBPjq9xvmDiji5I0OckB+YscinTZ+zUN+msGl6elEYokFIVxCypcmZ+11Shh2RJH
i9W75PMk3x8evrVvDvgnnihLScFKZf7hCahfsKffIGM/d6yK5CsLwMP1nVwyh4USj3VEvJHLDS6c
VrFYRTIIiiJsXOVhC2VPgiuTdsBKHU4TkBUdcIxw+Xinm/flqgIkPGnTySEyRgKePC+M4reDLU88
7TCqHiDcMwLyjzUVK8LenSX9t63k9rHhTLgN+iLaVp2wtEZkpBo+SYaKJ7SLQrXd9Klve0wUu93Y
EBic9zgxwgYH4WGFrXHI3ALqE/oVEC2i1qLCso+GwKedMjvaB/UZeyD1PPJmA9Gco4Okwy7zNJmZ
Ng3Sginv9mo40nrzZ3TuWHpcamnzOZTWOyB04UqIt70p4XzCOLO3JW1yIvQe27s9Bahz6ExSqEMw
sspR+eZ5A2O3hqVO3+TKKDkojW2FVYp9nIkLC8qQKC+dXX9K1KruBOqVHcb6WhkcpEUFwdnHHUqV
WIwqAwlpctqJqOXfrfEeBujPMWRj2LpLNNVBjwyYY2vznuqILX2CGbFzcWi6iYML0VSgu4GwQEGX
dHOEQJZN/rHGbQ6Fwrox0mnEZ/04Qdu6KBr1928QZqvWf2NczqiD96pHIsNGnDF8ID1yCXkuxnBK
Vv+B3mXh2K5YNreXrqnb1CASg4Mt3m3pthJvIukLR7DsQXYaMM2Z/o04PZZpWBnw/SOHNXmoSq3M
ihxqQchA1HUOvCHnyHComwyhXAj6+L6WIB5HdRvj9xQe09KPvgtx1PZefBrhwYDIFOY2vonrjKCX
Ota59yYDXUUt4c+mQgjzLjsH9JTg15XIEmVOtD/KBTmXWmMIawH1UWI+ggjnlqlvt/Upoh2SLTKI
3fhHinHeWawRTQ30YIno58sh2Dic9Gdo1GLO6LvlmcpHnnR9mxBgCPOTmx/DAka2yzuaD743pGBK
0Rz1+PYW3kj+maGwyv9L9qI7feavKce2+hsTzJGWv3NuzyUHpgq3iu+AwHyh3pSVTf35K3b0QgxW
Do1Ej+sGu4kLt4evoDWAfWjZzILf6DzfDPgcvHndu9uTOTryJNLeO/fHOSlaQ5VrPL/7eoAsbFOJ
Q4UK7apdrCAQxV1ygGlzkUx/xm7w6Oi72atJl+TpOzJyDkVrX2nt8vZmHafbWaTPDWYZ7bbeM9Hh
gZnbxO/EDZOc7BiguaFFfITM1yONwsK2ptCXVV8VIVBHlIMN6QRrpzCKRTQjVpUy+OF8NaEVdS1u
qvZBc8OFMu2P0MHNgWTMFbEGZ2jQkBkL9hSPdWdvaJMn+8W/eYWhdItCZiA/RKGPG2ICSCIl5wUs
ySpztJSx93h0g5mPUh4CtCEsgX9w7xQazgM+IQlTSoSzG+OF5nJCLaImPyMnBdJa4XWhDo47atcW
ZBqic7FQ7P78HGKq8h7jFovCUvCzVAx4Oq9JMDbr5X16Wt9/zpww1e7KUxujUvoKFg6NhsOcjNJ8
uHZlHqqi3r0MRi+O/9Zdy5qGYWb0ftccMt9l8AvE7/0IpcIys+4/yhxByxnlyz5LrCyzbPSSSFJJ
HOHEf0OpHcxGsQcH8QoJkyAdgI31JlLipfKKRKHp0oksHftdbz85yImCsDsD5AusC+ECniAcdbNH
Ert0hc7TM3pZOYZqCxbTKevcJeeiaW6eQT5XARjMicHrjIFdLdpGo7QhbkSNB5qe0j59vCLyEzMG
mHinHSMBXz8OIhYqy7gmgC8zRzFT2PJKYiZVqLa0OJk4MPhEEqCUd2O6LWPS9nEBGvrrXbpQqwuG
eKPJzc8mPg1Tqytoxx9wZTrdNrBSp8X6O5TkNI28SwYf26iDlpQQpQeKdUJNR2mhOlAW8+RCtq/R
ZtT5FGyVt7PC/p+WDPQka72Ote3LfMnEI/0jrJV3aBExCZ0MaiaQiGk+1BxA6IBqm/xdwdLNgQOy
YVB79OkxwOMqp3GwDxlEzok/G+gQxmLnXzlDUYtuMbCb0WyU5TMpkFUxhrsB1LnCtGcIC3W+GjQf
GhxARLRj4Lopb2WKXenb2DeokEGeaTGOmLIlsZjtDBU7OUVlCSXWp/rlAxRll172bELNelMN1Poa
2f24JH4HWdn+Lw664bPXQ5d3apbCRu8ER7/TOtsbVmkDu738bLvNPHAXSwG6JIHBrw3i+jeZsurg
ommPn9GGOXTEaYf/Jq4uYzh4/m5qJxXUvnhTyMH7r5lp91EWnghE4rSOpng+e1/IYS+T6e9aDyV2
DEKhyQEp9reb8Z5T53IsdToEVmcZkV+tqjepFkOMn1/x5H2Gz3O2+DSbtpmhtGyKt5XAKIg6jk/i
7Fy3ylzPAuf/nRMMAOr+QkOsC/EmTvNkIZ1wxzpeX++Z1854i9PvXnmz5YBLysQC2d3px1sicZgi
R30syju0oy+hwTcWFaO5B40wXA9fVSje1Bp+1EaaJRV5ZUYBcm5+B0paN2vOknMqGUS6as4Qxz8k
yW5iUzOSfLnNqfSBLrSrqyV3YnCQW2K/6pHDbtm93PcL2uKQhw9TIRRxAqTpAQmwdUwG2jxoW6oP
mirFc3Rl+sFXhZccdJ57CvtQqPYl7lMY0bFTEqRNlfSbAuwji6mw0oNWJEq7mpc99KBwVKcBaYNb
p8sJhy77rkv8yJGEZe9t3b7ggw9V2H4eD/ubeZ4p87fgQJYpdFuxBn9CqobtryCZ2CU6SgPMZS1n
kCzxkq7bPtpGWic5x5Ssc+tMEu4fWq9NPy5khuiPNSw2uYr7rCKPnPGbXi5tFp9Mmbv4neON/G7z
EavLe2aG/bCCfQYzYU7V31N7E80NlqlxOZNozJN0ak76PVrroVzfzegSL9gI6nRL/dJawMTdiJdm
rGMckM/Nks/feQyjbZiIoxX6511lj8xYewf9LmVpTUnjPTi0IjpPp+GNsyTTEJ3wMkiM7xYCoiss
7NRcPzIwAKM8vE2SRk3USXDe4878rLZpxNcAGwA/UoEBapn/AcDwy2fgE8sezDGXeH0RLQgo/mGa
kcS2ZD9Z9K6BXKegFCPHlwZQlrrpPm+J3nndzrN6ShYtewatNsChD9vkYKISlwPELb+uuxYgnX1K
smjzrxb7mUxr8uFuqgyv7hDWoOBCNIJHLwiM60D88NbJ2zZ36HAwNXwEcjKriTUAzXYBPfAhDkxe
RSNtBs/VTxsandfzM9u117ZIKB7EWvZakL0ilA5BWywp3PxPP841+gHwPTCiwiAc2F/eIEcnlfKG
0/VJaKQiWZXZjxZYtxGccIQKD1hnhLn0DrLNg8k0gJuqOpQWczqE8qWuRPyyULKI4ckWuioyMeMd
Dpk44Jc0xbEWMwfvPGY8ydFAZ4O+Q3Dr0qM+UlffiDY+cYzdi+v8x0PgAnH7M1NlxpynJMLf+Ba9
zQIVASACg+H+Wu0VWz59c0s8GlTSJ9PbWuje5lb+LJ9l50W6ZjZvb87HeTsrUTnpePPh93hpx74R
r3affg56u1KQ/bISJE6A8LRjmsiNFoxjmmkVZPWY8+w5g2Zw9sV3YCzGf14qbHP7Y6LxslXZSKdt
VO5YdLZW2xXwIcs0BLDPMlNWe8qIE6cqENLR8VqvFKscAntHBOUKgpeg4t4TzBt20jH2EVg8yMfc
epnnYiUAT+aNX2wwxsjYRTq9kLNHrKS2NpCeAyRo7pCCSNPRNhMIdPwGWTIlusbTR+96dSKQexl5
lR0nb7DRXiA3IH4jWMNnn5qCEg0lImdSP/rq4FfTGxx6zj0/7VXRZljhn2FXrSJkPP6/kU/+b7dT
bvfVvAYfyqGXWI4BPEiFznuYWrc2kWhMchCQ5igBFq/301BzEOYb6fsgyZWzhY/6Ma4DrN/Av29C
0L0ZUpEK6AGND9I7jwRCHvSaNrRhZnljzBgNHcZiAjcyOazKtOJnYYLc7YRZKj7B54cyG6dtXv10
E4kV/oKXUjaYEy8pnqY7ycr7bRRmBxTvWgKns9Dw4ZD4Od1ELPrZ2AueEkACJnJoefVnZDsjngqa
gU9EtpDE9PtuDLs4GrPBDJF3tqf48z0xrizqpyysnUWZQBP90F31f28WkdqkMe7T3Geon+VS/590
YnkNZvhcxM3rVrodLkh/qRwigdBP9tMBkBPl+9WA9T22W4cxg86QuClbIdyYccsV6V2mLvEb0CGv
pMmbtMpkReryM37ku47TScnj0rpgfGrQejIyEQSN2Yq63fGBGgiLxXLUIMpNzDFzcJBsfdwx9LLN
3xY4Zt6AxWwSKuwaY0MEOnT1gWlzt5bKBJdgM05VEg0k0+Kz6kdMMJGVTDxA4Wjih2uu1k43/jMF
6T5zvsZtDNAsFPO04MlZTB9HKp03o5q2ZOXVYUJGwyAy+6sykelKCB1CcuJGbCOdVqhqu5agAtWw
+bnZ6EAcNTzAI/xPSEs6XLmGKlaxvEekYCZo084ofgFliG/N0zntiYBEsePV4dPq3rJFpcEjwLT0
OfvZ9ThBsn/RJU+WjGGTMUCdIF/yvP5Zx7QA3JPMA2P1LdMvzm3ORsmZXLMOpbAd3gEnHQ33MlJv
/n9tzcw875fjF2OH3dGv881AXWdsNAbe+uA3t65uRl2UZUaFHDNQlgUfC1eOrW7nGtRNaLqAH7jq
TjZJbEomebXnEn6QM70Ug14tCvrkwrUyN4yzerJiMMGRL8NRuFSYVSyts3P1O9816q1bwhWNPdQa
F4tcM43TTChGclmgoC1dQ0o5yq1eq+Xtc2JBgIFx+nxdMrRkqYcr2mQ137I3h6Sz1XacPc0r96Pg
k+n1WdR1Bj1ElthUJkMS9RQdhxMf+cpreJCzX1WYdGHxQ6+XfALXIxaCgqXXEoRWpwI3wyDFNXA7
vSD6dNgvcKPTV5w5rZrnSVVeBgFNzIw2jj/1mJTBOBv8AO2PQ8BeULhFjN1+Jh+jayPeEg1EF8aR
jFwCrUsiTNGbd9FwAjzmVBiPYRmHeiqxaY1Q7+hyLvz8O3mcNsfiId1fKiox/0Qsb44AQgOy6SOH
L6f4QiBrGW3h73K5opqHhBSzr09Iuok3VwnY7sgafKd60cZX00oFMA8K3fYIN2Vhtir9eKTM7Mw6
UcpORfWOcfZv49JqZauhABhDCaHaQeIN17lhcqWDYWIi/sg2MRsnOsjkY3QpWUe0+8EBEuN+7WrT
oLrQVdq+aGREefCq1tTVMFVUuREApKawFQG/E68ljiayaHbYscJEUYJh9IQGEMx+jcWmMu4WtF9k
fcNiem3a/4hnmYM2OaDTtvZxGkqoKwGUnMyqUSH+vJKEnGWTro/oSfUmg6HK+lghYuqXKCR0izfq
/vBNmfWu2KE9jqy5SnP13dduDXPS1upo0PqnzBJ8J0tPJD6OHUApasMh7aHVNsbRHyYiwKt85fR5
wQnU7/JGk0jw407R4NMAvYO2YSAq+p8dgpo50H13H4i4+h/JMbx/6iHQ+u4Vm/oPhbiFfG6+sdin
ycbzQOdfdoZamro3PWO+79tTxvp4YllAnCnseyjS3v0VK3Re8cCIg361CgTeTRDann8ZA9HGJ/42
Wg0MXDiDoMhBWeVsMOLAAYo5//54DCSHfucjIoAMNkSgEGyUO1KNFZ7akR3iQG5gQPrHhH4pGvZR
6EsyGiUZfMPWH7RIgMpus3V+Gep5S0KqUqnhNlavC+ZdLb4ZYJTs7ekMYVaswH1MznIY7d74qJs/
COUSdqM2sJ8f2aoKddTSJZfo3Jr3yTsYs82AxJ/AcSBAKz/2KJOjTsbkiFbMibGxSZRD59u00q2c
o/I2wnSSZ+KDRtJn0YedQkQeqDsA2YI1N8UWqKamtgMln8XAjHehzSyh/8t+tocx64kwTSIzdqaZ
YU/9Ner1OHCjrFDne1TPPuWgl8M1bNDv6puAH0e/kxCaChKaQb7o/orYrFiQUEumaivcywpN5Gyd
delDCa/LGx8tkfs4Wi0xjMNHuJUeos1Opda80OMTrkPwZiaHHSKqDK6DgF6zuL0qaaksuLXnBOyG
SqlGOwDUYQ6YqbNgcD50EGqM4hCJEUROYp4F2wfLY8M4AcyFjRlK1hkwF1nQlpWRvW2HAChyMYCk
vYlNHZsiNQYdEneCr3EVWC/jjKtT6usT/rHJcyL46vR7xuCUZcloEcHcOv5h++qEljKGYkxwAl+u
T5+i2SCXYfWAzMDhgAzvL99eYJASvMmwwCudK2uqdZtIqvBU9BrvxhCd0bK3dXiU7PLcaMrfC87o
aRpCgcj6VJTs/nipNOTzqgr07sQfCDqc65B+/+jyJm9wRat2da1/Z0QMcpWSro7T3qZsLIOrlVJI
RS2BwEC1sBNDSr77G3vPPGbhrkANDOjjgBYft5eMHw/fa7oPbstSuFnshSHR+OGsMIHDaL4qPvlH
1nHKLU9Wqt+CpAgqbOdqsdf4evGe66iN+pU4xFMLIZtHKYjgxAMSLFH95mSxHBxvSAsln77W3H6y
qyXate0zbOwhOPUwT5QrWbE2AsM2RhiM4Z9cQ42AhD9oV0arlCEpIo8TU8S+xadAtqttVbDIyEAQ
o88texw0IGeRfW5uL77zd6pba+Vs0B3tXARYAG5xMKKN4/AD2HvGZqQkc7w2zxAJhL638X9QE/Ih
YpVfeK2kTuyRwjW+K7Ucf2iW1ryNrHjBvr3t4r906RSjypFfXonao3aycbhsnvWEeINEOzzWNiYs
M5BidTGSnpR6hLuQSoorJJ1Qy3Up9ZKASn0EAgSA4kDWFVBgVzSIdXvo6cKfdVqrmWxhJiZf7NkE
se9G0zO5nWvqA3QSFSumKqZF8QoyO48Aoryf8ci22WTxAoEdzz20AKjFoxgkh0ByjGjFD8OXOOyc
h/Rz1GLY/4t1zWtz+uNfS/J8pm5GpnqpENQJz1oltFUd3Psfyowk/po5xtNG9ZllG+5dwxy18oO9
L+Mf2jKpwppHoHUvDxAg+q4Kst1FOv3l5dAYtko5lySVMQduAgS7MngRm0FqnkTgEy7xTTMerSBv
Dcb4NBft4fy/hpPTKccJf0wFcjBAweraLPtNTSKjJKScktFz0w4FzlqpKZ/Ur8jJ9TdFU3EICrSg
JgtMwODoVFlqwHIp9dsUHb4y+TAjiO8kV2laNGuCssBAR0vz1ebpj3AjV4FDS3VlKUZ5g0raDLlp
SmHgh1Q/JMHdUVLwcnZALxq4hBlUzEmyygiL9XOWNMSIFsyX7tkl0mMBeXgc/+EaYVPbda4e4Mc2
mffjcMyBch7xsxork3O38fO8HitMDKSvm/CAObMqec5Uq95coukYIvPv8C4zE9LdX1PTUdsqjYCK
9aw/yOHjxWPuOBdRdQDh/ZQEnbdJ82Z2f1x5EUpVomwgIIyeArPW/RuOnvqpEt5S2A1zc1lSBQXE
qdASI/HB8QZI4BZJw4osbfRZ+2Hwm1zMihQwt0ilPiePUOQ7ndIwezPDoE19mzVAXDAoXR8SbNvm
YiKb8YEylX5nIuVcD8WaqxJ2OEVGIXWMJseoxaLA+sup80udy3ex6yU/a5CgZPKDVPGVQeMFd3fZ
HSdPgSkU1hmetLMD0p9uhx2/m4PUZjsGsRo+MNPw7vcZc+/SbDbNwshi4P8/Nexb8AvWmUszx48G
3mHroAg+CZjzvdl8b3KtkXwPagyOXwkMHUsHAGlNoPwTm9uuH9C4Kx66n6vTxWk9bd51GMueI+vK
mxSgmRTAsR3Af1ljIBvAK6jzWMc1ECcIzo2GPUEI/VCptPKF2kNBmKRnjtfquHngFh50BhKInjRR
pB76LZfHWAD93jgo2DlX4XFxtA3V5eR9XeYS0NNWLomwuF+0C4afH93eXwVZ9zdp/o4aek2IA816
49p7ImNZU9x1t/PjL4LU55EZVCKXDwDHGNbwJoSGhsoU0SGOiyw2aJx1yLfRxRaMTB6mwySxy64H
4InfMuy5Oc0NiCyOzzxb0DjmFzlFC/K7/MrZDdFx/ouL6xELB8Y8BVdNlBwG/xWKjcCtrCy7Cz8Y
Dx0ydx3L/AUWOpTktX3bQ8b/qFaV/mqrlW+7uhxZPcq+QgmklKRqch98vKwJr4IPJFN3e9ZNHNHO
qANGQ6v6KDGrOptCRFQOFrkMFzKVdNK0ztlb+C/vMbI7nu2zylhZQGKDeCTIpF54BKLhzFXuSO7P
SpFUsljmSg88bDvwFUBnSR91bqvTkhb793TYgp7ZYNZdnRdbmC0lp3KoGKr04pDZpGABctiHVGCl
tK84JEsscD37Qu+nKNF6l4q/zmdjmk6vG7B2SgQCVaeu8py4aLDbYOuMPVvxxgyN7wKq94/WeDwt
9INKSBrLM+sEoYP7BTpCY39u9qgxGWMAD1RciVvWNgEHwmMu9hahHXmPcP2zg51DhCipI2aWtUoY
+EUIY0Yip8bI7VkEPQ7iTSffDg/st4XCAXAHFIZ07sBfQ6J6lG8tWef7Pog3W06gyrovoUVFofmS
E4jLhAhtkntTEjrrJXlr7FsoDwevEZVe8a74XEIpuE5es8wKGDqht1PYXTVN16Wdt/czieaRAE6h
YrQAq0mA1PFd1ESmhAZ9Xpu+jTNUH9jOcZn7C/dU5IxXbUv19D53uIKBUlZuD4Q2BSH3wAPae/S0
gffCKtM7+gtz+/H8F624Q2iAm5nsnDmKE1srqsPGHCEybXOXXV/o1uLIG4KjDu8VbpksnHSPPdE4
GBtw2TKnidk7c8lPZWhG3HfaP0w6jaHtU8grA6xVDU4NGisvi2VB5y0Nr1xGReITeypIXkTakCOY
B0I3MTuGWYhqsT7W+daQSkxdO/eWeyT8BVlKCZuXQ2IGWV4+2/3LY4qt7a/jVNqN5iW3ZfPrg9Wc
G5zNQFkwElhCAbPQEMGM2HqpcoVy8mV2hUMrE1dNkCR/jfgI8i6hx9vhzGqUW++vzlasIi3F714C
KBKYIHsHWWJBc6OFj4Lp2AT+ZJy6V3Mr+AT6C9RxoTaXygl5yG4OT00R8lm+6blWzvBDbC7620d9
p6LRLP0GzoZxnJ7yz0BwQh1q33k4OKRvU8lpBy1Ab/YYT9Yl7yREwPSFsujam7YXpHO9U/da2WaZ
Am49enV1cJKkSLl5cd3C94o0lrrw5aD6sJqo9Syn4OA3Q59SzTzrmf3LoW8T+luPJ2HBsX6u9jiN
pMdrKu6RxaLXtGXDRRBOTqp9R/5Z1HLo45e83rUYfrP6WHutw3si8gBvGBeCjM4riC+znNYQT4dB
Svz+ANlkCgRC0fgu/UTvZRTqhSwnvZ5Tw0GMCIcyLl/A1Da6BBVdPsDYVOyi7RT17nP1g6rSNnSG
iueyJOOZDR006C2CYvhQUnPHDJzNSUXBPhX1l8GdobSZJrMbFZWNA2CeX7nt7sqTMIV48pDAXiTp
fs9fyQha3xgBkWfsnpVHLRY8sDBb26A+ErZYLuoW2/VNxNO9KkBxiuu5Uu75hQi2cqx+6J5j8NE7
Z4tz+OJRNeq1Mh1cAjbm83GNNLyyxZHnawWnXjL3GtYc/lXHd4bHnRA/D0xQr08KiKrUtOPz3Ftt
ly1bsWxroSXRRewDZYLozqcRrHXCxoKDeBvhHrVurnjeUYL0nwopAn+JUe6m+VxSgLUzMmliR9dQ
Iq2MmVb1R2w7/sriec2ZrmLbvuaFq715RrdxiLGGHuAeTb1PkFqZKg1re9vLL+pVJn5LKEEVFyfv
dQrC9u6JleWGWfWVjnb3VYb5IDB33zuV5zRGM5hCoZfsMWsTzI27lUkc6uPixvMIu5Rizn5tELLr
RZyuS+Yfm6wTZ7v6u7NELwL7OVZczbwPaLWZ2yzIea5tVqA9pJ4s7lKc3CoUWqD/9EqOt3+CpYaJ
+Pyr2+3Sl1rZ63CtcJ9aKcDaKBu27hFgOnnoIAx2tfo+HBq3DPXVzAnq/OZ//k5KB617evAa9N1M
dWcPoCqLYEtOqE/9hCuqk6KSPCh0dCp1S26im89W3W1lhpXu/KtsjLoEuEg/gdhQHPQrYh4VFRUL
JGnoe5RqRHN2mlqPunc1GsYY9vkbn4Uexs0KCYmph+/POi8Xy2i9aV7fW9Zsa8uM8GmhMuulobNa
Xj3X3CTBaoE3P6kdXcEo4AxCSCpJTn+PzDKr6uaeqX3IgOFssj8NEIMphyiGSMK/UTSHNhzpfoWQ
Nzp8FtkJsDcb3BOXvcAgtm2zCIDL84ox6myqgCmOmEkzZeq9Aw6l3JjPm2onZfPR6VMeGIUQ19qY
doQ18LLX7oAxWrQRnoZ0Z/QBDmhrSiwaMH0jwG3VDWHvUXwKOogmeyozN5/zntp/zlg/OfLPppu+
ET/he/aykzDk6PgOq5T+ICnBmChdU6zmY3IdzLEDC5MYWOWyQrH1z/B3NALwFW+UXt+LM/cIBJ4u
zLH6+UHdKTLZlWPTs4qr8RnjFyvpx9eWEk971lUgvrJ4+kUamXRVL00RhEiavf/x+UtvA5KBuk/x
G4tDR4Vy9Y81Xxr3cN7kNZ4TZzYqJ6JoM1A7PAN2dvIRXA+bdjLjILS9HpyFlg8mJBz4Jysp94VL
ksg9rwxjPcJBmHIpUe9EtoYx9J6/HBgoeZdp8R+COkkJt8g529h+1EoNX+GpIMYyiM5lKJwz0SYC
EXNA6R7q60+JJmOsaCBLayX+aUcz8h1O7uA0D3PrROPeUQLBgjiKc7TXDx+wJpBPLmO6vazRaI++
iBJVRZzTR9Xzz24bP70f1OnAPtxjKfvIt4494exDkfhwqlY3OP+/xPXU+GXuuGWIGqGyoqkI3HPO
cq5WlneK+7jwmn9RM+vUIgvnht6k/ct094z5VofJCznYcEh6Q9Lu6UxrtQqdgfh1gXA5XHCkGLPp
H+PDaXqRlwwnL1a+CatQjZK+am9GaEVLaCoJ9NZQAQMahGw8nSgSNlNg8GI2UziBRleTcluZe46I
eeRLAAd/+3m9SjF2kCqg/EMq70zxNcIo3YWb54k3mkYn9bRs3SeSY3G8cGiFXXZrerOZaK47uHuU
KECG10kmqy+EKUryhu7UwrnMr+y+czBOj2rl0StjhF8IABs+SG40tnWR7tAFQ+orG8LmCjaJaq+F
rlWMlz0mqg5NVPeT4KiERe4ojyOzxB4+WdU/S4e0nHSF3hXiaOjEdUSuDtUABnpM/27w971S5IwK
gB1yE1Lr3JY4mPtbvp2bY++TOISJRhsCIzgj52bnjyIs8XuQyUPX1bbkmL/QJ0XtXWiRlEWoMeJB
W1zjqJ1f/x3QkPraS8POgnvlnz6lETSNSaM0C8Ai8Rar4sSWblU9DxPOmC3NEc7IrhZU99/HfPJs
KJTyB1aNsM5bHT2fCj2OAqRVvMNyaXgzKkJyq3wr2+KhAv8gDJW86VX9fDH0JEUAiNrpMFJxky7f
5Z+ed/biIPtV2+/tgjxhj0ZJa/L6OeNiQb2JxF5xrFSWyrgFDbGKh5YP16X9aTdLjPo9M1lSTu4V
LBIRh9wJXlQYi5IL+sowlfMCRvzzxwsJyZ3hJ87TtZfisJs7lsSBMi0cPIGSGGsWZpxgaTTGAqXP
HCMtOI/ID3ese5BxD+vH0HTx4EITWtKO0jv8MVZOgmLjgLxAoD12qAtMs1DRklJyDU6LQoHkvHI0
Y1TRmrXjIC7GYaCy0yiuhZwsA9pvseWmflUhD7jqO3aFEd5VAfWZjO6uhxx+JdhBdmsFECnZwYqe
IrzyvbmAXdsYhCTAflnrValz2sroimM1/VKNAfDj0zcMU7VvQ+p5NxMqdAUbPZEH1KE6gJu5O+s9
DbLhHcTd1PEDS3TRqIi1pC5Lcoqo/16X3KWNukk2AzBdCWH4ChK/rFag7A0ApHVHNfDV8b7bnmTz
+FPco9ZMEOSdv6QNxuRlsnqYooEsv4DMIwXg5yfc+IfiSFWyCMVlNbkNYCtR6IGiGyuFdR6valKB
57K881yGHEe8LP6TIR1dxxtu+tq1SyVY+FjlBdyXIovtSooqbe7hAqdnc86j5X/9ciQxlnwwaQ0i
vN+f/7zbQR2INSfz9DoOdpCBtwL+qezH6o+mKkF2jbrchpdxZNpGZA97G1D8s4ODaDplq/03WhhP
S5iI1KhpchRR949X4NjQ+FlK7Hcvl5gjVgBHXTqwX/Fhrlc5nfkhwRQXIn2UvGPdsLTEbk6XW0wU
twX0WYXTwZssktij0UyF5i85+oZx8LdFCR+b9XVrQwuzpan0ux4zaC7abXf1tOkD+vlu+ih9gEYR
njkfi817au1hAw6p911XO/NtusLqC0W5kAZYhcxQzFfYsoQkWs92bIUINPMajddic4JFGvUmu5hg
sjXlFIh2JH4l65HTVwju0n4VZf4SMGZK2C0TU+qYD5whwDo/J1O1mchJNqIYCaVxVHLV06jXOViO
v/TwE2i/soXhvp2dg6hy1NgoHbAKpoSAF2Jvhw6bk/e8MjMEn//xt4M6E/kckt7UnoDbobs4dg7f
IGeBAtRQhkvW3ck8wGchnowjtMB9yqwckwaV48lOLdRgqL25AWV3fzv4Pa8M2I8l+H/m2Xt/Uzn4
z9o3/0iAuHDt2NfuMoxyEYouTsip04QF+DyHtjKbXlepQ46dn48elgCLNpw6TXFx0hZaaw14k5QC
zCCKWci+HnbUUrgK6VJBUyf7MJxaufKwlz1sC/DJAVekYd4GkNQSj0rYPy7aYuQ7oZfYxA2io80h
POvbmQ5dzdSOMs3HDfVF3WspgNXti+53StOV6LYrRAde/D9wuc1XyhCOFQ7oM6+F39YPhqaoDj8i
Wrxj8j3IrxvhMNnQpIoEVCxcIDTBXFFiw/Q84hgUC/hCYkrevuKUOUuASkliBkd7uHuf8zKlxjnt
FPX18NHTl5H7xNh/eq+Faf07w1UJwIpV9TUjsUuJoF0PocAcPTnH/l0OOWONs5h+pIb0Z2EmZcRK
21BFimlwKZ3QOOELyvWBnEfWivU3fVGlH+4MKjIri2fVZ+bIoEeLA4Sg1YwsoDiRjEw4YMqbIkgz
apCeVqmYNKLuCtE1D7J+wBZAlRkyJHf2fc5pPl1kEXch4z7fysLJ2ntNSdyHc/kYf6ALnu1U+RHX
XRhTUF8O4/9zmRjegE1VLTaE1ymdWhNXS3gRPKd/3S0UnIrlZ9kYCl3N+X612Vd4CVCLFSBRczdC
ZztVWR6GUdul2QrV4CQeCtg6RG4HtP+Qcgvwqw2EsROOkkIWLQ/hvhRwzwQUnrsGCQZHcsJm0xNi
Sv3EMUlcG9X9EqeGI1fx6cuwvb2wp04nrMNQjTbmkWkJ7+WmQwN6WYOYhFfmATRtspvwjjBsEIWk
uJGmJuUAcnxlHgJw5ATO7mWXCdgUOlRrJSjlGsRm04SuAXqNsiFgavZfQiPRbwIRulGmcRFTBYfj
zI089baeo1yqIaPYhJtAFr3lsu6tXuFz/7V9bmWivHKI/Qu7JUaSBylU4ElV3wXYducnSwBkMqYl
uNUUeIBKODaWF3uxAA7J/99BEtyD1HZnDtqvrHYZBIShw9X7/3lkM7NYzmsnXG1Be3MEpIT/gjNK
QESqJ1Uw2H8DAyt+aEf7eISGmgj/V6+CcbfkEmzqqYIDQDHB1nwVQeuqeOHNJTS+qzTSRjRnuzfg
I/nT2PWq0wGuE5az1LazjTZnn3FOfBzEJXnpiSnJYYmBlKSH7M/SUhreY7qJyoUxS2DBhEUTo0r2
YDDdx/gxjsiFfJss47Vl0+N9IbbljbSYwTqPS87kWn6acoLM74K+VgdUl4RRzqqYa5yKOIvoy/KX
irEX2WqsrSi0Ww5BgEzqsVqa7074AETFYBY4ERP/CNOa0J2bRJ1siDqhc+P4aAaruusgXUEAtOk+
xPIqhINpTFPVA3V/lmkjdYvEb3zwEjknTdq9DzvzIkFqKjjlk3Oy/IXKFr/lHTDJadHfn0SvJuL6
wPh052cmy6/YpZr39lYJUiaXOYCa16bFZMjPGthLWi6I1NeQFxs+3IYiOnzrB+1oe3IK8ivCFNJ9
Uvlw07FFK93+vc2hQ7B7XrnNmLzC00FgJ1HcDy+2U2iTOVqUISmaZe6WsxlOULsCRzIP6UlNfSoK
aKaoLIUN/lRIya6pyEfLDLC99y75WUBJBK6SBuE1hWtP5jHdnzKVinhVHLoAbK3zCAXPs8+g2Mip
9ZlRt5ufgQw265s+9lqJZrlmu3z7eb4smsvoGICrLbWFxDkZJjqu7vPDX5aAmcrNGOoF9gTZ/3QG
BFEvF1XvgeppinFkHw5LvuVtdk5NDCQfWgwZvgkeqMBBVC94uxaKp+rMzqE1HgHIqLNWQvDsRtTr
LTvIVWLEHksRFdeU7dvI08OzO2Spw2dNtDEuVIOObb5MLGNqvjlvms5LbAjlcYq3apRzH2p0X3gH
kOerp9EhWLHXtfKVxuV8SUzMXa3NBoiWkjNfciyVTn8vCvZt5YFmJKg2Xnqc5nmg5Gdj8dk+WV+j
3qdQWkDhk5u3VfcMt52MLYq+TZLojiEZTiP7YF7l+KLshHxex3HmgZ2uVzfD6gNtf6y73QXWtzbW
6OZyT2yF8oDjWDCpNjx36KgrGu/E7wk6R2D46s9zDjyb+b/iTjZwo6sS/sJZhtQkmFOS8bMUNf+u
FGv717W9hB3wlKMKTFdEKh+fxcvlB8ERCjmbWKD2j4gKadsJ2GbBm6mf26NkTXj1U5BHv0SGUEwD
RKfeFNyUp4xXlxrkwYPkyVFZ5/yNIic4faXEtRW8dSd0bjFKbhLic4pH4IB89HMPjI+KMrkuxjkE
CZbo21wcqg0nWXgbwe7dNvBDphI07z7iqKYceXuP5Aa+DD3RlqjE4+tbyXAnrVxRaqoHR2gBE+Zk
3ndbP0CEW4HNADk0YUQN+2Ib+3vXzdvFGkdpTmY4DQAUlfEb6ty3AXjcV4Pcicqcc9pynjDbvOCR
7zNEHK/WUh4vdtaY8MRaQBiUaDRIye9in5DwHBTh9vPpdVi97HW5hJWD/6YezMwgcdQJUChezsk6
b/OOr+V23j+s1A4Tykdn1w4Pyao/RagB/50+mSRidPk6+zoyH4PIv+gn2Iyxv+ODdTmMRkFZ3fOK
bEsNgeH7+YPc4m9k+vbnQf70kRCDpLZi16oj3Ou0aNNYwo95zZ228oxr2UpbaA8JLDw7vCkioZNf
3gq/foRTruRPWjQSIdaaCd1dcJxOMbJuiKVG8qoRUh73xtgPcTVH0bbRjrIELe2glbLX8AeVX9yM
ST3lfhSyxdm0B2m7zrhR1QTsZollSXHAtSdrCwRmzjXVUpZukjK1Rwq+6VHHk5Mpg7f2g2dVWgdn
Y5GQ8hBGomNFLkYUl53+ryDcmi0YcighujczIHWL9PfA+opbjcWvVP/t16IIZq+QQAvq5HgqCkMW
HsWqJZar/PwwiedrySz/siOdzUAJ2x+/PLRFzwxkIS2XSnpVcJkdPBuwrfoTQkqDBB8eAbUwk23L
6GYodpxUY+ZT4QjlW+wsxwKLrY8van4UpM/gSxXwDUoAYmTOyJb5hxyQX5U81tNqDXgulGC8pqTH
zB3m4LJoW2OTNW9WRLOsPPECPaIFOuZ8Xulq0I64/An2nWh+hI6I02zZGV70eXiZwmJjs05vpHCM
7eqRa7L6AYPL4tYT+bYkeBsRrhWd0cmRm41ktJvINE81AS1KecwoqYSXqDoSgiGSr2npt4rdebGu
2epkvFU2wqUuH0l91frVhwq11RqTc+UTgjzkXnoAA4nrgAOuVUQVPtENAC8Re5INSs5JpJcxqoU+
iFS07iLtLNlr7bDkyjE2ZhtnZFTaXPn9sRxuksxah2k0R/HuXgb5rHxVAmv7aE1O4XG8IQnarXLv
thaltXQOnzSuyDDcyHbc+Gf5qcWWK/QGvlp/aL4HMJp2OiqE4fTYNqIKFAEJyLaL2OByQOC8JkV0
6pgLKMK/XxES7BJ6ntqScdPmaT2dqkQwCm0hPjm2KaI9Zz5lpiVyvT1WNCc2icEQXloU8nDS3C4L
RZ4A9xfQ3WmCpBj79gdlZvanAfuRvItejrap+08DhzZA4URKeJwMUKAiPtSREmuHXpyiIvj6OyC2
3kzpUlD+ZqLHzjm1LnVWcOEuw7G8x5pgM4Kwm+q6qW9Uv6ow2UM2dCtxNagwAoLx9eUirujpG7Af
jClU7e57plYM4dY0SIuFPHp2tiukHevTKdVm0ulA96EUaSlJ6z0e19mjmsK0vGyhtFdrJzN2maHd
uj4hiU6GjLGmTtljKoyhkdBUpEIGyTduk4ZqCzLYuXA9X5P8FVVw06mScPWKq7nX3p51T7nBcH97
S1g189LgbGu4hO7foGLKfacoCrvGMzM539IpP/DaFGX7SH1sA6Ge7FrEsXguUDXzWua2wlByrfgL
wpV3M1QKLkUfLTyG7oWHRoqfjPf70b57KL9K2KzPxh6fb1biSIP1QivIY//3JZ8AWrIpYxHHajdo
BXF4a8sq/nR0hyEU0p83YtnrwTkNa0ZhktD4+UPLb4jlu0/uhPB+oVfQai5Oi05iV/x9Y/uckhAJ
l8HY434riT4VkbNdAa21A6oTQQiIwFmQBTIfE0R+KsZsmq8DraE/R4CMBCS8N2hVLBmIgSAKBr9+
9/A/O5xu/Mk6Qpdnm0jCXyOYRJVFDimnsC3mdWKDQF+nBd1dXThHlFfLLECcko3MEZbr8oTW8djO
bN1yVNY/Ot91PONl4VbTV5KG5wUeDkf8oRlC4jYhNnWqCZKXR8nUrKQajv6Kh0zjdjaEvTfTnKP7
G2DTlfDStzB95nImnYXTNOsX9O8UOw3ieJgrUYtthXJTY++gcw4PGJJEzbDFtul8955+hUw3Nk8n
kMl8uPvg/iVD9ZktC+OEaX7vNQErRSriZzu4kvLK3LPt5fT6mMvVZqTNuKA0wD3h4o2I0teKN5sy
KtoAfxKThGjrAbZhT8uIKUYNe0x47gIQuS32Eku9KVA1LC5EarJeEzZ5dTqMaNNF2ngsCE1VYBDs
XRzJQhkf46cP+vHTEB/AJT4e3D7yuXJXDhC7UicsTL8X4ChY6+K+hsAUbkdL41V2+0aaxHC3Wb6L
BIfRnCJjNryPO1t/w7N6F6SSv+ircq/USQqyGIfxCwIRDoCHHLyh3EEltpE22UCPbE/c+ieq4i+c
v7FtHUMYH07gxozGCoSLAm/uaHKo5K3iPR3/svHK0fdqqUCOvaoT0KxRXcedc/MfuYnJTFluwDhm
/5egk+COKg7sarPUVhFmzy5oCNmcjFdEIz9z8Rt/WOKHOJdDgtzcUjgeCOnu+GMs59OFgrADGNdz
X1COOvMhOxwya804d83NwBi6hqgj2wbnTVT9RRHP+CdeHgVAsa4UgejzPgLWVukMasH6M+tfGdTF
Dt7ltPOc2D1Y7/7/yVohs1ELJxTxsXx9z6e76G+hqheJC+OmXDOrcPxXpZvb1vUe5xB5G2gQEulF
sntquJD82/xS5b0TA5Ns5wRtyZTYDe/USdosC0ZaK4RJAeAJ9qBKGt5uFyoC4GoQND28SIG7kd/B
Yzl8EyyLJLtcWBZXXbWx5LV26oyBoBC47YO6Di0TeiIb9R4RbVuCRcsIH+5yFfWXV272a+NIzRQQ
yMg3JirksFIsUd8EfU8WaCfWV/Z42ZzC/QjsBHqZlUmE2T46CD7UGDN8Bx7WvHF2NUIkv6VOSdqE
4RAnuyMx2cE/HPkvpr0jDjW+sjl/1ESakScw7fUWZ8GUVsxxapqk0gC+ZXGHoSdz8oXMg/YAb2OT
Z7usNDImeMLFj9rxEH6YW1xsfhq8q3xLdD0+9iMne8B8LwuaqOKLwpXHcuv8rbQUxyXIkYhPAs0g
PEovUSUmcmHGjawUzy3IPtj5p2/kbQMGB+mtpKNtK0p9XSYeEqNcQJb8rgHTjz+3+EL/z6ZSEr/Q
vqD6vB5RZQ5PHhH8wWhklzed7XCwRZBTSZxAeEzNNrCEVImNZ8MhcJ3AkB3Cd+DPxgOInXlRPIDd
q2eCBA3AX+kpnja6QSacAYq3PdMVKf+n+shabPbcXqpu+TJ5lzY0qLhENVBBoxI6MdDGrsUlJQun
Wy72XfeySlBsmaTuWuS80nvap0s+t331yXFGR9A7Jg18NL+iLmOkbE+fAeAsliZv8SQ5bybDe2AW
ocjuBC12CXY7FLJ8zFDDaWxCL2iWxLp0pnMhN05zQJmHhvF5msztz7JUFlloQA/ZUki4Y9FkyzeA
kTgl8gDN8/RYFTyTYOt6tPOVaHkLfDUDVSHX1BEwZOz3oWwkJ2nPKR5lmBF1waaDQt70loNVME9s
Oatw2xMVF4yDWrfesB2snxteqts5WtDlWcqphbdQd5X+oX0O7K6zhO+QoZsO3x7ZR9FeggiOhUIP
KCJg1pmjWXPfdsZcyrgu3ukFE8ZCkM1lYSlyI8g65LqBBCF2Rhj4buqvsf8+M7oJYTzyFr3AtgmQ
MM/toFaD0rPYhYZLnag1O/RGsFzcJgDKyLx5VuOYkNXghwE83VbJI8hM+O3Z3XV/EAD9jZwShdC0
ZFT76SLTuIri3+8AcHmw7iveesqln5dyMXmVaQ93iTK1GdNfuph/eMpk2nCURVVHTpl1BjnclnGt
rpnRnLFbBbluJao30/30U8CSglr76bwivZsAOBC0PA/uwuffuBTYZatqo7XLXL2ieN4kFdEeGbzB
m6SFWGK7NZYoiZbS/ItRCfcsgPXJxkgqLM+TUP8o46uj1Hg2wO+bbC9fPALC9r/ewA6J9cbYe7ut
wFOS3gDf6Am2YP6Q7vf8F5Uip5ayBGl7YzXqN2BmMaqcZQ0vNrOLDnlOupkLXEaxtkMUXk1nUAuc
I6ki0CmpOBkI7Ov4DuDaUuT50FB8Z+Ty7niYl2BEV61gUVBvH8awSXtK0FBe5BOIT0rE0x70ULOq
h4vq1YD2VmK4xnjRx3INe+c6uAtIRkp9sdwTHO9aQZW6Lu8owbCBZD4B7JASZnRXCkESiz0G7I8p
o4azDan22xka6DNWz6wcZgOu1X4kYjgphDBSU3JKlEcHEipPxM18VRsTMXNP/XI6B6vlULIw5PqJ
WMYBDw5coQgwztlg5urVXYxGbvbxYeUKnPlNJF049xIjKSGUxfZTJXN+F63J/PQ8M9DVgaBucyDd
OvavZ/enrdFoGhGKFojp/mk2FuAal+Zdy55EUMQD5Lf7QFgwjzj/7jyxsRCHS15j12aVE4RKHq9j
jckqAPMYkzz2sim3Y0QSeheBRUNq1eiPxpKlJF5QNmGT3btJCHcrQ50u38kXdHse4ddYiHl3Yx9y
GkXrSDGZ+oqC575GAZZR7HlK2Hv5v58mt0DYQqfBO1t1lG0Uj/HXgkjdB/KKbY+5zUIkbEettt8u
T2f/4BE6v0ZN8PxElsjzy1RWX6XZfKbX7vsS6yJ4RNKzmrpspBh1zjYua3zvse9tyNmt/S/qyhsl
89UNCKNfebPNODFCxg7eV7qz+XpBPp8Ard/5SoZf2DMuDQbJgSgrbRzy5Qw1/EYWXsqVbIzQGnX8
IgKJQReejrhswJ6h+v1mL0cni1LOqfzaZSqiC1hSFRDTJfVMaTYDtTmS8HzzVzIkuw8zU3xZih7a
RIjEFFzPJT4Tv8BXO6emDyapjyEUrg/rmfA2spclmRzbcG9aMsXHl95TVJeAB9Oqnbb60rkYhlRg
VboSKf+P87P+N5u/KVZMR2IYFj9Fvc8maIOot3MY0IQGYpKaa1NBA72LdLWZWJGAptxvQJ1LHDP4
WKQUGLrGyFQJUT458X0jBxg29HinfVC7Y6qI9dlk9c0/1hdjDzIjF5Z7mzdz+a8rsXvwLV0I0jYX
LMiz6FVfzoyi9RHKmXVE5pXMIjmUsTsW06yHYmfvcLVSTzu+vi/vpgpZLFHfhlO9bnmYnZ/xY0lD
7+UoJ9zPD4qejSHEnvqMLItMADhqtyqUqIkZgIByOZwE158zjKXDFoerDmv9vl+KXIqvbYdYAYqP
0nRIXszxGLz4OiMXtfuoxymLahjBMhd9gjxRnmurI27lc7Zv4Mxi6r5NIASmmpV+DN8Wo0Vbf6GB
hqaxk18E0xPYg+Fcm/FH0bBb5t4RsmonXL3w9QteQfAYqWhc7kDwfvJnC1W3k7lwFq4w06IhQSWP
JZEV9yvBO+fdMnet+6LUMH1iVcJjmU4bsYu/spYaBdgCVwoUDPY5YCbj3PRPiqwU0sICg1VJEm+m
MAp7m+O0JIqwD4jATjd0mkHpkQqdEg3RikomEojoecxZ6o+EqEzPGarWfKXLO7cL1496wUQi6x+A
VGwyL4EDkxKar/kT4S3ILW/ei7Lw7h/dUZ6D2MqEKMCEN0JQnUTL4JvP0nc5TlwZuSfb1FQSivot
S+NaXu2eVecZpoxWN2m8S6HtdrEtnejYnhiFp0/I64syWaKZeFNvk9z+63epJO9PRxnKos/BvRWp
5PjRVS8GAwMdxALPaivtEM6sTDqYh0nnoUr0NvYmbDJKpLaYJs+tRaNGD+/+pv2mewEtxi0Yj1dL
QvyYiwkBGMTSFynqhC4HSD6MZSL+sBzvIk8tbUE7PZxS4+O3xaG0hXukRIIgYDu5m8Z/8xNf5iWX
1c1rd8K2nCWDF5GVByrE6sfoA449Ogpyyyvpya6Pj+g4M3J4TiBy68+yoJ2EHhG129OPX34GkOJP
hfO5KoHUU6pu4UVET24JHt1a5C4hU888YDBbIhP+JsCUsnWo0tv87Q/rtyHHAr3fRGq3JX27ZPvr
Jj/xB5QfPCH4WFzE0oM7eS9Y4DpDseNJD7iAZMLadooFyZpyGoklRKjHY9Gs1qfbfTyDgwzWDv+n
CCaVJCDkBo3Sv3Uk08fEruIhjzwxyzsuF1gH+4c2/lMIeUwqkbbJ16V7opb+RlM3BVn1KRQ4Ud4R
hgNz7be96dNsdjEPB9TxOU9CY7pqC38/I5xarR1H2qTE8jq6bNJo+38q6RUdHvRpbmIjz11aasP+
xriSBYS5FGyPRu1ii2laWjzyz42BwuzJCBTxup7dtWH3o7PwtOtWdUW/FXevcCVasTf7WMAD93fb
xZFKTlZZxgshSKkRzsna2RPBfZDjw2crXn5TsvNDpASEFSt+tnQ6bJNjwveLpK7N33I09Wqnszqx
ryQA+CaqG21GjKoHZI+/pCEwi0KZNGjkWLMYNgXUjQVxmsTZNPsFC7QvVtA5F70k3HqNFOmrLokK
gz6fn5OLnY0G+q1DCQ6u24rwf+5qQsaXxh4Bu2hAf6fAYx4UJYHjyi+85s6TpFr3zJrWHp3UpOaE
SF0l8FLvkb98A+I5kXEY3FTTtX6mBfWpawQH3c9A73RtcqKGDbTsFI4B/Lvxdwl1X08FYCz9/OI2
G/LyXM4ySGP4hUakZviv//H7xIrYZej9H9QS66lkwOrxA7RRNA0v3HEoMU7sjx/hofvPyIfhgWYF
lWkFvQifDTnpRBOH3p6sh44DwxXvq4TnK4HjsaiWVQFip0SJwtqxkpiMQpsigs/I7nuFRV8xX82j
ciu88YwIKoCFJtOa2eRRL2/ZuowdlJ2FCT9Ax5Twn4SMalX2fkIuFbjlHDTiBjwLoxMWSNKTKNuz
DvpAiA5uofc1yH+I1HQmnmyF+KPCT972bFOeLbMpxYK7jOqSfDs6E+Nm+lXLUyi1FUGa7iVuOsPT
ZqHNF71mWgYSQqsZ9+gVkzj07MiTiaFbAQlOGLRW1Qgo0dM5ax/uuuFBASTt/xdFIEAFp4Z03mke
a7gkbPXWVbdV9sQNf7Aj2gZkzd5fVe81oWGrc25lk8HyIZwHCvAahbq6H8PbK7/q4+PqfPbN9j00
e9a94eGxcrKHxfzzbsCCCIshHzQs/dNnhTaP0iQ9t1BvJ6CuEPCbGfYtgSiPLyODmjdMogmeoXZ7
TgTco72v1IeNFvPJrLl3ckQZPOhhREo1F8eO+HmjvEEsFG+oytTKWTc5cCFGLBt8GHaU8zrBA7BS
v7EEFZXJTqAdIiLQFFGhXwLLghKHVpFgGvbBC6tJOC6ovATkQLBYoz4Hkf+v/IgSWZIu6X/mIc0E
3xVVF5AY1e57S8mryB7sKQYgJRXqlOmUJ0O6EtHgo4TUyKYtiiTTXVidEgL874O87tmx7VELIUwy
YeLqxmeDtOjvRT3ALoNF5fYovahgevXEcuaX2t76rCtJWBctMeOQ7ICSVTSESkyqu+oi3Fp+vSIP
z74aI+SCW4zHwVxmeg9vMXDO2dxP3Zhvc/qYgSPMYEfOOY4FnrFKADIeA1wq49t3EUO+yjqujCAe
Uopwwd8UILb1vgHSy+3ZvOOMZJi4qhgkvNLxifJmsPVmlEa6lfK+u35zRmjSUnt7Z4vk3QZvWfgE
RLnZQVLaqANMft5opZ8bS9IJDsBYLy2r+XUQd9cA1RigQ7tlyLKgCCBde2Bjl+gh/La0i08SzIMT
T4ZSfd6mhALK8jvkvYUyHNC+cG5cS/GpybSYqWRhxyAC+DNy6YBcNuBfdOz9j+amJ0V1QeEAuyJr
J6I4iyDNGLogi3cBftyYYKdh479fHDUuxK4LBkdLglttPqoxFWi1O5lT+vbCgWyRrJ6Rn3qH4Pqr
e+T45SxRxqo7dShkGu50+50j3O4ulqqu8GP80fEoDnuLoaNLQgAlHIa1Hva0JF7S6wQhqI/yePok
bL+MIYWoqlL+ecJ2bISHky7zLkcQOJ2JRXkisbutEF8p67EpzDpQVC7aTupNPg1kterJCk8lohF9
uoZ/WQl4HTIwfGwmlu5XVQCDy/T0U2p8Y0nWSkNzSHQG4rqUpq8xeds3jucwq+v+MOqpvEp8BcWc
XJxOQfIkNT3KOfPzJqAKXHZk5GvOgpt02cgic8lKaGjAxpLoE6ZnFyl2u7qaA4q8pV1+yy5RtGqO
g9aDcsUFNU6uWr6ba8CkOyVHDdyJf7MzLPYrvaJeN1vmdVqyvx8HE9jhAuRXI0M5et7bQ52TtXDr
TYp0aO7hMEA0fbPkR8uK+yr3QV9Ob3o9zvmNPEBQTZ9FXENe0I/RtxV+1wwogecRjIp11Kz6oifb
mjuEa6mKLek3qtLUbSPdiB/jaCgQaKo1lLaFwMyqpwOwfJgqnZZHJS8DVcAvnoMVZzW1TsI4okiA
p+nES4RRLyzAnQFmHD1q3ONiISRlL6ikuBO7loK7DP9DRAkfh8YQDdoC2LMJ52PV08xUz/VkWMkV
1UwJ/Ei+5JU1loV1r31JemzvaHJjE/Ufbkvo7LwJQjOHFpeyAFleAbZwC2IAIJr+EPlBlBdCO1Jn
tf7EwZ8PE+2cqchAbNw/9pf5o9nNAs900rb/kpIZoWdZU/T/lgYjQJVuLFTnBxPW8HVfMJKYqH7o
JMH5TcPirhr9jYPcdGP6dysZ2DOu7gtANnUzXc4ahSTxNx2+Gx+43PltgvfP425QGZUb8CiFFvi4
Vuwa+8hpaFwu6iJ4HhGcS5I/smVJP2J++1pxm2v6v+5MHI7xiwQsTpAtjwn58qlELIzupQnqpCQW
Ie65/937q89X+a/p5gL1X7Td8BR9rmu60DJX2nXsT5MxNUKmcYUqjDtWwkICnAds0fkaOS36Whzl
ReB0x01WAjg6OB+YkPyRx3cBtQbeY5yGdcCrMEPG+XfRMNEIFqekQ8oSlkp1G5ZcrBi1yWckWAo9
7BPaDuz7c8/gAEPxxA2NkqtT0xW/gsKGYufNsUnu5Ot3h+Fn+n6cYA/1Vef4eezzhRYE110KQPek
kxaL4eA8ALz24ldv2u1cInshQbyOdaANI/A+XOmpv+J64hyvAOq5VpspqTvF0V9KunCfrEJytMTE
Vnurgi8gjZx8xmtWOn0GJmf4gxJWS/U+oBdoqitRkLJB7qShe3q8xk3xXzA679uqPKf2oiE0Dq7L
0PbCr+BFL9KBxBhb/NgoStlORXO9Q8ppfRyMfncJsoVn7nGzRApblCZUE6qWHrch6uF/UTElIgrW
qWLQGSm/Lzi/6K2OpNpBgeBX3hOJCL4SedN38n0H3Y7rCjzWjiVBI/RGn8DxCi/J6t+FCFpMukpd
WpQiVXqJ9vcZtl5TWSZ6KRw1gyOy0NkNnhUUBER1d2eyvHviG60z1kPuKM1STsD/osKAhgFy80UK
hDz3eVyFugvUyI0wRaWmoVdsw6LG3vEpkCvboLevBVUw+l2+RI4Ie7Mx2JLUpdkYYCVRUYzkYiP0
75AbL1Yao+mW3OdiI0QeiEmh7TNPnwetichyo+CDcD460+z4Kf6I4AB+ay53vdNvIXcOwzeHYS7T
ZA8UF/fmt8m2IhVxWNv6xW4nqmH6pSVaryU36B2IouzyDwDn1V9U9NVwUZV5l8ZPauvNoQ1e3gRD
2coaYpUGxKJQ4SOigTZHR36jq7yQdDYkrKRQEmVnVqGaDYfHdZqguChQWHQex7CHct7anN3W5+iH
sKv18byCMXwKlEtG8pGt+hKJ7mJqkvka2Rt5oeRFPNDKGdOcabfqfEPHJEe69fYKNhaWk9grQz92
PxbH23MU9yINlFXjBhJlZ6610z8SPNcDaqDYjZPC7AqEtz02uTfFehSem+zHaFkQDaoXb4dYZ7on
ui8Xym5roqhBVFTN40C72a2B4EhVHkHxwzytrhp6sjWqlrFvZOUW9Cz1s3BKtQxXrKNXvsMmqpgQ
bMjRyoI9FyWeHKHh1XeRGUcPERe198EproSuViGgQ6a7Rr9zCDOH0oYY67A0yAmZ4XDNn9UcIOM7
ncTzOnEhd3khtrQfelzjSO0/5AhtWtRPbtE96sp/KTzpNh9ZM4Ryk/Cd53CkWdQ/Mpj2VMRdff7B
4/0Tp26n1lLjrWz7JCuyuKkFjNmZT3xxqfBVc4acZZZ9t1fJDQuPzJylKOmz8IXUmyl1oBc6AAIO
oWWFw+A0ul3iBxlOf+zBJMXDVp84pMswCAqUPkDLL4rhlf8HSGjp77HYGOQm3CMvGyTZodeITtmS
qhPVrZ1MsbmPhK9VhzfUcZFUv2uUs7H1k4zF8gi/sF0DZ4p/To3Izs8IcgFXclBlI8L2NelxRG5m
PTfPi8tih3q+nUs65Ru6XkvYTmAeE4vPU3dQFTLUVx/v0oVWMiopvaLJPZ/TO3fQcvgxHPYT1hI8
cix1P0H6uA2zhNyxA63EOs5qfiiTGpDowCV6tfX1wPQXn+WGumoZht5Vuzgq5cQpGcOhZLlYPtme
RHTgomA7h9G9nve5vAYO3NaGxf6JSOtjXkfD72pZywXFD57A2spTfl2nYv5PNnNAScXzC8RFvRmw
/WwV57ygkS/DRrIxsbwmQP3JzwDZad5tuDO2CiWxn/GBcyMm6dghoSJL6v0sMgp55srt1SCyGdoN
Asq9Yrwf2F2brOXWV34KLsd4BHNOUowf95opGNcvZ6svTtolMtrJfyv1dZbPVtr2ZXHY9ESHNsFH
YtRKO0J5j50sBr5VvXnk7JQ3GPGaVSRZs43c9AxiGsXWSL4jvVlQuxr5Uc9XQiswvTD35TXDGhOd
wc9FU4tu1PJn/3uecTx3grMSGPvS/4rxAYIZkNtzNcxuKFm5/ychxs3s1hLDECKqtvpAmV6//gQp
MBjsX9lUSpGETbFbroRiJK6tgZ0o8uZJI5lwLc0b9b+zYDRYW1p/8adtnqHNfP7TIJe+zMnUWVD/
DM6cMa11R+O+20BUzzUqWd7pT7y7Ublso8HTE0f+LAdCtVFaWs2B7IE9G6EZctEmlK6gajtBW6TR
2KBejNeqYY/pNz0HnyAowZUMsa7SaGKBbnO335v4/TSUlwgSk7KMvexyo6DkHILfZqUe+nR/y1xY
bkFi7SCxFkVWge5jtRxq0LDdxD8j1aq0Oqa5BdXDOmEJ/aKaYHbPWI+xEg89LEqWv04GSkZDKZFH
94L4rvQkJaYAmMCL9SN+LDY+yxi2C8BCssjX1MZIAJiGPamVBtgY9eQqRu5mQf5UjYOoP47U7Vu2
TccVBUkdMlKlJrbo7OTBwyYLnvDmO/LBQ8RZxtBAivZ1V3zmpUrMZUuyk/HnRDhRfH8wwmHLxq4Q
1Aea3lgQUlHsYFvRxo+5b6/Uhydacdz/Cnp3ZQt4InVkOuIGuU9kKXnVfHy7KbxW8wBzgl2wQu0v
sI+EEQ6DrVG/9vMl8JNWtNeL3osNuWcr5PV+KdYR2o3IRE+Ao8ew/6PRvmjxCXCG1vYU+38i256+
fy8b+Q+0tTnzxJDxMjKSgIgvQOhf2F6ltBSgbRV6ErIE9uIpDdfjoPPMXqy47Xrr+9B3PXgEglYx
c58IgLKAn/lcPuPkEp8GizXQEF+XFKn5S8iG6j6exTPjmrIwcm6CiW2gO6SDubGfscGbzLgSL9Lr
w8z48+6dtF3OY96D98FB85l5KCQYTcQrfvXRoxmsXEg2CyhKO42gUzOcxU4FfI85eRbcGfEPOnro
B7FMEt6Pq9WQVQ2PwqiPd7stDq81LdKNH+iZjZ3hrSPsbYq0ZOE+WOMhN2XJaQ7VCxBGOmMfKPlB
HwRfuq5/VD42WBAjmdaqU0vE5iC2nvN1E7WNp0A5D33Pc/vOsttqbZ3EUiWGqGeo9IIOT9CspsLQ
mgLL2/a4813otYcQI70I33lIuH/kF2OZ/rbwXFrGdgt4N5h9jxbSKuAGVSVpKa8I8eka2wOHjjtD
Xcx1HnZZowPvj9sWSIWw0OPbokqedo5kCL9K61SmB7mFVKKr3TQGz5GayD9ys+pxbK/JMnBCijwS
5oahI3MulpMAf1crDJc+IcgjSlMoCWbqZOtwz8Z6jVvkwmAmJPSXsxtjq9qRK63pue4ISBMGse0L
lX1KXMI48FXt5cyt0U5CvznJy0MLbt5j/8gzYgfLbgAgghiKpn/oLcx5xLd5EKwbKQ/RSGfM5VNi
NzNqz0h2HNa8jyWRZxCu6xt9+h5kFsR1PRkxZEixu6+ZrDWEX3W1lOfNZgsk372Xrjfma/5e+Rz6
E3SwQqYjl/KQgNt7sjqbIXioF0nD6H9dfl856O8VeQopvoram9kuat1eug4OLiXMnetOSIywtHgY
6t3ge1ajS6P5gTU4jswG1yy5hUfprGs/jpr+5dZD8pIzAov0xCVGBSRVnwK9GzAOWLNRwztgmqep
Ujy6Qz2gPHk3HJEgJJVIWFD5NJhhRQTUrCxqZKu6kCI1zSeQUDiIEUhVs5nCkXljEz5neGXFhaZM
S8LotHMJQLG4VOTzi+B8Ifr5hrVLeLnPCpnicaU8oHDm74b3BbpKmJdlfwqoVZrpanGA8AKGDAAk
o/sn6Zg0DMDqReUmpDuMFg6egG1GM9ZO2UmpzV/z61/srK6Ktni+00gfmowVo+RZ/jUMaL5qcOgA
hLMbGV8sa1ZYnTVveZY57ZgtUeAJCqTdO5ze6laTefyrj3d23J/xNOlVDHWRc8gEz6R7FZ/Mojgg
yPuyDmlmB2ULNgkb6f6KfDQxVywseJhVouT+mX8bjBXX8HRS67Yb1xW/ZCyAzEC8V49R45GLyCvV
4ece0nieCJAbx+ZGc7coRVZX478kPTY6QyKa8QVVoLfWUdWdWEfzRQS5JkUMP5NA+aYuJyZ4yxsA
moerzeUAXP7oG6Zf8zuDCBtES4dvMRHk+VgVDlKjGbbcPvXqifyg/UXPtlqUxJvA/xNE8GWJVctv
vv36W3qALcclQoSC7zu21AqY7fgnV6oW3HW2wAEGfTXmNuSO/+udPogpqaa+n3/OBOjR0HDO2cEW
v6o4yAwholv4PbBAUEg8bjvBzJyJuvieaG6VEvozBRCaHUaQe12DPpENzDMy1telrkAe2d7TmRMv
h/S3C/viltXFyciCy/yIsanIL+b4/Xp2GWPLdbrtuo4FQ0FtvYVYfnz13pWD0NSldGG4KXPvmLns
ncq5HHYzIt7UZJeF77GirskAVEFx/PWhxmeKd/9ZIOivETZcO9OoCOn70elpk5XQCci4uSR65t8H
NbaHLSpBd5k0wtrhrzDcELKOSYl/RJJULf7HD5FtreBqugRv3LsjPlY1Z/t3tSimzH1RnwT1nfva
XtLHe7bN70jtvRPC5IJSkf4iGjHDMXX2etJpcsMIQXQ8gRtc5KU3J1j2B0ryE+R8ZlgsplL/t4Lh
UECue3xSq8eFw3V9/WDS7pTn/KWUVxx6KTo0lqCOOY3xpd3GDEfESKgrPdeUUNkgy963KtsG++uW
0fue3yZqmZLLCp+8KsiXs6OxYcj/gOuUv9JUKJu83PIzEG0lxJVbW2I8RnwVRM0iMfoMK3Xnes1k
LvdK7Yay+jZPC7qvsS06p7I+RwBeMZ3r1tgw0YClT+SYqvGpjgpWBLcfArWHLCqmvPc8agiAl0Mj
ZpXMXgn2zKYHUOPy1tePIKe1aUmtz6tLdhG7CNlJd69K4nhncKvvEbnqyTUtLlJayWPiYiHvvHvy
jWg2lCaahz26Gz/Yfjglj76DjzXzJUy76H4d4iCxm8vdgKDf0Pw9HFALJiAYWIFRo3HOjihskYvS
32Dx+Y3UcJkPnd9zFYn81bWbS5YnQUmdmbxfIehK1fqyOHI92rtqGGdvixqgqZU9s+iU385qvXXq
xK9lTcncJXSXZwD7v7UFe/l5T3Mv9Co5V3QVT7bn/WSIbYtMQinDEx1yWckG/B3Ja2K/Y4Ys2klZ
K7y8BNy/D79GceL6nLPzNRWuqak05StDVQapnwB8L7lt16e/vQH8XmFUBz7ew6LsnNTSN9uYoao7
BJoq5E2oZ8Za/1if8lqZcv1DQxaviFnVBfZRQt9yJOZS0h9r7jdvd45r78jymOaavh0mgkXNNZTe
20yoPwZTo6AtXUPMPrAVZMfMVMxifnSRvRPOQih3GHab/tWwHUHdPO1DTwxWd3p+WdGUY2ovcCqM
6F37iudBnZyXvwoZZ+vEg5+qyAmPrNB+orbg6DjOpoSbhUFTb1YVGR/3l+1W0hYC7PgDTYQDc4mX
PHKPOF1RcemRlUu4wSpnIPfqfPdJAIMcust+e3BVfCTOKgcTDjrydA+g/owTsq+VVlwsWi28huvs
iDKnMlJKCcg476T7Na2hFNz+AOcshJkSwBCioM8jBZijkgTS7WTEgJk5AmPi7VU+T3RiEaGLR5Ro
6Z0gDSHTjO5ojEivRAGk32uQurBo6TfA9DzIEMYxTPTpXrak+R9JgHZxpEr06FoQterIhlLuhaDi
/mS0elT0uu91AzwTrP0c84YRdoOHRYREPmwIJaq3XyZf06S6dD8J3+0iFp4PlGSqw0G6XOMfHzk6
Q2R3oX6sluPR1dBlTtVQ5kKDYJY0yk83kmsGsTKO7x8nqJeO7K4rX7WMwQqvj+hK0vHod5qJSqzb
vP6qM+TnfXajRwZbxDKFoV+YgbLaZfraOVWsw1o0O172aMtQvFtKhLikVUuua4t788KXA9UT0CUu
iLi/P7vvxFg4BOleC78vdj3D3dQl/6Y+mxqtr33cgd/sjvVNAKE6eeQSh/I3TGae/vPnOKrwy26R
yUDGizwwJQew7Y3ogQC0PjXXERagwVZeNb83G8YIVEm99ElIECXLEJRPhzujcFt9SyZwSBh/Z4s9
YK0KEa/T3euhA56Tfbrb1WhwMBxNV81od8/lOK/g671+grrNmlNlZLP0VdA+4TaJ3e3uUtBupPqE
LL7rmviq5JZOna9to/64MP9TlcuodBv6AJ04JIlo5k3nSnFuGM5hm5rVMpsQ06jJD1n8N4r+Sgyv
k7hPM7OkJPADRK/SWdtAZMQK9bjZXNquEm1keV1hIC49DKAaBZCUE9ihXOeuuAfu/NvEfeNRp1zh
5b22pCL4DeT5uoKrgxsCMNm8k6vlYj4nh1+FFtpu6dOGeyONqs0K0aCcdz60j6juqvgRXitadCHB
LU2P6UfgIU/jR2/IpYFyKBgDDyBVKyesyLvUd575Q4+dKr4uh/ZrUlWIZZi/gUnoZ7y+iWDRIiVf
6i0d1623xSITnPKVEUqQNiWzEUBhqPNP62hyhm8qCECXY6NPy3njczDx5D74rRymhduBhfjldsxM
NKq5+bSH2K2XoJXHKH1mqEXcv6vd7kqI09cQYAC9rUAqE/N3X0FKqDEm2IOh64PGg6jXEI7gum9B
ZyYXe2vLtNQ2fNZAA7GbKCjaZJz+9rOPFQLbtS758b16iyyWqHwmUA8oTVwAUJBkSsRap1+hbda0
5oR1AaJPszufFo9Tg9WqSYbzLDGDYOgQnCHWkLtok3nNWX9mI9XLRdCcG4wK5riNeN5nMvMsEv32
QNVqFNuLVQCxP+XZDdvGSfMcjPTm/yOM7Cso1OmnmwBBPQxwLkcPFjP03qcZHwQQWRPRpJc4yCWd
frfqk6+9f5At4arUT/8QNUND4CnOlP1xnYXC1QXSgyBaZ7KFuGGgScSb9In1kkuKhXVGEf7rKO3d
H768YAF6kKOmoFOt3h1mEt5dO5fe2Tqbi2MA6uezCdRtQ4mUnoHIF9fL1bDGoGTyUcN6xJYfHcbe
3Fwbp8BZiwaj6rXnKdjvUEd7XipCy5L385s5yGzmJuFaSmnzgiEvqI6pa7OgB5+Tg2QLZSewOh1f
UC36wrDZkq00nr5RRQ6d6+B7bV9IUc6XNtjVAziL4pJqnUp6+TzIuWvgJX8TraDuSE8eYcq9TwiY
2pBNrQgR5BNSJF2P837FfAmld2ovQOFweBZrR0pVYCDlzad38Su8hWNn/3TcS6tour8XQAIx1YVJ
5A65Mp5LnV+NzySiaAhjQyH22z1I9EjkTifMJ+rKK5dChP/P6rHmLhTB8DROb0nrrkBn08C2ZL83
pqBtt7BOveU6xnaSmkzMrndTDqMdlnO00FajZobYSnBv/LrK+sw41c2MgFKJG3A3l6Wgc65xlo/l
xIx9IFI5mEfkbX4JYjmyEQ/AQaQClfWB7Ap/zdwQmdD3ZlYy1smU9HpF2waHJsUuWkbTxjAkUoou
53yWzTDM/433Zj2vvMERRgy7V9RiI9YBrZVi/fgjI5KpHcCft/bc7YsuBz11DTvcGBeIkbB1QywT
xWzytD6j9BGEzC3cXBDQ8q+MuBluWhMVaR59oUIgSXt6qiU7CS4ajks+wfzjivrtb0TN2cK9V+Mm
yBMjFbdjxedUeSM+OH/iOenyHrkwcGLWh4XokEZub9BozkQm25vAYBH7dK2DggHn+FZwMiTgC6wC
Okuat2QveV7RFj6o3sgMI2EDyF11Hl7q1uMmudl663j5kt1tyLsgjABcXLXTjTOnJMT5ZqmEPVBf
F6kPEspWjBO0E0pUFu/bnBael+r0qtRdCWZOePdkxd64ESXSIMqTZJEo4GPUQ8LQKmZxWyDie8Cn
fhA3kTj8mnobkvoTPA60ZtJQu7lQaSESPxoKzDhTZyxoPp/R+x42JviU/KwZ4qNoySNoTDVRG4fR
ndI3aOmTnIPqPB4ido9dSRDQZ/VgrMTGAoGSlaef9wdrYMtg/jyxHvETDIlQ+SSrzcWT+dgN3kRE
Nok8xXkxhrltJNePkzd7UM/y/LZViB7UduoLzPs/VoZafd16shlDSLQGKlMGGcr73Cw1T18BZ4eu
BRQLIvZ56qzD6plbEFhUreuMCiko2FO0ggasY4KuJ+OsB5JFoABA3YLAJOdTV2uMRdaSkJxhzg1+
u/2ENu9oYWHJdfUZSQ7OVIqVAq4o8NmOT5QNMmySYhKQqlLTpyHhisO74eR5t1MFIuHUQgBPULez
YECi0hBsNW7T7+aZSXOoQ42+3mBQLiBlbNv6A9SBcq+VL0e3EcjE6FX86jwmpQqfVhJ8An6dkWlQ
EXeJQ0g/DTK03cpL4NTUN3H41jQX5dXiK+QM68bO5YHWnIuWD9U+X3kc55OKT85RZUWswyKk6grb
R6qVBV32mgmwxeFqadwxAF2DY5uY9KzsEADeSPQvxlCrfBTwxBG9OJCZnb3OoFsFl5MW236NIJZ9
3/I6OLnXeO08HzfzPWET9vfWDVYBOUYym8j+s4Qfu4V5gmGx8OlNeAh7YqpI25lltBlqTN+014iK
XowU10xxX1zG+vsFuvZ5IV9TV4kaFo/n4AeW1GX/2qhzt0jb/+dQAwGlkuBfkgftvoOpR/vPdkHr
Qx4GHiCtCOOsQdUwBkA3Xv7tTN4GtKrmZXToLonHI6MCJFtx6+ffwPLQzH1btomUREg5a8cd/Dde
2hz/odBZ7ZV8gSiHRk/yGnasy4NOE16WUi0+QkkB3AfA0mNi2u5e+uGqB1FRWiSKhe9lQnR2cvQ2
r599Pt2wPe6zgAL5WAfFKCmK4NfzheLDOfU+WdohxI0qDeE1Oj3ucaT7XG0VoksdppiOMK7nuhQE
LXDtqMcbBYrzCZXW2Jxv/ib0++bwHM80xinA/esL2vsC8yeZwstikZZ0NuePnEf34teyNEdwQKzY
HsqL2Reskm34XvDUAvJZZIT2+J1EbY8sI27jgth/0I4Rt81DTAnKQE76YJM7t6InLx2bm6b6ErBv
+u7OyNMGhDsk2uGvI4SR1UzbHFBxmhINTAAWat78uNBg8N+KjTdLexId4ant1E5saWagfiMA/0Lr
IBQBw67Fd1f647/e8c/0QgJ1oqx8DmRyXbj/TRDvdsKu8uqaq/5FzghJIWaJq2WGPgktpemW4N5i
XTbsNNRJFXicCwQ+5i74y5QmAX1lvLGWqzo1TVb42qITJ5xRz9d6UbXmoaRQ0gEEcW3CU/2LMOh9
5FvwyqxkDfvuIghVTPIMo5WlREWpTzUyjLdKIyYkGTRlDlWVK4USuX+SehzLPKCu0ruHIGdvxelb
6TVOZabA+jUIX2BDzDWOGg5KMMSoClrmtTSXU0+12jolg2Bs6f4lOTxanr8870Q0bTnvecCzJsA/
H423fsTsrk+GlGfOsqMhYA9WpO6r2a1EdRLLf2xqrIpf1t22VoHzW0mcDmm5AuZp1HWJrApvfsZw
nLwmZms8VjIkZw9ddZvYU+rowpziHHRV//cASuFiADkLY0OZEtvbp1A+Dq7r1OoclQAG5oN4Lj5U
VMUdXXLrDFoS51YEPmO4Xa/ye0FuVHA2kH69d6sq1/JOyQQKKnBM0VkvZmGVc30omENOzjLECwPR
dcJIqMACR1yTT5KDug0KMW2xGwjgm7uNXkkfB/DkrY7gVbTKjzNZ3uWlATV0OIQH3bHb2hBEdzCT
NAPwFuBpPkBEchsMJnhtdG1g4/jeNR0LUTvORHmxb1aTLTgoHRXFVpl87aq1Y1vqTLgI57aKEO2t
/Cd8oomS3kp4NC+iN+fTq4ub5xzvsmXnQAtCESJjxlTXUYrFVTL2DboFxk9Fw8Ro6+ALiyIaqIzm
5CvtiVzTAw9g43f+TUVePYUbRiX750NmyiKPq2RXP2Qv3QlZbqli4dikGakIXqaVuCw49Yalydrh
FWTVtKEIPGi/uAibBXd5j/hZmthACbiEWlMRNOyE/sHZk3exUlK/gVaYF6SGBfWrc3TzS6+Z64+L
naoVtuPHJoFOun/mIDqI4cQw2upSCuOdbhcEIkBvRKhiZYs4I+olx1L1Mp//yVjEppAMxwDgn7fA
DO411KLJ6u3Z/+b8FF7/bp0d1sU1Fowc6A9Tz8j7iq1C2WPyhpwq2LmqiMgnGzn7L6uFWYLM7VIB
7mqPX/ADY+2WqPY/erRPFI5njpssxxYoFYyJWPgAp5i2S1fe3uEMx0Awl5cBzfesTDad9hduGvEt
qwVw0/c9TnoBeoVoZJfsEnIkFYw6nJcbH6efJGucOaU5FTNp9v8+M9etq7rm1zdmHeJRMk32/7YY
1MDpRelBbDIXpiBJFuSO0iZXFCCr6fm2o5fQZ3sbXS1TQiDgAz0sa1r8pIo2zfpFKrenCt/2MNQD
mZWe5cmgaO91EAzp6sI83n0X7nQgvt+A041pRctxY2bL8yPgvy0ZWLcZtTB0f5FyA5Yaaf8XD1h8
pKKuACsEO8WvyKX0dRVWL2DIxyDl1yfUwTzbPaBLYp7MIRltr3fJ0bYF4f7RTMcsyaJWl/Y8AtNc
hwA8efIfz4wnUftr3gmrCcl/DaixJlhlcdZacBU/U8lme8jtjWWVrvmb+7r9+cr5Nv2+E6wcX1MJ
3D7AR0K2g+0HpycmQSstkel1SM2B3zjhoAPykL/hsX344CZD82KL3QDew/1JQ9vmwA8dQKUhUo2W
CjmnGXrhjr5PrTWW3xXSxOiV3zdN/J3B09eF82cKkA3EcH7xsbGIw9hLXpJnx1LsBGwBFN8KEcLz
gDMcj5XMfk7OLkqJnLkpIPHLNq0zJbGmxUTZkHZodrAqgdL8Su7MAzVE7a7Qv4nL6Kg4S+TAaLdz
NhJaEBQuH3ecs62pX2A9nNXKj5o7DdzvUrxEsPd7fTqKJdy6Aj0AO/YTcH6STn/So8NghW/rreUu
YXtSFtrHb8ISxjSuoBBCQ9NfRpDTz25pNy1JNvxsSfOF16asO1mABzJ2+vNlGhpolCr0zomFR2vo
+0FdGwxiQyLvhIIMcTGYsM+Teefy8QDVW3SjNl8+08WYXqMYyJqmclMZTmmPxQsDaQR2eWOoxXq3
tq8k/SDLuAfcbkBr2lTbskS4wX+b+6SXTn0qlbpyj1WE/bgT66J6xJGdyMvOR9IQc5oNhcYbaIRk
KYwOvMO7Fe8mif1pJ5MsYLDCvdg9Qu1eXLz4EG00g0vJ34O99dhwk+ECJ1rPYMaKIL0hnHfJOd9V
EkJNKPFbelJsQQXIof5rYHlY6pk0AXRZstRGSNekVjHuJjMMFa7ZOTD7fA0+PhBy7PpqvBYKx5YK
phdai4lw/pBwb+v+Osl9YfTbwo/pLPd7vOkJs7wL52/zDffSl8iRF4aR8A/G4zHyKdf+d9Kq5DoW
iQOHLS4Bvu2N+SLfHBJm6IPujlPlGNqgC6L035vqtsMIxgnsW3p0bUilOMtxoZ9zI7eDd4Png4Tz
5h+DQeB3EwjGRl41ClNK6++IxK1k9HsyiueJfaGG7S+uCL/zklaG6/coIzdTDJua0DCfPKc7l330
FYW3cvwAVtgNOubWcGMRGt+MNS8S8MClxiYuIW+aaeSTfoBJvQ1v4UEgvzGzM3Bx/Oyl/34RT/rU
xLPS6vvIeICuWNmOo1kYvW/GmwNlhfWx1Ag8F7bUIP8i904x92AgEhD7I3ajAx5ix8s4MnzVjvOd
8ubrrG80js2qdwrMZQcdz+/+ElhQVmwxU9yLbk7ubWMI9vjAXIGuXiZiA9ci2L5ccP2I/vFKTOnC
+28KfRlwwtTk1mOepFvnQTXCXfiqZtCFbBerL0j9oOiKp2XORQIGwhT2ZhttbM3R39vVGViEnu1V
pqbdMcvuxGIa0TWyTOrBGuBOUe8sQHU6jtPbqjIJuQB5mQX7dZ2efj79SUybTsVEW8I9KBg4BzXm
HDXqqVa5bZeQZzVGopFwHZ9SzzfNMnUatCFJjU2/xL56+rnm4P5kwHE59yhS90FyEKOcezAZyPZ/
m8VGqyPp6lE2/kl9PtlpBTcqyePqGD9wDCI/u3joYSoVgm3ZGPnhbU2KKQ+zUou2UMdNS5BFSOhk
s7jygdgNQmcFS7PpiTdQrfH0yDwczUBmu887zjq4EdY76Tv5x3AJDiLkENa8la+Tl3E4DE06q0gZ
uxMrYpZltbK37H4Ex7RvwqJ2MBzAjyTERPTV8TO1OZ+l386V+tlc9dt42FEjNfpVEZGKzrTQ1OJN
6uxMI/+f6a4IXa9mktsAGjDOtkaQF2etKPrq+Mndj5AoTK8fahnuEoZPJHkGK9Wy9iJFoWavgsCe
onTCOvnnnt5/fOTy3mcddd5drYyF3N9oXjBksRECsRoXC08t50OQA5aWTwexNTODVbqNTlUW9v9L
vyZAfj6/K1noypp2zo82D3NqrGhx6afUsFZEfFfl9qxm1anDdhpXFRg2XMvhs4pxo0hrMlpYQOUx
tpvkOAyej25vp+i+ngqsi1eXFPE1K5IZ1fNaSKm36+JHdsvYT6uFV33RdUR4aXpapSpYTTZ25Ni7
EfzrCNCaKz+D1yf8hAzmR4P7IvEglaxKzscVI0ZCFFuwaw8j2Egf62zV5PUSA6MpgLpvfsWI7gho
1V3WF8LGdXyaHKQsvTr2twFcQkVaX7cYJ5wF/lL/GMTHE+ItXosZz2phm4Ssu34eU11SCheXkvXF
4zMhuTYgEtQetXXWG11KELsddo6xJSGJK3lNxWAPERJ+eNA8EW51+bDH/mrAah1IkHH71amSoArf
rKOSusyX5wwU48/II4JFVCtiQ3I5Xiw5evBJbjjSR6EMrym7stP3Jzt4LqX0+qlK+jm1c3NhXrIc
ZPkUyhqQzvrz3JUJ1va0+S9c2a2C5xfFVqxwmv0mthIjnLBYa3at/Ns/h+91jD+hrMaGDyvoc0cC
Je79+Hxv5RL+Ofg8W6oxqbPJlwCgpqBm9EVyqS4YzXjZOGhhWlo6CBqL2bRS6Aqvp8uJOUF+gMhU
7o9TkdRndh6/Niw2Jvy6u1SKH9E0QZ+fLaUiOWA1y+NF1BbL0jVEDO+I5ViKQr26EtVI+q0zWsKv
DrQYcYkPmtHfklsWB96YapM4uIKoFKLH+Nnj0qGByntWtVAA+58hozn/QrgvJ872y1UTfYsBmO65
0DWPiF5Wf7DoO/Lf09opE/kkPEieE5H2LdnOm3jCIpZT68vCtgGNN2vr3xnajJrrevYFAHKffuk4
eEDmJUVxCVXavLOgqBuZrgVec6EOBASUkIoZdpwbiiX3zL+RV1f/SeOkQw/S5KdPFUV8lUuOMG4n
1KhBRFcs0bLz2013hpZq55MUWOwS6SfBIs9rsdiF6ncyG0fn2IC1u1b6CdBXGw2RGhW4Yvo1tykH
lR8ElBItVPI8QbjVoxHYen4kZaTt1uPNErC/QMbKiWaY3xPaMGOZgevLSUTh+YsklEBHni9rWEXW
c+Z2VLhCFd2x/ZZqfQmKDuJxnFcgpFWvFYl9jKIrkvUJnhv37aWb1AqKWoVgJ4BYrSRH6S032X6C
JaRqIxRSzoCaZnG6QCBI9vLR0v9afp5SdX/wX1o/M9b/SiET3gy1dcX4PX+nOM9Q58E8xl+wiRCE
FmK0IwptSMusHqJh5TC2d/iBoSBl2NX4MFhWOh8KBaBQToiveY5xF7IQtESJcKer1Mb4jgSdjNBa
yoFDqP6pavHJyRHjodOWLKDGtQ7UP6tAD1LvWRIs49VukYEVllRMsRWA/14i6ED28P/9RBk/c+XC
LF7w8kdwOqxire6gXyTKn2/K1WA9uau0rwgflAG79iCoucEi/ewlirAZ472HGcam6PrjJQTHcfNY
YnYMAWZhvp+l4N++vynKiTu/hOQb3TWLcH+YTzv3nU/JXffb1kPLpdPHOB+eGhQix2yk/qfqi3lG
muidKT1VppL8LFupO1Ji70wkk5xBDbbZSPPbBkfQjB9tgQn1OC8DG2V4XbYuP28BDgV2Giko1XA2
fZ8Mni4QO3R/VFTFz12ZWUtmbjrDmO9cfpdl1u5wd2eUXeikmc6wi38fTNdZs5KQHy4yd0lsDP5a
Ui7fakxwXy6oxcfuadXiY3CxSALzPzYWkxIH0ncV7eHzzBwizgzn3H4fyPPNqJq/NlqN33H5tETD
+SPCdv+VbVZBJHIs+23bxdkRuXuls1EPILETcgyYU148FI6FYmA0VN49OAVonX3PDGfuHZ9xH9Fd
huX+2RffK2iDz+lObGTVwG7/ykivisEJOZ1w1Qi0aPtZub1idNga4TgkwyqImzVmwuTECe6qGXps
+RCFQyLIjqpCNtAVkS7UEBkg01I9I4XGsPEbR+1qOg8zZNZBEHb2O34vV9mkQ8edVr7Udzw2qg4M
CNO61iWwkpKopQZSBtPYE0J1EcFA8ewrbA0uPhPk+qufzvHRRCf2PLu3fJ9UBg+ex2iLzVBntLQ3
HpCZ+IuUwbLvEnVcDX6PA88w4cBQmkHM68kQklH41dCVFONCghZBbLon8YMDjxrBbflIpLDRfQmN
4pOxKFeiUGyzwCwadNeh9Kp9OQ1TDxio/qCyU02fUpM/ieCeMiG3xPhMxPfKZGStWJwbcqj7V5ed
g6Y7P0YaWLzeYFXvJaEG7vGmUPXidZhcKYd6I9jdSxNPBiKux3EFGolDQGReqa+xEWk99PNL/Dl9
vzDoi9ws8t4H+gvX7fuqf/03s/7i7v/MwkoY4F+QHG8dqzgOXtqnZI4ywoD+4+Qli45A8bSmcWc2
tPufroSQIl3BSLhcIWtZiDfY4o30NiryBD/Uz2GjIhr9Xj/wWzTa6gc7mhdbLyR8/0KMg4q9DFYJ
DFEW7EguEcshn5hYKXMIyuTAtKdWoZ+pqu9PR1hLR2u5wtUjPjYlZ/jy4UNCTLP2zJ4KAtq5Whyn
IYUXj2ppa3KrHSwtDd/DAKRC6m8NOEVtTX1uPdXW0JS5l0mATxyu1KLe9BP3YmUomJc56mDvrOmt
s6TyA2JKe392GXqyLzR0LZ9J69HoDjiq7LOXUOtY4tdvNll0l+WqyINu3A1f8i8KHE8wyxt6Qlra
EMIXZzPHyaCJV/nt09RUazE83ZLrbJ/Ed11DvcJSfPVy0dVpZJxwViolXJwSfBKtMPlGp0ZTNOVn
Y8qa28uZtra7TXkdUg/p25Qq275rC/nygUjUytQ3MeFFLLGwP5mUDAbNb7m+gTT78BXmpx1D+fbW
nz1OLwO23T/s5n4CCnrLquED/WTSj5b6zpfejwh+pgMxLGwnXWd9jbNUvjM2cbiYv3hq0ghyfVq1
kRCZYKnmyg8iglERJP04xMt6xpFjXoN2nZnyd9+8JOc0AXOQOic/KFrgvyHDWoM5vRaULZljFPV4
Xc4tIoM6TLA87xEIQJR0N1eAqoiURNiTKlcreAgoMG9GhMTVOHE4aBazkSvXXvbkz6r9W0gbQ9m9
sV+mIKiYIXrywa/vBEVrJUVCFfAZVrrLRTUouvoT+GK65eNBPhEcFJIl+VIZY0tkEuuckzvRQtBh
lOY+i3h1eUcrq6DDU3EMVCMmXsGr90l95c90Zt/E5yJBWhV1ON9myzX8P/bKfcHHWR+0ANbpv3/b
Ffp0uKt2VkPQ85fitP779ubZkbSf0N4uEeQK+wOxPimG96vTBBuWiDnAyVZQsMNax2dcVzWSYYkg
M3DA8ekSTewyM2EszgwLmCB02x3w2U8ZXrOjazBp6NurGtR0bXgTkLP8emOtZyBhGx0Kc8vFJObw
evhyJWC0ncdFrKx4ic0GUyk8LrXH+eWLXSRyxQOtkvlowJtF1tsD3RA0CvMaPiSOQxFyPXw3Y1+Z
ShZ7KAnhakYJPBMtrIZoaaK013Yywae2BvNMVD2pVCKX4kvjOw+8hzd+TgfK1pE6YLpTlRw2rnPG
E+2k8jrxCPfPi2CT1aU6rC7Hr5/c+PKXhRxZAH5Xn5LEBIenrcksEuhZ8/rv70p/05siXQb7E3Im
AHBf6GVznHKHfEqfRC2+HOBwEwN1+JR+zfx3TbX9Lvey+T2NcpGZY6rsQilmOb3pzvILdqrCEHua
fjhrHB0mRrITpQuYXSZn1QcRwJ3okC8OiQXKNC/j3SVRSjx5AyeA8UfhfnUYAZ+I0duu51Y6lR+S
fWpXBkVla4IupF6zteHbZM15XcFaca1fibrjMRT8OuqcTOWkZpo+LnJzHnepgczPf//BJk+xv94e
3MYz+yP1SLLVRk/N+0xJPtmp+X3d2AT1N86jgAvsC1v/qFs0b8WxOqk8+Ra3paevL+ZDff1WLRjd
9eaT9vtJmRxj36cFobQLyajNguY//Z3DSKTDwDFAoXVUNFjZmrkrLL1VsEHNF1hCQN7r1VXdYXns
ADU37jyj3BTjNUahlpIdEfMe7mXP8HZlw5u1ODjEVUarge5gCwcvsLRJFXSyEwX/gvr6uUqxSEQM
er/kNxckfslRweevf6KBH9UXBFhI/P2QzFF4gGf7e2a2IJ1fj1pkZiRb3sjkp220ycrMV3QXR13b
MW6jAPL8vTrhLLOXbR/HvNM609gDeC+977AtOFPV7RQTGc2bPFUBH9cqv5fZPlCes0QAjldZREAD
ZYNw01GBXuSaV1G5Xqpfpuose0sgFHjLsrlpqSDxbrKWUYDn11vwYahwZ4Qc0ShjIsCtxg0MBpS2
dKuSnOOJEY+40t2Tu0v4XmShFrJ12yeCOzyswGgU6LWqCGjsK2i4rIZHkOjonSNE5O4GCTgDPrJt
CLgdpcmrlJObJQJkIA7PV4oxw4GWmicaz9YAaHxFNXRL6wV01+8cesqgY0COE7pj3aVs3u44uV57
2At8qcUUsMk9oAh58DBpsAGEcXzTMbDetScHCmarB5Fzv2+zh9XZgw0GqSmzKW2BUSl8vaBKyzE7
w3YZir0PBWm88QW4yumIWjT7zyd08KEonevRJXtnd8C0ilo6kF3nwseyz+zMRPCfeeZbU04n2nfM
8Xqyya6f9SQySzZKXzHfUjSs5FA9COeADC1RxYQNAZVXIn8yRgb2MbY1h7zKj0fEfmhbxiB7Ye9L
O///DfgIp5yC7xk/P3zr4voSlKekFDkcoa7Io+5PxOyN+jA2IF5yOUn3DTt5xSAbkqPzUCS6mR+L
K3yi1W14g7LGDa5jglT1V5lT0w3kmqtvp5i6Iz+NiddXXqVfpv2Oh0l812zIOh9Jxk6MTYC+HA0i
XN1f3g8R3KNrqaJoAIa2UhUB20oAWIRSqnpAbvVgkPETQRZ/y+zJc2/VwGAK5lR3hmneEs81dNBB
xEd3rt7/EUOWWplU/l40CEM7AbfUi/jL6Fs+MXmz6iP0BiBN/ONWV7uUOKre1ypUpbXQKgvFwfbT
sLR22UEK2RnhEMzVkWRhqpzwtq0Nri5zP7oE1UF7m+niDkIAJGicxZkhYhK4vQUnp5MbRXl7sv8m
cMJ3RR5XQYk/AGqVnl6Z6cjnivzbQypj9R2uFWiYyBT3CacyJtBq1ToDD6lULJTLrQdRWEvQQREr
vn20TyS41reRhRpP8Jd7tD9idb4oH8TITXH4f+GkdTJ28ZNQjwU2JrZiquADuUcWPz2xaPKWkzHV
EM7YNkkcfYMH188FmAlcLuRl/lpcuxzPu5wCZcDC8XdrPXHKOUzSrpd8sR9fW3tIOPHw6k0dxji7
05GSv/7P7sIssuiv7UCujgCrn7FML9htehDR9MansM2K4PlzA/1V37ugdypJWVL7OpEnAK6S+Y0g
9fwWLeXyC0R8weW2CIJAjyoSpH6iMmNWa4PEBRLyNVwXMCzav1CYvsuly2CA+w+51zJupYkEcLT6
J6ngOD42ZX2YWuK6FWm4EaCQ4wcaN4d8X0159kpC+qmK8Pv44rjj4K5t7zOBNLXDykb+IQcZM9qL
GUC+ZhB19KDxDQU7iE2pxTEgtRQoelb/hzUQiB3B5LdRuz4apYBCzOV5fhnmI0HUDZkDb5mScDuh
tfWFhf0LPzLyAKdB6A3XdCdNMaZzJkOroLR9JvIKfvpp2XHZ4BQWiK2BWXHZN6YECsmwvH5e6QCB
6vSONN4nCbjfBdA726MzAJCLcs+ycXAbyjipImCqyvuWw4crqcTHkJFY8Ld3xSGarWHlGCA8zG2a
cXsQdZlsDWPp4HX2JDAqR67Sb0xGHqVwx6sP/UE/X7GajX8DisfrG7GG4/y9XrlyM6vwu43A3DsL
Kb/1b2pVjfLEW/I0ZJvMx0RcnhO3jqV+pT4Y6E+Lf2AQHzeBEVTN0zimlBG4SuxzlpE17Hgi4h/d
jyyfgq5221CXBhgZlRXwGvacM222ogW0xr5bDpgQ7/fHwuCqqoWHWIjdMl1Wl4AntG4r18ZaHdPX
fbPTJ2lKv7hSFROOcLVq4IGeqmX16lt4HHHWtXSnY4upAqBjebCuOm1nkGlhLot1Bxw0grI2kz2L
aRF6o0eS1Mva6GALhhBqQq2fEN6suxnQezRLZlfyj0cMDQC/jO/U7Rh6IfDPzxMT6R9ZdCzHpfq6
nEa9tRGcgMZoUYAE7tb1N9g8Zd+/pajlDdZuUOeSNBRsZAG+e3tuehro16x8exQPkNXFdeP8bMXG
xRodjirY8jLQ1cz99Hou5dr/2p99oajJYKkt/I4hrhjS+6xSkw04fIAMIYzHfOeHpusCTxqHiM3X
IG3uapD5clcU+sgueqlJ4+jvbYtDkuAcm8bw2d/RpAMBoRm6w6Oc9BToy/YQGPlyEiyhHg5HJoAx
+QnCZqlloCF3nJYxeJzJzmF5VA9TT+NbO4psKFy+8BfooOppNLcvASOlpnDxwRPsvQ8MKQ+B1NTp
4LGd2YnJ0vkTxmWlyYcpi5PjjiwD1Fn3M7UnV7afnLY5Od+A6JP9jgg5X56cJD6ueUoF4W+R2Q3K
3g0rb5kRv+yJb+iT/onP1J2JvH30JbDS99sPrGJZycjCI23ge4A6vhUG80nfDcmf7dYGW4AS5mkW
tChm7iTtKfFNK5hegqddeII12rG3emzvmso6C2n7Csd/QQUHymNaUQOscca+OjATpb58G/cPqApF
4wQOHnfztk7qAADGwtlah8pGH5wgIVQtWgNpoQ0Xy6b9FlC/X0crUa5xrwxQ6lGJkqHheFva8TOf
nIhiYksjfpqI2R8IkmSnYZWCtukvJAm2gsVw7orWVdtbXR4anVpjgLT0G+gDgz8IVxYkOsb9z+Kj
9c0YPniI9Qp+eUg1NGlijg1YDNB4adV4ZNrbC2UPAlGYwM92FEcN1p7rcE7CJsBExGQAS7TRH66+
xbEx/KkXgnfclGZc3wBMTZIlax5ie0mPfD43zTD52xqzakgzCuFZHgzBxJxQTj+nLpaQhivstmbb
E92/OlgydXkV2qnykCEAJnnGj+IksVroyTNRQomkMntFLZ4i7CeHcDxfowsHA/XZh3ggZC6Wg0L/
cRtCb1ANu4XdtK/fFPWK6pj16D7QwTdtFhNBiIwxfZ4hNpnpaJ4VC+rVjelbBx6dlx68C4kbt1tL
ceitXIxcPaAk5DkADpj55XfLDaDGdR+sXiiaFz2t8qFTQYs0Y6YbmwqgDLouKVvAC4SNkzREBH9L
j7AUNuXyWRwblE/p+hjYoaVU/2XGVZ9CsTIkLzMKRrsijB/+Y46XGrumgC4nxtmCZVI/cyXGRx8H
NlNPBxbQi5YvXVIMqF5Lu77VDU5/dl5yCES4kyjinhx0SNlMu4e78DZO5DFkT3m+Y5SEsB0uUfFN
MWnTpVDbhcodCh7yq/M5VOR/TR+yl8r7mPo1NqM7qwu/Dk6wK97uwY9/XEtFatcFAlQeb5UmiR7O
crLnVRMTjkdTPLXIpT1VqGNp6tkSCje+FDZwXsZ0kSvtkc+gCF0MNP5bGUSLCfP5tt9h8b8RJO6k
7lTOH3vzyPZvNQfsEfCq/nDRI+eA3HZxw7GE++GCRf7RvM8LxAP89xfXGFmctJtkHTw/NDDSA95E
IgdB56uCAhFSRzgMX1Vwgkp8qvvjHi8xyRa2rNeZGce6Rwih3bTZURt0ieEbfc3YR8vzHAbrpmis
sLevm8Rfmr+poFedgmLf3pPdiJPCyO4DbdV3XnnN9ab36IIF9i9/KTPM0CTG6aVJB492De3AtShz
QyUmt4FJemUt6mCWjRdo3Nv/TpQudt3MRgsZHz9c+xrdN28nnLa0hhGoz4Lpat/IMIngSDbl8D7U
rMTT/HcGIsXnUXmX33nJkxt3Qp1p9/3oOaGpMKYZaEKeDW/HLI7qOTvhotUILVH1xQodTXy2EfSS
+NJm+rl2jMWbvKOUTGL/O8BnjgcvnEi7rwUygGOXG3+jONiZL5aXRA4Xj/DY8IlHHcAFYxWsAVKi
esI0J35eH7cVEor1vY9yjqU/Do1r6EaiRDFaB1/k4qdz0I7alceXrHj9h4yTuWFbo57PyCURgdtQ
h9NqNwhrcePAchmyHQ2OjZFd523XIc1+tlyAAq+TJOtGjwfunMUS5PdcOr/k2jyi2viaysMvXW3Q
vAXE859lMPr2e1NW8SeMvHSS+AQzcOnRFDajzz8JYcz8BWuQ5g5tiaB+Vx9++teqPsufOt7kRgt6
zPENwNE3Zo8woJwKRAYXrGaDtfDGdEWLnU6OnY58yX0cTbjzEUw5FK0CEX6WiMlhZHZBblLAtUpR
m5xoyY7jopyoNB3Tyimc6W3SFoEcUaQrEzhiT5w/HiM4xg0pd8F2a99oXNkT6xxFNeB3Ivggs5p5
3gMYs1h+zFVrZ0/tkOBb27KINGpP5vbUF9bnviQerBQ/hbbiqgYIKnzsoxj3N1HQfcaV2+ziZIgI
wwKqZu6u8FnAJHKQYFuPWZJ8NNpzO2g60YNCV3gARlOS+XAXXfRGyxiiEfRjeKPZUU/3XpM1303A
+xB1xV+EVfRJcA+1rTbjut1Fgv06lp2vKTKSH3xjGQvPKPnVobuBX0CpemN2FYdnkRD/dINtbWWz
3uqDnJcGOMO16yBbLbWsEgNvJKhel9W6lNTduwp/LPDR+O7pXK9m6GZFJmqBr2ehWPQrEqxGQs9t
KAFm1MsGI7/DmolB75sWOudJRt+ofWhwqdZ4pV9ugDScpdxHi2u0v8wXDXN1cMEJLxW83H/t5Gcn
bibgrLB7RBtz+AyAOIWsR3vKaD4X9tms2riZzTdDfTZ5QvtYp+MgpFeFZcFh+S99zGIkFsq8qeqf
B2CPUsjUBDkYFtn6TAOzIyblM+kO1jIabJLdFbCLT4s1jw1en9zG4Lxb6NAPwRcn1gjG8qAYesVD
of0GweWnWojExb6umaVUgCXLJcRrkEPv+3WGNqlFNOFmBLMReJJgzNtH29zBU06rP5RbrkGtexcn
cou5JC9AWXzfBVRZjUCkBVjxshupQ3fEP3HIcVLhNNZ3xMFYq7/iRav8jP5Duds9vj34jfTsWM3r
liQTUWyqpj9nHenwTYitKDnZJB9EdumtDB4JX3TVx9MpnC0ObuDN2GQdsCTakhwUEdfsjHubRdSC
6BZikKK4hDG5FsGmxuLzI/8giWpRsEsBhWIWNJXhjnCDM6GoaDxCFQEHHoP0lYpqZSVcv13dAdSL
MEQ2mOVAaddTTmAvTiAGm53wGyQDfNT73FQ513tmDdB2LiSXUZgsQB1gbMHScwJBOdK2Og88ezcl
vZetrreya5VVnmbTc3u7NpNLirOc+i+ym2fRH51hCMdpX09naAoS3SzKKrI+gEeg3eWd1ARAv+W7
QLhlMkKOlQGr+FGRR2R6CMOkb3LiktnMJCqVnasnOPAisjlGN7MgvULyPQzNADixJbPIDcfJi+Bu
ALJeOJtl3Vq32yEonI2ixMnF1kM3hUTGfUkBIgDLnKNJ2cXWwsKIrrOO0WYfp2v9RR44YL+2m55C
J6wyQhbcC8hcaROnBzxiIf+blKY7t5DGIO4+zSaoWMEskR50EkyoXW8Nd9JLkyKO6h8PpXAZvo5D
wE9OR+1NsDdrLMp5lWspgoCyCyOG3KEMuUgllNnedzH06CpOgsOoulLUfFTwn2qpQ6UvT8BPdDLZ
KrXESwAkwB0RlXrCraO8TFpJoq6L2WmE486BgQoAgIYWdrrqS104ffSphALzZtwI7IXWe9gLg5bK
uHZaLC2NLZTLBMGb6I/byPvYSVUMcIGQzBomAhpM/xC3FF4NHO9c7VmP6pCsJbsaMVHMtxtpgTPZ
nSRtzRLHYn4XE+WAQMyBmRfg+zBYYavnaAtC15HMeI8QBHYKy5n4Y9SS+AEX34IeSu8y1wy6EEdu
UB0pGESpwSoYBtpPPwL35QG9aOQH3GUw1Z0AF3qdLcIiK4BQUzg469wx/KlGPE1vmYSeU2J1OBU7
Rxr3L2ge8SwDgEYW0u/i56UtjAoKOQ5EdGkh0ljhiAk5Cg2yymWtEAsO1zzc267D8UT/K2PXKbJR
MT2VMikqlXnlyZjLSsl55xUdzV12yYs8M3nhuvjJi93UkuEzRVkJeqK4CT20bv1ArvMGGiRh//Wz
75Lpvoh1BChJRMlA9bkTFYPiFdUFWzxc/34samvGaUpKAbX35Fz0MiSjzRNs3/2RdIqu2CFpG3s6
39vlz9XohZJVel1l6YYMwdK+v64wrmcM5vClzObsLxs/yFhRW2XTIFjvKQwgvUFvkzOrRdIMJMOe
LzrehUdiIXfQBZkg/NAI152jAmWyRXHcClQ4/oL0PcXFnq/I1IFZooflPzwZV8k0h+hs+Utgpp7O
FbK3jOlWJSNm2ek2Ucf9oSy/xZvyFj75QfRhfvJ0aB/TRdu3RVMivhRpp/Tk6T2OBLeE/42QoGn6
JBcoOZ1plx7I+3TiIE2oNwOA7xd1hwKKefdbsCeZm4ZacybaJnjxyXMnHzVRLlWe9waVGvCFGLF2
ggqWvzPl4eruZUBHyClI6eO+jYakqEH8Ue99EkD5do2Ea8785maYC76v1JmxTJVcGrFnAKnmu0ty
39PQVxmjBeKTzykeCEpsOb0o0nMLitdojvFgaqWpZUO76UpVrHAg6ehzyu/Pv6oaItfGe55JN8Sd
f4eSDP0GzEmeAMDoFf1vIbl2LWfYqS59zdx0fTXl2x9EiYRHx+V/fiy2OwqtBVXDvDE8B59Hq5at
PJxnK0rrzaOA/eeskRSeS1HSf9vmo+dAuQqKaOWAyp//w9juhxW7UeqlWStrUQXtOuePaf/0U+1L
LIlK5BweTD7XRpRqzdAHWypej78xx30IQ4LhzWsOJI7GaAlDj1qCOL6fFZSfpvHiBY8Peef59Aso
u8OghgJEfXlObTm7MmByjO8iJep5Gdg5w1hOOMtidTybFzqK5Gvet4A5a1W2VbI//duRqrgsADbz
USH2I4p1B1Q7AyC7ZSy1aMyu0VGbiB1oCnTKdBOpqHFzAhZSgS6BDFJomO/KcZHzUo1dYhH0Mc27
MH+v+yZlxfenNkTcTE8rJgtOHZtN+EoOsPtAFe00XnBRkaOjXjIVg9hHjo2OwR70+hlrmliD7akG
SkLu2D0Hi+mS9O59DX51IwEEsXYOqfgQcvNszWg+73LjPe1xUSRsWNl0tJH+mC8zBTV6Fb2HSAQ9
Q07hKJy9/gjvlrjNaiqbRJEcId+ILTylGYbT+vGtR+noYZzVwhQurgSIL0QV0hcM+UzmtEyXZjA2
ZxpX4bDpbCZvfCW5TjAx4snroNnXvih361FGe5kyRN3TtQOcv68uybHWtEtmtSu79VYMh3eOQvVD
ye7iH61G5arEpGnLElDVdAWBA2DlaPRIF/m7jxGr5tzParbB/CTgrXThIHGcTW+RUtB7FQni95Ur
1+jz/pvEoECCX69H4+IyRehS/Oll0V7YaXJ3Uh9mEubchXAswZWeLg7GvemLn6yHeswLDk2aCKUs
1/r30svGW40z7Wl/ltRjac+AEokgCr2dIHfYAGXglvhO2qiFWU5htaN/KjRUqXpi+cF1PXiVbuJG
bsjKTZPMSGzYcCsSdyDEfqC1WDez/k9lmFIagwLFVSi4CKZ86VjyYbbxhHGHAu+pxkvqf1rE9tOJ
65foDTqlnphcZFTdUTb85xTIdTpp6zZaxWA5DnpaHROnUs8IcaoWOJFbxUJOU0bIdyVNtmV1Zct7
9xNiQ52eWrvQOV7W+3W0BayhTuvxQM1ooGgKEKq231qw/0HDQGohf/CUVPpeuSDOtwfSfQ0o/F2y
qpEpCTRKJ2R4HGpTLz2msuY734tklA4YZpuBNDlp3uUSFx7oUfxbvFq5+1hRMRmk16QYmqzJiiU/
alakWHJIpypl+qWSEW3FZ9NB78AqUXaKNY6X7h5Mk/LE39T2L2A64hUJI/RUQoUgBF6RoKS3gym2
Xb1nbQlMeEtWevUGTJem2/xemx8YhvB7//XNaFJhcYvKYIZiyjBi3oigTQPhyKZ/FDuJPL1vJZSJ
yrBOjJGNcILCwax5CSl2pm9gNP7pGpi20hZqrRKjoEi1/u5V4Lw5kxbOgh3gwoD8j03AVHlLo6KN
2b79R0Y0qCdJs1JVFUfu1Y7Ot6eHa9A6KjUyqZ/qYvhrWyDRFgp4h+FOBcPo3wl70WhtkqNg6zir
J5043cX9yScrbrnUoObnJ3c65g4hr/Vmt6ZC4suHOZI5oxmD8s8o72EVzrIwmdDl4Rd0RsjvG7ub
9j2Rt6Amxj8TbZ4YalCXa1hNW5c/2ShXLKSAApOsNNJ7+1PjAS/JD66sZQNeYFoP8NgvA9/uIPcD
HLTmDq/rxiRBVMrz4PYtqyQ7zXH0qxBwplutAflhSouYJINXV8/wi8zc4sMWqLKyxXujxdCtuQUq
pkO9CwyCDSxZF77n62ATu/5o0pjb7wPFECYrCBpKIAJwXDpihHBS7nScBSebZc089SghG05djQD7
+XxsZx+5gt83QJm4WnG0kJtD3MLPoVy8G+CVaq5EmMOVCnaawELA75vxMCFqBF9+LRQgzpMO+QEH
id03XA87+H+Uvndp/8z9/pCV2xFjqoX3E2yGTus+0uCdOSPLed1IjugDHu+idR5WQHi0w3QVY1VQ
SmuPjV4SrOy93+NA7X97lq2SMtffd+6svA9NruIBmzoduMajtfTY4PoiNUGH1PX/ksEehHi2LSAJ
BH5slevpaNXYWU64l6vGTbejmYXB4HTkdRc7vsAwVKO+Lmsf5TCTz2SOYUGndswEzelXZu5Pd+dc
cIxEadWAQGH0HoztFTnSBS+8tkvrryE+g+7BshfyScLBpHYzzZj8NCIaxeBx9+IqQnhuczaJXoBA
d/HKj/rXT6wvPb3LvBLyjPg4kJPuKqQDYfWYCun3/ck5BTLNatX6QzZSWHf5Kcm5kFfb3+yPGO6x
QFGquRvYSReiB3l6RluTA5TVig8KsQcARWuxL+mDHCixZxkWKhsbGVOXquL9H6bfXJ/IvebABmfI
ssJHIUFqaCv4f1RgrmTJ6YW4Z4hLugbfxtCXXTUm/jmMYH1RLu0Mgtaa3ueLAVzHB2ZlnohNt8j0
8e5Nle0HlE0torjvpSbvjxkV6djhtnWpjk1g0XKgVXx1V+3bpBuLPBIFIMz4XBn24ARAxO02sLBO
NOh+oE1GuRRk2En04NLX+rKEYxSiNVtQlVPdWG/qOMKZlp69ZJRphPw0QBk1sY3AOF9hRcm8zars
xGxSStS8cv1qvSdXFofyc4tKr2pIi0ZLt8MebKB4PspuUeQfwezpxEWq3+cIHI2sZz59kp0BvWQJ
s2HA9XZH0rrrBH614OuD7OPwoTLSpj5Wu/t+YMarmLb6ys4g6+ClPiWMaPvCwbAvjEQGDlE/EIxp
Nl9ldSun7cLY58aKJQCAL7eu7/4mdi1b8/H9axGQiGYOUygPM8I6WRPH0pKoFnheFaO66lp3EJ7/
qdu43b3wq+zNcIqiD+ntrVk16W/V6xhWvxNMjgqSAPAtXz7IfJdHuxG69BnJIB/UMKks4krK+KrG
aBA2tSSUNMMUY22RdiFImWai7UmH4Xp8cDHV8ACKBiIyR2RR6rbZu+C7gaIk35Mn6RGkP/7oD8hX
xDBrnGyE21DgfkMDjAxF4WcZTkIaxtGaSS82lCYEcmbwpOMnt9D/6Q64kSbPzABT308cU9j6RoJi
6WIty/hzmIT5XvIVDnLOKO6iRs4eaQQiIEZVYNmNwSCt28hWqFVoM8YtagY0uND+NLii4dRFwQH3
ihlnGXyMdTq/GzXyEt53UhrOeAfJ51zlZ/V+cTn7vOta/WHn36C87J6yKSJnjqYAHQNfv5Tur8iD
H0rd2mVtfYQC7jwFdXajRWt78yjf/KHcNEfrTMTLr7nnn+VpdOvOozewprk199D+CugglwneASTg
mOr4G2Sm1uRiiZkhPbyHBQ1DSRGQLWJRtsTLs3k6ABBP6NqilY3BdTGOq9yogFawCzWvRaKuI/FS
YWdib2nyyd5GvhaYIki5gyIAu0Ptu0EA071SlRg6WjjjH+7j+Twhpf3IzrKTkU8/sstqZ8WQOCGz
+VI1r/SwdK5WPVelRzccGEk//CYZ1knG6xbsUIwIByOSzCPwUwp14saO/7Exi0tiuKGaoulibfi4
es0BIAHF2+0B4cuhXbDQnc3XkZ0+DDH+CqItLAud/fNz86xegBFEFI472UqoS+nhJ8pnuH61dKlY
FbB+4s9jWUnSxM2Y3XSqfwEI8H+LTd8+mfO5AWPZ2a+9zcttaNjBCUhPEUOcpCHz6bJjuT78MR6K
Nlh1vaNEDDrS4cxeJQpNZJfh1UyBmYJZ01M6dPm9fBL3x9UXuYKAg2wFYqVkay27TbpSHwzym1v2
z2q9CP5LcP02NYJ8BBo0IcA29948/sGs68IwI9aA65kV5WoPcTR65jXdY+0VR+H+P2pJsPLYJkYB
/sJ2c01+JxSs1gkFI0cqvDDpUWQrn2T1RKe+FKZmHaiYsaP/+WgSw+hD50s/1FPrPiblEzk1/xlp
NohylxFYTbaLivLkHUIAsL/ekCSqwumT668v7wuuZolQZmQdbQ/ppySQN2Yw2uDoAs68KlJWdj5W
YxygPVkRyXaW1ftwzp+5vkPQ/QNzMKfyYE+5Q9jtY1SBIqr5gOOYC6QBEVWi/n2sJc6pTwJpHHgf
VwWrfgpY0zPU/6pHiFg+fOuF6xfTfz3865y14/EXr+WCkwR7l2rKQpjDvRO2owylRk/RsOzez76P
Vff3hoF+ukgn0QXjE0Fc3ikUJg5gweAlPVw2asyQ7TF9ZeyVG2/q4xY+rMNwjdIacT6eHoJqVNfv
pUVcfAuTeJtzC5b1ukb2EoWebYKKlyPl5SSKN/+O7jJ2IflhI+OYmXpzYYxG775BgD2NOa24gQ4U
8FwKTasYiWhCNQIPNuMeZfqKcyQQqDHZ/MjyJ0Hp26bo6LIH+ghF3IyQPXinVymb3p2tOFrtJxJw
32mMwnb/QUKZtkloKkuKB5gtkx/cypVT0lgPcWhRO+GrUQL3uS0xg3erdeySZB2yv4KpeI5QNC+P
gggkPSlntyAHrazVkRu9DvwIoBbqqFhpTWbR1uiqA+p5+BLfSMiVUvCyck2Vle0BSm4AI+fXKaAq
EFBu+PzhgAPJZSIXB8YuybX1oT5lTOJ7Mtp5OV4PYaJhITm+QpGOHlwmJGGEgFkjkFd00WJ2jr5b
6ipm8WFkR+x1HyNltCLK3abhn6UcRSw4g9GRaor70LxWpXAhkWRZ/HtQOkYYjtuqR7UaA8VKPQUP
nFp5KzLavWnnVaA6R7s1EcO7ebMz2TtFxAMquQ2sDL3rOI+bo2Hq/xQwM5WyCfOUUqm4iTe6HXAN
ogGE3ZkzWOC0OffpjgivB1ImHiU6lIF/F4fY3V2qsJnaRd4RmLQBTtVBxJ0Rw6gfroBOIvy0IR/b
S6g2ViEl834ZwfsfXscQ6VIZ1vwCBGvsutKIO2O6wR+CxmCBxaTZrTcZYFeYgESmpu8JgyWXKLnd
DPmc8upX55NKoI2lPQvMgBgyAhKiNf6UxIT3n3U7VnX+ikpHS6X2zBZeMiDm64b3ZU7KZGH3ozOr
xUpICOTS5OSmOgxLpzgza2naD7uZsfrCONtzpOiHPYdjHzPO4Gv6BN+p2nFfYmZ7raNCDUFX2E7/
iGs0+0oL8Rth38Bj7KAt45DgXOgupgWsU3ajcAwtU0nTnZIdEIBrBscfABbKwxGi5IwOAf+C7kNs
D938lgc56o2oOG8qB9djBrnaKTmyK0iFOejpEWc7lh+2inszVGzpQEX8QL93FCFVqG4IIFjmWajF
vZxQVufrDP/LVU+ovOOodbT3zSzkgBfpThZEfrO0+/UyJTOr5LAmSe40qznIVw18Rycd9StsfLTn
njJg7cLqgeuZhlYoe5GH7hXCrI/9toOE5wa4JWANq5OITC6UY+PQSNNuDJgi8l0DRmBu1LWF5P/t
0Zh19kGhRPvMCNB+DSNxbMHitjNBjlYzSbNg/dmMYPoDcRGXZg0PqYZLJzf2xn2LsJYiMpJP2+z2
ZnUJwW2wtKErSDcQTibNwuxmGqioBIjogLM47mEb9xf9H4VFVMNlYScgDEUqNkyNDpGb941vo+GY
AewW2rXCH7b6eatcFBuOhOrT6J+8maGgIMg5BAZvOCfXizOyw6G9+Ikr2SbCLUv/iQ/6Lp/aU2cl
CCOhOZsaQwHJJDygLyi7pKeFbuTPeEE2amgm80mJalzySywvive/VybtNfSlnHYrdlm0TmSqyH1i
h3c6tBh7YYjvRpIkXuJ8XoTQ+K5eY7qn/lJBl4ELE+gFdfGo2Bd2Lt+q68ZOP8j+UpqgmE5HHxqd
AAVN3czCxr7HnKQQQqmNUVlh+pt+UMCIpV9bbbHpTXzlmVkHGIDtulMlGphzoByOd9bfagFHXef5
DmVIZwU/xjdcyfCGqSbyQrlZmYS5ZWMB/CsiT3kVhk0W1qy9eSSUgIr1A4mmtgwteivdLeVyE6Jp
uUSco56+2RTqUss4Lo5pFQW20nVg81Pm4hwJ9q+kMb9KBsyZLgIxBhRf0q+2dED/XX3hXr7F8btm
D4FE4+Z+qQqa2kr8dU34xfa7g6kPr3ex/N/d2iHE1rDglAdQQYpjGzAy31M6xBsQfnhcHeIOdNJT
B8fYbrsGaKJ0vf3xlOKkZLs2SYGuL3r11taRoCbaNqnfLS5zLcechtyaO3fGIKwYjoUn8cxfByaM
6f+XTXVG1WhZ24ObCGjTdm0O2QpuMnqa39ly++s3gbllaSANEF7HxM6k+/1XUqhYOtLOttckPOG0
DVIZRSMDYCNPrwAS6PVG2x9yVokfzDpR8iEJ8UCxX35Xd3cI7G5xR1ppk/uYlSHbiX36M+OJeCmb
Q+qT8cFk164A6n2Fm2/UnYiXWyiwrkx36NwKEgDJm3MisV/ceC+0pHuG1BUBAv1/ntTC1fp8OpqK
CavxvQMA9S7UmoVq/8W1GxhHspGdxp6tjhgazRT8WHFjv/PPJnDGBT2PvyBZ0dGYARajDUDPiWnB
WzMONSHL4P/O4mPKECXqZPVMgZ/8pQxQ+H3zrckg01CCn7euXb9hgt0COZzuwEK2yYQmuwt4wMxW
6ZrUSZbI6ETo0JWgqMiFgs6J45mjgx8DD/YjFRNAoYw/lLyO2bfqYMpY5JYvNc+EVNwxbRFCVRUj
mNY0dnYNj72vJvfZz7HO2JSUFI41DZ0n+pTdkP7IMr+8PoPEVTmohHVPkWZqqeWDnY3C/6kpkCJd
EgOaboK2/BDXykb/Mgft/lQyLRoy06cTHrhSanYtveiz6xFDDNjo3VmgpqFiyRiUQhWgZ4SNdDwk
Q4Q4OHNoMJ6JjCW53mkl24H7oEIX6s5SOhCArSbl477l+bswMw7OZ1+J0AZ78n4vagyIwZRb7UXB
dGwUlj8GMGuoiy/TQEZV4Z3jfV9Zjs6m2cEZyDgMreFDTtkLbJARFe9zR56qIOsa80RBfykZnlf9
5VZFJsbn9/A4g/Q4sSVeD7VWgVKcXQRByYUE74Q6al5u6NhdipPxFojmNmtz2aZkQ04h9iAt3jpU
eZx2kuKcvXqn0fmTMdIJ5UUenCpYzcsLhNr2jJ1KRfrstcKWrAjdrJGLTRYXGOVq8XFk3naXtWbt
rS6cXJUiyyKaUjXRb9jeUuFZoHeRqOq/xqpcDIlFecpf7KjuRoMrPWbjZE9SOlLIapktb8h3D2h6
0PAC9FxGW/OovTwlnw78Ccxk100fesafjIzzU2OCJYQ6DyEzoyEkakxGvQT7uogOZKPEis+scOj9
XCEzutWo+7yxekVYQDSCPF+AeNwCRUF4AIgLVt8ylhgYkMjDSmn/T2lPlqnIIi4epJmF+BoC0tDv
W0qJHL+cZ73Dolw4Pm7vJdOLKOM7xgeNxJgzWnUnT2YBm7DQQ8LWr91S5/N1EumFc9SyWJodqCQ4
PWuY68zYDD9477y9uHGXpkXeZ+1GhFfb5sIb1SNcUrZncBloONhBbfyHdzQ+IfNr9QFIBu/dFOoU
3rXEa+4ZWHJB4q3OUqBvXdQLem6VOPilZP+hhOh4lOd4UyUiDPcWyF3WIvyEanF83GHAY9k34JuK
z4zF86Vf81NoKE0X1G+RUIuRwjhw9ERoIYRascrGPFpIKPoZO0oO4GpH4SpCPc2LRhdEA6fYs7a2
7M5wF5RP92UledVyrYeur7yfFT30jIsHZX0WgwiqiknTA7w28Vy1i4oltiYQFJHSN/1tX46F7vaX
C8/E5vHitF0JEu8egdnfanUquwTCxauZ96Bliwds4amdvlwZB+OQp4OSGqrByimO7A7+lJYhKWIr
Lk5r37PDgb5zA79+XOm0D1eleLlgseEnvByLuycC1GUUi3L1xm1/+SYS+vW/tHUj+J0oI8jWjDvR
2P/ScK/918j5fXzZgZIaGr7kJ+LhUIqQ2FmKtKZzZwTviIF0DBjZrtc1b/zWfBC8H06gOdAvusO0
Apd8xzMHdbj/glXx5Tm7w28hdggxbQ0avxUERmjGby32PMFWMZTwkUv5gB0mB+qtkaL7/I12OYPn
X1f2wvRVChm6Znrg06RaVb2y+nSgr/ob/dnTH335bqABEKDzwFS0GupTGi5DGBQwAXCggKvcm47X
ZxxS1v2tCLeqq00imkB86Nz1kDvd4lJAOqbDQ6oaOEDHLgIccSIAZ21hcH64iK8M9BtKfzpdf9oF
OXY6prfdGRYJ7sHqbZMZAYoawYrpiZnG1Vr9DW0HBG//LfQ1LcuyHnO1brCly7ecpVVUv/ui6qYp
vPfu0JkQH3ee3MAbi7Zv7N/6wokQy/vklrowFrliM4LJfbynk/RNmcFGrsygxzsHh4Hg2NV5+++s
+35Mfk19TTF5u7qST2YlcPxxY0EaUmyKGvVjZ3Lxd5qQ/DQ52jgsqF/rb2IiMU8Z30xXI8LlGzbp
u8RV0X8jnNJ8Mo74G0hZygXNouoEQMJMCUKwPcdrwK0vq8U1pkkPEImbjoq5Ji1Zx4tJXs09eRw+
iDBzHk7A9mhQzGGkD1ZAiid+xs0We7UCCzD7sxe/qdT8owuIo8PVG/qK3bfmN9bTOhGZqMqbheWp
1stjBoo3gx7a0lUyOnpyj4LfiEdiqm3K6TWZ0fGA+4QYg8ysgek9tJW/isDDnnJziXAuV9gL3cbO
/ttCZLaGfLq3viUkMctu4+LAkGbE8dbIfbd28eCKfyn6j4JDPdNIXxjS1xyWRC6W/9Nz7Gy81uuf
JpVNVwVR+638zGGbtO2CAgANqfA88sA5z3R4+rPzbvrVbBAco7f3S7AQSP2K+Rxro2cHWdGq93mT
VDsxytA5tLLkkjceY7lM+L9Lwjrt8yedATOSmSWgg3Qux5OIAkM1uxB3VsWLOr4JQL4OLb/SDKt5
gVFTcshx/JzXr++QZ5orwNSRjtNSTz1zh8ouJpBRGdBkwVm9fFayvqBR5dSeTwzcfAk16xExzRXZ
FG4dHZ5BWIE0N+w3i2SSBGaEaIUNcgU/DAeF5sfmj5GzlQXSWWYbE3Fdv3v6LN0SOsxU5XWRdUkS
jVV95ChpICBWKwNoGOBjfyaV58mNYTsvt8XQLWEpctvXagFMX3XsJc5SNJL3CcwyfKWhwYGniZDX
aeVtbtY29voVIJ2vWL493SeT2cZwi4U4IrZcinbPidhmd86YMMDAPEp+Jb3ZIF7Aw9tPJGQKgAU+
RzhZlX3vG0nemU7CPO8XgjRACPoXe8bf9PZVf2caeIWOMrJPT0LrPwpfDhd19BkVlUgK3FJoJxKw
PPsYo3h8bF7PP5ynHONKtE4XWKxCUHXx+n/rmQnr2XCUHcxYBCJGfaJZpvE96mLcNdA/xV0eODvZ
C0DZbUzmPUNR32lvkCUjAMEqPuKqM5qTnEr8Nk/MBHB2N+Wn/uve6EQwLCx8AcRNKyrOHLvtiPqc
cV1xeTgkCU5sxhygAVAuRud0VdaolvlfF+IGODJBKrCof1Vfs60zDj8+O/oONEATm1dNlrxexbIE
jPthN7dOyF9KPiSMrP6hI7byQQHPnh0lCWjk2nhZFWZ2/eFb39jD5tQnD3QF3EVayLz/VVN7ako4
N6kBV9yAAj+qF3stA2UilD41BR7sNUQMuT9cvj7+fxoS6vKBEr2BZc2snJkH5H0uyqWl7GMnJENq
TQu1IGyGo/mOGBKGUAd2XcLvCjhsxVaUk7KfAix7W4yIRcgp3jPeV0HTfm2sJ24RuH6s7LOzo2y7
CX8Soc1ft/DbIS/u9YFJSGAYICinwRheLtRRzHroY5hPg7d04AUXyoj5kkymI99Qu9P8APRJekg4
u9y/G5nVn6VSPMwppmLWMv0S/25wHjKiS/VgVA0kwIG0czERatkDTtFMoSyFGgPk33t1uFiySZI2
hIJBSmmRA2Mvsp+NPbSOIZRNrNji2GgIqSLpd2aSe5/OqvG1lbCC08oRKyB+H4KKhhinXGdTD2ms
8Njh5Y9r2jOk8FOMg7MZeSa0wYEIm5nICff3yBD09G+/YupWiw8o5242FLYIpMlZRNAq+imbYku0
O7oxTw0/7Umgj3Tp1KqXRMyXVifNhxKR3ijyQuNxINxP05YMDmXU8q4EXNv20mfXPSI8fsSSzG7y
XLDMLIdsk1LZe0YXkppf/btdgSesnnF0MInoOtx2PO/7EQLdGsQiqoLb35Gjvk3P7FQ+QhXZlHvP
Xn4sHNNI+AOWn2IdEP2zkQEumVRrpNlp/QcqjJaXHNXbuoA13Y5+nkNM7P7wxXCQ7ocYIakUGicP
1r4GYLexl07dQ3k11G2Is4hwWpkurIv77j1DXCv2Et0uIhT56IICx/OSxvsbUIOyotMd60wVHlp/
gM47sh3gQGYKCorm0FiKg8MBSw2nIybRRbtfxFJIa4bJa5Ar+HX6Dn4HWOyYWFhfNDz2q7+WKVQW
GIZY9+tIVBFAR5x/0pDY6A2AOCct52AVHIw+yTDWToyzcA2nn5q3UcpIDGXLM8lsC/CuQfdJ6RAJ
qbTZzfJeKJOTkSDRD85+vRo/vW6MTKNWWBFWPsoLa0lbVpHMJTu2uyBX6PyUUO1Lh5ENhyTJT/rc
0ci+EleJJqsM/dps+mQUwSi8g/V+QA4DnVqp86XHDAYfVCrFxr8JcF44B24+IPdcJLL8HfmODygN
973DCNylG8olpdCZPiQmrlhMiWovvJsiV60wDQIGnFeKpvCcSRtF3cflX/vajCODpfRoNJl6lS8g
V+QVWX8wM6O9oG0wOEzuITkYYSO20Qktc0ezEHAMWPcAcHlZT+CmwG4nSdVL8ebCaKR8u3kHSzCk
7n1f017+pOaGFVpgsp84O43FTkXkE7rkff1lOklsvWIixraA/l3vSm/3ecvT4TwDYgRqSKRU5F7A
6L9VQqqpR9jcL1Omkx2IJmjVntV2bZIfizz2GLGkPeqP3Yex2WthXcOyRlMWLWQEuPyB3obDA0Aj
xh5Vz/shhwYj54RtQyHE/5S/YIiKoHWvsMGqB2goj9BFCcYGnBUOz/VtI77ImGOyFXOp/AKe1W0F
MRS0xpThzacT+fcFB3T6xmdHr58iUGhl+EGgCkh4SDtSX0/sVTrEc+CkE3JObRXQFyIeliRL7QoB
0WqJaYQq69yh3XciDGcx0oIvvwklTJ/21+2Zk7i9oDoloudVUVJLnzqQwXve3OsOXIXFfdrShtVW
Gl/UXxy1zl0Almn2uDtNvceP3N07/PbIhQ7wHDql5fI2Vu4H2op20cnyNwr/EER4I1i9opdNu2WY
p9qjCE11eAaKX299fHnt41PUiegVWbsrKDo9UaitF98Fk0AhrX6vY/zBoBJ2KdkSOBngqrwnyBq9
lvuSaEfWEN4MKFgYW1yylI2eJOqGfcEKQGxfl2g5Srpf9V4XCijPLhnqBm+irBXuKWYhQ7PPLWAN
e0TPJWQ+HB6wEuYoPixv8imjbS7zq9FusVHyxJgr1Y0QRkmfQME0e0KBfIQ0z85xf5uvOrAamHKQ
LRbqKNn6AG17Xv0lfFzEkask1p55xKIG2Kwm9nfgpy42LZRyRsauH2Oin3H3osMxYCy0J9iospxg
AhjroMef5sYQheCTHzI4B18Ct84ZpnXhva4KdL6qw02kn65djQPQhbLv6eSUcTs7DNMovVfvv7v0
/pgN4mSp27iwZSo/KWm/PmUwd1sc6fj58HPRqjsznk75XWTuLYpDKA0Giw4ge2898JTZCvqCpSvY
g2tyJrozN2cq3+7wx1DBo4K9t6CbrS1s1mAgyHeSednsil4dEwQ6lmPYJXo9LsTTySO8JnAkQyfz
FJKV/+Qoj6I9XjLRv/E4IbmVHjWu1Egid7JL+IvH/EvtvYNCiP4V74Ol/iCbF/+ooVvuyRLRICok
BHJJrOiU07QWwhTiAnhr9w+OxtSbkcHqV2Gq711tMl6Q8/PkkvpXJOyinXhWs6wScPtyHRSJmAWg
H79phjmB6kjDKxrzyZ+KYlqU/dBdagVXltBzuzeRl/Fys9zj4ALYYj4d2fUtqMAsvec8hOnzkHRE
TuEpJEKTzXg+bvdMRDbMsQakqDWNS6hofV6qNBIZ88Z4EFfURqjQR3rtvS0yRyN7L++/fvOGJrn1
3wcdXV3LUc3DuTXZPrITWSyBPdBvaNEh+lGSKD2/3ylRglERhSoHmuxiwgHEkEPUUMes62WBC0i+
CKYC5kYXL4LLxnjepAs9fsCCyNv4BL5Hmp+tKYf0c7F6AVeVLf42o0WKMNRxH5wqOUFXkUNpxNuU
METOlDjw9AeRMFjbtZBkaSQdjmg3xfPUI9q4Ayp+iV0MiEmE+Ti3Ef41XgvVnKMFnhifPF5ShxY5
3w2c5ImxCM+5vCQGujrQOqgSx7g8G1/ZfqenWYnsp6hXXVxFtiGpm/mLyOEtcIWeX2VRaRV3tCXq
/ANVTy+DG6TJ/3nv2YgXZDFSa2TgePefDLN//xJhYkOJ6UC7913LZdedzDC08gHWnF5ITyFAVubp
1ottdz5j8tU9B/6yZi/1nbFqOmKNGF7CqNbHmMtIZ/VylRFBYAxBv8SCXpTP3qZh79edORLaYeCb
ZuRO9+TR/LBQ+rEb0IKf9SjrjU4hS6VNfJEBa2FR7hMl8nVnY8XJPAmYyK1EkfWcgSo18itZAnAI
HeOgx8T9Nni/IQDlIoObw1SCkrYkdUV3XL/rr+mHLFKfNGIT23GGcwMqV3FEUgNxIxZ5tmOepW66
blDOi9vSTd7KN7S+zsFbuk8DXRN2BOx5aJwXGJryGtFiIEz5dII1B0ME1fjHgdb1Wj/HgEi5a3eN
3oiAW8gz1idOWBhdrKExnYOeveJ9tXPT9GrA818SAmrqPv6REtdFv/PEDuVdRYrFh6+kiUUJISwQ
SmlWVEIVIpx/YhnOn56bbrt3LWms52mq7zxSgjFTUI2qynB7pv2AM64fC9LKFo2jQQZ59SOhcwAx
IAv7Usqyi7PXpW6UdY/ooxX/J7cCHV81GcLAu7yzqH3+24jMkTXU/S/j54XfGtvpdN3FRjxLZUA8
6GBgqlju6yEgFBsfpXo1lPwSOUcCniDVv40HETO5Y9Hv3Vc+ioe5KKxk3uQ3g2O81cMDmIEimcH4
fadzljrhUYfG9vG1jeyhSoCUAsOLkrcCnLYdS/QE/FHmfFeRz/dpT0bSYVWvgCnmnULcdYce123p
IMbuO4bqVHxORunJ/SJjQ5Q9YDn715d0I2VlgbHK96ybJFrpQAcjN6ekbKtpBzPcK7sgNKztGELL
LmNjKgeiCudY0yYgqfkUU8PMPQyrO2Sk9Rxy6L3mcqIzchb//8G/mapiprcmJ32tgO5+Ia+98cDR
trLl5NouU9y4pcONxBhAZkNeNJfh2gQk0xND/pc1QWkPGcybjInTS38IevakheTnq5zzgtxVhTQG
Yhoxxu4KX5w6gmwgXl26DTAvf+wsyuu+he3g1UGql7ZbVVi53DFXmch31gWJZtSJCmP9byfU/rJW
vYELjGIU3YcqjkfWt8wCBpGyjiP4hmxzw8NJxJ29Md9lzhivGOVlMeXumkE5fqzCRGBXxRw8DNef
Pcek+2FaTF7rz1Usifnhgeq3XLIKNYrqVGxLvqptylAzFbpTGUK8dTB6iPslUAN0f0por45NdekN
6HptIkS+/QVWbcYtIBLMZsYyirTvsX9NYkEytpcKJ8Nm+Tfy7svyoGqcm2YFT5fQYsdjkvHfuvEf
ug6+7fD0yWqsGU61q9VIgeOe2mo43XvK26cntyfDzsGVPbA1SiaI5WfjUW/xBmjxVzez+JMlqhm7
YsLi6pCC/6yF2x47nguScCAatpyjYkUB2zAXyYBEze9sQPDObyXjs8AiJpLcn3rs+ARj/UNDfjmF
uIMW3UCzbHt5jacn11pGaZF5gnxPn876OzTpGscsy6kDEpp41vzYd8r1MEw+3nhRTIjDd6uGkbxl
t9qvmJXR64lnzoD9IBr+onlKOIT6o/Zrb3hf9XAE9t5ONocV7i7KoY7bH6KhxH088p2/rd6lZYB8
ISjYYFZKomC41gzdlGaPEB3u7XEg+3kolLtf7uEftE5rJ5pX1PsmxlqlnM9MsFPovML7UWNg831A
7UDKk4JM1fFeH+d3tAF2IZVt0WI2o1Qcb+t1Vlfbfjb/JTccgvzM/03rLULbmSp24rbN47AAMzWF
zFsmE5d/fBzugx4L9R5sDLMiUhGEVBUOsyxKoFx2ZpnsPzZDbrHycidDLJQsPpIA/DGVkEsvptkv
Xvju6BAFLS2b74YVaaXMSgpNogVXz5nJK9OVH/kZxEBA4WvVQ7JeETDqxM+frWRhhw9uoMor6LpP
u4nT0ii+XBrr2Ij9Cx5bLREoatWl+7/30gmyZKNot3gHTiEW8JTqcin0DcWvfgCX6M0vqttoz6i2
dwriGP3h2OVM2lhIM+OUdo0rByQaiflJS3IqnZRCQ5OoI6vRyjHiI6Hws/5o/n7kvpppQxfDn2qT
Sw/dfWYmp9SIvEo4nY5B2989g4eLxZKjDTATpBHDrT3p+nN0YomU5xArnrldsyrvNrZXJhvJ2lzs
pHW+FVrhkyL1pgWzzSrHLH7TrzSSKkN+Zv6wFj2EuX53Tng5pWrtp7EVrjaaz0jrWKMoDNCyDhws
HOEFEDmmFYQGV8DNU8GwJB4S68AHx2+pz0BRuM2trfm/xWlHF+kP5Is9S+KBdQTTVXTKYe6UW0qI
RaI3wx/Cvc7Q1AbxAkdRFEaYPU5Axnl7HCbPhV8O+IrDWTTSls93ts3Me4IHGbHQdyN025wZBabV
j6EuG+M6K/c+tmPkk1iL7qY01HxkXWjZI8p7OfvwCNSdb0Ybu5tr7ynScHOpNyDPgbUF5mLZQq99
X4/14UHlS9T2COhVU8C04cjvciDb9VOU1b45vkOSYeycPux4RVGgdhDtElCNHA+zRZhLjopy4vxg
w29d/CAa80Rr4b8L//YfCnTSgr1ZVgVetanZnJETBZo83sF6huImQISY9XT54C2SikmUGIA351eC
Em8P80ckcY1BY3gDHba3h4m9xY5SRPVIDZ3RjuqbqVLkM5T/eZdRrAFrbV2q/W5UKiiEYNhuIwZR
31EBayJiaL9l0WXTm118YFCWk8Cy6nTv8tGhdlSGjPZvxvqZT8GfHJWBhYKcOmTL1Pgsomww7VnQ
buBj79GGSLS/vAWR6KrgbSA9jOfpeoVYs7CXxzPWd2XSCfBlo/c9Rrksqr/PhE5Yh2uFvpcBRxVQ
6q+jvCuVVCNMtLfiAMITl7uuiYYhtZAOOH8sXVVCyeQiKs2G5IyQjUVky4ywRCts/j/gVpd/52+a
bz+PoFw6oh8QNhNjA9Y1wSF60ssPBXWjHuSBvW1pmyP0oizw+lMzCblDPP/aO5c7Z6K0iuFbW7gD
tOfJtSLHRE3O9loGb9sc+1UjKh1bo5BHvjJnatQUavXAWmyfwWvWI5PBuv9Yh7Tq6Yb0+VVTLiZb
PjSgOmON0zYUvFQhK/fMynR/m2uMF5xiEYteOAgAqc1szBAg5bg6+Ia4avEWE0CkAAR5EYw7BVhE
lyx1+P7XjOEaK8owRUyGPlhkWHMOC138B/U6pyQvYTFOKHpGeC9ttPxdnoBhweIfJDFMRleiK0/h
r8RCfvwZUacropaYfTWcaccdR+PdI0VpCTJS2CQHUWtwGVlXhrgW99GjWJ8fHCIF7NW2btOiRfYU
H6TaSSBWoPRIZu/RSHYX73IByXQllvbQX2tZbBijlfLJ0tFyjkIGU+G9zFuRIj4FfRGKlVhP3rqG
V5G8he/nZukmUIOwSKnbJYmgQAC9BesiBr03ZTazw/jY4sfIgRwd3/F5wJSV2sHVoTCe346o4PM4
TrrfaHmg9AoIegnSQ9RmCOyZLVWkH2YpPVJAWxUS9HMgmINZ+wFErtH9TmmEOKrogll93MAZHB1Z
d0OTRUgVebOpIXC0M6qb0M4EAxZ7n1JQVsxyXEJ0n8lRCPeiOYmG5bVWpN3DzaDIo2qYPvj7DelV
aZW3LuASyXVGVnevENrR395D6rEBsBkGVsq3zJeIEkBdmX4vJQiLTyrZv3xsBFbIL0vUXuNaN7oZ
By16ZneSq5CnCw0ZuJoD7ywN/51DbbPaxmv6Rxw0T13YbGa/K56G8gQshj37mrx8CMWSiJabTg2o
nS6Fmu1dIVrijv8GSXE7vytmYkkUadqzHlQw+L/ORxCIvlRMGzcut2hPfSaAUAKyw5owbuiPwpQe
s3ISLqYDOzseX5lw2Belkb4o5stXlnGbovvTjREgA2Uf4IgNRw6ruLITUpiNwYr1f5cUmZpLeT3V
/VprppumrTo5t3yC3x8OScUinVitFTEVks/3L1n3/WfZnwez6cH06C1B+xJkLRzXZptKsv7cOqTz
mNvt1UZIPPWL4d850d3CyGgXBOv8SJ+u9WVMGhY6k7TwO8ZTN56jDil/w4Obr1P9ECP/9LZBu8c+
cmpmvg5bJeWU14Ll3mFeFv/SNgKUcjX40DicVDdLDTgU1TtNCOMRnoDe1pkS5Ex3dLdnm9PYjTJ7
WokUHQx+Ku58ZqM36gsHXiFcSE0PTMHQGeaHBSIS1hpU+APYIpmzx9lnOH73GERszBRWcYuO+8jV
Gfc4L4mnpj6P2hnpo08NwZYbifaiHppZ6lzB3lPQbi26gV+RgQFY8yZ4PAEElX9VAsTPBKZjBRZb
LXIwDDFW6ysU99VpzyZrv0xjpH65FNoOpwPc6VFeRIStoyaDZEUpJWyBy/fk5EGoVZBFZIYCueyv
OJuLQJSJbwlhN/Fk67Zg4F0uIRik47TgWYvmZu5dYcqRyhgk5Rric0fEQDx0OGWRs6u3L+CVkCP1
ooSQeBSjaTerPLxLUaRNt7JCI+aUPPaXj30HdDz7/X/cD4+biJ6nB807VXSzjNAsx9rMjG41dT4s
I0jPkLEQ5wW2apyDgtMPcHOIrTMKxjvreyB+fpIDQ8MLb/nSX5++1xvjmnP/JieAUWBz85fo5Q57
9xx+uABOzZhiKAsOOX3yLNrh4oLPYbz+/lUEyD1CdvBtPx36R7fIE1bZgoojiMdHtUwMtk2jKYi+
7olvvnOSqMHbplx3mWg6qL5u95TQ9hf7XgIztUYRHRJ39Esq+B075aaXJEClG88TDSgdGCrz3j7Z
bCyH46Ub1p0RXUrQk14D8LLT7jQjx+9akeLwVLoQ0wrpz1SRWA4W84bbaUZ/RkvIRylfoNdny8PG
kYIchaly7PAUoAZKFgqR0O1GHtfSfHP8krliOQQn7hlG6KrmH9pIlnElQM1mGRc8KZb+exaQKsqC
g+yi2VwVyxv+czesLKDSexC5qySB+6XVUZIvdObe8yxcRkOI9Nccl0XdmVD0cjBMIsmxnzds+Jr5
30quHnlda/Eks91X7ZbalR//nYVCYsRQedZgD/vcqgcpcbc2yFtjImpWCN/e/7jj1PTrdmHKiWun
/aWEt4WpMAAcjvRYbpbIJj5siRy/c7pwoPFGbgnxXjAGhmf53EEuJOxZcCZ+owRle+JHjNsG5CmU
zMlwQdozZklkglRIc9yanNcF3Pi1vbYmbEmxH5MtwUaUFuJGD4xp5ENHEmiTraxscllFJFQxSiUx
ll9wzDpPfKWhjgu//MO6rRSr3llslz0xmmFWRq0OjBaMtqsezrADBOh1Ekq4kkL+13oXhnC/WOPX
KiodfryFgWeev8gff58iqn9yGI6nQRhBQdEuqyTIzjpG8FnfR29QCYrnbIbR0g8FeEbl68PfLyQA
kiADQO3S2yZzxFrrqcxMg7bgsM0VGXkjsPeVvG5fgPcRESGLLuYLdnT76h/+yjmS+FuFP5+EMb/V
tLD9MHbwT11LY4+lsQu751U35ZRdYPeoO/5uN5YwN82ZSM62gY6l9rWex9tBpHNZZI+iS4RJLIZ1
hEI+/8xUlbsidWfuNcL6/AV2wlaJj3KKBPscy/vfFHlSypT8tC20jQATl7ENKSA0HQ4Jf2jiP3BT
jRYO0hSrmDIiabPVCobRN/PeYqoLNwCywKYr5je/RVRXVdhGJXhnXjeNH8NNi7sIdOgBKE+zYwA8
yH9A9gL+IYShhVWfbD89Cwl7mBVMFZqHzNnjqh37IKWHlG7a6UgcAU3sIVYJInGTkunmi4HKb0d0
IPipuo0e7VOZPqqbIcWCYTMmaKqW0am1sucUHK6/EqwHVbQWMXAcL8wcFwhJi4geUNgEvjfDnxES
mm5tJpBVkXYjwAhRV/MeqyXgPXlrJj8PaRmlB/S+GqAEa8GbdCe7V4iqSnIHGITC8iUcXzOI+i8Y
dPQx1S1rbAd/d1ZjZ+UaHLdxhGtFNGp4Y3OV/UA3hltptsT5zyToo8Jq9TtjZy83X6xB98DF4YH2
Vid9eydFLesxla0jKP/7eoXKoR1QC8yeEhUJXdwnyxxRDIxkLWoHom8ALgC56GYscrwT8rZvVz1h
TTKNotl14OX8Ij4N+vfnrpB0cetjo0o0Cp720lMTZQP12on8v3V89e52mAyfwNl3n79UDm22RbYe
qCHkcBIi8MBKQCiunApZuZ3m6aRZczEsu7sFv4sRb3nHM2z0AF+QCxvswgp/ycjhjCgPPzKv9LR7
ziCZ9u1WhOTfvfiit9oKitm9iFbU/Igl63CqXpnRqQFvnw1jFxO1RFAYpyfnG/SZyTAh0G217gB5
tqOqiFmvCtMPKK0ezP9g8XyXSja8HqjB2ITy+Vw8c3AGc8jRZ7jVzrSe4Lhfgu+LuETu0tvV7hGB
qqH+goEP+Bv/RbRP1J3MirDAHyXZo+t5FdZvNDpVjaLjTPEXl/VJwkKPJSJv2YDzr+rbPZJzWhed
pgXzd+jcAfdX51DctnCUUQI3DUNFrdNM3xfH0MvU+kkqRT0s3Dsx0BV2c61mKVxjYkF8xL95aSlX
h1GzU7OOaRfdnccBkqLLHs/qlOf1T7rwnvey+XvKZt4VenWt7ZX1ud9XGvq82NTmtYjjOWzoQjdV
27LI3Bo3GSCxXRIGxKlshqO+VDk6bVSakzD6XtS2WffBRCRwyBohNfVu75rkHincIDj8a6aKikzb
6ZTdHs2ItqyfZMIB1frdWH+gORHMqSTzrWckprQATdW4cJYBoX3G215uUSE4vz0tSK0ZNLhl8EOI
ja5IsvdUj7eDOmmDDwj/Fovw1tfla/nNj9w0EDbVxAyvOL9Y8IyjIUKgnlLZtEJ8MCXjEDarG9i0
1e+qqLCCss+h5ff9KYKFLikzdW3lboJ8f0BfrWpi1qwfTx1RdVg8Oshwmy2Tlp/IkHakaPfAszpD
FMg3N39rANJLhHPM/GP5FM0ypwSqMylI5+pIea4pGeqQkgR+PHd46Jdbf8KFX4KIJ+yfPhSEYP+v
ZxFq3xEPLdZhfv02BkHl6bvHLNZmYq6rmlNFDXQ0pCVbog7ygmPL5L0JFCfyFdo6xQyRukK/t6mF
STx9WNMiqCCj8KZzlzpqM+33D8h5UYB+Ipl6iel21Cu5s6KeOsCSlfCCmnnm72DJjzXEvyhUGPMv
qHWlRqSXDArE6IO/WMgcngRQ/5DouVrz08KmQ2oKz9pvhZdVhnfulLSf0MYwLDWPiFy/0anHEjVJ
cjEli5uWFP1cjJ5vDBs3FIGjZeYhW81HO5ZmVWZtkpndtae5kzQ0Eb/gV5Q3oLHQFt7DSt5JVNul
bt6VLArZIQXnNieS4VqrBZclJUobUEj+FdcBsoitUBWsE85O7//YJCISu9NJgoWy+9aASGJ5Mecm
ZLJhPadwwiePz2Vu372aMwolPi5X+tPcyGAimcTuHIDvCu0506rdaT2QmtNo8ZFM97U8WJ+Ponzm
39QO3GrJBcZ0ngRxKU47n8tYa4gduyzPzm3vFASmzyV0LKv7BBVoj+1jtZ/nxQg+kFLYIBPlW0VI
6cg3Kt72mAafVIZsqFxdjN6xHMU5dsEp4EBCDZjNj2G2Aviw/EQXrfXIEb+aLUPQK2I2TbNvvzfs
gGgMF2BXmqSnhgPub/FbPww4wLGfL+TsBkgp+cxLW+CoGK8R1Vy80aBg4JWr5zaCpKBZrvflxVsr
A/Whdnj7nnMpcQIyeD+wUaw+dQgzi5W4YCURhtvjCp/neRDAIH/npxZLGVoyliSgBs9QUysEZyD1
geKYIjOkwkXRK5BHNT38sE3PJvS5ZB2U+ZZFeVphoJwLNgCR4cDJEjsZSTg096gOzi9eovUlQirs
VHXF8YBRTeyp8iElg9CFPVygofqHChIn9t0hjCmL+MLZltAWm4iYPJfB1Zo6PfwaJqNCrwCcGpcF
Tu4B2NHYIiELNA0EojAuCFEqGvvDkI3gGitpYuDTmY3qX1ZDTLcGT53Xhq26G6GSk3i8Ynrf+2+y
thmKlQASBRHL7eJaQ3BTDs4thXXQwGSZydEBK4QPpbkXOMwFRnVCfrcA8J/YLHv8cdkrOEgyYnuB
eh9ZZ29qhcKr6tNvyh8VsqXk8EA9VDqrhBGtxF/yJyVoNoENQ50XSXtzJpVIFOla5I5ZfAtfBC9w
QwEAzo7n19eqQJLF1Mcsp/Sh6TVNAnT9Dc9VIT33mOfXwjtYshkwNGkZX9PxvpBTnmREXSaGjiHT
z3zk66i3Kosi4y5qgVUCjBh89bfDfGp4VvW/Y+zRbkcrujd+7BJdP2zZospGHuDeeyHnYK4bzUpG
GeE9utE5ShF4cY6VSGSdPPIeml0vcHF1rUW3FRmKQh3eUSVZpkf4h+AZExKFa3bz+aI9QkiYtk40
Qbvn4xofzdAkA+3REYd+rOoGzc2q6VoyGlkJQ1uNf7hREwm5fenyLV4AyOE4VIIfLrb7SN6eKIe8
01pWu5aSfOCzq/+SU79X2IOzj0iZHCTIHybs57WJG5JxbfXiX4kr7nRHPerq+BBetn559Sgyo3Nu
UhPqymAGTaYaGbpHpz+8UqRrsGMC90CKPj9uLQZteEQCdEJG/Pxd1/9plWvBAuv/6UZdPvAulWrb
VxBPX8FseGzBhmEK74OXoV8B/GvctjBjapc497KeHaxt1kDo7+D485g9LDCkl2LRn+kRKLCAL371
vR6hyKK3Lf0YRDN31fvLlGg3kSid1gOk7PuOtZ6L6l365NuiKIW3aMjQc+b+SHc6cg1ih8PV9xA0
BhvRe+g8uoBr+oKyEYMkt8wk7IgddJ/V9L3OhhDPJ9TJLMfeE3iZNpds6RSYT5R3wOHeGgDGmiyA
Akhu+eUBaK5OqVVGdZWn8lUToRp8S6J9ZlucI9yM8yRQ/naMmDaSQ0UqBbTOa8TmTHX7Hy+fVp8W
kyYzQsoo2YDJNsCyTxpp89hWchE6VG2LZZTFESC2tMKxuWqIrS04DAX5ibz8OhWGvi8zaN9m1XVg
ZrsziYnKPVKvJCDxxcjgKyTBiyCNb7D3lPvmT2za4JdDoBLGCT6Oc8gz7FSfF9vlsFamaskosbIt
vSM7NZOheyFykzxFVColwc5Dos8/tw8mLbZ+Hh6Ph7p8j/ku7qNitiimdsU98Nt4+NwiZuKvo7Mg
EGfhEkfjWLK/3ECu5I5TUghfSvMTCOHAlEZOFO4ZvYpKv5eTAUrjw5wybbi86CIAoOoHEm8R4uv0
LYuOF5leYN0OzQPwGJ61UfVN3o4ViItz+WpqLAB3xRRQTIZlTy7IAXTFrn6VMzTxr5LBqfknDK3Y
34VykMDxC//uRMvLMI/1TG1gmeQbYhffCg+p7/Cjy899+kHm8l8uzVkmXZqeeyIWqF3IRclXx7ph
lrzGf2/Ibp0BahvRRLzH9AvrkugiTOBAzmwjGajdSv8Gjk44P/8CKj5+WTQFQzRDLSbZumVEokMg
k4n+vUOH07GcBja9AyXNM/nODREhOGjX40PjczIEvPVX59/fZpHI3+mIISNkaTYBWa95ulIRQvc0
XvtaK/rgVa8l5LRIqgaa5j97aUlsXfm4rZ3KiRXAqQzvyk8vET/smy/bh2Pvvv/CcXGwlCOPKB+F
8PEyA+/uCNuPMldVA2yCEt91KbTBxSm47j8C9IRso9Pj+ehFiu9twXj7OU+Sw/iSQauybbMOFYR7
+K0DtXn9IaqowM/TExSsb4AT3gJDHLezkYW9VRC5H0LyMV9x5y56rM73/9jBLXDPY93Fpc36fezv
pV309oLBXLCrmow99fQumkdwWGOJdVQqJZQL/GlhOxLFHWLZ/CUr5kbhlxK4ULo9Ylz2/7nfxpnW
bzceAJqWtMptp/1O3YYe7cYCyby8g1nXzRIBH03HOygxpV1hGNswuJVMDd0IawX539uiQbE6nXjK
mZi1RIGpOV0vgRXPKJ6uMUGXdCTm0wrk7dvaIfuR2fZe5jDnfluWtLbEjZR+BHsNC+/vnNLDDa9G
CGHwgRf154DgLZK/9j2ww5oBzCtPSZVeq6XlcWfO6glMnUoz7TMay7clPKMtE5dmweoGivNW/cV1
lF2pwvFlbTwaWOPVzaGm8byScW83QJmjZ0JmyGapETUo2VxZurbRB3Dq+iyOPipnYLReTv5gOc4p
/TgwwVk5lluwiwVFPeOT2U75oWQoLqIQ4Qse9PcARJKlZjaOhJWq+ZgAKqZHgq9nXgqOS4b7e8Zq
WGzCVlJddrJHOgFQnSJUO44XRtMyNAbxS/GcLY8aTNh7/m0RgqGtmBX/kNDx28oPg/hORLaSY+Fg
8ptK1KhmVUb2U7R04IJvyBk2Fj3sPGBoWtgr9mfsXxOMnOVwV0duIUKp38HYBSEE4p8k+uV85FOh
H9zBDsWDvz6WlMLYf3NmOEBdUorQ293QaHnVFzpczsPrIY3wn/caZn/fZo9DxiSU4OK8UKqOLeKF
2//HLPwE02HyzW1CZwOSJzrjuz87Y3Bw5TqKZ3tJoTP+6XCgPYHNuHzRE+2YGTrdbLwdzGclac1C
7Ce5Bnym4XjJltyrvq7qazTm6mnukDIv1Ddq3D4URIE1ZYyXpF6KZjkLAe6dhRsy/h9pLzTlVHJc
jB7vG1lpdukQJ2wNtr3K3AbqAAinvSjDirHYxbq24ceb2Llpaz8gMyKzl+/chnXHc+rNPm5AnUN4
oV9xtGucinoJLxifCbmkWtalPyvPY+fqWX9Gqz9GdQvGbBgaGyQv2r9EekoESZzagJv/FDX4FeP/
JwMIMmj0Ty9MVEeG7L/uyhqZ/ZESPkcPIfJ8UPpCMhLmF0Pv6AkYsVVA5Dfu+E3pTq8JTOy328nQ
chdYgus3xy8Dl0XvzkV+dMUHeP5Qgjo6/4EOWi8Vvtr17TBXO3tpTy/OfPU2OYq86ySxK4feYgIv
B+b3UDftuWjzZ+CWoNPpSEpeAzOs6RWB+YTdZZtNc0XIOvEEomPILaeGYpN18aAa83jpHyoTpaBG
8lAWZggoFlbpN4lWbqceXxXU5Rtv5JrCS/f66PypijG89ba0GZuLe1wzadIQuXB8AqxXwaIEb2Jy
lVGGxxEqH4ZX2TF/Wd0Q+ahIiBS1+NIAVXzobdmRcfZaTjFgpOxN++7/3L6k3xKduSb588iyvq9a
DXBJrgXMiYECNgT8z/UfsE/MGByiR5tUSuwwLRjuZAlYuvCG04azUSf2JBWsnd9zYXUs+l2o7TQL
gU9I5Ho3tbXfC3h8Cmtc0P9C9xkwU5sbyxaRqgeurQCPPOpP5QW+mdxEd6RIZVHW4hNuB0xi3Vte
atNXIfxMl6u08R7V1BvB78G3GmJO2FnK76gh+Gqad1Gj/wrKhuP6FpqYOrfEdrAy88igEhKqRwkm
35PuJmWpEJ/mNtTck7uv7YM5XHqAjZMglWp5YlU9RVlbuW2z7hN8wemnQxiu6vFICmDduQMYKe/+
zrHPqav60hjSBQMH9t9FSyLP22clp58oy7wFQQxDvuMGHujIm0ydDd5bsR2xZ+H2kLqpWe1Bz/WM
IZA6Ei4IZiPhfcUVThscx/LBHE7Zm2UAnTGgdLPq9ACYVPDa4UaE/ZHKY4tB56ACnRwUGf25xAw0
YhgD/FOztQFOSccFvS9S51OSSYtvcVL+UzwUqofzpJIprv12ZVY2VwikZD+x9czhmXAZ/yrW7uIF
qlj5YaUgxx6iL9bpEoTTX3Padr6jozWpGjJCDNR0tWUqMu9Cv7UOwjlDWFxUye7GbQ/RgMKbUr11
Zqs2phjrKEZzE2PeEmxZZd/rmfY568zxbBqy0KVn+BtTXemSftboRVD0kGiZQ1JgbXX5vyN3abpl
VhnAXgov6Cx91z/b5l5fT5Y/NnMVEUJZlW1yY6vPcoR3hF3jWuFjTpaXk2fWctKwzbqL1hVkUm7y
jwqnERbv87NpFB7rcjzAsKSBxTs4c1Yr6sjYucfTWFk6UIWaopVkO9dBZfwvitAleORwtVPPYe+T
uhLw6t1Wh2kvyBl5kzp4a4oxwOrNmYiTy9gRXT/HQa9op8EKsIiRbZi3XR9W22eU8WFeSrw0ldxu
BAOoNrnwhTXpYFWm/5KIWlW7LSmCgvhyq1XJVgvftwL6lL3wp3NRNUqYA/VteH797jGnpK8+cWGf
iQuaqS7MedGWxnbnqqBh6jUNmzgk2g7wJF05iXTew2l4i+SqTvMHE4og8Y5nYq3uYQBp0vxOBqoF
a7vbxu2YLce4HNsMOIQpGoIk51I/ukFuMYp2kMkgO6WVwBmOwsCesk2l3FNhZml2OAOBRtf0t+XN
sny6dzNB96XtTF9Vm3gz4filZtfJTJkXJ3d88yOPd4lN6UlT4GoJN18XijUxWwokBednH3raGVG6
TVLoxCtIC5yAkJQGA6Aw189K99sFmo/B2cxACJnFYtGd22rax49JGuK9DVNcZWQEOtTYLfEJXTrz
/u0BQC6vcyL3riEtsWBjk6+aoRYxxLnB2ybzxl6UlPnuIU30smggj8PDzEmuGNUfBQ2ZUR5leWqI
KIXmhqMyt7L2MsJbGIYwvFCcj2GIHrwlEOhI19puJS0D36ZC0jGoGJ9p3+4y4Z42bFprSZJHCBGJ
4Amrdo+9ibULfbDayVQRZ+vONeizLl+lSxJKqyTWsvH5zDyAtbbI8VHeMLyTy82oUMM2Fkxsh8ti
k3KwazdXSkdeK2ByqNOM8AUZngmgLdM1iwS+6+v1x9aQhYF6A638zNckAMaRf8+1ZZG4EkD6fkqy
BHGt1SaqlzhBN2uTh72lX7g52r1evKHEHq5RMniurfOT1PH4e7hWiZTP3TriNN7VAW8jd0pS31lN
RiRgIDMgXx4f65dR1fZPcSqTz9Njfhzw5btp2mS15Hz3VakHhGHOqBuNQB43UrB9yo+3sUlTb23f
+yDIllliXY7wqBEkoCTeMPJIMWyapoyE4Q2tdNnfV4j5eZkulyCP8FXbGMOhxxmAboEj+7PCGVNA
D1qlEW1Jj1rKqE8EavPd3aJfe1VZk2wll/1KeNnfKkIRdEtfytnXdl59+QNL0KTxpPOKe4CjeH0G
M2/CzyTZkC+ur37F/07976bOaV+wzSE/n8I8iFHQB2NgmlvbIWjzafRWICKFuxXF+QgqVD7tMqo4
DXdV/ea69g5r9wSOyTWnCmpeFbUCq6ZfsHYwbS4WE09C6sB96BjSKaRYCg3G0CPBrofquBq7wB8D
eQpvceUtSr3GnHuXGO+1jlyEhSi/1bZWOLHv3Y1pcDELEmoDY75XOX8GRAB4BulFE1xrCFeZhCNj
Q+9JHotoghXj0eCI4iU9TVaYIUZbvgUiQqO2tWRklSOdfTu4rn/lCZqdtZJ7Y4DREr3INjlLzPSy
xj13ePM4mNSFopFaZL3oouD/j0N3KVVrf7EtLCB29zMkbu3eQcCQVxBHaJK82pKUu2SHZp4HW/aF
8HM+mI5JrVuZmipifKSWJFg+yQf7ZcTRc4I/VPUYfLGLr8+/OPypByHiFmflnZoNbt8d/tjexwr9
YjviCZLo7uUdeTr1AHoLWtE6tAWDrwoyxLSOoWp9bJ/35MDRWnoFyBI7ig450rZK6u4HsAbr/xjs
z8LyFegFpZ12oaVND2c4iPgV8o3qgXOEatfPKmAKerBdtxuOd1za0T3PcQNp1a+zm+3eki+zVN5y
3+/12mxYXT/SttTqAGcwuPvIK87iWLJt2ror/WJRKhA+zZfmJUbPHHmSVlQUlYkc0aj8p8v8rRIe
2M61NYsG+bGXHxE9WKI+iFLXHWw7awC4jXih4V7sZquLJIjrgbL82Nm80BbhtAz7Q2UpUj7i6N8U
1YI/6Y4ayK/PlnItE/v4kLnhE7RrDxnkBPCbI5O+dvEdaTop5I0o9PF15jxIj3S/goEATjwMvGQx
eLrWl0vtSiqQCM/VaMvLmAuzO7KEXZAPhy4nhccYKhpSxD0ocC7Ip9CE+wFu0+Lw/qJnZPDy3F96
JmkrCLvJjljyWujenhoKEqF53ty1T0Re1eXslg1rskH+Obrbr3SjfVzuds5RtZ5xNIk/1YWsqlLE
YZFTiZk5w//uytKlq3ph54So8NQUxtkp3+t2RrskDJfloVTFkcVruGMWfcn48irJ/kNnuTJYl8Fl
/x17lJcvVnvP98Scg1ZxkDufXxen83X4milCcb9jji9waeKa4khF+MSgGNhoPXeVqAwCym4NF7NK
BRuQamd9X6GP7oOWt5I51+cTuHtI25ldZ07XLoCFwGH2KWZUf6MXdmCME/jZdBBatkrKVlUk1YEU
fFrzgHKE5ne8NhLWDasW3Brd/vM+lUGivtOIXYSKnE82CHJGb/iWZZow/pgqbhiPPEyd+8uiDD28
93AKEr2x+H0zlemXJk1IiHD8yVid0TgReT+VfBxi15vgwhhS6esexy5dd7UU3yFWOxovo+weLcrz
txE1xgk7gnyWg7pqhvW86h55PWPcHKb+gKHqNMi2JhQTigWwCpGkFoAaT5MzJhQRk9ET0P8CQ0W8
ezHZN5wNos526BjbpnuFh89K+cZoPXb0qm8WdRAsxCi1xXnqtT2eL59s+mIS6alW0RqspkaSSALd
inFp/W8jQX85G8UjCcDC9d1rLHb2Fz1E7M5tafrZXDfBtrkHPoCjZftKFRUKr8Nagg1Fo4M+gG19
gjPzWNDxwrK+WWe6ORnSza33yzW8kkb+xrrjqMeqSdXfiVrS2RLp361nQYtbAWghjbwPwLEAoUML
nLbxs0kejbV3u05OMJ90wztxElNUFMTSRiJ3XIa4kiiBT0E4OJPMUQTHUx5YRUb/ceQ4OqPyTCR+
MXQzqdIrq92swgrFskmjECT7qcbnc7Gq/FieXCW4T5DfJlSA6eSxBV16vYvgsaQD3EUaaetSJe0l
q3fDN1RY7Tc4Is+j2ML583gsqs3TRq/hD3avBvkTwcS5OX7MQFzQvilCuV+y4/KITs++MAkWPW81
alrc6kX6TVCi2mnV7dcQzEtCi8rDICEEZZr07ut3iIkPjIojdOY4sY1F25xUFpNOma4PFgCB0O+q
0nxaffaci4EgSA0zU70iJUpXu4eFse8DDMGd5tfUDhQIBXGJjVIVLGVMHgoJCfcdBhsvvw/I1KUv
JNjsPLFFWgwW1p4OWT3MfuQ9fwjrwWn2BKK+s0SmoJ7feooXxzRxUx80xbk3QNtLWz22LM0v6QC7
pINh2C3KKMBUyALK08XEs1hbe6LHU9DyH8QhrThduME+BX52SDXoX8iuHvFAFSyP+MRrwgAn/g0I
bJBQa44SvXIf2i1RWHrii/zOj1edXowKReZEgw9k+vZeV50cq5DRu+Gqy4Uw0ZbdBaykneSuSjKa
Q0Qy9kw/v5+U+G9ss4z7mpIQSbP4tToswXR+4gTW04FqeUyv+TcbUfdfrhGnsVionGhrp04wOD2z
GKb1gs/f04DHhww1SX5Mm2IBPcL6HXB8V3QuqgJmK9Fe7jUOYVLxJnYz3zf0Z0EKrXBCliwc3DwD
R7mJ6a2Uc/ABcEU16XuZcJ17Do31SCS9l2k4NnkUX6c0j+zAGpPqhdPtKZeybrXSsiizykkrTJ/n
ZfcQVysHWVmDExPTlK+nY7w5DXnH2fcOLbo5OqmUe/CeosbwccBQWkhC2ZUZPJuEYiPwuGA1FpYV
F215Y8OpiX0h3HeTQo7OxWe5N1N5gIUfPAD8TUTsDOX5QyJRwLsBSgKHGi6Xm/eDu6CaXS/5CZKx
yexpDtZJmYgwhVlaDSWDyzWpYE+6DJ3YAcDkvwNAz2KDFX1ZU7URgFgjwtY0fIN+fCebnzuk9QHr
ZZikAG6hwHpuOeKEVFeNS3MfISgk3Ju9qfBC+f5QDsSoe4Q8cMBTJ0r3fm0Ru0XOddF62TvocWw1
TjBZ7xLzXo5nsnsg6z+38ciwcA4l5AR5fs3bhFoIE1xkqf3ojwrWAWlR3kETB8znB7TujSwmFnVa
ZWP9iwmliVY70oyMv+V3ZlwwINKS83voslHFPWso1isXNOUpLjJbwI6rXfrwTHG3EXGNDnWDKnQn
ptNGMxwz/7fvBXvugNcKztGPNRCNmO9iQk3NVaGuYBER+mbuPNI7NMgs41IrFXGH1vB0VSPuHd0U
hp9rEmBvaJsFk4V9wDg9lf9d+7YQ8089zqXW5mYGT1ef+DQkUKAjNkBkmWy90H3ENjX6SSf0hR+u
m5/d2zSnRa98lgSdvTDbLxdbPWOM1CuZtS0geJ0lv/glolAijFBOVsrPrjBwMCffWVig8tuPkJja
7q4KvaAHwSV/NaZLb+R7Oo9ZkuyZ8N74YrgJx3Jep1bF6HU+BvgLC4/yrswHAZnYcZCV1Mtky+kh
9FB8VfDSlr/e34j4/fqPkaai5wfFjN6CG9LVDMD8Q/0wEH7uDUg6GaUktodhsmT5oCqMnlyYcvIG
3fvLEm8arP7i2PpGF5NrgYrcizHCfCWUvUtJzVPWQ/fopWHup/+M/DOMg6YUDhQvaf1sm41FdGUT
mENa5uVRqWqEGdhy5sAotIztRDJ4LWSD0vflkP6FReOLPrQSQs8GBT07kSt49gK9r+VRKlwSLMcA
drq2UDQY2mFmxxJaZBWhwHKk1gVzxY5Qfa8id0DfPTg2ohq1nVITKAgbMVrGbxxP924nDqO+F9UP
Y6EVF6i/NMUPf+P6vuTOrUskDs/r3n+qiol/PZ+HCzKEMy2nBYRrs7igiZ7Qw8nuXOppZEyprGeg
Pau5nmAxDNIiaBc1sZP2dxa1BLfFZryXq75sphyDM80SDK6cL215gWmJ8D77JIr50g+pnmlc6P+n
14TbhHXoW7S7yuXD3sMPjT1ky7DY4+NDhH1cL4wdoe+VF1L40rB9fQ9dRLzJ/L5YsAV4B/+PZA+u
ToLR71x+O1mumlSA1blt8BayMZwerFO2h9oTDrQz1U/uLr2sTajanoR/cs/Ny6qTBP7Hlq/KSrKG
4Tv5BGBJD1UgFBconFCbN+2OXGHcLB6GJtBoY+cpoKskGhHNPdk4uEG4nzDozaXDK7RQvaPlq9c5
/shdbZ/tnXYNpfqVNIc7wy1a3iiJzaJx833hanGO5UijuDsFccjsiWjkHHXf4mAO1CE1HLy9v6rF
JYd0oRP7qsRWGOCUkruwGzTFLF3h4USmoidxtqvDOyoKIZWHQ/71ppbKr86WHRLF2V/wYwM/MI6F
GWHxAf4s0lHV6lLVUS1uVYu9xblaeIZxX8Ub01nvwdnE3iKK4sFmDcy67FeysaOdGIxaGfbmpSmI
CGDuTmZv0NcmK/2C9BDaoosxMtdQZOvM8NMYBgtczvz0oBg4JzTwlyZkvXaMJKFSHfTb/LTEtBLj
MPO0ajZI/pDUz/tEr5R138oBwLEBdS4d20w5uuU1MIhnmnFT3D5O4NTr6dPtdvb3MRVdNv7nR0q+
sBrrK/UXJSSPHquPLFwQmTgBWaKlhaXFw7iOTS24nTXugG+clJNxcrqxrYZAyc75hQ3p5oM7CVbA
vYLZuzy/EgNH1uOA2MR2kiDwcCFz9AP2K5kmScJuIkFQmcZsdcAFVTE1dM7TS99MXP1k3YOPydwx
st9GyWbgi6E+BssCyxmCs+H3hDsoS8qz32mPEKUHZ00McgGPM7K1Wk6GtEqBH5P+BOtPfI6HJLKJ
uIvpLwegXIZ3JPT/EJtJhvfq6zABcZbRoBHTkAxuqmilCXDjOLwaa59WRUQu1M1hn32t/o8mKxjB
LjjqaSh5NHZKbOWElS3oRRecifTchDPmFh1tNHokXOE6afi1UUvXNHMF7cnjulD2clOvesJWUnM8
CkEUIDeTs72fQ8weynsemqDyC2zJEBClpy4oE5vb6zHkhVf64pn/h58U2olgP+arrroePjaZ52FV
+L+3IX3aMNEhFXi1vWYa+Tatkyev+GzdIhFYBNb5pDItW1OMArj3NsjI2uKvoY7pjeN2QpdGLWQ/
UDgH5o97pZ+7mbxgp9y0CdM+yYpBPwsFBRHWUFlHcsVRZJ/t9GJ/zqFftFZRqcmvk6NnBk7oKlYS
pR+N9PqYqdPXweagL2DgSG9CLtbIuSIS9vYc/TmO/Rdc6eBWz+pqYw9JI573mM6+P4SIowpprwmf
5cn7ewISYFB4XsVXvkVNT36du9edRbk3hGsSJ7oVW7HPQtwV8v7COawNaq7hyb0/e6hmJM8tDXLy
msFhk/FrgpG96bmptxp1HCcvAxqqkyBy6RHyeeAZELpRVUTrDYl3i98LUZFLnoCX7jV575Zh6y4W
VghHkZjkW0ruXsM30w642ShFRovEHz5MHpKZQfqoSC2unK+rszf5tFuSo/cadKrTD8bqv0Gi0Tlw
8Ap9+k3IuU12xURTntMgUQfbmmPxLM2Xb2hTTmDlguCWlBwx68dYVbQZZyI9VtSDAThxXFDx/7n/
PfLqGNUUTWqaD2Qk9XYleoZ8kVvaZCtzi4wafsfca3OhmH/MAMgfZ6KFEq50A/Do+b83K9+Xcuxh
KabzPVBAPgIkcJUcLJAxqNyFByISgxTk/5RNwA54OYvnJWcVZ3Z/wcbdKHMeuIugtayDtGOBhUBW
4YMh3M5c0bD5Tp47il1aspGxk5T9wGXUyvcLYucAxt+aj891ksOKKShBsiambGRqhDB8SdBxDgWg
9bNsyUcq/7GBK8oEcllNe7iXNPDv7NljRhOlbjRnkZzxJUPiKAMSbBbIJrENw8eAPazuhykc42kv
noHXD1PUeR+Bj+T4lc7o+FIggOlOR/p1bgLBrr8VTMrIKOXccLIk5A86NY9o3tgQf75AV8e2lFBZ
oB8njhpK2wo6msEVy39ToTX+Hz000c2JMeo0lTE20AZ4+435+wBiNaw2fVyxVjRlYeL8doZC8KKH
Is2uVK0B7+OEIAKTOErHfoAAdb9hD8FCJIasdO21hXR57zIJApvJfpiWLEebzOkFgoh5WpWVjTtz
4RqLtdtCddQCuSno5uNauMfSQAUD4YID+z1rKBQXNymR7P77gDmsnzvDkCqYzgJcVnHkKpODxlcl
eXVnIhY02L467WGI0xq9oeHGWMonR0FXjQMpDD+oMNDEtcrXZQFgQ4iqdgHMo+16a+PwEIaLoqoY
Zff4oi0fKIidrL6vZWcpl4Aw5PykCJjMrwXMGbritKpgmMdI7aVWr7nSDv99Du3q0QAGqfplL+14
DZDglD3zh1bLCK/DAor8qtWqH/zrQ30LFZ3shlEGCOPINHll1plorhXAtyn34QoW43dDcwhZeBjV
cWMfMrtr2QUTAdGg1cBj3HkI/Jg3ewe+8ggF2Doq4KBZ82otNRO1f/otsK/uLvue+oFGIm3/D6Jr
ltm58+6yqKUK1gsq/EW+6Gwo/vOuKsL9FIK1RySuNBrguxbNZ0+l1tVMKbrkcV1NMhH/ESplIs/q
oCS68n8jDuAprdFdrrjpbaz/gZQFseExdKa4aTsewju5BMHryDs/gMPHuqg2R/WtKJ5avFzGLB8+
+5oAiFOE+OHEIDOZKWFXhIJ2+1D843BvQE5gITHN2DnpqPmk72Hs9cpE9aIqG/iSlbMvLetQ8Czw
hBEi19wVPeeyNCbORa/0mOXhZRG9b0oS1FilNVr9f7i8cXpd/fr9988erCE1WNCCZukiuXZHKHaU
LIejOXDeuZTq8vtG45xD182AtQ8CVcjgaIOBITaNHYVcYk21W+ln/P8145+07HLtKMpU0XjoXLFu
t7bEQuP7vZfWb/7Lhd/ccRVW74Do9OgnUgsXhl7iOZxHEXwK9H5K0ylWRVwv6oapcm/aXy2YxtNO
DZH6xmrP6OdR67WjOJNscdTKGdWm8dXcDaoaWNOYD7G/XJUrCnS3tmdgoiBaPWHj1fIgVr8WmQsh
pQAQtO3aGRlkBL9oY+i5h8i0KBr2nds/fFQQt7Mfd241yD8l26r6vDGz3gypc/+W4VELKD65uheW
B8xj8OP5X88FVyhHfiCeQs0qyftkF9dhG62bCB/wtAW322qy2x55IAY6q+kKrfbm8NcxMrp6naNY
Cz1vn8JEsIZhMpgHF30cEDWZTuj7APMomwzGjzme2UR8aU2vBS7WANpGCTxZ0leg+5qkXi+tmeiW
DhB7Xog0gx1Sauy9YblBCGKoPuoq9X1cYVMvbCproOL+xskHpj7NCZLrpBzPuLMs8x5L2NKPkTUC
xGTJX1E8pfMmJCN6qXsB5wZQkxakpCiF7INxgIIZZwORO+hzn6dpmI8AT/zXW50X7ppoQwWdo+Zc
QnHZoqnzCreFM0eKKZ5a0qEK3RSZHul2qKm0+wKWvUDBNWlH2/+kbx9ETKjzNHe9iG7igp+reO6b
Tpa+QMY7At34UT0hzoYn5UOS/28/QVchVLPr9x54zLEv8Vo64WtWxPmJSwvbdWEHasME8E9b+Mfu
OsHSmExb23nHC5Z+2WsZmganj6qy+daIvUVJhU7EJber6gPwPS5baSbs/oV2VCbGUBtTIK5agUdX
1vE4yjMJjQrA8+Rq+lswg5Z+OAaEM6IUT/F3nOR88rJjKUix10PiOcRb6RV5AyFkLwS6cpbomoB4
02y5P4pzqFCud1JZJ7WWHaoOk4EVjGTMuPuWm89wvUznAvZTonRV/b8HX+fp5l8IQ5p4jliRtx2B
BZzGPEWdbNyFPcaLeZR3RsB7CA2PXGaohshaWCEjILXbc+iPqn8uytCagU3weMug2U2kfdLCNikK
PCygxq9uWFAdDoPKBwgn2SDZtUfvu74mS9CpP4VHMcXyXim6G0JicBK84F8x0anMDDM36Dwv6/Lc
ws7mG9rmtgLv38DusLh+xRZGOVbIpFUGfhV3jIJpPl7hjrms3khl0bcnea/Fbh9hN7WvyQg3vqc6
+dXURJHEqk1Fnib0ijZjnaTydBjBOPSPaTYQs81Pj8baIqIBQpjIOk3n1chf/ediOleCrEgRhRVI
O9Fc2jLNlXnt8Za8JyazeEr5dQ3YNRz2GcB8zIwnbxwbcr88LXqFwqp5+OIpB1JgaBLjJMzzeEX9
RHFV3cGUGtcxriJe8erZw0Y3hpnHURizJL9sbWnB8B/RDdLAb+OfxOQEowLvea5NKcasaBc+tbRM
68vqNWe+/8gynpRgt+/gz1VmsY2KyCyuxEKAIMmGx+lVZx3zM7gKaU/irzT+RC/FMiVCWXFS3++q
OJid5/I8P0pfDVTpgQlWRvEhVIY0AzW96Qfam5qG4+EG+3Bsc2gi8m+cR21JUg37PCru8RuAqjlU
XGvzTwGES4ezsqFEH4s7sF6GuR1TssESICY8sgMz4kEyv6fK/HM3zC+AA5TlGFdJSr1SsV4enF6/
4o0Oh/yF5ccEv8stQeTeKR2juyQ55f42azgaxo77WTxKGD7kFTLciSYSE98vu+i9fkSVgMNzDvZN
GPp5e44zhIaZ/7icUCmaH3WgKqmHDuEJgQzh3iwbEwOtr8a46GtJhZaKzCEfBH1nkcnzDC6o65Hi
y48CVSmEZ5TDiR/4I9t1wxdZAx7NpFBbDbIfdWi4kI1WLo9l9BIftX4L5TiTmBCe/kYudI2xQ15t
IYqARaIGrgNbR5I5JbtxNU0q1K9azXD4t0r1nXkPUlNdSbE+r0yzscahaaMvpDLVLqJpl88z7Y21
cqqqPeyW/YzmlCYY1vP9O9ymRoZYStpk1mt7UfBjPjSWJI8RGJK1kLO77EyrrREFMh0HmgrU5ZwE
o9jsTdOY0/5aWOOfIn7ctotjT0IFZNZiy7hPq6jRKwIRY5bpg40OpxlvT5ATuLK2rTdGLYer5DAc
hE8lL5RuG4KGKwt+RBBPuadBwya1/IKjMkKmU16bLJCDrRqXX/vDvNu6bGm8fRvaez5V4m5FyOCv
N/NKqADiiKwOGYOd0KRoDMVZ5pYPdKCk+tUQFyN4IM5xn/EdjMOdpgL+alWOJCRlLCaLeVLsQcKc
aQVXSPwBriX2575QtikXDN8dUyEy7eguKd3yNMnAY/tBRGk18GIBOK9+bvXwGqaTaM9eTMLzR3dT
J3BN0XQgB9HFPzfkwc6hMVLDj5fyP3sLS1L0DzpUAaO9CgepPwTgNbBU8WOj5QpPDIlbrx+sR5Df
ZlorrjP7zuCgEHuqrOhBgE6AhMAqezGAJnFSkK3TYY9A1oJKPKBx4YB1NnVDU7hkPuEcZ72roB/g
G6nwKw1XygW/pF4CT9PWq3nZYv8TN+ry+LTxpZwrL3BSWXjE0rRX934RWJP7Pys44AKZ2s9vL4b1
y0n2DknIGXxrWg6QvnRNwJEsHb6cKrHwIalE/jg0LfJz9DvGuQAkTXFUAlhzF49Ajoc9An9ruf7p
eUZ7vChimyt4ADOptv4t1drfj9dh6Kh9RWkU9W1aoY+xlAEzvNJDcYpZhBataYV2k0/S8ceKzF5g
jFiPBfU/KCPZ3Xlye4XCqUOR0zVUJsDFhdsPBjfZFVqpmHuYkD7EItRxtYNLX8Wf4OVU4DmVGk5A
cCbXQM8Xqka8gM1T/3BSAGRVonJXTehwf036xGSlEtYzVp8QKl6WjbJU5JDCo0chv5g1hwlKhy6P
uH+MkIeSWxy15q3pWW7p3ES40D7KgLPWfgGrwhg3IsoiysVe3jkTS1QlVTfp8qSNuYK/tEpsxTC6
8jZM/dkZ44wGf0Cs91SBCFLl5jlJCMe7zs5W5pWMS7evpETIa+SVeEzHBXoGpXHQuua3iP8dm/o5
8sJyKwP1xW5/R0n0bO3uBb6wGlHX9cm3IiUf/foQlMh0ujn0mFDo9qv4WPEg6YlcI0q33OZ1oazc
fUEuHmSAGbERb3xAWIiX+BCCq1S5e66jmYhGMAZjHfWtzPj6g1egiXZuQsSQ1t3Oxnl3R3mlnH5R
EA4RQ2kXqpQdV9CYxy9JPOygbrq+ePoqqRW33JLrcKDQcTkOCSzQaVNZfTl9KIZ9zqO3Y7u85CiT
mxqvLLl5PUjoO10JEZmKI0O49DEYC2ifWD719vDcG/O3+oE7H1YRbRXGbIQXDWmLvV1dnLzSZYm5
0vjHWOfOGGFH8pDstI4d0xYGrTbqM+RiEJm2P4HgpvGRi4C1RFRB6Jltvh94J3X3o0bJn5Bs9c9c
vkSv1lr/5yZOlyFW6eidWKsP1SoNom0cbEtRgOo0t5mWycw1jhXXdPHrV0dN9vN0hOpGVR7oVeLo
vHRg0p7n3XGgN3xAQXI1OLlFOlDoUz1E/ubETx/arxaS+mc3RFzpvaS1K6HoeEn0BUs9KgBuUMxG
25WZvt53VoMcp8e47lPfYk8GyUb6cRD9dK+MYfQ0k6un4CPp4OXL2/3ZYP/7H0E8XC2kw24GQsYv
1ZVW2qZ1+TH1h/cjj/5oVa2/GXbmBGyGDANooRQgyQHstLx3/67i/f42pnIfe991F4NZpPDKTd0d
8lZnYz77zVD4PD34IRVMfu7Zsx4KWvyYHnHWW5YHnVDsoiKVXCcRt2yz+ufFb1H1riH44Ma4bhqq
BOVY94zoeUIjIUscQIEPuhiS6tKwKypk4y48teUEpvKPOwtC1fyQV5TnW2zSBtynEYsErCH+5RfO
NNQTWOpwlS2W7pk5xCXyckpOuuBFTLyksjNVje8hOZHh9H4QfxBPI/X7v4pompuH6MPaWsMrvG2m
9z7H3huScCw+qh+hu38sDyafTB/jHlwMjvuTe5mQooPUTj73LMsOoXc8sMiQqI28dZKQvfil0eyH
h9DOJC2vmuc4hFkZqInOyPdp6BuxjsICWRff+0l1Cb7/gWRmkUc3Y0YqzYvpRciw6ueD4n9UdBSJ
Mz66eYbbC4s4ctU4PdT+bldM56BRDOtPhUhdJnC81vx+J6/50r9XQmRrNPI0EjtFMML4+kzpxXsf
OmP+3o2twqLwBUv1rJ3XLiBHluI+61gFMRUlYJijdFyvCJlcl3NkayMIlSaSxYCtXoaVOvVaoo37
MwQSFtgxgDfZtIF81CpJjBj2KrF76BpPpirgb6/WskJa2JdtnEUTKlf+Nqf/wp68Ds6skXjFIFE6
U4HrtbSU5x0FotaJwzA3pVTKD+1Oo7Ooi0D6GVbIp+6X2mcOjCR5JtOD9A4cNc1NrqzS5IbfrbbD
kc1f07MGaF6H4RyUuK/q7d81QLWDmlwp2yQkYaEYCyGmVqftagUyGA9x6OFr0Ihv4Al23ouL3kee
0BKg4h7+yGEQhuIPdwGh2QXd3pmcul2a4fWy/Dj0ggarKHTL4rpF8v0TkK72X6a74WjXhKxJLG6M
EJ8sDkRxOqGl31LaLH4tJKYTEiCmLcqMW6hwynKV4mpsIa1egdoEx4bfjX0utkrfOaHUdWQFQzl/
y5J1bN4JtLOHEn2qmxb9e5ASl7Vo4rHuc79MVfT9V/eFunKXmW9fqQLfgAnmLFn0eMqBdOQb/MXg
C/h9vcViUN4XLvgn0N0OLh8nIIlZP6jcyuQGkZSoen/0eftXayt5QCDtD7SDXKmn6vCgZVSqjPwW
HP2TLNYgICepp04KZjnXVcy8biqUsbadLd27w7vMKYI1f1p136Hl5gA/mhO+Kdt++0vLGnNb4gjH
t7xF5+JOYIauyn1zljU5b0ftIibXBnUOg+9S5+MvZA3m76LBdX6/c1Xv3+Rrdpp1Nh1SQ2nBYehQ
ooa0QymKh1RFgEQYhNb0epae7SwlxRp8KMdoBSJKAK1xOgiSxNT3paYvb8zz8JDQN5TdvKmscd8o
l5JiPtPmbseS1ZZ76qMbe54LzPrEZh/V7sIM8UErur3xviXlN6hrVW/hLZZh4Q7yzpIZjJeAowxD
HYOeCtGDgH+xuk38NRmhVoibtnQy50gc53x1BKmDwEiGFUUnjUBOOK60pZuKMaVMTUsPHHPitn5f
ydfR0oes0r2HF15XguRo8Dj72bZpbsT+sMT1l1LTQcnkd4S9Q4dCI5lyn3BmyK7pWN5DzczpXOwI
x6r3vCcTfVkpdXguxyjxBkvOuF33Vn/jq4ZR4XDf2RKMGsEREozWd2iRL/TL6DrcOHgTMaEgSIrP
c/qM6EzUOioj83Iw4PEqn4eXHe+a2Fm42OZtMITWXExWyKOit1bcElcjwBdTBU9UdCJia/EDmIWv
VKMZUWi8MFiwDgQG0PNf+Ijb4zT6DuJGCNrtdpzCwMc9KQve3+Mi4pId8cmN5GtwOxm0RFZkpcAD
qilJ6sqUUbxzn6P3s8wxm+vWJdQ5POTxqTJyDmL/3HQ2N8dhr51fiyQxk1dWtDSgs7aTqtaBuJOu
9HWb5Z9J0S3xRxdKn/DVZc4gXC8LN71QnuIRLsFHSxsuDETTEZPx5dIc2GNRsD9EnpC7FTSGh89Q
3btCLsHJyJ5GUo/oKgXe05qm8PceX2lPwTWptZTzPsgplRjF336Q9JBefA7ENRj6EYgouwYr7ue/
4MbVdRn4jMtB3qDFSrBooufII9RtE9fZKkd3qckKz2o6SgtZFERg9vEUeMEyhXON442/0vOfs+Z1
kX6+O46ECxbTj6atUNwwsxXTDq4RYTHLT7y3mfW/ak9hQwMAAcwH4i5LkwnQHOXCuIuyWYED24UE
x1d8zo4NsbMhnXAsTIIWSCc0LgNBiAqOhBxdhvPYAE1V1Y0DQowz8MdbOnr40FRWupyKBTfKCl1Q
ZnZme7WaECbKTkctnwhNfEZ0McsJkmL5+60X7IIeGt4X6psvNTZGL1a+6YjARV9dSJnZpuIJjjfw
PRxpINCRCpegM8t1DP52018MU1koKZDERCvaxqx0g5xhyXbO4KMEUWJ2551htvCAEsa2kVeMHa/H
EmlezKIGAOu0etP4HN3NzNeXYCyvh2zVFdYCaRqOGg04IJGqy/8CjFAVQ+lMQ1CtqxP3GAsgi9Z7
H1CIlwp47S76cIFoKsOXUC/ZUQuTCmmMmiBNPXoqx8xn5mG6uEG9SD3swrDtMsDRistLO0JI6N25
EcoVGpk6YZJEpmKtcaooVoEnLWlGQXG0P1dYlN6kZb41zWWfd4VQ7QsEQNCWjSOojTkbmX/SYMMj
0nGH3C20/9egB2NFi2bv9mTipJcq8/Hif5SoNf2fQbiu8VzzK6KZ61UImXEhaYIjb4ZRlqPoHVUg
3VeX7yms2/aSYaQcjcB+M6qS6s/3l/MMXQAmz/gKtS822Ji6nnz7qgOVPt4bhSyZ2jv5vao84ZYZ
0ByuCUgf0RMPPXVsWsKHEixqB7iL6XGUU84w3bHbssWvkRX9xWtshtsUsUgf1Q9R/wJ2z7Pfsin9
1h2gJEda8XqLYqXYgU9W1UgiAyuitgINuW3XjITXwbiX11YLZ5nbFdUQOb/k9dk6JGpD/8gpYL3o
MlAhc8w4lKbt1LbEPyi90vkidgIRcf4cuSfKIr6TudMp1Rmm+pE0stNq0AqQgRTC1rKiIWgxaiZC
ifvi9UsvpOdu7vA6JrjcUeL2fSl4cH3bTUrYiIneG2h9eAOkS7t2L7/dWGtfXx+TULVasYopVsl+
Fw9Oyd/C0kEDF0bAk52Q5WMumUjegg76HkEzwfrCUDowLYthWA+e7w315wNXvgeqn17BEX9hgnKo
7kUfFL5y7hTpvolmsxFidPa0Mq7sO5PEusbbElgOl57/mbV5yDiWbt5wuxLfn7UQo6mpd3WxDHSM
tb4VCMx5Ra+L21b5vcY0k74U/73uabfdmnR/02gXM34sMSO3NFsUVRrw4O0TP/BjGG62g6DKomt5
dY+SrWhYjviSIc42vd7LREilBqRnByJcgr/w8swbag58J/9hUvY7mTAGwpXjEF1g8scvXJQaXNJF
Ve2k8Qrv3/AEx3Gt0106hnsQadxGf5jFxmS0BbiKQjtgTnR94hNe+hKV7IeRQzIOqzm8D1giKdmL
AALDsC9xxVJuy42b8WttWiO0v+quXibYQrsGVduVFqJQvwmNwJeBqaR7tpyAKOTWOKM4cGdKGDM8
7GWlqE8NdUZ6HYYbl6Kkqn/p+uDgmz/cj+45aKLdN0xZVrHagXi9tCfkKoU6hAF7q0vzdItsLBgZ
kEXyDvR2VuXebI5tNEr8+iBLcXUapaZjzFMTKnwcOPJqpFMrexilv45iZwfbcJC9J7Mj90HjbE8w
tFCre73Iom4hTJSlDJWjPrweFWvt6EE5ctP+3qCtsVSaqFQMSDBAxEhZC28cv7qrTlxR4DHJxs5H
utbunWW8ozN9N9SYEUBwlPU/44Rce3eler/0HuW/zD3rfot4IlJ7Lq6qtW6hq7JOlRQlz4Qw4IVy
LYVOSEzh4TejgK3eg8B7vcBsNg/p3gm7+WIUIkxBMmNmxPPMHz0fC3cNaE3zDTGw129k+Vh+NsDx
kvi0+U+ItdUfoX+VMCnZqc0Dg9m/TW/F/boxcq+KuW/ooVxY/ENhQkq0yIh3nNMtVY2/rY/2zIqL
p2CfovvJnQmgaYixF5mVi6k5UXwnRzNt+pDZWeliuepbKFOfBvMJQSbxKmUY7Lubw5NPfrGuCBlB
5LgmHwuKYTF3TbRWSnOK79xCTNXezQR924d+jPjMcghH/Np8Jxp8/13dw8jrzSvB9SwJR90ZJWYo
YF+SMiahgOtsnESZxZEpl7RdqnospJ4ctqBQqzdWFhNyBt7YBaGB5+99DwhsxZLz/OiWdNaHK+fu
nAH08OUVfdOGdzYExXoAccw7JZ2DQs/D8hgquIQBj5qqT+jbu48QhkrJUNsUXgUKrOsmVSvoJI5C
KsYdjJLAhdaySF2rEHQYO7Gi6RkKA+FWft5ekv1fBfwI80Qcq3AuxxMpNZp91reXnMVwFOG96sjU
5+jFyylpOt1On1sWehFX+V0jDrb5VLxC2KA4wpzIkchTcFeNCtyflbDs0CVSKuea7CH0M/W+yc3D
if4uczn2S2XW7Api3mOhyv3PhmDjng6uH97y/lKKHMEly4G/J/97BBqGuM07jqTL5QwVMZjccM4Z
9M058phfwZ3Y/wGKbNHRVCYXCoKimtzb86VTNoWruE/IEkkICbfZMDrPw8aQYk79Jfuu5SjqO9Sq
TxMc7ge7sNvfvd/Ke7IpejRdsiH/Z5qBgYz1/92PjSgrSO0kdXFbOsCZWFEAZ22JMHq6uXNqoo0f
Pehgp798BEZFF0ClX24vPTK3WQ0OuacgYtbT0DAIoaasaUHj3sCN0qPYyaS5CnwRH21P733fWUbe
B5CLDC5+MdQaUEwGEGqS1+7UuL3V3qyc3S7qOAqHRFEtGKHxc0lxseOlt+VDCazbpRClk+DiOhCm
l62fTdxNdMd18jX2qnRZvn1gH5jG1AqJqim4zWcYvstFzyOgC/4MOf+8MBte7znEbJrtUE75oA8t
0pbUvdy1w9QCON8A0gS4iZWzcN7iBS9liYOXoajNz87tiFYUgODLzO8CQhoSN9bOK/ExbuQizhor
5AMDPBtprYXu6chQHj+ugl3nuWq2oB6P9dGkBh80ToGth6FuJsJuNP2Db5xnnzeA1eBmQQrz2aTz
dD2M9YRzeeGNLjqptPA5+qmujtDG2sOZyCUw+XyMKcf0FIvVo54or40jqfbV7yRk1Ef4HEaW5+Wf
6OKkBXagUJyfwjNGdjRgOmsSeW9m8h0HEgFgGn0WLqell2Fw11hFuiYaDPWSY0EwHzeogQUk/zV8
BoO+0I5k9YaNpW5qHFdddlXG2wJpgiNl3/Fi+XnoBPiG3hr8sN24kFBpHENM+mreHqdeD7wgR++P
w9OAKBKala7giWOv6UNADSo6wTIeO17Bk43n9fr/t75fiuHCLjKX3BBP16BoKIu8jr6aH+uBVtyd
rWE2T+IxlHg0o28yPU5w/oEms9ar5tNdcZ4UnrPey/Y2w+ZyhBuFPUciE8IYAcKKFUfNqP8+xSq0
/PAsmIR+OpSz3XAifM+gxab+4wVaWvHOyjtvRu6T9v4Rvp/hGfQBXN1mUVPVTPF7wkcXLzsVIXJ3
Rk3ZHv/8ETNTfSEj8D+Cpf1x7KKP29wEJM3lkxrxrZz7ocBJ0kWB6k95zBmx0iSuOQEBJR8uGHry
7bmEoSaAJIctuNZS2Bd6DGABNWUfzL2wZGoITSivdS4aOuc6N4Js8DQfyfFGK4t9FXFDvWCn8eYl
FxY5R8xFcwogSXmh7mtGRy/KDozC8pJFR9T9c2qwTfCs4Qq856xOquhn3pAmG3kuzrFLmeUQEk1k
8nBaUlh8mCVuRSeRth9ZEO8SrXHLguDeT2YZ6AAEkWaF9xr5iDlBjzgr8143gSDMknB/Nj4xCaZ2
qBg28Nk+c8JFkzOGFrWIxumZwsn0ea7kwnXNoProdqukZSF8mS/rYG2YUq3DZFL1rA8S7QIpTTKp
tIz8eMlGbrFXtElF7hWecdeKsi1JIxpPVJfGa83kCO0+9o/hmKocq4Ar83WMQGGzyMMoxdNkuUF7
3v+66AZQ1FZ8AH5QNzxtbjiPQGvhorIGn7cGAJRyZsp858VR0gGkfZGVLOafbW0EzaSqM2InM30N
MkL65/YYuHnVGGxFNK7bvfRcMnUWYNLOHx6wITuBwJt5r+Pbh5zcgKE8y9wHV6NTmlufpmM9Lrqz
mnXtYud/xtslpyFR7pHpMQ+Z71L8eRSkR0nrRJ1XJJyQY5nlPNOQnMEn0egVwRe7XCmBxwPtXh6N
+qiShD+bMYkRTUM5VjF8JHCgxtIhE/AEBc+UqvvWPCrBVgMTA5R6w4hETB2pZzJaattxbsrESQJ+
DZmRW0g7p1CnBtYtTh82HHj09Tct2RwsxYl95HmUZHzMtvMN4SSXPntPPtCdeMz1Ckxc+m7jtKwO
/w6n3wtS2mti+7qgFZhjEOXmGW89zFpHPdlFTtBz8w8NcafiSsNCfO7a4qWrkwSdlWcTvInc7DNP
+YhxrwJgUYOSuXeBYoOws2qswKvaA1CV4Y8HxASOlGqhDdD9mczdZ8GDCxQYDKbfZ9UFu1i8YqDF
N9ityqOYHf3gJmJ/8i3mRE//Nozlzt8GVT5wnokAV8Gc5CgwKfcVsbIhKtOGS6dBPxo48CJQHcth
dQ+KofP8Ri/Dq9HTkYbv7sEVBgLmvtNq4sN9ykhRYcu5M2vnl2yIZbpSzL2nhxikdexFlUdQNwn1
28qPTbg+AkyQVqKlYoDor3JixqXWQkvM2pTcuvT7W0PLu+HwWYQDxlqR7rpoee7AhdRyCSqnyvJu
AdYAeH7qA38tsuKg8p5Mc/sIC5W88jbeI0ZCpRSpxRY3woN/nIKvthEoKM0olnYLFBU1CA5ktnWp
KMTQSrkVAnwaVKU3ZBbl11+dCeuq05NZvDaeQ6NuxnYxLKQERjjYkaETwYX4aFMP+W6S/Mc2m8db
hDR+pRWUIiDUes6aFWi/dNJWSRqoDRFRIioHd4PX93qOzZfkk+mtWKWpceB+9lTzu+7ihZv2AY4j
3k797QqeFZH63UMdr4zDKWraW8t4lrTuhheCVuq8r5GWNPmUfOEDAjzXFG+A3lUmp5TWlloW7NWx
Fv+V/TKt0NMP7Ml4jOzdJM+fprFN9QVlUyBLuZ2h1/4Rc0Oct+Qy4oerXFlBIO6PSYz+NBM+Wg3V
kZIN0/+HX12eCfM/nav6xh3yURC/za69X9L8I9MU4O2q/QBgA9JqvOf1qTq3PnK1kqIwrXxrGZiD
bPAU4wyclrStoES8G/NQSneX3ZONOMpqLJjnajnbNXEF69YB2kL/DaEtOG9iJBxl5C57lEG5KQDT
ps53bXac0OnNMxrzOsVyKhjAQjdLCvk34ex/Z6pQSDrWHLw7jfGyLB1tCoX1GqlBJ66+Fft4fiiV
WZOrVjQA+B4s0Q/E8XY5XfYr+UHqMJxAa1cPyndofcKQWVusMcuyM2T9D779vIu00bCoYI/juFQ4
IQHtKiHbs/08fI6JP5aRDrqABTWSchZSQCDEv174aF//OVWOSvOtGs8KP2tmFu1aICaDlGBoW8PC
xTjx/MPWfOv3/sZcmOveekRBnnk4fwAnl09a7lrJi4IfGGXbriL0jrjiduIMsYQIMd/Xk3UbkBzW
94Q3CNi00OkmZKAFJyKhpTQyXBffVIUKvR3aRAbWt8saw4utPhgG15DNZWleG4SLmyR0RLsqe+BG
Xp3fz3IqWN1cYjKyg2Djowmkt5sXji+ntO1NYgDqKlcYMy/U0N7mJbjqBbEnhNyMzNVogmJBFKi7
bQigIDfHgvj6ranszi9FlDUsYZlhmqf7RcYFYQIvHyO5RHRbbo4l+S/OdOWUMDv5hYnK0a5iAl+y
8npz5eVXccqW9HkE+j0T2WoMq1L7cLeiIW3H8DsmSpPRj/Xrs/wGNZLH4ZJAaM2IRg0lt6Dji7sB
N/GBow4mh1FD9AifczXJlJxulrr7GngOXCUAlcHqjJS7Nq7nDm2I/tse91oBE4p41BP0MjgXlkxB
YN6Z3vqeV9Mj2SjMCQ2i/RkdB578aoRUy2Ldi9vfUXGbKy6dMyN0jn0uoxqFH272K8McIsM5fwbi
PnudfwmXhxRajnb/nuln9QPNPjo+/+MYEsa84MLS5P/nJhVquX2PFvQoXs19D5spaR5vqRPqcyqv
91EF4444BcJ3KiSsZRX6dZSwbrbZ+JPjpKk19DEJ755nzPYNaWWDRHT+YR6CtAaSieA5l8MdI1JS
R8fLBEa3UNMQAOKyb9AMuBn+vayweu4c2TS/+2bIIkUyyP68zc+BAJYTQSL7wgJj0tnaoukMRtg/
4N/7Pv0gf2zUtqkQ1cg60GhMxfFL8ACxkkPMybrETxcYvL6pN6YKu8gpv90665e9433Ej0L+vJNa
91zFcjAJ30Y1hstYgx8tJOPAqcnAXCmYyDXCyP+AucgVyj+0ptv0A7Jj6u4cy/yPWtV2+Ec0VM5m
xL2MoaXsGOtbk6MQz0uw5Ky4YhH9ylenjzxOLADwMXPaxBOnkgNDoyKaaH1XOPeFRMWEMJfaeaIV
io/Gb4J0F89OGJKaSer4WP3dmm4xYFkkWwr+abCxtYea2qP+3y+DeHsQ32ZbkTg0q6DBRgU9ym1i
ZY0lef7NCoL3xhtm6xuyGooGcjDmNvW1tgB4vCN36rWbbgHEHZD6FZUNkv0PZHySlkcH8XKwBPkP
hAUwp52mAzSDefkNmiLuSslMri1v/S2TNeCkO4caA5rahSnEu7/BBZvfqHq4qXvK3rtbj85rTVHb
FBjqrVIkoPJf2IVUQ+4Wu3wBzzfRS7ELFff3KzOBiGsOwRQiGg5AHh9q+kdUr7S8jPJHjMIB6tcT
WfQQZLOtRhuKbNnxUsDtLW4jd59jWqEjslWCFu1nAIEh/6532OdjZ5PXn075Q+UNPxJpCKav3Wdk
OQSz3hF+2skvSQkDJTFDeJex4MOmEcTZo5sAEY9Kde7181VASJtXb3nKjpgLXBrdcsdw3PsIVsnt
Rtdn7rPt/pksiuPrUydm9t/VWnXx9SwUDDE1/e8qlSIqtg7T//gkqj2w0rm+YjSNararGmvF/O1l
A6Vwz3bbS4Y+QYhxVqREqokmsRhS3CBfvQbLApUthovVNZhoQJLnL8SR0rUfiQAypjnt1CyU72J/
DnZ0v6AbRoz9QtnA35/531UNtiJOSudmhJ1Zn99jHFHiZDXwmuDkSzdWspi+B2MNLhWJV7ZmJnHq
TVMvieKVliUw0atTv36F+wA4Axov3j9/N+WyHSD9BfcdrerdJh1kMxA5yWQtLzs4KENbehzFa4qK
c+I+WwFRT8sOYMgnms57uwHjAFxg0IBBtsWYXYDtqUwWlCLMjKfQ3Dt9OtUbAKgEdZKNJIFFZaAg
BHlSZIWYyfAXL73b4m7yNUbjUbTeLR+8l6h76AwIQ+zEHa/nl2biQfkCIKj1JozqkmX9BU3zE25y
QmYbFXc2PmfY3Ps/lzj1Lx2Nx1YQNBU2c7eBbXlIgvuYLvf/gcpILMzbr13kkrEmXH2wfIdCiwGj
cHcP5UFdguSROPxFGQ7k4nQtxcfPCxfpEBjdZ3LbKaObi8dJcoRtiMt9uksDvwfzwFR9sEj0yBhv
uEdLnPJWZIMJ02c8oogq9PqPG91N7AdskrZ1Hy3IVXvmm/1J+8xNDbQeYYlU8R7sIspzWl2CgUFb
v5DGnmkOicyWAvWAuDltr5cUL/z2L+iiR2KmcG7bnv5cb38wGoQ+ayJvdmQ8dcVN6WMji8+xvR7y
OqUSCvCRnsbJ6Ke4Jx3YWPrBFH5O9Dx8tT5bPb4fi5FXKRscMIcsBJSvg3AxVn03He7uGvg1i0pN
vqYjR0p6Y0a/ZGduhQTwEvhw20uuVVsZxsIEYE11FvVvcC8lyB2IUtalOTkowDopakw4DK3zYRGe
mjGyytYEPqtOS31wCBp6kw6stgxQJKNi5BQp9vXbtn2W9LZZfQeqPRl//h/qHfZaGbMQXVXKVnT4
XUGYA9CIO69XwuAlBoxCxXJyIlWnSTsHqwAwhoQePfKHL5h8nVyP0aswjWIbNCKBInUmi9CeNPz1
RQkG4zmUazNPg4iVkcWUwk+zG+oa7OG25p3+EUJh6nY/1EShmXlKpSYPVIwz3GdHSqnr9NXh7kWh
cz/XRHvsrS0pV7AmozK+qhRuWe6dF2QI4MCPeOfp7p5bsyxE0QmTF8hl4glcx//SWw+nGfD05mHI
jyG6Gb439vRuDKHhrFrIcOfPNCPaOSfvRuh7/GKAQrFtZhN35EbZ6rWDN6KWsEaIymAj8OYNNqcz
e9BZjfbVWTWFvWGB2xWgjQM/Y3BtlhzrvxQExweSB6+7/5jyg3MRGHvc4rlpo/ipfEi2QqesNGhF
NBmpshhHLESKPb73qDJlsxlY7KO9mezaUbwBdlKxNdZdTt9jX6nYOd1iQN4W9hTisxEntnR2thRU
ZWoWwpMOge5oaLiF9pYIlrJJI/W+4L1ae0c96fvY2ivdtaKb18Db9eqoE2upl2aTDXquo93w++6I
BQ+ui3GMcFpz+LIYu7YiRomt6kSNYDewXaWr855JxCd0y7HWAzUGAMrl3oPR+3OswwlYBwiYgYhy
oGCakPHzYbNk/STxAUGv7FIXl+jn7DEmM8eOr3IxuHyU65Wpb0Ec+yQU7JLMeiIfmkdC0Yxvq1wx
FuEayEv+5qT1/K2RPHncJe4AuMcBCPcntmwmQY35pBm67nOhccNmSntR0QIh0UICqJdEPnYA8BCb
rvy4ipQT/J3UmJUWQF6RBph6Gg0OEO9gV9oBPF+cRIQD68MKipb87wLMaTz8VwnwrKeVZI9ROp2Z
crjT6zMbQ33I50z6mA8xkhoQ2Vvp87rh5sM8R4u3QoN5G6Eg7u2NUn1GFyzpXEi6GazP7fbg80h/
wncevG/mk2CgYhWBlQq1aCTKAeQOq9QsFNgCD7uFrXsmkrjYOgGRZFKzobJCGFxnmn5u0miS7KSE
UKjg/6w7brzUElsMchZYM2Yb0yu8ho59QzuC5fNNQlKDqxSgIi+X0fStA+JUBRICD5WGEO7A7ERi
rCAg2l/oznr7Qpr4/TcdMyyIg3zQo6meqZzpk4d26Dbp/9IkgJnNrWCMMWQ6jvQ7dyB9Mgo8OH2j
+z6XoDB18Ubg/YdJQulplts26F29M6MnibNstLaNOSbdHEpMy6nN113iHOq9JB+CIuM9aN6xQnB4
vesNRA1wNVjehlqMTDg9Fg1HIe1CkNOdCBBoA3HvoMuEABjhRTMTrNka0u4eyexNjHs+LJwixMV+
zb1spkeFAj3/0K/jK6jPWe96b0A/S7GTXZOikcDB6sDyuNf/Fu/O93wAFjIi3lvsAqY3XsnDzsp2
zIlORLgKaETCJrdr2LTlhqIuZtriWJg7yTLjm9O0sQ/vnpt4q95GlwCEDozZ7ywsiPMc1abTsW1X
x8Y22SVQqDamXjcrj7ZwVQKAOall/Lo2vLTradMBQembsHpfPh0rV29B6gB9xejylxFOJkUq/pBa
EHdcJ1yfJzjxroL86ZS15toMH2N25v64SHduqLFU0xfJUIenrV83oXpOJeVleNvJLqsRRL4ydanF
fh3DvOb3eWSRgziGCqr37JBeuXe35SVDwHMUGCWNRuYN6A7lQ25mbAhtbB4dflqRqHpQg3LbIRHK
d5FLZ1PjKErHu4EB+8rFb/dGGK4mZjgLonmdqvi2G2eDrzD736orDCc/Qvhzdko71MOcpwRdCA1N
qs4uuiCh17Rw19vHiic1TWbBfCahhGXU8VnTicSkxl+C14SiBCa1qc2575Ix+ekAZ91L5lWI0Bvo
V5fkkUdTVutWdIJ69+rJc9tnC94Ot8f2JDIjsZ2Ut8tawiUBHLfNEw9A7DkOTlfJKRDUOJl5Wfxb
siT1N14kXfddBVOole35pu+krWYOtv8n6wlI/gFKnwhkdm/+vU1JW2T3sdbBATuayBd+dDx6QlT/
OqzWTIwoXnvUZEodYdG9BszUSfKLRmjZCMOh24UbrNEfVSkaz8mtjzIxyZ6WdtgRgPpPU+WPMSBB
+cTwhPH6sIgxh1vZQdmaV+h58Nzg5/y557dTNypTLKSmjs9Z0PfRrXW20ViL/0UhsM324er3pS6r
f0juJTBXTC5cSvi0K+UAgOW5hZTOFrLQj3GDScy23MoTYjG32EnDD9nh+AQBLkOKwj8pVdUOi4qf
gjKUFIZeF+0SkoQ50Rn4Y254UGVWW5jrn2qT6lfxhbkdBc6X0OhgaCkXzcgRwWyACu2ZvDjOIugs
G1o5+9obVtMTLEeXqe9PcqUeGSadnccIGvYY9dpaBVU2yzwOorcIzvkZW7IB8BEOXrc/fV5rUBN+
Fpk9KBHlKd1SVivuV+XMwIegPdWacgjqYnX5Cgcg3v4v4yoEj0LHC3ezicn2AuSo0cm86J9V+J/d
S4OCo+m4pd7T65sWgxRk6LETdh72Nd4vwWehDZx1dHZItahPgg36J50PHnwPSySHj6bFC4fZrMA5
IGHEoLc2T/9F2YbGxvhDyw7ghN9RpiCcOqjPTS7TcKzujppMmWTMJgwiYNK5U9djXLykkEv9Dgc5
tBwGN644uFHvgWxZUInI89S6sRaHkrAxs1ORDBDCrchUbJgJO1y505p2dCjYTlEDJncioz7FSt/1
yzaiYdCtdzIMPXyEgci8QZVuI+j2Ch5KMdRpoHo/pUUbm6B1XbNnle2FSQxUCOGIUpecyeaoUSTR
CkznFyZyhJ1e8pROLthPKvwdxA/rezviufJkp1eFKnlRgd14IKISkWjsZIlDvrrs6p278lgcd5F5
pF0uZrQ+nyqQ6TOgLK01rCNc55xFjh9EUgDIYaVymUdVlVphGBstt2+XgUgYb9lxUrOxgPMSMBy2
nl/sC8Lv9EAzKqp5uWIh5LncVHR3x2dfqHyxN/iy7Dxbs+rA4cTdxhz0YAnU4V3L5cPT07ABv9WX
rMM9WUGU34P5T1v0veIxNIAq1dCVxaHJQiJ1BQ04OBhpkqiF+gDvtkTmFL7iXvkGaO/Nru9wZREk
dQ4ErWqd9aX9rkB8iTUnZMta7Mmcyk7mlqiU6AAzH8A5Z7/5iCNHUX3gHZuUyidX+EexrQHAli5B
c1gduGtgO+pMr/URIiKsJMGer91Cd2HJOSlMW1+35JK725lK6Ju5APHyafLSL2S8SAo5hOc1tYsV
Qx+pkBPtVTPuTr8hm2BrNCt9lKvFVdBLzObLOa3y8vCG8NaWuVJ9IJOzEdx4d6sW3Oc4qL2YsjrZ
egtvzLtuK2ezCTj89YM2LAnxrYMbjKKR+a26YgfleNdlz8gN37IxlWdiposG1ERtWoxyC12VB4oe
5yy4iyFBE4iBsLi5bovT6MB0ZbcuvzrPfxNhMeoDK80lAY3BsyHGFfREjv2AcBxj/Txp/jeUmhRi
lxpcjkjodhs3kVyUJny036sb4DlOUzysDZMXnAYtd/3B2gyWipX8veHAVAeBbuXAg++pinQLuuUs
wAQZNChNbxeg8sEhYtlVqTzEwhcigJjHBvc/pGsRgY+pomCfAZ5b9XznHi40WsP9bqD/mWx9Jcx+
XAlmt17w3Z5J1qiAg2fwLXt0ucP2CLcD7EdhXr0Mh/zxDO90AiThHeZ/Qwl/JqsYK6m1U/XeL6sy
2/XXE6yAnKTdZUKjVI6ujH8y19QRp0J3YmBVcRWqQP8YSL+ibln0kDH+XJjNb0Qxz30cLuYd5uqA
pMsOm8NMyOgAJLalXcAmyvp1pSinPhqhe06IiNurGqdYLVw45jyEEfWNSLvd9U04GQGVjgbCapxC
SLOWI2vfmNyseF+hBjMniXZ6elEWYxM0jebxYhVq15YSPAKuvlpNa3BWaHNq+Ge3Q/tHwDNmwFKS
y+h8cHLc2iZqfEjXG57ERDSNLvNn70UR9DlMNqBrnzi5WBU1rla3kWaLUSwQoQU4Hwcdfhsx+K8H
sAPtTOLGhNgb4QwotY/9jGNkQBMcTkQ6kOiAE50ee46Lpd/FxDTbuGH85/JzoOop+3aTaatV5SaS
3Kr7QxJGoF4bbe4WZOeBhjISpLpSq7eBkyunh9vgdHug+Obwr483ZlXBSQ4CJyJPWAtgn9EC/i53
AJHeOYqV0Rk5sRkb0aq50yg3sZbkFuiuLr1ErZ9H265gts9WhoHAIG0oe5mZsJv/EF0mewx3rNvH
DLbbM4CG9YdNcmWe1AyOxpUEAxhMrd7Zh8e6p3YDZqu3R653D9lA0Tm1HSddhH2F0H3feH3pNVdV
MEAZjIRAyWoB/k94yXB0m5hJ2us6nGAiJGmQuGbMWy45c9hSJ2sqcsJjv9PGIWtDrcduDi+g198e
9sB9oQqKJ1u6JDsxf5QtH233Gj+xn80E/F5afjGtYPaRfySqWv++YuN/fENfllEnht9hjTkwtvMX
yw5hbNX+qVXLHjXkgo8frdvvNpTjyAbR/exhChQyqt0kr+33mJdHSvKh/OTO0ry9aa+evhtEx4p/
z3PH0ReK0DcXAqGANoAlPJuvtHS3IwqDwVkWwgYIYGDlsFTe+doNFaQCRQ7W8QeJr0KvWNfxjMDQ
+3ZVAj9jfx6M6YtrlH/VNgpny/LnX+npJl7KotODaeKATiJ+fwNoAO61ZAzfYY8kfWyLEvJr1Lh6
qRIM0Tt5WGb30o0wQQTXcQETWAbKqSXMyirOong2kCjY8vin5k/5hwDZX8tek3YKs68JcIoIRRt0
nroaYXzKhSWqDvW2d4QzF/vKrHzvVc/pqMJaD5EyVDqMbEj8qEQgpBtXd9ruF4CvWdSxZCxpKUqp
CKb84bJIyA5oNePhhaGqFAJ/EF47aFGRzRK0knXhDxnN3KUTy78eRqpBx9V2dSGylQsBkZnBoHC5
bey2D49qpq/wNPo4/joh5IaxUd42AR5ZFeWQMgVISBBdsv6dheXAuCM+BGIJmlxZU8JbtEeDcXxb
FRu2CTEccNuRSC9jnpU5y+uj+zZmvBxmaWcAcPcK2FKSASkDxcX1+uBMTriwu4U6Z9y425EdpbGI
axwNPIZ986bxgHsRFLSaVriIihvCzHpxWyxK7g3QRbZuvmIXebOnJS5sYD7WUMGD9ZoxO/OBKgk+
D/jcaT/2eSMg/TzAizJRcwPVg+jVLVFzNpBk1lT/dzYG8xhOH569k9/PQNOPsxsL+aYRe/btrPoJ
5FY4Ow4uJQgVMECS4iaVSY5LyLJjawkoYs6QSamEwU19XfoqbB9PYxwrarxNE0e615glSDJOB/n/
5UmJLtGIROrGGdfx9xsk4AMMZNZfVJjzy+0JJXuH+6X7pkK9V6BeN6YtLMYrj4qxh0OxbWEx2IIx
UHrztWrMuglfP9k7CbsVYn96SrAT+ILCN69+iQ48HynMKexeHnyxsCJ9iaYQUHgP1yC+xmD49JAk
Ln5AqtPHV5KQTyyafeTmSUoNyv9C+LzSsA7jCWcFZyrDlpWIQ50CXdB4SrwpbQqAigo3+nY6TUnK
qWnd+YC8bRTsXW/8z3IPWP29y0ywkkl73tPzgwokfgJo/TY/wIHKjSMYlqTDtTiz2HNCLLqWGmnc
0I2ETOUCdYaQCzWAJyCbcQR3VtH9QP3pfDVpCCUMfkuECTmKsiWUuU52HS65NrbzkQZ8kH8xo/4s
IDMmErWfMJSLTR//R+4wMd3Dwjv7vNWQ5dQ/Fb8zirsPEPRFQKltyNp0xerGYn2tE0dmwT9eErVq
5LTpbgDKS2UdbUtICjOXIo/eCV9Bo5ISfqOB0QHSbFulG9+1TmdTzCLIVd4gfKGKjdVqBLZDmGCc
4/nOEyvZPp8EptBhZqW1uGZVIeLVdSm1WxUIThlqLPQ/F66fMlTQjZT93kWi+h0ky1H1f6s7MBVs
6EBviZu3ZZJ5s5ZzJIgsrQV9jqevVK5IzEVucZOmPk/jy6glNEBFyGhOnNWUqctN1lUOcfsp/lzp
28hbvklRElmbvm6iMgVKh8ha/EnWjVuu2sECvKSM9IazqzyKMKYNtvqp+KIHuf3FPjhbYA8QknhG
IyZ1iltZU9kw+v8anXV70BTe+qYWzqdsBxJUujcIBsGP9Qz/4ONOyG9uV7p05BRNf9BBusohN+9Q
oCCFj9sSMsIE7JSEcibpWXkjPZ45DHZw7nkBy3kvMFwFDA3/lZu/VMGNlSB/LIjPeRVuWFDIARfV
ORaMDVknanFTV6eENbYuYp6gY5m1nHl2k8iDsqP7W2EM+qOMsrXlK8ai99cmxUOXpbmKIP6ASo2L
gATYUXEf4uOwGqURct1k/ibpT18dPNTlvklVNvh4VAECkcBwp4Cbd4So5j4sB7a1SxcY23nxQBba
8Wr5yoyrRjQ5oK87tkNUSDxPogOQa7i/qLu+O3jOGkNfc2G4s0Ro/6HbNIa01KNDBqwKU0U4P+pE
bw8djPcG5ZpQRM+cUsi+lhPQwkgmlkE5NiUJedfTZ3bKr07c21mzRkQ6A8olda3x/GVQGVwEPNH/
qwen9JD2jGhsHAUiOTW/yhw58u1d/P93JMludI5E0CDHMgvJBIo/A6/b5c2ngpjhWXepJGOGGrfL
yvK03sBd7Y/mmT/0c2jHOwPu6CrT7ox88iaUxl0X2wxb0PX7jznB/mX8bTgdQEd8zoZin6dj//Uy
yUZXK+oVKB48K4zcSWsLPNMIsPsXjt2uGnz3aFh/7vPa6ZxNJpjWvfZvTzIGeK4lUmLuTjuwXM8R
1m/Tm0DeDsXGWrX1u+i6dUFh6FtTj8CEv7ntw6iLUJEMDkX+ykgCsCHYHgw+JniYavgR/LjYy/ZK
q7HmBWa49uC5tnlu413HfSJsvFv0EhQ/SYU7QCG4YuiwC+naobnAxk7P2z9hct4Lr50t5dayyFbx
8ly7P49/L1pPl7pcOhXbUcvqvxbrgKXq+wu2tCkmeF9UvGGWTgO2zUP3m65xdB+YhzyxyQww0gyf
yEl9bjule+7FTULI7Cgi+2QAE0yh9Rzb15ww3LeHykWE8rrqvi7ZBJGXMQUNvTgrK7/c6+IFPlxH
A+h+Os3tCamE9WElDZnHI4RuHiQiQuxcRWjXSU3mkqTd0Q6qfIiV9yzdSw70Hcv5tHSB+PzbQr/c
DbmcBtmPKnnxe5dWcKtYrkZGRBapsLszTFSiw6PLkHXFFP1YYHNZsphI8Mc6g5vax37RnxlRqXWs
IPH9Qq9dQruFPQp3SCKap6afUnMjU+S2egJnm7j3xgs2IsrhArBxmdffP2hBzY6J1qNxXtEMDdMs
cCR6oOhPp2hNACKnv94IAKBVE4h3iYQ2mHsvtoDzyts/wTh+6j3XQcZNot/QljMcy6lHwlvT++XI
VRB3mYP74gP1ZmXaYieSnXMLCpeUBrT4DDuaUTizagL5xVX43gQbPT6nZovzo+s/WInZ7gnFkRn7
3tZ6TLtHlkZjqfJCA7V6arGH0VVx61WlUusufl3ndRdzKjvP0LXs7Cx3HJawKKINon/c4HYslUEK
xCkp15VBFFBdx8obDETs9ztejjIs82k/FgCz8/FxESlk0B6EUwosF7gKuxnWeSOjp5rTZnXucPAH
6NWOF7t4tH6dlUYmoA/OuWPHLaO6YOVItk8xGwGFC9mpz9DatTkA3oc286N6SNahV+lJH1ZzdvXD
8b4TT0gmrGpgYjREnIGOEJ+c/6weoZfmsYhuVr2wJu8Vsl9QTwnvfuoA+79Mlqy27wVNDJwlcPRQ
ySNmEbs99ooT9SMgbAdVqbYrZ0T2Em1ukOPk0829Krcnn+ZqLi7cx0bhktC2+d3sInj//d+p3xOI
zvFyhuqyjug3dnJf0WcOokm49XLoZd1iVYnLgeBd//0yFjRsDdXwKuoq7wzB35u5ySvb0Gg8cSGf
J2LHJLxZydIbHvlcSAKpBJUWw7syfDTmn6DArAo6VPxTPsikCxWplrUEfWCK1eF0wZoxpnELK0eh
+nM90czNg6LSEow0MSZ0tNyV1Srg6OiGr7PFqbpJsskKh0+Rxxfp6IuNiYwtW+iGbllrtyoP91Nr
8Yq5MkQVT0enEi144v3ZkX/PhbdMtmWRVAuLVOkxo6H3xHBb7U6piLtX6jO5hspiikdz07NGngOI
IDGQQZvFxy4Vzz5xnXudyfh5gwrLlAS3HzSwS1VI/xkyhHLzEL0jBvGgEBnjrOwO1dBtMFagAnJc
3UFoa3cNCy8HCnB1RR1HmjdYDI7RbhN5mt5OZnJ+/xgIKYFUwlhkWKHV4luHMMK5Pu0QZNb39Ii4
2SDPECk2VWNK7bPF7xY8acVRlcQL6GlsEdHH5edX5I+aeFpM8r4fYp7bIJxICOLzhZPEKsLbrSBx
bxrx4GmqkZ6mLUVwSEDbKoPxjdKA0/UVebkxlHF/kXLJ5OZc7lwcDvjVDKHx3E2M8LdR1PeJeeSc
f3iWvtUN4VubdU2DCcDLlJK5zaZhw6MGe7p2wy5eKqwOD1GvzocbYy2if6lCVkxG8BFsd7zVxzsA
wphSJGxSWnHrE+NRoI4Xyy/tIYC40fMA7LaxJ0juLwIf0u+nf2voVIQPJQo+1sBHgtIosMEmbwAf
PVX64UgOus1jsf6G2QKq52uQGCRPoNlKMSVGlXw3pJ7pQmHDlyH/HX0i+PXnPS3WRFEuGiZpt49U
giomK0aCpf+I08H21Yebonc3GiwM+jUQQqacmqIwbXrcK0xHb7jDeLWjyojOvg5Fp7Ct7k+A0/yc
c36XP3yRK5vfd/jJMJvF/Ka1DNpEyOUGFhqL8AGLPmx25RK7oarGb3FETsARhADYTLUonTfn0NKA
r9an1z9Q5D0u/6j+4Fcmm1DuLr4K7xknCJDsnx09teFiJQ/p51HsJ8AmIHPMfvAtWd9RW+LXRPPp
LiH9D+SuY3LLg/E0jxjhlbHF+bQ5BZXSyAl4p+SF3/k1u+LXNwhJoZYQvJpcBBh6YB5dgqCEaBZ5
6TYvN1u4DRzqI4SnG7XEZir67ui1qy0kSnb8XRJpwF8Y2GUiNYvyn/eXMgJY4t8A8DDFEOn8GHe8
ZQO55fk0lPvkKYM4MtpjchwxJ0O4jk3unBu/yANe6EQzSQNdX8l16aIBv+kPQXOEUf+mCBSJUx7m
1Y1Q7huAxOJkml3iSNY9wfBHOGVQK8/byYqMV/HViJ1I6ySyW0GxwNqdGkoxiz6mD2oUyh87oEpH
fK1Sln02jNVkvmqKjHnFpOePpekmAbVp52SH+ItWJPJE1RNRq6QxIQAE1D39yiIYr/D+ZG4GzWzh
nw0QEF5u1sTQQs6XgyE4eNVQWnBS02QhpRW5HRpV6G5d2IXrFyTvcG3RPOQcFIeS17jdX1j+W0jS
YAXCKVLoZ97JGxWYhlD30f4geXGo0cwKNp6heevLsne9F5oB6u1c6p1dGMyvoXAf1toE5/4PxTu2
ZzgXRF7b46z2/YjmRh2UvSuqtCANHvTD9uvlq0Tm/OQylxVDyy1WsQ74Bq4lBSBe9HtTXbl/ClM/
W83+ImEBCV9/lbAIeNMvI1bCmsgwE8RNK8yOm95C/D5dnizRX21YfP09vVY8AC8KFPYcYWFWHZLC
+OEqtobq5KuGKTY4ABew9BxxfSLm8m20+mUhv18koMXNLOuEBQrSKlI2ehN8+X08vAKRjSPL3ZxR
KHA7SDkJcSVj5TJewmAvaVo1MDwfH3MJQ1Fya5Buc08eWWMzwDw5LiuSSkqe725jl4IuBKq7ZxSe
kmpLcvzc7UippvePJlcquBApEC3PKBYnQ3VoRo13Acn8jAt9wgl79Er29wrCxumfWoXR03U+8riK
TDXI9xuf+Fd2osEIHBVx3pbEXqxtgFhejdvgLbRzxs+Rh8qNXi+J+dn1CAm0+bOqpGFL7j5ajr5F
2sz9zcMM9hmochsPu/1m2eRCh3ynV93nAq2SvrP9CL16528tj4PPqreANh3z5KCjXTkobpTecSmI
2MM45sjKJaXdv8SAIsCdahvZmA/gNIQ6IlZQxgAV1jgIKIe0JLyaBw9dZAKFqMdR2brkaWT/0E+S
QHXy0YBNYaDg/oMg9MxsO1eLbR2eB66x9TdBinL3wOvCliy5wbmxl9PgphPZTZiijq/DGX0a11H9
UYSR+hXcz8hCaAcxb1B6z9A/UwioFeXMYU5R7aYkgwStBpyT9MFN4Y10FFulw5/IVCHiCH32nDx7
vUOyzws4kT3i0JMW0q0cJWLDjksDNrNjkAYNXjfxH88fMsSGNePMJSJMMHNzUFl1GgFarbmVH7V2
axg3YKX43bvrQWzIgsY1+3Jvv2zIsQm70C9X4oouN0F4xbDmQwv0CVnazRl0APWpYJZuX0RVPKwr
/jJjMW0Satury6lmQ6E2G5sAq4IvHNcpm+lUeeFOdoz8/wsiJcyV3TeObbdQ1o/jsxfapcB2faot
a0qoKGdCSVoUe/MDTH878FlxtQxHhjF9XFiKzxpTGYikc8vvWkZPJ+U0nvu4Ro84BXxTbboBzM8I
QrB2UPcX+hP3enuUNnH8hQ/hOo+rchU9r/bBX0hqRV10CSd2Uc7DLzeyDDk0mX638jRjwOamZpcz
tTzdU7es1L1ovAQhs1rnIYmFUzsDegBaZWAe4pfRwt4Fv9NXfbVnJiAoyET8ToyBEbeu2ZoZkHZF
77RnSsdJZgIKzTi0zHLawYPISr2c/YvBBbVbCF3iV1GvgNd3V0ocivmrBMII9cOMVWWJ8b9tPqb3
wf3nsmw+r7k3anTjM+vtMnTGcjZ/FiJq0mKvIAx8g1Ruyq/Ctfm5G7nQENKHm0fHmyPsPRUGjJZG
cTIWyLL0nqFRSzEtrAR9CO+BbBowbc0BDdqc4fqMCUWXF5ClD1XYJdXMb7t/MMzYP856H7cLYLCp
zYOXDQLA1v3Uojm991GMbhMJRTCwVw6H/GbMBEZkCkI7DLNk/4397VCaMi7a1O/AzUOAOnsa669k
fQBiGc1xNkQc/XKmoD9qAz2uZqAS5pNisbo40sAg4A/Uyu7IRWCmYtNvqvT2uSSbnBVYlZFR4ndh
rtUYMrQBmhLwC3oMvYqkPbWSQislOq1/mqrus3H/9OVJgM0oo9Sk5toRjSzLX3XQM2lA9mpVFmLU
CW6nrRCjhHAMdtyCzCDqYrHFyQdIqguoF6liOAzl+KrXi79b391LdOq+dCaE899p3EKMUS/smTj4
h3Odu2qwqMQqNvqlXwWIV9EQofs0oP8r1jO/fggCPu6oCr81X/JWkHBMvGsQPL6U0EsMWSta1nZg
b5X8HuzLlN+td6tIkUIFzpjb8XhFtPISgN1XbwZ3CprnJEEuyRt1Wl04vuyB+vQUllO2+hreLppp
o0ud+O9yS+AtNcLlP4GOQ3ofjVe0jndgiIiE1as8R2+ma3LiUUYadxPYCIAR3vzm7kY5A+NDOYjW
fAPfQD7tGWcUHFOz/W3guypcZvmwWnTrt8WQPWqj/RdAIbt4tj6wvh7Ke1cewP71wsLGVWSA2PUJ
WHVPTedfHGd6sxMu7OUOqXQJZIOtdH0RyBFqfUiNspievzzJbJlTQW7wHgvz1lpw3+Z3sDhAXiar
X8lAYNxnyiA7ZLe14SMkEI4DsjAGZWhH1uuJIqQbSbWuTRm+X1HU4OtWUxeBTa5u9hD3j8tcj13f
CI4ZR6jzJAXAKz4LnOQ7oNCHXGKo2Gf6YjNTBMyspW7cM6jnq6EFcN/Dq2VPFvGhRqeiWmXFvTZB
EcpMcmFvEM4AE0D6jSJGwObAJfaaWNACcnmR0H97Jz2gpA2mEZKnkp6frQPjJEsgbmDrd/pdtVF6
+hmKW3w65UcIlcu0Oj5vJIjJmGqzFVWzjmPbz0QbWQcDYJXnIj83pUaPHzqBExkwjVIGj0LCjBr3
gkzWyMTkG2uvVNfKHpkLZTZWkQrtnj+3wWvFCdanI/sSpYjIYvFzeJ5mAxXv4YJQjGqasgRF8Doa
AMWq6edcgpNbozq3kBZbUDbQhz0ytpgdU/YiLNSDVSuUfzLhKf2HYuXI7VOtUmZIBn1jpT5MnnQG
qoN63wVZ8fVZolIuFxazgw/4AVqiB2Lgy2Sokt5ij0YOQGlr5qbCF69+i0+7ke+0ve4QGA9aeZPh
NjxTLUJkaN+ZpBFwankE2Mq4sJNCJb/iRjtrcH35aZU+dK48zhlqVrLN8U3uK+/RKmw/LzG/Ez6T
OFZNktB+wta/X7tyRK3FLdvFwjuw9GZzPhQXT2M6iSUOFwj0rMDdbUiSPhzNakPySvNXv1mJHHGe
37JiHahYdWztizZfy8MAXOEyolaCrVq3MOXRWl+pwt9HLCHniiZGOU1rx4bnS2PWeTweo6sKudyY
whrNvFLGhPsmAy8FO/tAynilKLX2lhh761qQkuIaHLxUgAm1aUDsbD3Q7IlePxlhsHkOIh134vTT
mZ5kCo7gY3aJTyj2r5heZmLFXfvoOUrKMLbrC2dEYUuhbLr2ERrxS4lcoU5+X+z4rk7isrVS0MdH
4eBOAIW/LziYqQaBMznDse9yKjm07cqRTstHnblVZ1OWi5zxrQH0m2BzNJCslOi6N6l3dnjVEO56
oVlBe1sE0tVbCMwDgJDu++alE0EyOfGV2jX+jMRjc77XW1TM7gKhyHATpg9SkfE9c7rI6epyDcP3
3ZlfmizRrejFfzd+0OZyYRazyFLdgOIqo5YDYs7n2Vjob9MUPEMmqIYzZiC3SErQkEaSrsLEH1Kf
dzMcDWJWSLhqF5ODShdcmTtgsNZpGdvuLSPocANO2EvIj9xApPCkk5OVmBfYogeVRDxMMGdg4ib1
Qt4dYLXaMeYdIP5UliBJZ9UNRc3gXzSLxyxmA5Ezw9Y02u74dQkKCg6XT3GJxbW6UvsXsX1aXP0u
R98VICUpVPVep4nSz0STHsUHRovh/KytCWIeK9r/SLb01vGGjd58M6SocG9chGi3Roe9b3uNetkx
s9252M21Ph/xbNsC3WLlCO6DkwFE304nNPzviobPQ3HaIvGWLzBcHwLQzQj9uDhFontTUROkjLPI
ZrtmuWpQmYF4bPr2Z/wZJlGdnUUOYRdJQ9uGvYFbXobglhZhEIwbS/tM6X71WtshtQUK4RvhGHPw
7HMmCPWZNvByXzkQEaIWsYf5PJb5gfwO5GyUX0VC4DzfZcs8jfZMkbXfMkmBYu09I76jc6tW31S/
CrA4KLzXm+BD28GSA5ZLQ8495CR5UXpWAmjLCE23YSYiDW6mbi7Ql5gSX4lUqHAkGMFWwmEg06kK
ZPskqCvsz6quB/WUbCSHrYwKC5LGEkDEIrQoE5IstJv47+/89S4eD8Z2ZGzYKfwqow8H89S+mn3b
ACE3MUywfZQhDBY1PWy5w4bJpYRneaEYqYYxldB1EMOhTtHgt95TS06M0o01tJSBZIXALnO5k6oI
XCzXK2iJnen5eD0vwz5dTKfn4W1PxbLTLhXXFUo1hlTzm0xTLX3i2BQTWrTMbxmQ3QQcEj/zx6zv
/kEFM2iKngK/fLsRtVezBv+XE3DKw4xFiDTOPc7J8jQhmtqYNXwe61kR2cJ9ALo6pbbpRD/ZhY6E
KQcso0r2dwi6niKaAgEkJf4myHo01e0CLuakZ2TsR4HBls3Z/nUMOxWjtC7m58vr5HgiOejL3/m3
evQWerqwGV/VqygL7+r6SZh0U2jEa56C/RIs68vC8tJD7G/GzaQ/1ff8oMvqb2Lavfx9bAuAmNEj
7NFZKVUsuPHpBsqPWKspztkBORfX6rEjPCZWHvWrS5WrZMCPU1uKGNDFV7YtG96orpasngfuzEC0
d5ktEKtaT3IkwfkahOXNM7mx5h4bMHOMQ+at4FWmKdm03xEr8msD/G5+Cz1IgQ5SLIz3KGyGO5qK
6z9zV/MhO0cTJ1XDUdYwR6ijVIScdXQMKxzEj5gw2xNHd+rsE3fh+aA2LhfQ5PxoSp5iFTVd1+FE
181CCGU5yhBxh8hiLM9rVnyysNzHxpz34ukReOKR78G3HCQvp3gPwf8jk27Zki3zNW60vyuUp7O8
GYsGI0EMsDgsi+QUub9ALxBDuwcB6H62x86WbYH2zVC1mARwsrQsN9IFLcWN2B22aXIW0qWBMg4+
wvDdKM1yZj/Cip2Dhw0wMStfssG2t3HXuiGrVBbz/cPHVH84NobuQatIlcmrIy9Ra4WzuC7brYQu
dMVWvvHaq3HRC3Ws7YpUauqA6mKfEnq7QXg2d7fptQHQW2U2/ja3FDRRORS6d1Frd5/qVWfhkGj7
XYcNoaZLW9Ib2xY/rNRF1+U0tEQh0S5RzrFsaniJU6FdtzG6HzZZD+AxoVgdndbDWCpIAcdxdQV+
5FZpx7yK683Vmb0FCwnC9kYHhRRZU3XLT2CmRXMx6+12/o+o3ufmiutG1jBWzYx00M1YIr9Lq7P/
q5meVDaFpN/vFTYDaRs6HggCqtcW2xeGJNamcsIiyVp8TnOfCfGjPsJX8ASw0ZH/Ej5zsQn3jcVU
zC5MZtzYdmi58ffc9Gux0rZlPBpASD1LFxUdhGUamVAJkbjYsag02SBzFLguP31yuKg7sSg0QrIv
nBNGBcDSrQWRblamSjLWizkyhPGVachqzL+CfEqZBx9U+8iIg/n2c46mxIZZm2tFjBZX8JHi8Qxq
kvizf8rP5xURDwDvynE2A/XHgV1vHbpO46I3n0Aw/5Z4fll2szfaAOUctyR/sqljjsaiJYSsDnyp
DRtzqKhobLNc5qqpi2lChlJJ4rF2cQERvar9+bDBfqiLzrwR79EiIOA384Zo9O8kA/WQ649v0ZKb
+QjqYZjGhTrO6TeLu7PSwR2Pk7IiYCTlJOd8GsMG2sxTSYLQxR71VTiRKMzHvo0gdorcvDRX4gqz
0x30kXwf8jkhAMhxrUIBuU+SLd8Ug/1XiRzQ4KFU7POhK4rQNcVDFNIz80DDxtpO8aciSeuTIl+P
jsOTZOaryG6pypcOxe7ubGRIK/f3zOa0rfQcSFi7D3U6jZYeKjtoSda8+UbXoC7l7MKAOQtXEOXi
MszjNBdkmltTJNISRWRjOmRYqk5frTeK9gdFnYsX9a01i00ISB5s/GUN6xrX/gfJ0cG4JsVKGRP5
72JnAZnUlLrpawKVZCy2dkH6TSU2DF1TP/DWlLMqadjmlROrBDczp+KfOm7tNHOf4JJHcXMpDTvF
K8u0KoksKuOhhNKaHlyKtLZ8LDsTQw3QRYR1BKPUqB21PVh9cTtRigznneB02fw8calL/srlGKKO
gIJjeE0eKKKfAeB+4TT6n/FYOYuMtUmQrdqVc3zLiMIjb2lhch9Wp5l974diUgjIy3cn+lEyc8rf
pX4CSeJolfDJDKhUBOZ3XEK3XbZwc0z/xija7RONqd2FtuGmokE8Aoa/jF8S5LdExdAYoKbLO9Tj
RQ5rQMnM+g2n0W8BvJEB2XAzVnkZSSR3d2bjCQ3M4bh3Cqn5we3Pnxebpda8lXiALIUd6grhmkuC
jAylT5ZQSPK8t5qzGmd14i3D30W+m0UpetKTy7Iy6al48LYhaLA112Rx8sTuOTalpIJ7HJpNXVgW
HDCdFYwHG4pTSZFdCPv4x3x28v0VHV/em0CUqiZ9BtbiX86M0faAI09TRlT2lGS6qjTbEZRlRUub
ducLSUx3OfM81cangFsD33S8OOpF3QIIxP/aI++skf7hKmfs4JLzLSvEE/dZ6TCGb3lHDiB+dcFW
wf4r/iqUgofQnrFQaNuq93rBQ8gsF6KmmBL5L8qvuJqoovXBM1w7Myl4s1D1YD8iMgEnjS9Fa1Sp
MBNgtvVQlIyNyMiIOcSPnuqaUScz+pViBf5tcxTV+GrNjPL14xbbJpvIpzKQ3YNZzNFEZGdY3BsH
W9VzWZGRiECbUL+ucVy8jJRj+KL/IbhLgjegqM+CiLrSgj7LGQb+3LweNu7n5MMBz/tD1nUg/fiT
n9lUym2pTzMKmRo/aEeIabpqHKknOo9BVj88bYKljHvPLsq20RsOmynHxHiVcsLzfNrdFG5u2IRH
+F+y4DEZJDqGLIfPTbKjVjz9X000A+Tms5kgCBKIufG9ED3OY7Ftfk2J0WTMe7YGqSqdNRB6K8VX
M6IkhbLT4akfjZzb4hH3ESFOcZ6HC7nefWsN75xf8/aePvP1OcO900H+FcH4aEiPXw+Ved8Prk7U
XwHaWZmoU8a7B//ZznAr4Ypt3C4CPQYOE/5nNw19dPZcQ2/1NKUhxqHMDhXm3x6/FVMNI1x0QUkp
V7rkC8+lJvwnTyR8fEb53CvNy+Q3ky7ydE6ynteVbB0VeSUBThgacpY63bq239bXEH5cwu32Xp1W
fCcgwalx2Wx26QvmCak+bgOHALHs3sZuqEhnbfqjKb1a7l2GKhvBLIdJGH99fsuGi56VNEaAEmpV
2GcMEt8ySx78cibz7ea2KDk5CEvwbdLKMADoSp4aDYMvpPSQhXTILTBqmjwTXCYfqnfe4zEeNvLs
U87SZDKFcKCSdmK6rIdjzb7BEu3hwC8LwWd/fhnN7CWcIkqVlE5zvxWJm14op0u+wGXegOxXEBDS
kcSlOgFkkfgZ+qZizXHRsiHa4A5v/aNPBa/sfZ1KdAuIBHpBUaY/hYUfIkcp1QlyLTyZmpPJqz/x
s1DpACxmROFGibA/AUVDuxvIMgctBTHuq1l9tFWJsYDXh0w0Qk1T4uhgbZpOPAW+SLNc/jIdz5QT
ILFRe9ve9w0Y+ycKfIRt0sXycUhlvvVsrWgEjgiQhKJPAqY4M1wegFRKGPW+aApUsorUWri++Bxk
NtzBrZKCcimHQD/cLOfT9BINVXD5E7UWkOIBv15R7loDlgo4mlcAP62wOQln0zMK2uBSsIzchS7/
kGzje32sX7AfCXct+jw1UrJNQjA42fq3N8dRK9J/TMPmAuRF2lbwpaYCJB/hsqO2SUOqjDt+AhBr
CsAHleM1AhI1TMxZxcrjXO32b0cJeQfMPb24FtoOvkvUU24i3h12lDebXO5GeKNbxB+BHUuv9Sw1
X9SGXmun/HpXeIHRhEr/r2dMs7pwEsHa883gyAhDnyz7rwpsl1jGRCgtyB90lR9lGgGOdEqDNiaZ
4wiZ/tJoxhVtp2tTfBmqP6tsPNmAPUp+pNSjicHcB3kpPFFF2MlUGWzaHDtB1LYlfoYrxh0BHUIl
TcGFvEWhQgOpuFf/IQs4C2LNxe3VbZFEmHQ2asPVadmbKaTeB6u04428cc0vEB/sDkMBRbD8BYNU
4hn/kJBBrCmVKD2fs4DPwuA5TyXhq54poKGcl2IcrirDZpKMmGkZl2bmxUDAUk1Xd3OhdYzqWbcJ
rxRirKfwZ+Jc8rZab2pPixEgxHlxNLNiI3uKiWLK0WpESw1iZwNBSc66o+LB1omdJbxfeipzWS9J
LfyEWy++6cfjM6fUCisnvMOZQtjg0SNixDCx/HfKJ+dZFLV726ksKuoC1qd2pRvL9PO8NxYXxavR
mDWa5nTicNX8WrvcdVkM9TwBLSlCNDuWSThL4vpO+TO0GAIHrro5u76KpFYIZJYR8Mjj32p4vSSL
N5Yn1rlpzoTXIzTP7vet45riiKsEFPus0hn0vrHNkx2lCBS9ZrzHTXnOe27o9ymeQIzfWDLXvn4K
AMK+7jcKnf5rATE5tJsoP4UmcEwKGTE3Lq6ruypXuRR7pqN8aVhxLxJYYpA3R2zIvfB2Wo/+K/uE
8uogA5ke9BJtFlUq/juarAWNw1/6CbecjQCTRXtULNUE3IGKS3w2NJok9JgWsnwLFbqSULZTZFq2
33uMtGtYXffHLROcYjsoPGeFMpuV8DNBmpd8IE9hRFzVTo1/ZkGI3QdjrclOyfRWe1mH/kQkBNDa
oQlKeg7hBHwcLMVV8DKv5lQ0AW5nh0LppjvYgzuFHpHj22m8k183RUeDGy9+8chk4ktRSBXYq/y1
5nxgSGhAFTdzRhQV/Ga1Cwgj+zQ8mbqC+68L9xK0AkbOIKBctq2wiYEjm1GBgT2j2HkEbMab1cPN
ZUBpKz2Kmj+1bQl+zBzWdcYrhkDxiIXm9q9jjsrjTswWHW8nCXeDYbrYg8pWnN+SHsNc23fULkc1
2aWEeXzsvY+swpEE3og4gWfR69nbuqHsLxNFUsVM97miVT1VBPxMSAePQ3hJ34I1ZzssAd1gJbN1
TZWYJag8cumNbb1ehf2ET67jhalOpNW9TAH/sizJGDKukJ+5uiWDjoJ3wrYMTqRSBZ71kkIxX8/i
tFX7hMlYMghccaODMsFAe6C5tE/YimXDO7Uf3MgkPYGetaZBhMIp74FIV3kr0Wx6qAujTYuCZKDg
2ycMq65UorYaFDINbjBzcBPmsETXZeFJHQql4CxPNXQOgZLpXRfX+dhcbBrqBkMc44iWD7g+xiJp
4zRt+M1Zoou09GbFNShA8znCUt/IxFEmgpWFTXJfbvt5OsNWlSP0D+GbrH1zn9PhDmo6yH1Uk4+l
oyIlAjWnrwwEOIu9UTxI+goLaVXa2k6+giYT8Buy3w2CeytFOUmJ8X5SV8xlUpTfEGziz1xiEiq2
LYvKLRb50jn0zbr2Qg40hXuSAJPDmHh9+zlP1zOwHCP7KJcsgTPRs+1Vil15iFnyeR4IrVYarWEP
/yBpYwQ9aT2VmUZbBe2JQY2grHRZFZIbfQx7sY2UvqIWDSFfECUSU7AKAgsE8pjxjCITbCyp9Keg
ObXdgBKzzUWmm0Co+sCm4p29Gby/nolMawJd+SAEj4L1rh6TSJXDEYi0qIUkhZD3VxEYS8YzK4RP
a9DOjv0IItdouJ8A9dcuznOegs7Rr1KjvpYpX1XSp2Mn4CPyFYV6lWalwwClu+67BFdnhK2jv0Nn
W3owM0EhnInq/lTA9QtoCTTnBzbO5qImVRtfm7xWIKOEFnpg86/B9ee9bXnGnY6rVmrEBaENtzTi
ry0UDpusefKr0mBSjeg9F/3vVeFKX6HXuF7mKuYm06554IuVXarZR1cAoov0JzHFRM2x/MYC26Du
iI+uU/PJkqF0RRtbiTJC4DKj6CN1IigDitc3ecTaFCWOG+Gfu3VscrgY37phDD6VxKKVn+YoDP6u
91kYTbZuyzymNBzH+AOmOz6PUcONB8YMEN5pZFLVEpIZSCyV24DXDqUEY+LGUoIaDGFSAgEoNcKm
YQVW5LR+zq/osz5nxoc3WljPYnfhJd60lu7WMgENU095DOIur5VdUE8pUuEN2O/RtVDUUXEP/nZ4
PMMXzp3xbpdR8BoQPQypvgpfK1Z7HbHQ4bS6YuHs0Y1fEWqFUvoiuBzQnq4UVKt4piqS09v2vkHP
NkeO/vII6yd/wlSi2BxNGBBEXKBEmwc4y4MiwK9y5EZAmPv+gqVVY3WT+Qn0zUgIe/OR2GxD9Zcr
Q/qX2KWGHZ/yOYraEJVC2GPOAHn8vDTemsCZcZn5t6ubuVTfSQYHJM4/F/q3x+KWTbv3dp7RPM0J
bXsGCG3uwjpERmKIK3doQ7aWSAJ+DQP8WlE/xmRjAitfRYqtDjnOpJdeqbi5agiSgPK+xqJ5KArj
cVTr8aomJ8FNeQBkczXnwhlgRjlauQu6uDu43GHz4xz3+gK0PsDAzSiv+lRukt8QGO6N1vWGZkB4
roD9yxL52huUGWrxXAnGXRLcz77X/z5GucL4oFJECajbdVEm9o2sUmRjh1iH4xfjMbZ3elyKWTeF
4LMpXPoGwVnKmEq2+FFg+qEhtxQqPKfeBxISokWLxubxzbm06elP5KXCcYR9jLvCbyykXvELnd6N
4nreqxG6Ib+8nXrAM1ndlLTZxpA98Hwb5S2783bds/mSZ4jJkbCh3eFr+RDiP3Wkogw61qDGwpqT
xqEB2+WE3+6ks3jk7GyfCY6IJDtHvqKLaR1aFvC/hAKfrcQibTuhVd3bmXPQQOgouy98d7KQn+Wd
/nxDGDzye79sQFBRjp+OB8BWvNtUHGV/noofngAcyL+vGyOGFQq55Nodbcj1tqfV19TdbQW0xtkR
uUus1Ct9mowRoulpTOjuqjXKkwYLxjBGPmWAI/YnCYMLdTKxXRSBjduv9R1z+cJKj59cKQ6iBAmj
qLz/FBSTQjq16DufxcDSQYyCWcrsH5RTPLgmwl+jM0qwBX5qL8xyWy1GKqFv3BR3T/17jXFJC8u5
/YPtuBxNTYBzCnjX0w8cW6Ty4Nc+fQ6rnSbaTDrj2ymY6mkf/BQcmFewbTDQlCH/Qm2gJzpVnVMV
PEbvQ4Pj5iV4Y9RMEp57qRp1eNnrHyiQHpAQqu2/dIPtxllp3YyIgFE+Mf+1JlLDOYZ58QrEnLud
DusqZgcebU9hmxHzUJUgbdgGBn6SqdZgOn7Y97gQwy+NfJ/e6LVYCLeS0+QmgBofQVFiU6UbamU4
/l9sVwPbxVqIbZ6CZx3GorwEM8OMqOHrIzKHb7q/j38L8gL81OSxgCjZI9aNPB4641lWcktic/EJ
HUO3+jjTiYj58kF/DwrTbtvMlHqWMFZx5wZkYECQOYq4MizW5BEUTrml0aIjEQYWYGVGyFWguuaf
N/qdNsBYG059V1G6cxM34YUEHQBbSN/d8gZaxU9Vd094I/ob0CX3vuOlZqCCtCRHhv8A4KbxzW2S
9uiC97uf+Pfxpr72r1mJGJlnvMBIgDzbBfw1heAUZ4T3/xEjOdAIW8OKm4K5hrnGRWRfIzk6JCs7
AJQXVDBW2O0gfte6mS1q5xq5QLkB4TyPdcGkqS1JmQdLDdW8CW6oc647xKuzExTq1G4S+2wAoTpO
bZR4ztz18HaWHhmT6TQhfodJZaOGIDByXq9Wg9zyxk6XFb7Np7/QBnORWs2SgynjfV8/7uo3JySa
gx98E3FIOCNBzwxM3ZORylFfcF69FXkEdJWlW9IF7RIhFjce6ubGtsK54stxxlkxfdXug6Xv7p8I
xoTTpN//L1VjtWsD/whae3fSy0c8r4CWXWO5ZnoEFvDG8D6jyKugORE2gFdq9CNaKqD+wHqG+3aQ
680vRxjPfVV82s5sSck6th71kzPkLNN0d0AXslsHuBvoMTZUXDo1mZ0NGozFEMwHGzl3xmd2MpXe
9eFqHl+8UgUOqb3R+fdSZEidHm9qlKuVJorXdeTmfECu6ZLAqlnqmGb3xg1Zi3OMLt+jcM4X2F/n
jDhhcaFh458gs/zwxExx5q86miM2uluJVd4l9KjK+x2l8St+O24pbbytQD7hGVozo7PR7Mhzq9Y8
lHcHGC2FRmBrzxCLdM3CWpV898Jio56xvP9wBkofyLRFmICEcDyt2MMmhn5937QeeD9ctbYFpCRe
61O/402y1AJaMQFJw9XZov29L1uYgi32vZJZvCLNXjhb9qQyks3ULqpeGlbJ+clY9SlntFypVK1J
l3uHON7VWrj3WOk2QQADSFUn08u845SWuNIm1MM9dxajkjljn4djREgmelEqUrqtHH6Mhu8hS4q8
Qg3F9NwGVacvg3InPbKQxKFTCgTHL5S1PQAK2hIZD9ee8/kLb6674JnVttWqjpnWren/kS5vgxQb
a3/6Z2VkqdPPqTEBlwzy7yPR/2pxcXb89OxomcEsqWCXsrdKkxW2Z0XmbJBTkoiMtnOKak0e/hGn
VABg/BSpz2UcFd+978+fXqscgibX1L1vxAqYw19YLCDU3NX4+41tW5eAkN53X3HAMimntNhigeW9
a9uVHIVcK9MZ+yj2ItztG7RJvpJxn0KnC45HKH0Y4CdOGVUYSzjtnHj7zo2+EKcPIRntaJN9+v2w
Ks7+fC9eSWpBiiEJGxssmA7VI83ZnyLxqjo/LPiA/mXNWIEbLnzRa6ljolib+Ad8vyAPg4JD6W6p
s4rkpUdVk6v9A1TUG7BUYgyn5vy0FHFtAJuSHYJKgB9k/fzQ0sKHa8OUPwDudv6Inf+egqZxffiI
lYx3INjVH58h4imF1iv+vF7D79cKzJpiK0Zdv+5iGtyALX0mXIzC7uSebhWS9QQ2PKkp9OBsG07/
eabE4jvBLnemgDsEB/xz2cb8QpYiVlGn6D0FDx6Wdc9jC7jQc5K1Kut+zJmHX+2B/H6UU6tr6NzG
I4oRW5icB6E2AIAAWRdYR83J1lhNQr5833NrkOnzaogMaZc4CivOyScDlavCpPeJpMEXlRQph6vQ
EJm+QBrZSJjG+NT9yxzqy2axo8TkOyPWhLf6XFgmLf0PC0FaLeidL5nGvh2PSVIrd8m7T7HeV4G6
9GytgoVDTgXsJEMASpRcETm9QMxskFuiC0as2ODLGrawxyml7VJUU3miSmkmLZEE9UIH1soLUb67
OMGyxq4IBmM5I7btaexsruz3rcQoYXDQj0RbDTxOu/wYeIpsoPpHCaikLygZpQZcbX7aZ9YUjATo
9PCCNvgJ/z8m7jYwyWnDKi6dDYqzj5jk/rYCnr26QmT3G2NBrk4t8rQSivKxWEw3kgN2r7IOWaIG
nTeZp4Kh5zr4iKFnRVKbWCrl3yNJyZnpd44m6OBwMsriEcSAPR9GElXn1jV8ccC5xmS42eZ1Ma5J
hIQ5pY+ygO4rqyr8eyLBJQIDp4m/q7qyoZBNB6QUbFbhU4wHrZb9ME0Q+g7m1CzumJLSqZPPvbCf
XCe3bv+RAZLR7hHi6m66TvhDTudDedJWvDl8jxm3qTla+cvgrqltfT9/r2OV1o8r36f89mYhG3yN
/XyEHQknrxMktgOYI7KLzYm6BV/LK2fW1DDu5lWrhOotoIWMbsR4wzXtG7wcxfCzeBMkOkZ1OvA3
LLPL8XYwa7UFRI4VkTD38+n3xjp/qm6apXQtUSx2yA71v3N/UsyXjjZuzCTovAcH/vZ7nK0DoHNV
Y7lim0C5muuJEiCz2EaLCFfmvNp9nLKBSzHVJ8BuVi4VZBo1UQWL90cgqVw5WrUM72ePfKBnoedG
33uo/Uxe1HEtmmrEPHvHwIxpSo9A6FPeP2j46Rda9mdEELtx7yEjnqG7pcz8UI2phVB5ZyJl4ldJ
EJxA0CrKD2f9aKSmjPnKQRIf2/7b6a86SajWY8dFY58reFXvqfs0+1i+NLtEbB8+fOXSbSDmw7ax
uMDVu1qHDse/Hhu5gQn3JfAwN+oPrsmPTQ4hEL4Iw0EEIgbtiy6nbL2Ldagn6m6chtRdLaIJvi8L
7baP+WtGsWhHP3Pf3e6p6OA5HTY32jtIwBbUoqixn2CX7s5vfQ0u3546t8/W0rNny53J/VzNGckz
Qk7cb0R4XLOzg5MYgzScu1Y1psLdAWrXDZ6Ek3wKGA5gATS+blQAyyeH2AN3hFDsxPM3OzJUpDRH
IZ31lNC4UjNtMRp8zM48ZFVWz6cIlBh/DpjGqVd61sJ8pp6DaleLUUPYtfHqjnxEHBoG/RngrK4U
UaVR0A0/JY2w1tMRi3gwISYy+H9EQF4uFyoavDoiFpUEw366QIJZ6S2lb0zUrtkbzJpcGsHTBXQV
hwibNGQaygNupfHQ0uelQ/emYjFmBlscJ78LRxMYEMlafRN65vTN5QC3j8vZJJ8SYJPOhq5afJCT
J+z9IBue1juVnoIndaLbD3kTd8T4LVrpRYKQPmE//CPKGBWS/IWdC70aretGov5VH3oxYsnSQ3iX
DaKtnYtejlb2oYfEaP/ga0gybPD75b8A5AroWJ4qJ//4uT7WKVm+kVLvJCNY2C6+sMJjdmhDHh9E
b+LQ75GuD+giIHH2TW6Vuh4LNDIAsMFBBmiOu3ygzlSfwxlx3ODXFtkl+1OZvzaER8K5CDphHTAA
kUuGAdZ19YAEDJiIkrbq/x8EXz8DQcPr9aRwgqDHTUNX8UMKUrKEQH79PLeUCEGQZNd78cdd+nQs
MtTyfI/5lYrNlBnv5CBrhyRvkwLll5ukrQQtElnifdhL63rLuYDFD9UxtBqXF2B8EwohJTNnvMhg
Dx6oDyKNbKYNK37V7YhmcMOLfncR8RVtMk1mlV4VfXfVT/i/KFRyFv3DnJu56p4zzlDN/aMZyDZp
i5pwlpPHs/kwUNUKoQncXSa2L+giqseOpFhaRPDn+GUcXdsBFBnDG6wyEwMdkdkgpH7HDhrW2G4O
6JHzoUAM+1N55MtYXl10sCcgK1P/FARKm0GCefSBgRudAQyZwa1a5hgblAl5RqDQ8YPuEVNXiyay
t4Vvrk70lJ700wG73qkM/kMovjtekzIznmboHwpv6rlIPBDw44BnL3mSlSeY7U2ZWPnSSXknWksB
JWw0433FE434BGttM/H+AMYG0AT5ep8IBkI7IxQv73MW0lKxITPc2My44q4czG+FFA5f7lfjn0XC
Y44CT+SCEQd7XvF7cZZnR2LcWmWqkjkRLD21VfhZ5KhhVa69FJFnoJ5hNEQqWYFKNnROPsXMOQyV
ZVwwnV2SmdoEYYI6nzNNq3y5GoJQdaS9bc1DbJEzlBwwCjhFGWV7jc4guO8ti9nCcQoluuzDrm2p
yiJgr44GxMYZkPI5BC4meda4Nn2RDCmbGAfoI4JT8f//SCNdCU/gfg49W2Ug6ZCjrbFU5pjhiQ19
vSTOEEw5DnHLyRiZUeJ9iJ0mx2le+CCgTugoawKE2C9ma5bDja/+O69NdtmBkPT7LFPxYjTaevO7
jbj4eohG2n6zv9KHVIYr0rXZtR6TGU6m09alo9AFctTThPQgjinQAMY6uNnd5GXHicvuWdUD+LBg
LELlU9YN3ciypH8wmTP9K6j2UwZgOfOLqlACtPe1AbU7Y+0c4unxL5HJyMiRN5JqLpED/9fLog1V
QSr4Ue3fJhbBxXYQZJ1iMyHv7nB+VVV5de2N00K7PER8VFNpaJGS84WPBYqOhNA1XTri32SRPnFv
mDUQUZ4EOFFTlS1iblPoMIJbqdxgHzhymaYe8fHbZ764Jm2mXw9EyI+2RNCttnA13gdQgkwuzkw3
aN/Tcz5k9keOwatf1I4RWv/0auuAWPW6kyiE1iXLahjN1jU55wHlKnJDxyQLPms8zdxoHY7HvKnW
lJMAanPSaN337H9XfGKYY5QEuXMlsCVR6E6M7t1CzKjuWniH+QFSkxPdFGE4hi7UkEkmX0vp1w+p
XBhYeClz7FiHHrN/yeUNAGl00OD+lXLu4mno3qk3k++g7snmsadu0QfGC6bNimn/0bGbbVmRpRt6
/W1bIi17/i0uJ3y5EPgtgzSzwH5eDDl4GiMuyMveZphlKCMcam5jWAnhbvieYOY2VjI8zHhqMMPg
jjj6XQ8pknAZAm7RXUQFrE/triQV2Mh/lhYxfOfU+7xgQG0LIqG6mxOFVXeT5xmIkGFZaEx8hywI
UI0f3T2YPGROwlIZAPfHB6cKYj+jAckYalqB7Ur3d4VWI09fHKsNBIAddWyzh2htJR11e9k3c/H+
mPyZ8NxDXq3KmEr3y2n4bqkUteBaiBXrY2EFlkFj0Zz9UemeZRMCE8tPl3Xs+ZMVPwJXdTSXFEm3
aIxQrarucuWvxgM/eLoq+bLzAs5HEeSykElBoyADeZbYMFHnuVVxvTt4H7h85uScD+VuqymH0JQC
oyOYlllZ6DULg/j+1x1ps1JiKvu/hH72aF93G5l1b9pQ/UYnnaGQYgctzz+0qnvDb6lkC8T4dSOG
YoV2DUNc4vyZ7DA1WH772DLA+WQ0GsCj1DBho2WnGYwozwrEJ5mBlF93cXLij3JXMEK0h7hvoArS
H21DKjlCT0fANP6UhrBsROGdbNY6yM9RLUDs5glS6nk+KrYiJx+nEF75ZYyu6vTtIqJb4KM4mhHP
7hhBuIKFQktutVshmWWNKLJL4GD+MeP8iio5UbRuqnQMcQVEkAwZDuVn4e0Le6wT1I5ZEOYWiVPO
OF70GQrst7Kdp9v3ZJK0O6G/FBi0WJ+ddaxUGjKT+m03EX9DOqLmKPFsK9kv5fcpN24VrtIYduze
bPIMl4v7sKi2JzUaPVaO7qV3RRuI/Ge9zUmhu8HmZh4vcZNhiSQ8B2mYoVjKmgey0NQ8HRMA0nYy
htf6QWfB/HlowewXGEK87QEHKtqujL5YWE4BfmERpdPLZRZViEJSh4MSO8PNPvmB/33YnMrNfpig
rQkKaUnRJstRKNEBGMJWjae7uwSI3T7YddW/cRGYLz+NGmJF5nnP64VcyWmn0+kZy0awyaf8Nj+6
UqzjGUPYRD3TFpAJhSBUaAFLc1BL8F6eYbTKRiCSg6Vo7hZvBAB1MG1qlG7KAnS5d4gTJfdt4/i5
0NyTOcSElRsXgaEp9T652CkZuUCurx3AdD/2Uazx+J/+OI+ysBQWP0mftS0LC+p9CvhYAcZ+P0FH
DmZU91VHQmqQuXZkwTrD3w79Bym5zlKFK25fl5O0k2clDmzuA/YcAomRuC8ERq1knkhkKlJ2HimW
6LJvfe31fDfvQJGpCf42p5w7j0Gjc872fnwxYav/sTs0ffE76EMKkImO/jSnMJM2VgPt79UNK7xn
nD+qMAem9WLjTKBH9uC/bNGpgpyBnyiONneV9/EvuWZN9A4cTRyadUzLCF3ubZnQndS4UbNNOW4f
4v89v4vuLHBoWU0jh+ippK7k2cw8udkMJqPOS92qbRH6Z0ACAYx7YmwM2FrmYUClfKnHouAhK+9F
Je3R2UpfyhbXo6jXBBLT1CNjjm6QvzmzJ9gUdeOTkAJ8WefGVoNR7ks1VQeeFcqZJGtfvXZK7+j1
YMT3bUVRBpGMRojLrFVkfOSFPs7KcWHYd+/bBdaPTdqGMIUX/qyiGXyvMXD9k5jdgiMGbM77WlOT
Ykj98lUImGlDgiGl2WEHnMhoyeJqJAcAFI/8W5/KVvP7A4jeV9+wXwgX4Oxd672xAEitTcp763TT
JfLx8hk4pYjARByvw4NRgubJTq2qu04WWNfc4N67aO7gidLKXPqjHPEpsj22zFD/QGSSuw5UJbC5
gTpcEs6XkZTZAJsT3zqvxYngAVilMWo69wHwQCfx1PV94FNIvzRe9UTSbnJUpgIgjdkICEDNpLdA
OAdi0+DOe+JncrNZ0AIUXTEmi/iMHxnvvwMQ2oHENSbVbojBE4tIB/XtWhVJxvLc8Oy2CbR7Lp7a
TUaxFieR3guILo4py44htKwywAo9UUquWWq30uCp/Jp1HV6yMzb1SD31glO2SZu6xeh8p8iF8Sj8
3YPSflG+3z0sun3o7sfrrr3I2bjuZrdSklDdYnopcwriVb1RnBqLTK5eaLUhW2ASRxioCrvxJ9Hz
EhtTagSpxreZ0ZHOTAg3d4q6NiMYDXQ1xYKouvj967XpruamaMxrLR4HTQc1CGVMMqOViyBsQkAl
BacytXjq73a+rcBpyrPgyFP3qR9OUsw/JQ44GDJUJdmZ1/FXalyhq4aslyNaxYRwSRch1aCYRZ4+
4lr/sHxA+jTMk9w1s+R2ohm4mW6sr0qTHfcFTtb1wlFwjnrp3aIuckiIpUXDKlACakCHUwgoQqhh
h1CdE74pqv2PrXMWAhh54bN+fdn930XETHMTD3eN0E4eKZnWkeCFMAevnEBdkHo0iGVguNzKwz5a
pa0e4LgjOKBoPPGJRgX+hA9WLX+DbBlJTkHFWG7mqVcZCpl6+HQFQQbexEXcAkaRyxBrbxOismN0
ePStbV5X2eVPBnoCy4kxQFZ2LqdfQ26vkoxd4DPkOrU1KIFpaVe5gVCtcwwySbbhdElfbXb5VNb3
ZfB78P5maG9Sm/OIla0MhIyxV9WrGx8UgBBRH2P0GHiyp4aprTdVb9Oc1B3DubuBEEh0G2QQ7JIN
q4pUBddzJRcFosh5CDEtDwvEjuq/0kNmwHx3TF85fJ/zWca/9TI84SecsNYturMVoDxOG0Cgaw/U
sk9Gbmb2QqB8URJtTSpqPJ4cK0SIyZADTWl9ebf6K32OJscqWh3aWT+c0XzgA/Sr96MgymlMoAst
j7Z8+UVH+DUkH/twyk5KHQasdjOPSvPap4jJQFySjw3jW3KJdEnHr8NFu6yu4VoQj24Jk3wJPiLp
itO0VmkkS21WyxdJGRow9aadP8sZgF7tR8DRRj2G+StQVdQoU/tBkk05sKU9hpClj0gVXosy7rJa
dPZZv1v3i/gLhR2dVKJ4H7GNbuCKnLJdHeg9o+QrvZd54d5TYS/3Sy77W+p/XOvcp+U5jXXzpTay
73q5cHmRGwnqeSuDQRqLA4caUXTjxCCnhTCWn25V+ozgRGXrKR0uKBbwUNqka9J7LGhN/bPKhjWG
rzdk9rEePNcd567jQdMZdI5LCfHsQMvzhbGRsB0YIL9sMwt1BqLZjGzFdVG8mf9CEg66iB7qxrjS
CY1ZVJ4KJz62slUIbvDsQBFzj8HR6Uz/9unAu4XPdZ6P4OdY3CtkpmYkVRCAUEj6dzJk6u/4q3g1
e5dgR7QuioaK7u3x2Tqqqd5VEUQQ+GR8KVqHfHS5oVG1Ya0MbgGtDJnN8r4oSj6GIKqnMasq/B1V
fT09JyYP7p4b+8B789ywxQYP/b3iH0jW16/IuewqlA32hVEgWqBpDWerEBu9MMR2CAT01UCugii2
KzQUDD/mBorUBBDbYy6WOQ87cMI1Xk6qm4n/PZ2C9DKYxyV2fM/g/lRe5dEOPjrtk59F4GNWiJWU
x+sGGGjJVGv2+WY/b+EeSxysj1FeEPvuXLKCzFpB881NUA2WfFzPOTzTZ6+JZcfyeauZSG3LtBV+
mNeZc+U0ATS2357/9F6YRX7+oyP0ZP0YqTu1P7gMVw/ZnbIFcCUCidL1dbS6Db9C7lD64mSjMtGR
3H4E3PQxANBT5AyQAk4vfmxA6z3W+BRtJS5PB/LxTrFc7MCD7n8FGzILZ581vp7SJWOocVeaaUew
jXDIMqp/8+B4wj6yfOFwx6FpPkfe+QC8grMsNkTDE1o15PSkaa4yP67pWQirMCSkyOuRTUpkxp+c
ayucbOJI6Ta1HE8oc7SYnIQbo3GZ76ydrMcYbRd246mwMXz/J/NgcHXFKfWes2qxZAi1fzNczzxH
KZw/HBSBgvNgpi2+M5rihHALlpJao8fHuJ85wrAGRO0YIo3OdAqsOg7+vSi3Kk0EB6HF/SDbkiJh
0wAK8oig/H5cnuhPGr6RF3RmiW4wJWiSnYvmHf1x9iivlGkgn5jZn7cal2NO9HL5ypoKHBFLEjTX
/BWIXIOHuWhzTs453+VENMstzwDUIqzqknUL/01JY7Bks9IcqfzBtCAVRk67gxeqNtZbsqXpj0Ay
JNO38pXCPWq/Y+dvXQdrGGfkmxTNQiGWV7xuChEXgVEMKg3nBIN4eUwvfRXAZxRndvhB6qmv+n2J
qbP0ipUASa8us+NQZT0apppZGIcq3cathARULXtd57plTjD/+F9yX+703W61TvxsSGdORwkFaTjm
kpB1pCsMz+D9QSB2bCQdEd91QcgSDMi5V5M3yPOHe7PspP4IGdUXTUfBMJMD5cr8iH4qZ2ouLmVM
zrTpTC/GH77V+bmz5qn1NOjfGBbLAQ5lJsC6gxe9wwYpM0BeI8UKV7U8Ck3RwVfyZ3JOR9h1+Gvh
7FDZ3mIJZ6Q4XOWzF+Bx99HpW4dl6EDKmR3PW5vb2s4zEGJwR66u6p/TGGMYn2wXTC7jwBk+jNUs
sx/n+rJaK6pDxJ2Ghl3Ef+jqrjesuiuUOnNJcn95VTF3Quf1SLDC0skw/ofeIXGI6PKxczN2GzBR
/p3+6RgWuS1HgJv/bvltwcA0eEk1W7sQeO1tFvTcuQtLGwDlodUODks2okEJxZfBXfoIyemEUv7k
UOiL7NO+Cp+/vbD5VF3fccNemH2pKfIs3vIgSgpTLZS6+vbHnPjTanjfq0029KlS6mpQ7NRjRwXP
uQiuQfXyy5/x28nfT1Vk/8FipWAt3HfgxPnOdF8YmPDa1eWShADninQPHJNAK68+bAYq/tO5lwoX
4VfgedfPYZfgDDWs9G9FBFBaE0iocsvGvBBJNgsDY+2O0tejt0G4dfMMpQc2ahMatsgMekLXSibr
+COd0G5UyZPBUGmiqOfEsz1xfx7yqIi9erNGi5cJRck0yXD/Zr2kFrsBaLYozjrCS+9mpYtcgPse
Smc5RApl+EGxIIrCcxwFj8XFxLAU6Z9eXuN8pTLEryfF6rf1txK5c2soFEzNyzhVtZj3uieUWLhP
5ZPvur9Bv+iJpHS+TNTDzn5Sw1PEbs1VgnXkcd23dPgciVppRnzPqKIjV6Q0wPrY3IQ8XzZ+cEVa
paWu91cE5twbwYFXirSBY7GNoa+w6Z6qG64O4jlc8iCfKISjQfGA2ZfaXqUxquQNo6zk6Z6ijkgg
QIaf7pbkAd8hMJHwVQmqRs3cWcjXGQqSbIcidcsOasFsSZrVZ0UX03rLryp68UFuFOzvFKGtooR/
L6/FiZY+g1X9BjjKgFQI6pbiVzKw4h2XPIEDt7IrJa5LUi7SfvPxMMCwj91d9klLnWHy5KxiQwpa
rRLALsuRrMT/NSY40TjJaAAMl2ScupH344wxA/tUyLw8yer5iZbs84yFs05i3m+/tpArbWQ5LI/b
Tn2ycOzB8nR36qr0BMBjNAro+RTQW/YWGhmv4PJhwEfWTDwzwmLBaAE9wIkUYUo+ig9ne930lGZk
qB4OvEr1lGXLfRWJAVZB10Cd3LtA+dU5pzvIIRxTB+mdB50ja2o5Cm7V5qqokYNJOwjI8veJj2FJ
ehWiu0ojXQkJ+mD7pqogyF4mQYwzTRPU9snIwKaTokFcHeys/Ppf54+356sar3oe3GnBlbbvPcUc
ekvW3aD1qFaZVqdcVPiWys5HkhKMtIVgqWUxdBNQBNdKqoRIEd5QgDa6nK4ISJLHadriyOhJRlbo
DrI4DMCyFFTw10L2ixQL7+M9vyrr8aVaITVZ8aI4gkuoxCuQ5uE4BzXDAhVD5CgOrvkWcn+tNqCO
fwPF+esNET4dDndZYssSKOJ0IloKK/sDSt68js+HGBH/6mmhy4Hi/utQLunoq3Dr0JkBHEqNu/sF
cTydWM27yKqrrNXI6fYqPmglDBqmmb+Yb4uK7bkhq93iDdBFdR/8RVADJbfEQc/ZOpbWtyh9b11X
HojGQJGX8UWdzr0c2bDi1nWQIzZAXMYc9wX+3/x3XZqek/bz8ST4gXRBNofsu2iV2ziu0rHBamkO
CjeJ/LUMxjcDhXMoZ+DOQmptrMieIfA4FQzjBW0R8v/8N3QtnJP/+9CK0oVl0S0+kL985QBzs5SE
3nZIoN1BZgdY6h8EWSj1k11w2KOlootZdVSisfvR7BppOs0qjC+YsgcEpwGVhgNi+WbG8HYkJgXn
CiHN8Lh+RF1blt3AAIvzaQMToaMOf2vY6U9XFqOTYFBPyioQPrhnUKK21gppp9grhtla2ce0BQLW
5t9L7qt5yKunm0b7PGowjjD7Qk18hjMMmzRVNjA/0MY0AW350X4ECliUNPtKy2Ppwuo2G3USYEJQ
Cz/18ocFKCxpQLns2GU2z0TNo/h1t6hgbySiU8twhuAjidsv6KYmBpNFMJQVh+5VU62oQzXPXKlf
y9ZPOlGmsWgRDQ8PM9xfJw4PnMombpTZFtOIJmsMXyNhfDI3rSsXs7atHQ6SSTSophN7ZWR8nX6b
L7abv4lOpFCjsibgysGa764HP33uRB6FAqwU9VlGh7lyKFMIeSGqczCEh6ZFs3XCkAR9f/eAqXn2
jqevkStxB+i+7zRGJXFRBMcVeF2LSaLMmncTMGv3ViECVKX9TQ7zCFYfHCvfg2s0e3WwCGjPDE5e
OMkNjpuT85SNAvYmDvL1ZgGitjKxWmWRU/VticAkX/QaMN/snyYVulg18GZ3/fuCd4ea0wAk8ZKC
os77VSf82FKJE6XBW7PU+ZXE4mPe7uemtWNchtfD088nm0oDoDrGg0ngJ6+MCh6GYvw2/rY43y0B
uPT8li55C2acQAARzBJ0Ij0EmzN0QmMaQy+uXFlLxKmEhLSuqc9vlwLM9iEigwZNq46R4HAGwX43
4oZwvWms8jJ6GQISOkLIq4YCzIATtmzVGdSMqlYRYPJ4Wo7x0uG4W5KiIBhSwx1pleuacuskw+ME
sxeVnZC36xp+1R0KvjLE2CwwIuOOdFHoY1TH4KAQCSYs2iJU3PZ8Y7GNwactZ22mxZp3tE5/3uLa
A4vi+4Fl5bolfiIhYkFdkrRLcC1DlSHprAXEd5xTgukxW4V/cXscYvS0eRx9QdG1iyLLRchwzSp6
YXKMrg+S5QEtlYX5dwu9pbpG+Zc6ep3VojA5QU+5hnIACsGPcCtEvf+Fh2tcfRRglKg9qxWB/igM
H5fpId8kBmPAjTjmVnrrnHG+8F8ENGX8OrC5OQOKruNpmV5m3gvXKyjNfAgOFagIiTA9hmZovIwa
RAGUTMbwVHX9LjGO5J4c65baVHN937oX/sNRe/HCC81jlJcvf+86xwNAE5UDuKH7IJeg4VmUMLXs
2rrLzWrgK9yuNXbFyP1yxKcQw0lg3qzHQZAv68GkCFaYlWhgiAdsfKnIZIlGID1iJdwAgRxS/aO0
Gj2SWzRNgDpBTymrK+u0qhQbjJDyopEmUNXbBaqSRzVzLT6OwKWTgTIcVxyLLNLeW22jwwGjwGY0
wnOkkkXlYN1W1T0eJOOhwke/T2RmpkpDcRv51QqbUb6R0Bx2PykVxHWLJV2N91Wp+8a009OgZjEe
xM7I5T0CsVuXeTCSRJ/ezkwUmC5mSILsT/SQNRVHxVq42t8Ep6Jw0QFF7vDFn05jcW5o5X2ESlxb
jApelQj9kjBA3o1VtPGmMpBeckEBu2W6YU8fW97n4hySn4XdDt1B/Ly1eM0jV1yva06ZlVT0GvXp
fhnceM1XxWBU1qFwm9Y23j+Mi4bS/N20GfP4dS5FbUJmph6imppr+/XslxNU74icpIzVAa4xFedV
GUs6PyW44clOvO4chqDijKRDWcIh4Nh30A0wOKuXe9p9ZruuxtgnvRL1K2dNg3cBlpXhX/85KcgA
I/f5aerf2sh3lEWfQKBvm9G7olkH3+9I557w2FxMaqSlA0yVoVFiZxvnXpLqCRV30hNQv7N2IdoO
5SLOfdvBtceFikn7t7MrslQxdShx/K+VlyJxtSZIqhHHfdzX8HrwKaHndiyt+woECQjUW5fnkxps
WVvg/QhEaeB4mIDbCKgJCkThTtnASh3y9JTwZo5BoNc3Gi+oQMfHo941nYcP1srgw7voDW+NBTOG
L3lyOoCp4MAF/RTVlRyMbM/QGN85D6UbO+mo/icsALoIe4jpNvhLHkre/S5Dac0U/GNZDEfrc36f
1UlEUU9Xl1wqmWuGTkJ9dkff0W3dcHpAl39Xsu5gfXX+gOocfEdI2xqa4sN/QqOwSPAS3D7zO5Xr
8ALc94VMJwgkYIB+uzOkTKvUaq9lgupP7vN8DO+XLtRO3ercRbbLzc2nXgZpxYfh0Mrqa7SVgDMo
njlhxvH69CIbkeS3kY7FDhbTrghGBjeY/gbYn9ZK1K/iT3FVhJkZoAGc73qLJpIso11WgyA0Td0x
G5G45ugbebMq4BpYHi5Q+5+nn+WTx4N2/nw/RNjQVuUtZLF/UseCN+Dk5xHzjcqxWPfuykYpqMEO
ZWgnC7sEwj6qxudmmks6yBDD09RC5XJ+hjdQ7ciAi2QczpB6yal+zb4BPRXloZRIp3Y0B0LVxHbg
8lNo2evBjmvBgSX0Zh+Ucf6f1Ug7TH195XB4Jj1fWfN9NeuOUpAV3jHTLAlXfMcd/ByK1SqeLm7K
rUqVGpKKt7r2OV8PiRj4gOu5dlVQP3Od1i/O+pyPMljBdY+xV1UqL9mDsQy4e4npiUdeNUgKg07b
Eehx58YXGo9Xv6ljY5SCJrCX57wqhdTLfWeZNU1FZ/bLSHvYIzAjuIFLd2QcB6xUvM9t1nT878cG
cwZ1/+LTiFFWi8WY0snsTSP+aFIrdvZtuHTe076W9eC/RQba1p2yeJOwmug3JbC2ZwtYbCrnhLLv
Czz2vJFNc090CVbnqaP0NvyO+eF3I4WiKiEvr5KnErS2V7JdOja8LAmz1ss1fZ/3ee0NOD7u8yOk
Q/UV+CuH0TP+7K5+9DEJR64QItb2zve0ZdHZ7UpGXtBIm7NhEqpCGLra8Yp5dbtLGz4i4WfJt38p
5w0oPFX8gWXD60HMsk9msbcIXPWEkXx5o0gXk8MIQomaN+In0y/BnjBo87vmLQ9tcVz2lU6Vlc4e
CV95zS1YnWV7NLLPEGOGo3i0RNMBpYy9E6sRM66sObg/83fN467lMLHcjEJHrfHN9KS4gYTyr6nG
i9v/105hOjC4cgi7Q7EMkWol6VSVMDiBR+yk3GJTa8/ZLIxNSQstcVrB4H6CcffrSXAmKm8lDBPS
+IRCgQCdhvFT/dWPld+H8uFd2lcPIn4AjiAzPd8c2Sb8qwWslmG+p0hWYY8crXuCqCEHg99C3hbh
6BhdSiqhiQ8/yPlOPqYThTh9HQY1jGKGXguY3L/wABkRDQxYrE4zYAoSJWN2uURX88qOmvORtj/c
VSziffR9h9giguetcbsM2L8LG93n2DVdM0XXYL8VlpaD6uRXUbbAG3+ClQqULk3brOMGwxA/r0GY
COoXMMtoB1uRkBayQvA6spcujNLYv6XaCsB2Wg2ThvIHMb4DScCM/J6X249QAOtTb7oZ7GFEDuMD
L+fu1In0nxcp/QpFnSzHVqUg8fdNthgPcO5TuPBgbh/cuVP+MEu3+qelfB+A9992qu3IIyy495iH
FXy/yxXeMUivigd1FNwXpZicCtjB5oe1+ZCtyigc8ZpJe8UXo9OP6VaTecFju0hnKWJiD9YURets
xGfO9GKJqscOHQ4mT7Pa9LBAoiOKcRXeCUcloRlqvenoTeuRlv/Q9dwJ0vSFn9RSeER4FsOP+Vt3
Aoyyb58qMNqFRblc4EGs3s9re42brUhV+egQvcbX+KSzIT8sGfa91absRTMXQEMm5NIKJfrQeXCk
OE4bnkxDnk1P/pAw+ZASYp4kHQLJyOQixQK9pPJyo2RuLvw5acGMUanRVN7QIB+nx+70/1zUdng+
K92P08QbkGR2Oa7vlRXjUPL4Dvp08G2IhE/0412h4W6LkN33GHbLgRomcz1x057tdjHnZPW5ScXJ
Phf9wLPy9FLAEHPFEIvVpMo4MooEyTkUi8ttJap2pYfHhr1RltCnUamP5jZVUS2mNEBP+GMcSL5S
cU8j3lHWKa6uxN7VsXkvztEn5YvgI5LK3X4c23vBmmPggw4Dj5yrPJlkEio68vaysjHg5b5l38f6
DxDLIwEgb4W4Wzos/fGFfbB8+UxT3E58jyiQV/BtboPUtsSPz2efqvXy9o7Orx28BbEtUbAF7TBY
sZfInWuNI6ATaMDsRoREBbudUwqCr5BV4t5UtH0cCRn3mHVGzMOBa55QON2HvG1Z1kzbOEuOozgE
jyoAxrz2ZhI7/aMaDA7T2p0Xex4ojvocGOSQ9GOIAGAjhDNxj4tKU9q/gWkLlTva80KUczZECKYb
tzyTCimmLgsNZAT8Gj4AqWi9uRiTZVj2ds0LBInB1UeJe+us4kXAjmHcfW2K+IEYitfgfA0s8vrA
8hJlge5AUPL80lhhqjPLzmvpI/5GjE3pU2ualCarSzEyfrmY4hAyl7Tr4HI0xdl42HGGNfPtQRKf
yfrcL0irj8yqS/6DAMPZI07u3SiKkKo6Oj4rY88JglWqexCWWvtDUx+3EL//7PxQi2qK2+tuw7rx
dpWRVIYj8a0QXvy/iY6GGw2OSSIVS4IZouGXZQEwAFSKFEmerSpo3lnSqr+y19IQSKTfJDvfzLt/
YEDPSZBnJgGua+WDIlkAI1u+lvBcXAfbDqurBn2ZNIzragQ6GLQkYuMxW2GruiqmQIyrViN6zpuc
CwijcahtODRr2yPGMkHi80Ed3ulSOeCGGsvnKHB/p7FO6kmTnmd+bSnV1hnFLriBr5epahxqpDU0
2u6FrlM5gRQFu1D5X/G9YBd6T0Pk+2Rc5cQ+E1DWoJCl0ZyqYyr7eAN3e/Z+OWYsOwUyQgxx7adV
ygd4hAoZHIK1fCxAGKWpnbhAyE64YPqEt3YHwWKTjxmUew12QAr6FDIVpbD64wBet06zCJhSgqr0
8+xoZHMHpOERO1twzlwYsswTtZ9OMaiDsWEDw80UToHPsId0484K1hRePyHbcFsTXmPM4QbRXMrA
HAJDzMghmlFtHRnPp4bhrdrqRb8aqcv4ItVH6dFsGdm/OieIEbVwINJRgk2ji9TTi8ZYP40CF+SV
1GpTTxyzm3VotpE/xOtsH6iOcIehl+GvX8EHTZZmDKNA7p0ANdLtH9DgWBqJM8s0GFCQ3uf/Q0Ro
unNxeEOHj2jgVrvMlAAKHiAX4jEysWEAmOCi5ezNOrwM6pBl82XuWrzl+J4pGBkJCSm1kFfTYkPM
TilDY3mcBlIMvHu6nsssZPrM94A2xhYpnUWAXNCTlgt5IJuxE56I68kTuTS8Xu+q4EkjvLvFHfO6
U80zWbtXB1wy2xvPB8nWpmASALgF+Oy3LU0uL+OObxnbCDoOqEdPtrxHwHHX4E/NbUtJiHTMj/EU
z6QkxSVykKPWgR15rwLToPJUAS0xV6OEwxUQnpZ1xHi1j/C0eGB4ntXNJyDKdxNu06xDHhVIUMF+
oHwqs3E82lDKfqOaawRM2A+YU6fz8teyZ48leVsLg2oQo5Xeo7pvtuTGPU8vTwuDE77lxmjzHGyL
s+Rm2FP411TqATWQ8uOTgC2caqJhGATk1O7V43obcnIxMp9LXaYKdrM1giKONbe59kY2pd2Q0XcR
bZYCa5kAs1p07lBqPZCNU57Gx8GyNoHdO3MBBgEN6ov/wccD+72UfjYYv/xQrNmqeZOEesEXwCJW
gvi5HnD/NaCAMB+ZJfpKxwXu3mPbRX5fYCShAuUvnZ9kiS/WiYyOdC6Wer4Cb1KInnSEuzSjI/nr
2M1oiIkXVIn418L3Iv/BZm0enmbuJf8Y+08qokOzI9yBDKOFxK2Otd+NnQ34b22pOI3PhENdcU6H
GrcbxVSIxNHTRp2nK8q7Qqc183BQ8sfgzp8KErnn+uhYOM/2i5G6ytTojUyfUKX48oEU9H+PIyt2
b2VjKbP/tpLag1zMVIblx9auHI1W+iQdCsHNI4Ucor7lGDLiYRaOv7I3Qp7PKbYFD+0MpYk5xFC6
wrbFGwalYOzouhhtjP/kJb3uB1SMAANNoAgCnIgLKcBld2yZtXelXLsuHkTL6RHFIYYUQbhz8Wus
VFcW+7syjeph8DnDN7q16jEm408yQBbdNYetsMmh23JpDdyXKIMtkHwZzMMXemfrM5htbGR3zbfH
DtdHTLExI6bdC6N0ohE0SDbAvOgI4Ob0r/whXFPoL9ee4Zs5f1SNlrxHbk5/qykcyDKj04NqmFQo
AwsCBZWVU9zuETnARELQwkasbgAayrUgPfZoqgsj+prXDLn0aaMhxZAm+eLGgcojXGIhndCSWIha
y+dHXINvBYCn7mSbGpHGwBpJj8JqvomlcmKsTZyymX7gv2FSPN8iJQYYl10z6J2B9K64vz4580SD
SlrvBTMyXvfDcz+JJAfJSbThdnuaBucqS4B1bzurqHdr7eyQ6zoYkvN7AlinoyFu79HG+JkFC0ia
pY0xxSIblID9ByqdUH4EfHiajHmKVu8r21bmFARwmm27Ceqs/jZZJmYurIbLgzmKv3mLqZz4iKxX
HSJnLqpvajg3Juc5nT8WtOv1gA2Ww2fY+fvKk2NnTnBJm3ZsUWEPD8GFkYhXq1T3+4n1xPo4D41p
vdhsTyn2zb8JlY3cIIFwl61Q6EQFNH65vFFfv/T8x326q9GdcuuXKHJU+Kl9J3FZThA22UlqnocQ
MBEd3/dA13OtMd3r5LsorK7VrrFkXUJkFDoBhHZkUHE3iEtyYxK1oVo8WESgnEhtrs7wgWsX0TlE
9oSi/HhCzmXvaR/ixnMfOXlyDU8QceUN4lybxr6SIdPOTYx1Ni+MLDW+SXUa+j1otoJ8L2GYVUwU
SfFano7saeVeIw/apbTJfcR0vWxW0aYSGDiu4TYwaqaNgugD3P0aUOwNfUZgpjHVArxTLmFiXQ8T
jviCEIpR9ikVi6LwTpvFoWpGTHc7cvVVEbpog5Yeyi1KVncZhrAs54lFUR2QD21fTcctCaRX7O10
guSmVrC79/ZFz4tuBkAGzB3X9oPoKydqhqyEIKp9f52QTIuEW7KtKqLFII9azJrpBsPfuv54cOAd
SqpJn7ulwNvuzPCB0TthW7hTbIIz02FPeiV3j3en6DPPmtyxsxOEjpbw2L5URXNelzkAkgicJFVR
2SATIMch0iLvbZVWwOddlb0fTixY4pJip9XW6OBYyrZiPBISsbw5G/LxP6cbd/ijG/lZN2ZhLnzr
8SI8dxzrcEkhpr3giCFIqlL/7C9d8L5L3lMnhj+AmGdMJR5a1py5G1SSrWrKMdRcsFp/7F44FZ2B
J98VGNAhXSkRpFa1TWgDfFWv3zCDmZ/4MIqb21HfskivrOlrjlsxqRGX5i1iTCjIHVo/jkknoqPQ
Tf5JitNJHgW8PpdACbibQoU/M95KCYsvkMUBy8DIbYcqs0KVvQszmkBE7qn+zdshZ1C1MbcTqCuh
FFLBj6wV9sQBefsIDncQpqk2csaMEhZaf/MA/rjD5shFNsltY+uC2aUnEKrhE44OW8txJ1y7K85E
DIiOp4S+qBBLa2iJnOZn2VEtrhHKb/ZInr7LGl8FNBsUhz4zPMG4FKebe8U344xOnJrUnj5Ks57v
JRroIUlZspz1cVUVd2+gl2PWBi9jGgHp+0ihU38+q6cCj0XdmCE4Cso6+ZCUzflcAg7bXcxt5EP1
QdTEOFos1iLxE56TA/1yg+4TGpB6fi9uIhEskG8ae7MsTpL+7myFuEbB6y+uzWxm/XPq1A0eCXr8
qTkFZpH4LM637tFFI922kj+JXvT5noSNYEpUG48Eq6qXo9pbiIHfmozmxgq66a9Eb70TAeVPZOG/
GovvkI8gA/OehkhMuZ9wGj797yeDgInNNhDPMxy53TLi9R5RiVALvbmesnUyBlBChCBeJYPVttsX
SMqV3MZbI36yFcs078QbMLIk9/RbGEFhZXQHv+zYfJ9PTjkXEFUVXl/8Qg9DHzsEI/LlAfaIH9UP
Uws6SFtjWdqLD4liCZi+uP0NjEGtzwiHc5TCocQGM7dTLK0LnCDGgZif2rEI6u0A3Rtawn9gBjIp
TN9vVXoX0/eDQeyK3hdqXum0tK61H6rCa/1R3mnyGUJLaBu9hiV0Lh1STFP4bPHu47lLH4QS7QyE
wgF+e6KpklXGNK8cSsp9QHwJJoNtX19h0z0W2hAv4zR2NbKcp7w0Ul/l8HMpeSMDAEMs+ZpY9TaP
1WHswtEkoMIdFSYAJZDorbRAWA+LAK7c9mhH9nrq7q+GXU7ioU5y7oQIE9Dd1+VWrw6WF+52h9mL
5XYZLfY5xAyWUYp1bhsV269yij67gaZmposfnvWGYV0w1AQAOlkQGB+QdzfxUDYnyW5L5F00uhMS
vJpXxNoUxitSVOcLQ1nBOH7skXoeA5u2gpHsNoD3yE9aAjnkCYRG7Ybj6+JIOmFvdb+bqU+AIzhe
p2xIfhDp/Bz18cMqA4PoYcFvU9rjskKTjp/43MR3o/1gflzJ1G5qzgPEQkcBy1EoHV3DItZ/1EXo
yuWVQtGBQMeH29Ud+dcHZQF5BXJjPMQkn4GSIFgqn9aWWBgBp6uxeFmifYTEI1uqEmtF1Mr2LANK
kug02LKNFjcnrRo2/zPKIXfAp8lozbY82cHG67Gvip20eLXl9+I5J9p8Sd2KK1OvNV2xQmRTGnrx
lcHK78vMl21OpFBYuEqLSZXsQc+pZH+sUdD9bjhGkrvUDEAup1UmMQUXtJXqWgsu0PfgYDJHu6eo
vxtF3ycvNlyNEm1YAbrddFSIErKnm2vzzl0k1mV8EOBbiDOkbawF8lLhCYB0yseNUGgNWThlwVn2
CVBTQzsZHXkziV5+mJFNcDcrIbxbE81MFXGrxQI/l8OjtH+P1u1lJIKOTyk/8xFr8oho8++puOGb
mRI4PWMKRekN+8xMf1/TozVOOBPIhi1vI6ng0yP+XCWOfKqPvpmgBXIRmfMjl0dzMvRa5Ct7igVS
7Rt99o2fPieVMx5XsZQypNSzbPEVUvxmEqHZfiGIO1ke1HGTEFqaqYdJTCkbuSokc3iwhNSpibyv
EQ6tJtQGQxfgXSjVVDHZLGrRzSJ53SF+St8aXsEkWZJuK2CLAIgfmWdxnOWgpv1hZ1ylFGegFzPb
W88yeSxva+mUtzS2F0vFf0vhivuuoSrvtb4MLx74APn4iLen5ycUXsxvHW5wVi5mJwarslBwlsHv
7OftGqNcy7AK/R8mUh3cmooSFZc1qWauTXeEQmgjNy7Nq5KCXg+V10yaZRx37Ki85NXccuAU6WnU
e8/cWvly4tfAVoiaD91LphkUFJ5CAN/78vUt+kAZKXU6VHxy5V6biWUzmWVac79z4Z4fHgSj3Pat
4T9vfnkAlZpKY1XS1WzF2cXjwE7Y61hv56ekl9XPJ/7C8XWKcweZ26+Bl4dvf1EfHUMF6vZhmN4J
nErwbtplI5XsczDdemYn0+DlXYbXOP1ZCi3YErBfauL8aFVcf1lJpoYDAauUZSPQkw+3MQXYXuP4
YLgSfOH69420qUDVIQ3zSNAdLEu4+Y5dBIw0ltRVserfRik1RUBqvfe4dsSdYak0WCdmwibA3LmM
AuqAuW85MazD3Eweinw6VO4lw8d9MBurGqRAKr5cSbvSKe/g21N6E8b99SJSyMp5iw6KGptJ+LQb
nikSJTukQ1P/jrzNIFPa9CWnXbOQ9VjtdToez8AweBoH7pjGWteq3zgFhE+8Dwhr55D7/ReGMdgg
oucmcsYkwi0S8L+XrIKfIKStvKfj7/gwWQlG3vQyXrQmQyATYTtqkPh2QhUQkUV5/nkhWUT2aAmH
vs3UafJenVS4kX5fJjiESCiXVvXWvRazGbpwL437zLUUNBZzz3/EYKBrywR3H2r9zvF8VWzcDKR3
4Gnowxx5o7s8DKJKgtNxlp5EkY7BWG1BYPGwsJZ6OUlUSQ4NPxUTaC5/R++YGJ3LvRO9xlgeR8z2
8MpYGo2+5g55jpphnNIUZnczwsHDLhmK6WgmfncJJVoD6UCP+r9ZCGRz+CMOYOWiO69Z1BFicjE2
KxoE5rEH3W09c9MAXABPcDCep/DdVAvJwr4Nul23YX/SpFQzpnu1FVeSoFV43lhZgFKlfCSS9z3Q
GrIbC1YCroIDHEnzlEKWbkAhVCrJpN/L1b/nATSQc+JfcbWsN6mzJOgx96KCDPZuzH9Gcal1Mern
onhKO2CiOeg1xp7UoZJBeTQ+mN7kCk5lBdOX+uvBpTrg53qNpbNg1orv/3PrnNpHzL5dpCk32765
f+bYdVyocMBLO+3mODlHa7XklLUhW+Dsn9Q4Ls/k2thISB9dsJTFb0iib1YTYe2a5+PtoKDmFkZZ
vmKDnQaHl87WrpmFezATJcPm0Ca60ZUVnhT+T/G3atpf4jdeZYfi+zgITfmjwciKL7a8UY5TwUhO
pKEKrGGZbAojDnzqbS7pEKB4obYLapGOgbyhyAIFGHp8MUQgoWOBKDdQBJeHlS5qXfdfoKzgZ67B
yKgEBp1gKd+deyFjMUSceZzTyT+2pe/usxfs++qDqcA2d2FwQhFTpbwkDblkAj8IADSRZ4fQ+Gcc
VgcLHr55Qg2QcmPQYbp4dbXYyfF+FkayAqBgMzGUxmrEZUb2bxhWvRgUhicRf+dTk48AP8lEHJZ+
yfsWYbQofeXTHRuciDO+mzasmiIaRqiE+Q6c/EYJUPWfYp5RlP21rx97iP0eRTmIEOiB4J7o78qf
HM/GXOBlzrGSD1Wmqovl4Js1szZQBT3uo0HiD1iQA6gbiGTnHNVNoLtBnjL5eUtmpJgKMmNtuAfK
HnNx8tnTlYas6gqrjaGEA0U508vWAdpthsOi24dchx2B+T6c1hhoD6Gbz9T+SgL4yG6gkustrvGn
rr4dvWYIG5TpfMcqPu8OHgMoh9iDjiWVT93cagaW1713NuTS+DKFZFyyTZwTlLKAgfhOM10D6Gse
BPlGJRts1155UB9uQjeuhE5xnAd+V5vYmnIRtK+9ZhPytff1gkSs6Jk0aHkFfOrRVHYh7v/SjoY6
vV/jUDQWNsmVBDTG4F/aEvqtChOqCuhC+NUN5bh8L8adRiqeDxdc+M9G8hOpKLkFgzF0U8pUuOiU
UdoHwKmn9+BbEPUkM9vklHIVF8s+MYp8NZZFsn1/NV2at5ee8Aoo2qZDY851licoydUbAr7OlmtQ
c5UMEFbleU941K+ORewYqqRSkcB7CKQVyU73jeIJj7FP3ykOJgBwV4uMMaDtiKPsANZqLeDyUkK+
AKk4K3a5HLenHDSpCnLS2WLnA+Nzz5cZ1O7gTllasf50ZERKwOFJmeORzv81p0XWBKycvELzfC/2
crJ8QiEn8o4WbANK486ntrBgclA29RVb4DM5Z2efmkpN71n26k15+W43of+gO8rmYeg3ciGpMBXm
ifQJ/kY4dwD0Lc0eQXQqifjTNP+AVmulPlE+vHHHPE5mqMNNQCbeurghDFDg5OtQ9QK8Rtg5+CCc
HEmggdiO80uqgNenPNixckRbP1rZfeBqwCXDIaZwXqfNk1SOtEFs64uik8fVEV3VyXqcMN6ZngAa
GMxSx+hHWgZbsvo0rWAmfP6D6htzM5+NjaEUiCfIM20i8L/7V5XTHrSugN2Y8MIK7ySn7m80ZbC5
c965Sv7YcvMEfxe3S7NHJjqxTshjgsW05EIstOLzZ+iMvXJE4JhO29Gg+YHXRSn4feRhMI8pqOL4
ksbG4sHQBQ5ipsIDS3w+2A8YaaMWZVFlGtlVGJz3sCQ8NPJ7tfyftoNvs2iTK6BiCJSBV5+yRIKS
meyDT6qGD2XrESJFPpJaOj0KdlOWm1IVF54TG4m5s/QRav4IUbQC0aEKutKnCT3k8AT4GL6a0B9y
0buCNLUvbrwqOMyO86v2H/dsCJsAnryBFD+eHmh1oA66uWd5KzCilNudsnyOfclilACz4QcI4JlR
C7gW/7skuIaWKSbMrVyuITzXMqX/XKtllRwHNyMOnZKkmrVDhRRxkA7MBXgtpDy8vcJB03EFmEWW
R/7lzmMpnTibgu9p8KNh1eUdwSSUzHBGureu4BRLE2VUK/Q4BoMAFa3s7QeCsRbhxXGI/x/iEzOL
wSg2Pyi12IvhCIebztVnOHtTZ6HQTLkyBcaK485VpzAKwJcVShQTExx08ZdfS3z4gE1TswoxDYHX
svoE3nhF48OQ6kgQdfxuvE04vnyDdgRpktwBLHuuHyU60FectzFyEfMeATyE+XU9pYmJJcCzJcra
a+JEVtgrSFztS7sVkzEMzwEH+pQJU86gCaVE4Ym+1VKIUcDYxXKyaX5v0rhAtRbwtVDhBIRiM2t0
mqiUi929ybSey0G+Eehzx09k9tXXriAVxGWxi/JbkYNo/tx3Bpl/yVzACBWWrdzxYvwUlZZE5ro+
zxFnIlpsZbF14TFbFYCFqjBlRSW/IYzt40ohGxc8U2gPqFuGLhO2miAlcWAf7TZolQImZx+u56sm
qOCEepj6iJXD31pwZ/t5JCjOqZWwnLk5+Ibwq/TC07fszVWtZr3F6UXY7SeMx5sz7kouSG7s2IWQ
BM5dN2XcNl8LNlwkaKqx01x1qYqyLIb013zilwlHb9JE2doBrOM8zS0mzchUma+oz8gIlAWB+Jv3
nr+fWb6a+O0fBzyV2QdLuoBuHDL2O+LSuB7SyxCuOfLzB0i9tvFbq9DQvMu9dpTyPuoerN1sOttT
TxfuZtUmEaZZ/c4dKPW8A6g1c320J0+IMirfUVPWtdpnRwhjNb0c5YlNjlOATbbzhEVK/ZXR7gbo
YvfgkDr6UvZ92XJ0h0I0BcjXpK0/K+fZbyRaoYDSunmyjEVHjLdC4LEDNN4zYNxcAT/jLccKmHa/
gYE6SFQ+LJGy68ajMdioPPWkFv3sYdmUJenI4n4/Gpt6QtHnyZVTHb/TQDeSIYERbVXxFDW7Ld9m
AenMnVZUSA6e22SHuP6sgMJESgaz03ZCZqFrpND/o/Ue2huAH/WsGUQJCLZb0hA6zvtdwWTQjnYU
BfR/TRXk1p6BWKC/WSu9FxFu8Og4cfS6TD/SJ1WLXyQAc9zrOkZM2ImZfUhBgIy5jkUeAIwngS4x
pBrUMcgLmwWMwynfYUF4t8rz0yaH1b4+pe8mRHmInWnvsu7YI/niT2jXOFvI9GFI6S9PL1Br7Xd1
7sJcYOknCKlGh2IwEt/E50IBMovWsFa92oBAHUk0iDzVRLjOV66VE6iXV7CTZr1aj7uCCeBr0/n2
wgszHOHjnUHwvFGnAMC2JTQE270kgFqvWVb2BZU2/z/qXA8XFmf6SuN27xThoTaLFS2KRMv5cbwa
TP8NEFKLb3B2i7EIVcaNqN0C66yGIsikxUk5AzU/A/GbpTIgV3Vs1Qe74sQ7ZUDSP3GFD6mehUYv
HSvBAgzx8j95m3rVDfP8nMrtjPi7YY7wBxdjQBrw3jkfPaXM8k7/AYf1rlgs6RWTU19auEDqnv+E
i+XfBJr40f7emstTqTYblFP7h0fKCUcLPC+e9lUayqsrOJ9m0Cs+73irrxDkDCwa6kdcGe3aID+f
9XRyruRs/YsxblfReR6pVov70aSLhMsPKwUoreZpiIEY6mCqoZBgZdrtabhQC3Q/GKDvgDQJ2wzb
wh7kp2uJM/VWHWDlAZIaGf2dLetn6TKbM2rRjKlVLRNHbJKWBdrkGLpKNxx26OSjkBv9HrnFDXSU
hq3JxpURQvkq6cbJpIEyV1Aji4Yxs7j/PPU4igFEoJXYKQLbtXzQGiFZDLZx5E54xLekZk6l4LJq
EpG3mTvpmZE1VrVNT7lpM0YyRGXyj4iqE+SJXT7YS7U5lyC+6xm+tKR58pbR0jK0QUXS+A0Fj/0h
Rv5H/GTHoE/GZCu3F7ximGHc6MqBgqhliSVWfiWfokS8QjH8rvwCJsZfXDJS0Qze3sjSIUkShKvC
EOCU4j6F+dp/AW9QIO4POGI2rnWLO75NVTHinXKN3ijFis7U4xVRCBOkt87xwAhmzzMAnnGTMMa9
8lIPldw4Iv8b1EIBtTEamq9c5JJP/l29dZ/uv+BXvREnZ2UQLlx25U0RRlsitOGF1yx8eLXOeWnh
Krvx0SQ65bgW3Pb+wN97+07rXvTAg2OznXn3jN3H1VNkPTWojoqdDfu62hqiRU9VJ4mQZMswZJqg
RyMGrj42V3H1dUwrusdBJ49aO18goBUleSAOqpwSLC36spQbJ8VEToUAn522fnNNR3WZoUgV82LW
g9YZT9RgvDoNPHxsTKZxA6Bupia+aQbdyC8Kc8iy9ZXIDomHWcfhosoNmy25Oz/j6h94VdeTyLau
xg/fOqvsncDgxWSyTtulXDC8JwfZITxSxXlhgQZIl2G4edzu8PtC1gTQNoSgGESTXcXNVs5VKu3p
R8Lj+hxAWY7tr/eF7UO/J+WNA5QXlHUfHgkP0uMrm5MvK1+RmpqJm50d8Fknu43CedvV886iE49A
6zufA4jF6Auox7dmkTB44hG5GEu/MHoEn2+yL8xtx0iWP2oNNqD9Gvw4ORSwf/i6g3oA30nTJ2HZ
4YtoxbxRj5gW9/a26FWCXjOX+qIWva/WDeHpenCaf00QGUlCDKapFQGtdAte1sU4STpgz9QPM71l
+n93KVdVKI5PwNYPmHyah5VK7VwmEXAgKRTZzBs5LUAg2CflY4sxUdB70wRyaba0vDDpNuKrgbXm
zz3vuYrjytdFQT1P1MC0HLBRx1qrMLPAjNBAh2VVGqHPuW0jdkkQgD4qUEqQSpTLFgZxL84Iho8z
iR7ZaW3m/CyarU2D/v9CX3t+2MwiBPW5pzkPnp1M/B+Vg5sDszWqeBo9QSjX92zwQy0UgPneoEry
dzO8WOer0OCi/F2IkAvXxWGwWcZq9tXE06h6ZJZMi3jAPWRKO33ByyMAi1ET5jJB95E8xbKilI1u
fmHRtffndUgxf0zzxHAT3HHBWUuSWiEUSJazsicO53e2PHhQVxQzn3lpNorLyjqWugcLXmeba7s9
lGoech3stCDbJ0RmnR7lKN94/NLqaFz6FlMRwz8AGLo23Ttn1Ny7/hcRQ9jFWzSgeILuJaEBnUxO
noAAz8tYbK8BfEWi36i/1c6Ju6CGKb7OWBOYYBnJcYUSddRBUm5YdUk23szDHq7+cV3Kbxz0c5lZ
sDLmsFe4v8TDycr1G06vyd9eCtnxLWa3Agds6GaSzwKAirFv3WRWwF5YFtO7pnI00EugdzHPhnje
3ONYf0KIej/E1XFJyTIR6CO5hBOPv9pdgLAXuG0FuMERVzPUztCWMLNqg03z4OrIrQRcVLeYI03v
JBYRIOR9wSIcFfdB5ne8NgCOkqP4ImFZ4qUhE6F6FDfGCnyIjax9xRv8XYNpos+Wbq7jlYSh1PqY
qVtp87G1DwNEs3hgdcECBuah22c4VcZcS5OGFaP1Ic3aPRVE2RpdWS27Xoh80nGNm1aaiio+AZN3
5/iNzKRRxu1Bqq6/hP9/TKgGZ8628HfjRPkISy7mms2w9cw+PdBvXmkBeEDRy37N2BH5wf9swmNW
HJgydnD42nknuTiBW0XjalkHm+BtiglK9ZyV9Uca/mLlrraJQiq2DhGIU/TJKDWHFflJrRvFMSy5
pzUhCKU3k1OYFwu/x0tJ5Wh8GEcHdk8VhX31BCsmAtkPF9gkEFjq6v1quGJS5AW8vdUcCzoCIaDv
XK9hLaOW0iafk+XXHucM5/q6PckDq+4jJOxxeF00nXi2WYVFI2D+CyIc/cZtQHK79ZFUxHvFHyK4
rJFc4Q5OqjLS48rB8pxKK9y8anA2EdXMX1YNkW5d/L059rJ7ZEUqX3skBkdRPhXNlxN7XsKMfyQh
O3DO0biVhPJ3Z7jMYrjFNYWDrxvS2G+O8ipxB6vrPOrrrnmAGNI/N1MyKZfZLWWBq14eU0hmuXlj
IUI66NVG15CRy8nMxqreuYiZC9X4jsqTrYdNiK1u0qZzsm2ZFRgG1LoqBY5wS2bYlTkTFsXnKSrc
GNJUGXZaxROp/4qptq51i+wn7D+/uQeWtuAbNEW1AlTor4ag32K5VtK0mD1CHPTjmefjUMICpdGT
5Ktlg02UT4jNuhCESYponyBqqb+O8ppi1Q3M+8ca7vr/KR1ZMdeQc4fILVe6ygxFP0q0qw6iTllU
02ssZbODpP6UflD08Mo0Xnx7PlJ8ihWC0/TQOOYcYl0/55TVyaLMchvbv0cQz6QA5YTrvJTVDa53
ktAYOd9n+JpDe3wDaopQOrwvIyX4i8SEpzEuUayrEBHMcawKFPWKxXP6VT/hHpcGYRyNEnJh0ic0
Yofx9UJo70buAzZnmrK07ovBhanvIz2aItgeMXPxEHb3Nq6poKpcpssMlcQe15tfOv4meiQ24uDt
2X6waU7Uis3FLfWplvFjnWpHQ3E4DdUjMvl/kCndnA7G1gwtaWQDjz/J5E5sEgA/SC6YOuCRDe4m
z0cM48znzClBFpdNsV+1FwLc3OmK7YVb1PonFf4COCLAA8/MkwTHMJfuw3GZUhGIQCd0sACppVxd
S56/CLfNgI+eSSjJFVbQreOXo93vNaaRhnnDLt38INm5Ga1wqMzr/XAVkTRW4TOXiVp7l54mblOA
xSOc+7HDcHHtYN+m3eBPE9wL3wx3BjdibfTcxtJjDlJz7gfi/mlINBrmIvcy9R1beKm+JU0Tft66
jssOmjJC9E8CV8joZyrYZmDcTSKGseXMvQ6M76luXY1mnHzamse4Wq7GedXvAJmcOpn2Xuq1tew5
LRz9c810w7PZQZCWznL7rtqsLXQ+mP5ojStcrm34Mkye34SxUIAoWPgmPkwCUwg3k9cIn/Dk1cDR
1zcCQoDH5X3iDgQeBWaowGr6eqP2yVozLPK+YRiv8rqGr1y61y4Vd2n4JbhpEQ2wJX/nN78SO8Nn
1gq+40nLxMy+SFlM+79Hyq1Izv/MJk1DKmfa5i79N8kV2Ie+gBdB/9WyEEzu4Fld3Wt04+NPzoOm
qzfVydQBW9bXb0HEpm/DSGos49uzhem4Prm4tqtOt8C9U7+KVpo8JfXjDadhhuwqzb2cmjBb9xmV
GmX63p0Nnq+eCyRDEmu249ZFeuJYGxYPzVme9to7nbib5N8CbnqSZn7WJtMt1ZnNWwLRo+JpUsbx
GRciWGDdtohIkVL4yyeZ3pl5x89twO1nx5ZoQADs8g9m3+QIADWFq84/k7bJXS4pHEaWQRNErVLr
RrbsvCqhH2hyoePjxfrzFx8BhKzRAdL59zXgaC/yLPcnlQBNvZhBrnWO9PsrTFTEkO6g1FbKI84W
InsfTwGO6h2PbYHekAcU+wuyHyWuD6j1qvw4A3pQobtw8t3LT8lPVXbF9mEOHbkVsP+HsVO2S56D
kJVm/BFkRNj1iLiQ9RyURbOu972iPyx8eSImkekAy2Tu2O66OFTkMNl4bBf7OUzG4L/oH733L/L1
VKMDu1+ICuO0jqa/ozq0iGR5xlTnCPUrrcdXawT+YIz1ZqV5Fo3gUkaqWWXBwZH9sV0hE23OPwL6
sPM3gSRVci3MP8YK1SUPCVN3pSag2w+of5evoyNTmBW0jUWhgpji7vVylnb710TDJC2vl2fp6CMj
q4js1NjJUk27R1g/SGpTFZxrRqmcx3Hyb0RlUsoHO5KIWwIkmPziRLYW/ibfp8RfBEtreA9J0H0O
kknKIhnnBaW+c8yB+X/Ps3WaF924xNIHx+hVMfs417y7WfaMnS+oprdhlSlrqozLe0+PmJyIZAMk
rUBzb/PYW5H9+GMCtT2bPabrJGdWGQoQih7nhuAUFKmjN7u6KBuw8QRksqXBeQi5sAYFOHLKUhGe
nqUzdhlVR9oIUljmoNK7KGk2j3dzZL8ZzQjr8y5g6XeQZMZuN6/ZAI1oBUWo9k82gr3kRN2c9FNv
zs7l2KHhGa/NT6jWCHG3z1d2UPVNwPE0Cf4rzES/GFRprclZ9KnwgTCx26VBkDujgWt2SSpW4wJj
j2+e7VFng9Dz0zcis2GF2WQSt/0mYZZedJVoZLk+WeS3cPpxavG9qp2c+z4VATsuUy2gabzQggJ5
1Vr7l4ZyKosQIcwl4+RWNbwejPEMb6M9j5rrRL/KiNVaD5JWuIeCpcJefHLp9F8HZ3vy7FmvpM8/
Y7o66yx6zTz2Bq2Zdm7Zb82GzvGs3Rz6a2lL/NFIGippR/XnanElHMf6spXR7hUkJMqW5dIzYXus
8lKbXSVua04iU4AGAG2e7U6G77RSffq/4AjZytqqszYBRV/If+fAXv3xQIshn1ckJTiXr4FOnCzp
E4m0NEAD7JrmwjjoOX8PqbBqrZBjgcjykDDA5vaalJvmLzklj2UIBbjHRaEfvJwQeaZcLq7R+xgQ
mG0CvRmgg5J5VMgsZFuVQh93/8smwq2FmAuF4dgOeMd0mqEEUzjK+iJrBtBrnxAZUHOGlSiQ9GBY
RyNVHJqyTvZa2Tm2YL3IY8y5c0sbCTMN6C/o3qoJJ40UrnGm6tq5lFYN7cn+reZAymDo+kWdLc6l
v6FMFEkkrrqX1JEJkZIJrdzdHI9iR9Be9BxfXaeT2SifVxFzIJr/mTk5Mlw7H1eHzVkS7EZ165Z9
eKjOza2FPpO0hJp1Hj5LJ2LUhuQXwvzbV7VL1NWIbrncmyKqZuA2ixAJIyo8J0yYBWaFodxsjbqI
PEz4+yq/siTu5yvhFwPOFcPFyI2qHOGNvMtZwyMFoHLvd+oJridnXhyo8yoiaB5t+pehMI2FwHPX
YndGTsjQXwOmgyU8CdVwDYafhJS/WmZ4vqwo2n//054pYZfqVpAy6F4Z14pL4vg7oSFBZY5gate6
AaqVU2btX9rZhzid+qRBA0Ve63Kqv7V7pXXmpKRm2j2qICDxQqGH1OFhH1HKIcFJOkLWSj2wr98F
aITpfBfPptH90jsii9qAopkIvVi7tVdYI7vKGHQaflG7aO+q8ggh2NJ4+VNeQS/BKS/MsHlPOUE0
YPuvvdQec8tIwUv+IIfA8wd9fvzejdbTh7lJT2VTjkLL0aX3BmM2lQgVH3DImECw8U31nQa79lxW
bK4q8A2UVJs97qHJ6e3/gycnGErcqKbjWgUulApL/g/JMVIM9rRN0lgHaLWp9XDwy3Xj3pG9+ref
UvShJSgTuWbMXMnh3MXa+FLfwjf/gCQmEEjYu7Ep6BVlL2AJiUBUShq4VosB5rn4SX/5OcadCvTw
f7PD766Q3XCVHV3eythYHYMV7AedIrnmmeUxYJGdo6lP4+sGuywhNfPd9C33wd6HWA2D9p2ZUZac
w6DTIWEEFUisjZdHvxVaqN95Hcz5U3HKgCMn/619itxWlS91AO7R1w1A1XcwwlqioOCFr8CBqoo8
LDCfPi7Yd1OOrc13LzyEy/0A4zsmSIfIcXg9+e8yDfNAvdwcVwuqswquLYky7Mbg/2W+ZcB8X9TB
RGBop8QjNrgrWLbX/dd5HUIZXurcIAQhZKeyF3ZbaZeShRRWOdP85jR4ylglfZMItn7LY76sSDnW
JT1luWPwaxZq8sL7T9WPyP819eSzFLMfIEDMrBLb6fiWJ+z5PnB68jjt4F6CjzQVjlScJowkbI+B
yUsjcK7JcWa7+APUAB2w37Vr8hSPtGNIZsjL9BhC713u7Kxnvfw3S3vnPDt8H7OLOE/V0dnCySWd
1DVLvxByVT/Fn4OD+KlfbMJG7vVKX8EeCMsp767hss9iaQpvDb+06c9pmAmpZvSK7dy3DNqYXMjd
jgRPtZo3wBQprSnMGkotEjm48s93ovgAVNAwAEhPZq+9fjCe5WCFqzh8VQ2W9M570X+I9t9r3chA
jTrshwoGE0s59hR0wOB3JNUYLmm4GPodEF8zH/dG2UPc7GJMQ2zX7n6dNAr4yS0Y+SRksa8s7IP9
Nm+Gmo+XMXFAuiEPGk0SDGyB8m/lhA855doASuSP/psXDIgM06quDc0q6P3GmuP3cFY43F0oSuhG
1UZ899LCueyIRJoPLmzLo9GsTCqsT1xWyUxRzKN5Er25adbuNketqah8RkSclWxNDlVEdFhbyJZR
Kvk1l2OBAqtsKy/IgzX/HWHFlNjXkPAI8mpNvFD3NvC9mhuPBv3UZ0KR1PApHe0IeQXu1f2L/ojh
wpjnEhjjXNd/mCdLVxgz3ck/iyK13B3jQIjAGogAUaJylSBJDr+llT0PL1UWeqI9/35dp3a3dy9s
2OWTd22f/sne0QvCXPBZTlj1gEGmRreJMcbl/oMAWsAdHGs3AL9pnCb1rDUk9+m5M86w1di3BfDL
UWJli33eW2ANrAdrqaXbsRGiG7zjKcyrxwTtskcL/uc1aqVEig8rXHeXuiGLMwTtzpFtDO7e4MXF
xDLiJF662+TDFnVGzuezSm4rVRisMcJWYSba9nT55EYFtzHHhcRCHJGKmQiFuvVWTRQDjeZKDuuf
NtxMHt/bpyER+BAPXMHkKdbs55+mG5vslHBfv++i70LbinSEn5v97RjKvoS3QOPlnqpSZjZLG4tN
K+BOYO5JvIKsbv9zpA5C2hK6Kwv0N6/kKwF6FWGIGyM6BeKwTm0p/MIF7Zq/Flmlo2hO4mVcETA7
Fq6jHNHFKQ9SPWov7RObTc7VwuoAi6S/n9Tv/j9Mn7nynGfAGKRO9a01EWL9391X4V6qYf1D7z+m
1eJn8ldrTdvvQYv5NVgHaQl0k0oRYA40jaHvFXshMcMiuCrnWfw/967uu4RkwuYXePAJWhdUDEFk
IrhAnxDKGo0eNPY25FQGC5Mc9haUnR7iSrIDbksHbqA3klUaQx+VI3LLAuVaLUe9wkYOC0+1XNhA
ho4iB3Egu6EIiNfhXRpVXZdxmmTwlTcmCzDKaEKefteX3KNaLuSLt4Pb4XzmlJYkYIutrkiq/gtz
Q/MbgIdf37CqnltMRJJUOeDbp2Qx8bN+Z2zWfpj8m6keSlIuZJxD64YPXVNnZCky71dHf9rPXCPE
W/4xdT7ce4wv/OwH/VP6WUoKA1xt63NNUQ5f7c0PBz/hj3kub8KJEQEXTO2kKrZcSaXkPhTA2HxN
jQBgAUrlWtq/fnB+AcBojvyrkq5H1dSdXuUknjzEjN2EdmNy5pMfqbgLuYrnbWhAiZ3eNZDrW/SV
DWPG0PVzHHhDzEdH7dkQkv4JkbTodaXUWSTZ7e1e+wKxxIUx+GpCxI8LYJYobHBOkOkk4vQpc/lO
gsvwFuCZFNAtp4zXIbaTfCAltxPiLfL0yRaOXwdOEMYWcKkJvO1vQcsi3jnSpDBE5TWecW6heLZH
jxc44GD+BKAOhTLJKaarUXTfnKC090QMFdxw8Weaet30Qz6zBdh2Ffd2Uzs1oXEmCTeTYp8knNgy
bCPeMEn5brMk4BVPpwpEhSM77cuDjyhaOw+LusLRoOgfHKAq1zyekxilW4MDf5PPVxXMiYj/VmmN
uIKUy9UQvJMRDxQAVeetMNeriRXM5YCxS+ONqG4cnxMyqhmcecxMN0U6eBaGXwv5NM7rmJiOdznh
tXYVeQejyj/WBJWBGrmFfcxUxt9Mdy8uJa+Hc4JReZdkOhLvctuYmBVOCURy93mzvjqtcyLYH5vK
87zkAeazE1HJ9HlpulTGXF6i/awOn5iYIslgNDKw5AmQfui9QOOc7RRuvkH9BMVYAEWOOF7jTku9
CmK503Q/kgy1bqiie83p95up5X2PLWPjomQvtbIwLrSsTPNMB/WzpHAzLwj/PXbVd2bldemLP1Ws
64XlGcEFimr9iyyvmC/X4V7y5B+SJo4CELBp961LHKHI4RYpvgAPQvQEzDRy0ajVE+O2PKPZHDCZ
7k6oL84bdqNRgQqvV0kkeua8n7v59esg7+dP9ZwMd2PtXPqUQK2wWsCgvbXOcUCKo3hTsIPuF2aI
aa6nxPc3iatyE0K4nsCYvvqW9O/CHjx6olC253IZIjVry8Y8By6w0YVgVF9i5rC01uqD/L/wRBr+
5wE5WBbxLvvGUaFevvL+mAHCuvZh51p4FcJo2mEmQlDU9pwH8RRzgDtQAa4H3iFdqFqeH4LfUFVR
kZx9/9wB6q88AGn4ZSyeM51uyE4xzG854N2eZYdCC2SvhEUx7ooP8mKF+bawy78apGLP/ehO9HA1
EHwdWgf/brgcqo+NGGC9ut4vA1LGpI+5ynM0m0X3WRYt7Z0aFVRBl9hA4tAZftlgr5GVarkNe5Py
/QMDf36rNr61puqblTDwXM7ZohGP1qG+Ae023RvvLD/PqGYg/OTB19EOIXKZqQzDAbgkK+eqywLp
Dro9AY89myBM37hQpqImwDWZZoL+2ooPijxoo1hJvtXH0TWxIIqorbCq/LaQ+WTneyhEa4YVpKXv
/pXYcGhOEzFAGCBz2pqCbwowKuWV+AjFbikWulv/cHTD2l+qldeoWySWCH1JEuSJQydofpy6M2rC
aN15GDCJEactqqxFp9bukzs/RgOZ9CARRsJkg0rJlx4/j3iTqUSSw80Aor+UH3B8Qn8p7533rY4i
4iqZylVKeusA3A5JLb/kExlcchId7YJgenrqw9MwEarTUcIIdiGxg0pC2Izagsxy9EH5ZjodYBia
c8DP0pETCn88L5zKhKEX7p3EBs76/4uG28y3DAfneDSg+JKj3W4u8aJyLThka0+nfdFz8GEwr5l0
H0TaAdGmFUT4bOmK+71HpJNEWixTG2/nuV/UDbkyp2KftIfOg/iS8kSC0r3Oe0vKjdsLIQKoj5wJ
pKFJfK48Q2a+g+mgCFVi/60lC6UoB1U7ddYuAKBwLUJSeRgcOH0vs9UvJSzUJHQK6n86ZjZ/5/pD
xN2BhgVB8DnYadpkdb9vDBYdPj88befCSxYys0JV2tsEJhlorDGYmYpcZPBDWDeGzjuVGXMpEoWM
nbfaKthg1IfdRThLNSPVse/Q67acnHR1fc1ooxz8fEQkyGxslm3+uoNEbg9turX+KS1gegKz4L1g
eT64FZ7WsjYLenid6mJTY0q3sZNKexaubcDjJnfzXajRDnkHicoLEcGbqLj7yLSHqZ9bOzFVx1ie
ENWrOpizLp8qQVphFX5LD1cW7UVwgy2hhMrn5rzqnZcihjL0oGP2nwx31kxwLi1DFvF970weoAUe
GQwAkFOqq8/unm72ylVxukk6W4k2KAgqOiJuAEy3uney6APM8gImMKbC1bHlqs1rMbtlrh6wiunI
23bn//SweU+mTjjWAmOaAWBsrwdKBkekpiHO3ghkQTI9ZA4mWh14vFPxEuYodi9I5xrffUxQz1hC
njSy5K2J0UFySHDTKvikvjErZzAanKKYQDbBe5f9cMSrpMa4p+ueAzqv92IkSO5/usaLj6Q4HBcX
TI2oBOikHZ+aYQT0p3SMmqzW5OG54sy5wGGep7s4OrQvpaHzmTtUf5zWzn5XFwOemb6chu7cunux
olgj5krLkDwaqYK41v4GEKf8jEN7Y6eF5WSfuzpAQymiBhWus90KxzJVpbnEwvfeP431ZV9Rq1i1
Ma0M1XwtW4OmIQoESeIFg+WANmxbeaDbBc6xhyY7AXTwN/Y3SxpnEy4NkVJl78dQ1foUWuZP+iXP
S7IjSuP4/pJv5zxP9z6u8HKYULtbayJCxTs8wOX7ik1boaw3U31W8r4BWv33vaIiZ5kOZGkQyJtt
PQy+6SPwgZi7iCoeX9mGJalWK4luSamHSZ79Etk3thM3LuQObPQQxlhtW7TgFpkKWjC2z+2QZ59Y
Xq2CuOb4bhs/QAONh79dylBzJY4yvHJxV1Pw4Wtg7HZ01U59q1aHObwQSYrcwMHPXb8f6gEt2qhG
UNcq7XE/PH1Wm6hmmpHBgnuu/VxLI93RjJAab4IDw0UW7tZ+ACyDAxp7mfs6PPdtBv78KrsfPwyb
dton/TqrsRFCe/M7WEohP5CwmT9Tc6/7lX7sc+Afq3Sn3LfWHsFUpZ1t6lFelDWxj4Tp5lbcgnia
Y4WMVFyKNFq/zxGSAJjLayNKqNf5yhEjOjyK64YKoI/8fv6VECldVXvK1yeC4qSSrTL4j62RD64r
G7ctb0h9gnkdZUp9O/uq5+vFhgSHLV/iQK8cFVaLVHl/vLd9EjaZn/Nfono7lhTu01+1BVjJ9jGc
vfMNT9DjOLvFTxn//Q5sDdkMFbFlD2nMwxt9sPwBAVSWatn6btCy66ww0mNrX22EUT4AxReyW7qP
iJUA0lnZRY7n+u8aabZ8DRIymQhTf49F1USW+Gep8XQav4IU4sIOc2Wlu9T5G6KT3ertF2P6IjMe
RqthltZjZkfGGUDcylByJN1b21kK1H2hVlKvrJ10iRGWJK+bxsLDo8H16kkKP34LqVE149V9GIRC
A0CWvuJkvyJ8TQAhpehzGsTZdFxGEIj7nayh1lry9MYguk7069+aWFP5tyOyiKXaTU9eEVL5vzNG
PAq+sFchJIVdGJds2FZbnfN94BwbeFzOVzp3YHx4n9c8qZMFqNNKbmfHMdaRokmEcKdChuqbaWka
WUDrHHHkH51smgrqHQUCvxPty8nlDc3We8MQBMQaVbmhHmVzC8zfpIUjcbQuFazHOIfdXJqShXcK
lxQIzxtzNz3of3ycvRIGP6hENrO4F/FbsL0qhj5wk1Gx+nOz+Pe01DTPewrtYUE1yEZRe8vR6sYP
EOSoujiNHSKwTFnj/WD60hHfClEX5BAHo/aL6zvv9O7mTZFhjcxyKvomc1YjJWnHbme9oUj4qBcT
3f07o8PO3eTn+CPYEiB2/jhBUnwv+0psblORkQnAjK9a8gFC23Lu0ksD6HEzjOoBqY5WaLCpUvBa
J8itE6j3hu3vstWENYIRyn25ptq8E2MfhoeFYZPp0wayAZ6qQgKP+3byVNYNl75iOInm7rBJdrse
I1/ZB8rNk0VjScqa5AuVVsJ1vPOEoLG8w2d6Kou2EhVIAJdNtzLjyxTIh4QtEidDK7Hf3IYGZSXL
+iW0wW6nCNybZ8vh+N71n+XYd8Xqcx+hBsuWKsPwR6ykObCU1vy8ABsmDAe3E2Cg/geOwBrU1m5t
9zRamQVzRQrsDpq7y1wnX3D363q/Vzf7B0PqxkHFaWPU+A7w9veIM7uUCJdraOoj+S5b87vBYpOQ
tnFBK1F3HeytZLoHrgbOqknuW6Do6dvZ6IlT4hv8ZK8a+7UaF/tAZ4RvsDHNRqmm87HyNPOjwIZo
gErKJa9aG0uv7ef5Kzh3I0YJm3KWoOLDabE1ose+n1Ay6xytK2b1mcszaMmaSLJdYPNiWzGec/el
og86DopLIhHcmOLM24/rQEami3U6kBGa0p7OsJdwiCAqGiTMXvfx4RAj1p4zXUqUWJaRBxnOBD+8
y/dxut844EycWOo9griBpEPk0Ph/6MlgLkHW2ZAQ0AEi/a/GZlh2J4W3mDW3Yn40kUrUX/BCKPLC
Dhqp/oY8dE4mYXhQHRG+PZV/jUA79EpKVhzV/Fjit/SH36D5FXII/NG2Amry7GNJ7nmyA4t/fJM+
in6atB1ns0axvGuKf8w6U3pjRZjO3LKyFzJYdEkh1bbPjVnJyUdLVkBRD+O/cGRT18VRZUBQz2wy
upDrrkJYCw4SaBOcO+VRtUpwWtYTYciTH2CiScPvZxEwdu73xMO7ObXPldYo41Ew9mjc76xXAiUE
Q2rPe8rwLGfWK9PmWBJUFVB83SfdSHzaDGK+58CZNluTdNBMh7Pw0EcvNFn9yeBrObP4ypyo5q1H
dI6mJfFMHhhMT44DM3AWg6gtjp4jRZNoexEpzPueT9NcLbAmohY5Hy5P379m4OAHJXo409j7I3yQ
rpUUssRsMAkU62f96c9DzyIIuEvAEBR9SF4RUAFTUow2BmlSBQFiRlNe+ndGaISvoEmZyt9sg79t
m6Kwl9VYokEkn3hP4izXO/oZKwGLfxs+l14/BW1AowxvS/hDhlp2K2fMavXQ4QPe87J1RwOd6P4O
5KGRURdSG+O98nMurXUjm2olHse3hQw6c1b4sqaNAh3uTyaaOdVNW3IbfztG9s0gKgetez3O9Q/q
Ob/qonDmGpTQJJV/GT/g0pDSZfTyWAmoYOwb8QhxcPluEbDwr2zWuLe5nrqIjIkknl9iG/azuWsP
8Tc2aG0+iJKFlWW0hRvIJlgm/I05shHiO4hm47i/8rZNLGkYnSKbCFWEd3zvaaQ3iximOEH3Hyae
B9uUt5uDA4iLLVtkAyQO8sf3nVFl/rjCOENCRjbhPUcQ8YoLRwWOtUJ/Wk1a2P4n93PYZE/+l6YB
6WxrVxH9zwaN2MyZSf0LEd+5QU76wh3MDaQxQHiZGDcowW3xR0i0BSfesA+q68GDvMhF0yJsXgJh
2m95CSc5ecrYlrvAgChuXmBgXmd0AVJqBKmBNVtkYNOsNe/GOxh2MjFhZuwIHoBd7IJxwTJch878
9UFZqxJ7v9ejLDgmvTqS2TVURj3Te6/n2P2jQ9DDzHD5Yohg4DWSSFQyMTu8s4uvdFravHAagZUD
AefGSUUOGy8MT1/DsTWDsFzTDQ8MkY3ygoSq1LCYh9qBI2rD2qd8g9MBZAy5HzEYh3iqHdM7E0Ve
EtQvGleVSRf+LP3ztAES0k53+FG77ryoPO3eCn5vmpEtvGG7tF3+VZ2FXxoq6Mfyu5JrQwBekCko
4cJCNPsjN9gyvziHUNd4cVxNcfHH7Q57scZru5bAPZ5nBS1V/MuossVvGFVrey42n3t9ioexOH/2
EhFFQlWtRI/wlOa9kqf4ReHDLTx1LN/oGsSjO9YrIhwuDEIprrQIfbUEy8+bu/j1/JU0F6KwKuMo
eyXiMUy5ZbNyrO73PMIlDm3kj7it8oUhhKebZpbUtv6CucXGeZfb/SQt5BgCYmlyJHI2+/4RMVO4
k4L9/PhdLsnDuYcyDZGHJunEYAfmwPPoo9QrDnTpWPjqfreQcuUpoiz3CkG0H6LIwVb6JMN3UJYu
GYrpnEXV22xDZFE4psxI1hng42tcIL51mWBMueKoFx0NDzWrUYTuD3Cu7oUFLVw21MNg6cWolKZo
QErpO+gaEq6yVDOx6Rb1RGzoos15c7VT+qhA3JHPAbTqoZRV41eUv3ac+JKajvmSGy0PD+ir4xNa
EHsrjqz0MssiFr7O2Uf/S2vtoJ2qRRinBWFLlNAOqzyV6ZXgPsrWPlrRUsYmJXh8W95BwKUn4iyS
KoAFG/YRyvfooOHQnrzd0ggRiCwwZ5Sxsm+zkSRwixgI3Z6iDv2zafr4gQH9LSiMSTKkEUqNQ8Xn
uV4AjiqVXA4kuSEpEljyXvyq7L+z1xdWkDmK/YLQBNMbmc9OOA4LuhhUiAj5iriP0S3cXE3Q94ZW
kCXpECYKpNhcCOoBVSYgcUbFFAYIdD5k2CncEw+DRvUa9X5MFRLjxWDLujIWHEw4Z+pFUvtnh5Nl
tT3gc/TNcW+bVZbZriGlaMeq6zDoJVwYmuYQd+nRucCnJFAN4Z9Rglls/v+j7V+XvB/vESXDqln3
n8yKewSr0/zVwXbtcuihQ/5oOKtUULY5Brn6rW/AgF84yU6YrPsT9eoNMmvEYQIWlMoeuIsPhKMt
m95IhCxFYGgKxJv7yX0z9LhkchKItu1/4QHgFTI0BCYbphnGVkjzXKwz+djwNe6B78YrtYb0KPn8
aG81YNdbpZKxcT9TCf6Yk6eRvO4ngV93jY00YsGCfM61Bo1r4wkIX2+JlgFxbaocUrbM+rIRdGkO
ha3ZOSolAI8lg5l0NeGkSHP/JJeaVlM5xuJlSBj5aCMRVfB74xYy3wOI1ijz98VV1F1IUxawnCFj
Y9MQ+Aa/T2jQpCLczR9ovtHLDOuMqjpCiTqh1mD/vSGtZXDfh6efzt78+XeP4YejuDecuEKKQqL5
HO/v1ho6MDdy+/c06D9K+fbdsBLDTun9vMfHXPhKRzt/n9RGm883jG+pf6kQYrbX3Jh9gDkqmVR/
88wgffk2+Xv2aAREeJy1eh1NT072kFWPTmkTo5jmqopHv/WcUPIKSg0NXzbwjiKEi5qDAL70WXZj
OHURKxnCwtmpzYNTVWagJvqG0sa2XAcCKimrKPUrRNzinQHZfTxA0b6Ir2MJbKwxU9poQ6G5LrnF
OqWjZ+svXWjxkkqsEsn4Ivns+3MKnqgQhQEk3wRY4gvxKey9QqwFdcvH6LooG4Q7UlNDxT69sk9v
y4Dv3CAyx9tFn+n1L52fB9pdAKyHjQ34ul0i4WrYsastWa6/mBQZZb/IpNwGgB8Q8wKL/VykSlKR
B1oq107LfJF5nMKhkob7oP1/c2gtfRxX7YFcgzC7RoJxyRUCJ+bhKwjSd6UvA6tlg+n9iIQtp1Xy
FzA+8kW2HBq8oSY29w6h+FhZwPBE5SmjNjoA2zXnqRUGMZc0o3gqBLyYkz+5LqqpxQi6muPTThZv
xIJgojF9O3Xzgiqhw/ML5kj1u2sds4Ci0r+X9aO1EBqqgkI2d6QmtbUaLvrC5tAAhLlNQtRZinOw
kQnfIi/lI2r+7esFTzBpu/pjmjrvk8mton4hpNIbmS9nfFWq8J32FOn9m/4A/XDXOQlSom/kCAfh
oMJA65bnq2zZpYsGNyHHBezpBfFpQlW+DM5ZZowxqoZ0FRPTvWmoDZGN1haTiwNyMsq3OGTA57an
PwcuZfkyWxLuFGv+u28OHYnCw5jdhT71ClMa83/ZSbJeL4Hjb8AHC/rgjJR2Qs1xJI4xguy42SY+
dFOUiwrLnXtPh/MnOaVsbnXBqDwGam0+mx9yJ28Qrhfzi619A4eKfQmqpY7vdQnk1Itb5sWX2Zvv
L+KJnqTTnWwAAra8DqX337AHeG2J+NIEyG6ThLx7yfPLadKofBEEtbKcqbd+/d9S/uDCfYpJmQ+l
FAlNPVhb/f/O+YLsdVz8oxAfg/kJs7QQhLcTpIfPzSdqr/OndNyd6XPBcKpCIW8G3yWLysi6JQVW
7d1N+bAe7dz4Kfc/S8RNJFMvmWfutXTQ6WNo+FzFu0gr1G1889O55rl8NXlaxjsg8pMmspz3RtMQ
7ZeOSr7PGrMGQcKHH9uaQehjgCq2uTaezX60vNotVAcuJEYAb/h0kIV2hu+s5Oh9W/zWfup+QbOW
wnOSgmtlo6Tx4rjMtQ1v+0VkY9LZqBJnMG/zuBrYt9TlKB2+EPlhAnV6L3CLpQ0JFDBOfZTIy40J
XqlNw4ck86JMDnIel8qerxNMOQeR4zj05k+3gTNwYjkNYBj9Lj6yLktqmABX8zPcjwhNvES4dkkV
zjAb0T/OmJwRRwy8c9QJv/4rqUZ16iSKN9kvmPPcTtcQ1iaia/rCDnbwUDv0kMEVGklWAgeaq3ez
v7STP1ogMgqqS/Y4Yw7mfQELDfBXXNIw/Fxb5bwDZjPl/aOoXSFdnNp7TvvmMyhvMFkkHiyzFYIF
RdOrjuNAertLeiNLcLjCgHb/ynrDvzMv9Pru1Q/Ohq7Es0x/Onb+ZcVzsBZN/BR/688+LDXsk1hc
IIIHWmaqUzkaSsWyKGjVr432ft/oRgVud+g1DBTUG3V6qXTIhcZbA3L1/edpC0EJnkcin1C2toak
oTHDtrxxTT+4u2zE9fzR+RWZF7DnpNgw9jx/imzMLWNX7VbnZusQLptVFTMQ5HQZTSWUlSJONurk
sVaOzgy+IDYeJPsbZaaA+Ciyuuk69vUnrZzpniKIx+obGAaGAaB1DBsC6xlsyRTXpU3JEU28NDY3
Kq2MdXOfJkbRenUKcd1TKEibk2WwQ1/I+izMLzka0LKsmUsNXTvpDrojJUeW7xvNt2UCXdOrRcMk
t1T/0iHzetf6crqCASxwRJyZSpw/4ArVeGQbLkPXl+D6nsWfcKdSCFtrQWNrMSgEE2YOih/yv0cP
RUqAgbLWIVm0+i9i3G3bGsMDdufykxkES1ucewZbxmCchLljFIQJwJgIBSLS9I7GZWYf8qvXeOuX
txooWKaDHSGbfIHUJPVcpqheQ0ZW9FtdPeIhIYxQv0cKpwDScV4tjKpSs5CfQjvSHMM+lC5RDU4p
KgpXfdREZVh/Prn67Dk6dJVuexdimi6qQ3jPXac0wFQ4FksTkf70nEB4eNI+GnLCig48g+rpHjdC
wPWKFgAI45dAYIUaxQdaAnNtFbQJj43y93rx02xhGLEH5zBvMWWD1T7E5ug1Ji/vl0nPvb6UkVp0
BuYAhcZnookhf1knknEb30aA5WxP77TcrgQeI7tfTUkPUt6osZ7ZT8zGPxJ4pzRt6tU8Yc2Ex0dV
I0sp6eK698HkkKImu4nskRRAgIqK8R56ZzAnAo7RKxOeMbR7uwAGCWN2DWAlXEI8bhksAuCir5SN
YvJ46teS6QmBO+iMSOKyMh9UzMkezJjKfuyKve7n9/SHzHr3MRV2Ha8YogUEnzfcBhmPqE+66EN+
3pL3O8qCA5BR4RKALXn6qUArcpbkrdtiqExDnxsFIpSCgz3ZPz4rlv7VbSxRIHKhhypgKi10cXp0
ocZc1X6Qsp/llQooBcjblJEc5xo0qHtQ9RPh1woVuun4XaUM4RZgzuL/ob7hhWFcBSbKddI/u4su
pxf4+IVlMYUPBUpztnHNK9+n4cUAEVN3IsiB+kCS0IVmjYzOVi4GJSW3+wEhzJEh6B21ESczQ5TU
jILggcV7GzweP5JVqrG7q3C2ktot/7Thyy6Xbc70ktRN1xw36482hyBLqdVvUEpHp6Jtnjd7nfBL
HwTYERseKxTZTQh55u2U5pPh5T4uSW8QvTjaPyS617Kc/LbfS/gj6DgV8r94zeOsJY21U9WbIxuV
g7/g/1fCUlM6qfuFnTSVNhA617O3uL7ic/0QVamleZEd0BAV/Tj0NsYcG++1R9byVvK/QTa+Qx9+
UtJUdlAFfoLqfnfgcqhaOoVINuYws787iBqUspyrIuO7ta+d7OxY3anj2eguGQaB/+JuOuJBoXxY
8BlErMiSM/OsTZPSuuu0I2Ddqv6qR30ptJZZ+HHsgB5d+3Qhazfjyi5lsgSkjmd4aqVrKfBm5NY9
68TYabUtI2mbmxcJXD1NBPgVwA+ZNRSgI0OADa3WzLBQOFjCaOCU+7B/3QsEhMLCnCbCR7aSmjri
9itEuqkiUH7dJD5keX8hdSMNCb1in0zTgguj5xD9uHeJO6Lkf8hPT4wk4up2jZsiKDj/SezGCwuw
ITW6nqV5GdpqXuQQBhcMoTVWIb3rAgD4nEoM6vTtXEbOAFh3vLLoAFL8+JDQMOnQPS4PlDHZH3rI
yWloixs7eTe8sRyvPAtkbhBsWKnJkqL+gBygB7RD/b01GkkBJWxeu24InPk3HmlTcEcJK/O8DniQ
HTuvIitSWK4zO0grShTMLb7GQwgxSOspXXz2PeUEyxBr9DjenDtF1CPErYMVSqQKvbPEFDmXUG1r
Z63iEDASMT3f1zohaQxX8Jj1QddmvftOK9kputikriRbu/N5FVS/f/AchCsMw48wh39oqtykfClR
Kht4V2cW9BKB0Rzgp+NNMixTcKE3TGh2Jr9cPQJ4IVtpHtYnbDDCkfZz4UXp8sEHzM7eIQWkRRD+
68aPZS9r9/DOz93IzC117pXxyPgh/9+PepFuivQ6eQKAoWRbqbmkWkEZtMpnw+C63SQ2AfhcIo0q
4qCLq9LAEgKj4nvsO5i04Yx+pjDwrF2QSMzwkJcWdy+50czKweK3oQv7Ma4tp+SU7ZdyGr7Kp7hW
xMUyRC/HzZycfq/NMWym8/3DpekMOpXqmb1n0vi8+Gthsr/aRY2HadSkrVN1O3XNStISJB5c1ffO
59y+DtQFQxu4JDHDcBVwPrFSuwWooQ+WCimLjjPh4jwNTr/KEI+d30iNxCdb1Mza59jTbR/NZcdK
RXRYLGbKCZI6agSURcSL+TNqJfB6DTLJA6Codv0GRbRiGyboIqxH5DZIxZp4hrkVIb4Jcshl+V6h
ltLTwbmwMbhWakv0vjmvCR6fNwbftHUqCs7gN/GtfAXp7mYxnoXeltDtm9D8u6htLuRx6fvh94g1
V8y7ylADIyLZPVKPAkk1vQiDswBrb2ByVVQyhRSOCBQW+hdrTP2qKWBRQK3QgFn+RqhwMEBAu74K
PzBTBCkcnpzpLuep5kISv/YR7XbXF6U/Jrv5W6y2p2ZYPlJgt5oOdpr+4W01QRpQ+d+BlhCY9b6F
tL4xJm5GjIoOCG91WbIhtJUDnC0TmPwkLSlNsjeSTWNkoFswgFrElTmOa5WD+gqSUMVlcuBPf3sL
63hEu4BxTtJKz0SGRVVD6N+jZJwqG+m0vrHJBNHt7cskv/xCEt6hlsGW6w0pnj71R09GgZfpM1tU
aHdkiM5vrNmUUAkQUwXnrBFQaQXhxBvSDKa+Scv8MabGQS9X49UNWplWhcxMa0rm+32YUCYBYYYy
/mUSu/rKMqV4clrv+5fNuCUAxQ5yqmNO+k2FGQUK8/Mh1qXZBL8krQSHASHv49wpWaO1Mtep6rnB
hQ+cRUVTTsq5JOSL5vlJSdr0q3wQoZIzH8zAkjPVwgK109nXm/Nmaymb21CF5eAtR+npNJod290V
G/xyu5leeWw8iDnRF8M2P8ja8F0HFr4ifn7i7I7+CmFoRf41NT9vw1E7DmRgia11akynWYhP19wY
nxbIcD4wy4piKrVSSy7j+d3A6IgZmbCTd/rrKWg/eHR2gkRmCy3DOvs1SPekKFHgPXnNiTvsw1c4
iuzXVBEz4c4hjnF6ANwPBzFES2XXf0+OaF+KlWdcFGVowYmdGEMuDL/NwMiAkPW3SQHQfJjPPHgL
x5btAm7T+ZgjFLNhjfKCw+cH3RWA0GB9vr3rZOK5Zwtf/NXAbqjuzOyk4Sie2Rqpa9c0LvR5V3bq
JdqJ1cbbFi8JdRKK1i0cf5jHaBI/RJz9fXTsCFfE5r6lOYbrEFLOKH7adxFRw93GvxMdE4MmbZ5h
GQvDBCflbTCi1YR4vpS/maSk40FFHy7WRsJZ3V2BRlEWLtbr70E+4K9Y3C57qLIZbhlDlJjKO9xi
uXBNLAvl1TseZ81ZQwMsA0FRweJOiA8zwaUA8BwlkgmTnztcHlQhbCsOhSvapsfN0e3imhJACpX8
7WCHw9Znwan9/Yh3lXAfSO/qbg1+nnFsnKIfZpIPkFg0v5CLoHpON0SxBfKH49jdcT5FIWTa7aqq
lwqPA8nlRO4AInFVfELhoMeBoQZG/Bj3FgRsMpcGQdIq7lRlkBqn0id2b7TJf2ACdA1PyS3NnmwD
db9MEidLRzlaBKm3wniCjkueGAThB9plEL5vWWXgLcRlHZpAtsO5xNcdlCHgzhhUIjQPaV3Fgzlr
f5QCGgaEYTtOxtOP/+KbSE2pj58Y5+3PNK/Gi2v2ccB1ChNt1K0trg43v4z5nWg1TNrdBXTU9OY9
RGo9Pr6k4nfYegUef30hDAQ2QFp7A84fVuXhYKYyMzkD49IqR/X21PY7fpuUE6errqTwww0HTWQm
4vivHXye14wWqirqbffM8vmXyEgXTw8gstgPEc2zX6r5hUaXFLM8+t8+77Ac8lAKSDfpVrFgPUkh
bKXFm4u8l0l3cFGA23YH3mR0pQTmvE3RlwlYaVjGZJhxifZMpICitwe3HaQGBci164mi+Xqixuqu
gyJs+9+HiLBqRze7Tqbx0Mlfyshg7OyPJaNg1NukcwdGH8/wXB3hVKjeRF/e1hKOHMRSSEvbUaKz
jIu7kDNqzJyQdYR1XRl/hOb0jkcs7Q+Q4WRHGnlh50c7beRAcB60+L3p+jzlWoBpzMfabW3UcmMi
qCfE6x1WujQgNGoAs2BjyiD0S8tFqvyTBzuozUcPWk3jkQURHRzrLdxByWPYI+o8IS6VufXtVQop
Gq/yC4mxCHxRYjaQDkGOHz5NNjMTZbAAfLTiomRGPOTBwf00UDkUjxXXuyQI2Qy2pbi079ETWT6K
Q1OCe/NRgBD5cl2e832iO7L/9sBM64h3Gk5E4F4ztQkYoDPkyfc72q5XnxUV2R/8F67ALOagW4w5
kVuqTCpQibDrbteK/KmNSg/8wEsUh3TFefCm60O4NsUFlxMETAPSYL7zvA6IXbv/VZslCG+7YDHw
+mA0I/vKUh5jaui1bBuedl62856Uh+n2ILOBP5vvQbhMUuB4tpiFvOLjmUCMZBUrOUbAv5KXnBkJ
JgUgOM9LMMQuGtvtWmXLfLvy/BbkRvAmGMbZCjB6wItkX+LVkwwlM+R7fGri4xMsrvun31nQ581n
5JT0/k9FW5lkJ9U7jJ74fpgu1EVhQLj3CJHrQDIRoj02CpYIO3rQaxTED7gDxzpTcwZreYHVBkKG
5OcHAHt6O+BJbNC+Ile7qoB+F2ZikwqdBbfbvRps1/v5ti45Sf4TDIlqvSR3QinnvaBOtPUjJ223
tfNKmg1831Od6ntVQO31IKB1KrgKBsmvs6q1+Kc/mmtAh0CMmweKSAbz083VB2ADyLboiieyuBJf
kiCWUdkgRzui8mpTnF8uQ7LtEe8yaiku7UkIARi34ATn8Au/rcBdG5gPhU+hA7IHwAn4gADGvUUc
EBTQ66LEqgQA792q27aDRHXQEyn4A4KqG8A4aw8woudZaZfa4uu4SmAOXdo7ISPiRFj2A4h2x58p
YalT51yngiBsoyN5SCP6XPYgYBdKQHaNArZSVpVbvdSUV6Aj3fcKLpv6/6cgKdQuFZQFgVs5g9E1
PrOEicNmsIm1V5cGXdStTUUxEngD0gMan4M7QmaFwwsCfiRgfwIs9y2/DCxkEA+mPUcPMGBPB5vP
/5xtE3vSG0O7RZqwUXgYjvuHf/eOZLY6jUAHID5f1Ib4BHQ8G2OYQ177UhgcqtspQdNM7XsFbCXw
z6g8Ouv5R2gAt+XXbzr1chmM7MelMvl10XNkf52NDOhOLxjRfZ4MQlx3dh++waTJ521d8WDjOewb
EU7nrFTqHkrgG5kRbZlovKO7neQoWOA2JGP2Ii4xSL7xwIBSV5+/sPeIySqwbQ10b9kslA8Jr/bX
RRmYpxww+/sTZcIVAc0/YFLpCLTwtvbZegK1GSFz7JYfhkJB7553zLcF5jL6c7T3bumODZ1d0CRm
9z9hRGkT4+91pqLfmVqGLEIXAkEIHwspkudjWk5GVeXzepN/ZSBoodl4SYkllC56Bkbe2BqvF6qa
E1B55LFKkKuQKK416C/3uz8O5TYsOazLNrBF7UvWoKk9Gg9BwM9sJ5NR1fD/rj4okwwQsYzSrqAT
MvfvGo5EFJz4CM2yVnc+kKRB/lpxlkVt3tcm3o0pOExYqGybejrsGUz41hVSJu0we0sGXk31yOJA
EpuR1QZwwjR3HbiE26IJLAZUz5AdPpCwm7NvmF9CoChWu31FerM+pu7UVMPc3+2DimHS2qcO48Bm
pB+2x5UDap0Rn2AkztsHrWUxccmwjw/319PhIx5BD1J7Thgw7G5EJ245+5B0oh3j2+jdVhnfK/DO
acbcRpjpdfBn1co+XZlW8vx0zPW/k0uFTv/ZTlf7cQP/4+bqD/MrnqtpgJ9vbvjVHGNo9Os0dltp
g2Qpou7aFfqmkM5pX7DprjX5bZG5Pz0Bows9XamUs3C1rWtCBHczYoLpOWBMbYXB5inqMTJMgQzM
dZ4+vbnEkNwtlfeMwdetSY2FTWR+t+yGD+miMFdnZu/f6cfnZrM4JL7fqPtTaHuIJUCUCu2r1Wtu
IV5IR1cvdnmg52IaZ6SPvmKKOsVZqLzfe+NJrK3JdYV1HrQDDQTNtq2aKxDCQ7IjK4B9190Ytt8A
PucFUTaeJlvfcyu+qiCRvDQN5OfFQw0jTn8vp07bocWNdUn9OQWsnmonP5bc895FS0lL2Ojv+k9L
l0iA/yEE0UE3t/FxopAYoHvJo5YH8BvnToBoQYPGInbsFs2J9JeV+kS5AyjALNcjirA78LfpPTTZ
hFrAEOtbpU76H1G0rifwCTxW4Splxp9hiB7K6RI23Ej3+z3eUjdTp2JVMbkwrGcKtePcvk9mYcyl
kMKZNLL3NY07NWRrqqw2av9cW5HlewgAjRwR78AW341f4QdVf+ETZhZJXDKhSwxd4XXm6VqBpbpk
86esWylNLWE6hll/gd3V5+fQDRcQjD3ALMuM3h6w1tG9j2B5g/LE/DRNtYMrMkLurHS+SEeDodNt
pmb6dsGi4qHCX0gYnOUiPHTNTmL+53rdRLRLg5ThpHlePmAde9JWTIoe/8agldVUipE432Dtq2Tl
3BP737VdcdkNG6kA4egcUIwERyGD91j6t9Z/Qp2Qk7RU0y6iljyR5GqB5lbZO+QNf+eLSqcHOj85
YA39jn61XdU9XTWPTruoi3r/r3ZYLDbllP3k6UumcsqMsR7oD4ovR+wFnDE5X514vXHOrrywqYQZ
EeY7kIXlUtISAqNziu1sCVXSk8zCScsW+F7nLmsyY+CBOjjdQTA/IZ8O6DwC5npVcxkNE2PGBp07
C4nC5xD9zUSZOLIJoXpjv1YjGqAxcKg6ca+zwDDocXnNmY+GhHZq/DLWCSmSUSRiS52w+5gZseje
1cEV2UkvwK5ahj1AV+WoGT2I4yO1qEeerI0xZlmT1E12rXxrb42JM5bXEvq5n1UJn8CA9p0FUY9k
B26b/Z3/Ac9nAtQEN+cvAP3AVyoGuImTZIFb4vkoSUu1P4D64uGZx/yplZiULu33aMLGZXJ5l+RJ
g9lEtWkWjE+FvozL7GCyBw0AKRXfXDI+ZHM2Z/j0Ey5bcLENgZe3o2aUqXvAHmBeLl3CeEfjBJ1T
o92UnX6UW8WApkqJX63EJP1Iw2o+GTxENT/Sw5QGkcB9u7FsB0m1EwZjVhDP4iQtaPxrjmiI8Xz/
TjqY2H3qzL4a1+fNHEZ1j+cgWALxZ5mq3wdlItWwHMNxA80dsJ+y+0H2aCpxoKWEMmtk6hu7Kdbu
jOasSS7v/1iY5Wm7xeJqLKSVHPoCBz+qE3+TXQZwo60Q9vsv2WTtN1ZPEsHg2svCBbBZmW8p2Tz9
LnxIxHo4Wl02qMZx44vx/gbu8tN/2Jl4zcQMycdUvl2HsDdBMMiuTgD9AQISf5A4NQo3J8L3/+FV
rtL06ddIBOV42MkgezIGHDjjB+LnI+Yf2eZmBvzaZRHpyIIe2NyUO9ftnQDSlHQL+yurqPDHU7xC
SFN6NWXQDbH3Y5OvXINKcNMVMj43zhU2VQkTsa3/ZX7gmCogl4H1PQgI5cXCDmJ966aBUGjLTE/H
caCSZ/kV8pdT1h6Rz0o39lc3x2pA4fSuDPIe6mTlnLjwSjkfROqknhB1/LezHI8D6syppzThm8cc
xOKJ4ZiOh0DdrhF4FXDlagilvozkI7UXgGAzF0qKwojSstccZXJzgvXS/K//gu9xWM/rzbL41EBW
QXI53c8lpt9GUgCLGxnUWL1GaKsEc2Y5JnrL2Y64fOTcVQY1+goypRYWIsRmL8OdDb926i0RD+/6
C8AF61jETNQS/7gKXINuhESr7B3oj3eCA3SX9tYR15nEUjLfA0HFqcAWjzRqxtVCWB6FHSYpFrqt
/S9s/9JJMEG0Zlgn1JmGMXmkBkzSxDX17j7F1dqnHny2iPH75BU5ExOag2tXdHAlR8KOcKaARdPw
pyg6imPCmqPcCPn2Rx49OOaSQD+1SyeUMAGSd72zi9CLbKB6CeEcHPuMc0H2s+nUANjkkAmSJmma
POLlIKjOKoIcURPYNB4rm/9gj6xuZwXr7LYFmTvG6GQf59hznt3QdW1uWBkJJNQLQNs0NEwUkfbN
xlPF1QWDWbo2G6AflyWBFvXwjQyIklibly2T+cYjN8CRUpYjoaxdSRGTn8P5ah7o38yVJlaUt8wq
FqSwHZ5mJRQoT51PSxXVgWiKtudOBUmVsiirGAVa685RrnePyPdXvCA/T4rD57JsjCCQxzR9JMXc
Y/MEqKsKM15rUiNRyjgTO7vqw5ATE/RKGWDuSUB5exNTqV3l86Do1/JZNxCmDNQPXam3J8fYACfM
wuAy0FxlBfMwZd6qf3fHx1Ps4NOCHoSpLuaQvOzXbi+ERaFGF4T6cfZziOT1k8+hC1qf4EAaXnPz
hi7c1fBiFMGG91bvaKVeAx6GHFPKkQorVQG3Gg4x9wMJ5VAClXgIAigsB7TW5qVS2xwUnrM4M8Z7
0T36dLpwXjSJXn2ZiAc7V5caCseOjBZL6DwhuCAPleCaUn58/o+1H2Wq5BvvWxlGfkCocssRW7RH
pPXWX/WbOc1XRGHX9cSb5BQs3U/pBsEd40Ao6X9BZAMz+0VSs0ID8CcBzakb8wM02uEbrPO0zzHk
tUfRvZqZeJ6d+mVP2fOJYVTSD9D/AAFpuedQmOfGwvaTxp/70SpcGz7/jZO1tIfYSGsYKSqoPihU
UQUpG9ZF28+qClgaqbWXf4ZaRNgmNaDqSTWth6iSughvDLZNdSiHOkZ7r+hkvY49vWhvMrrMXTWD
K5IEJHrl2O8/P8NoSP/C3qtjCp2DljeY+i0iD9ecMrSdiDgMrUaz4JoKoD4oFBdV/8In25vWyNfV
8T4Gv6OpTDhphmM4/fzoL69aZFTQ7d4tG6yiWr9sCL3AQ2UQlxOfXgq24T6/mcSCr9qotJYa4abX
p60j4TOPEIA/6JP4IZqMD5IFoAs9WxkDy6ppo5lk2MngW1KiZ497mnUS+PevEqkr1hdXpaIv66BA
iTye/8k4DDuQFHn2kR0Jrwp/ipdy/b3nt04nE4jrg+cgcclQPH5Vkayy+JeSHZ0JwCV2QdStiCnJ
gD2xWEt+lQ7gi997qeBcoXQxtslE1qK9apRGlhWO7lQnC5SjVeU2lyBm0oVvFCa5hfa3Uc2C9chW
Bqk70Ry4y6guSLXlxSv3eudPvQObYocX4nEAdI22z2rMmzjIoG9rr64n0ZEvU8QoxmP+g4RefyDA
D930ch/5QDjSvPUfBhV8+kNFQZRKfm3FhmW0065o56lXuCbZAdwGSAxTXHBICvdWa4iQR0smKQk1
eEw7iMtu/e7QLwedP4bF2sDFmHEecaNuCcaSO+0EFReij08lNvG+OfV4XMdgmkoi7HVyvg7MRaLU
mYGn1w8y/6cwSBXmdFd/DPmSa3EjZUz+JxjjuZr6z7wmPCTFgVDtxZfrm56/i+skFZXa2xifotcY
zVlKpYZ5sds4w+7s7dMzAGEyug2Bn+GAK1amuShlEtO5pAa82qzR4fxeafuM4EM2i40iYZNaRRSg
MLByTVi68ZBecrzMF8ZL3udt7721XUA6WuU3vGCOkFI5CEp57h6SrRlID2ywVyfhizrSHwtuSMBW
kubYGI0wJaxxVWO86HJ3uFjADrI1nAfTIclZJpikcAExp6DYaWwyzAlzWX1+mQaC8S6HYbMSKMG7
icyKkTaCf3hjldvGtlDUyIyw3LIX9XpiaExOhIAj8j2U5b9LyFWtKOkco4daMOmovpRUG/LECb8A
PBQ9uIjwMPysGS9Sxthw+7BTHsg0GYKF38359w9iLd8dmzMJ3OuHEs9neTsqHegLSrMasPQUmt/J
DKw0B+R1jFCuB/CTOemyvuKoQmrItlbQGVf6KzInETCUExdufhbDhWnQVihp92f0oKHkqGNLFQQw
sTgSTFapvPmq8Hy9Y6UDN/nMJlDBq4YuUoEGXgXJSGUS6dEt0gK9d0CZbdna7aV8BWldTGpvAbMa
Lm2y7dn9N6vUEyH7gSEpC0fk+O/GJci8GldvKUmrstpQ4+vM1Z4F9bxo5wck9tgB+lP9SsjajCc3
57k5JwnkBq759DRYsAgR/5cbPgGxlgA7XHS1DbkeqwfFcaKRKf4Oau15PO5zSjJvMjLO3eFxJZmv
JMdQtufVo/7ix6K9WohyUlOCHGP4y2sv2GgJ0khAdakdqxKqUHTOQyShe3E4IZYvQNjHnelRFOa1
c4HrKk0z1gZ2z6+mZP+rXjX2JV72j11RlE/k4hqPbfMvZHbCv6Kx01MtI9p4C+0+PHNokL4zSJSN
sZTIq3yuC63N2kzxJUYN6xn9yNGc/Lnhq/S6Lna1wZUryY93mRNVr/ieYmoHWebm2LzO60BFk+OT
eKqweWfGs33OG4BwhxtgvftjllAFF/7Jg7mblRAcNuh6fc5/K+yKNrtQFPKOicMRFIfholyYFp0G
S7ZEAqFncrfXPKJv3JgGK314eBa5WyWisvbRV8Z7LAWylPJV0Xv3qRAnh6308vW6EnsT5MV7dRo7
4nyRFx3ybj4dwOkuAu85+suaI19GcALIhxTmGUsW3aJSmvvMnZZ3TjepyOi1IP1KKy/86SyhLyHU
RyGJjnOoyZQLPZQOfj64d32aekCHNpX8tRz01q3pPvEn3GsGpMAUXL4kxQh1PzRQhALfEUYv7Zbq
hRZvNP3gQIFNBqAqaJExBtZCVBgoRZmo/wQJYuTVb6ReRT+dTcqjUyHUU56bjpCHflCD16TSwkh6
GwndBa6ZvXnQ4VGfgjqcffgeS5h2KMmkXzGphtcKS03L/W0H3yLCDQk3FDCLDGPhKz7pFj0PA4Vn
AcsASaMdhwaRoA0fqsbmnM+j+BUQZ5Vp/O1IdIhTBmVO2kHRmyV2QkOyVNMUwSMUMGYrrSjTnloW
/XCYire72dGewGlKaYgN7Y5/QYUlKOCEl+Wv1QOjn3SymDJkQwdXxG/Qb1SFQ13gNNA5QeXydBkK
dfDTLdtM3oeYgOOK6NtZElZOb3NWY/e9ugO6rdZyAAFNIWvqsIRHhy0OEEE9XRvpaKMTZegGuJ+z
91xqC0WTS7FkKi7cl6hrBwZpbSj8T6jmCWCV0dFDHq7FX4DYs9tfgLBR27tPsDM7oOn1hfInjwtp
53F/BxjbBvPy6vTolDTk/HlNtZPBCUCkY7HMa69bElsjtf2rWHRtqTMXWVzaIoBoZy1mAymYXn1e
nPDsbsWxkRmc9xOMudcrpxtctWMPUcw3wvw0s+P59KnKm6lcAkp6bm4Dcnti4vgv+RWD6RItHqsu
mBmxeJ7YnzVBYdNtkOK+5+a+60L/nymQBv3HMCPAM2UdM/U2VoO3JuWQm+f/yt/QPFucaCfIDibx
l9K97vLpdqm1elNCijowWXm4OfpVhP3s0jp6ZD3HJoxHUm9dudFDcNYzJ9nW5G3lx8u5ZAhR/1vx
59kPilBh1xutUgcuTejHH0ShCtJ4DByJ+3dDDKhIqctXanbED84pMFZlj/qt6OxdO7gcdYh6kAQE
z9MQxR6u4yGzihzA6W2VDMwTPdTE3vqroTuD5jpdFH6ru3nuCKi1PWIAX/h6RAFe+Viz6Sepc/o0
RcRDeIpmymNeAkkt17H9KwzSroy96ntO21y21iXzmX9O9ufDMvvUJBfxMUVAJBq07bU4z07tj9a6
vvgLYmwvHTWKbF5/WLltuCQlW6EQ1a81I5TkJflAGCyrBTImZT4uh9Y3pUK2Q58e0CckT8hU3SA1
TOPKCkSNSpQU2vduCvDO+LIzx0CU2QCCk80moq1N9XM8EQ53dMJ836F+uzlIp77JbL7/rh4dsbz1
+w2FreTZfqaF4st+Jy3HcsC9vUucLn9U9/YiGbn3M7F/BzSva+RyAbFr6HlOCVWBFOe4b8zyx0Gk
Ic79bN9mv+hUPaX3kKrUHkKdEwdY7r+kfI2E0T8Z/3be3opVzWT9ZzSsj7E8qQDlTlbqTQk9H7LV
qADtx+iJK2Csz57FSWDQNQqCMXnrUG/WTPST2qmNlEG1P8vhTGjV5T61PIn0B3Qw62ZLGR7HnNUp
ALmEElML3l7I/AyUEIJwFSUHySpJdgHrb/OlvdmOx57gFq5v1v7E8FtF5MSrbxOrT5uYjdNOCxjl
Mh4NJmMnPKTocv2H+oHF0DqpA7RSrrve8umqR91EvWpbY1IT1ocxmvDKHE0liYz16ECOb1zZx0jE
zvNv7LouN8hpnHP9otZ2TxFUwvw6QpWuE8Pi9KQpz0Oxa/Wb98sKMc+cNroJpW5yR1SWFV6DO4iE
Yp/H5kTogdHmon0Dp/Hxj19wbeDIEuS4vO3K28sNaAFRK8BPH+cicMntVBxxAEc0yG6wU0GZs2ul
LwPqtK4nRzIaJeoacKY+xMc9rbWiwBJ8qE8k241PvQZsnhkzwHnIoLjW7xVjCqmOyQlvih4/9DHN
ahc1/WetxIc7GXsOB/vQnK5j97S9+V1opulosumAucqJpMkLEZ4OSGUzoTaNKxe1HewnNoHruyu3
whT5oafuGFLWp/Xb3mnNu3QoaIbdzEtbkXsTUZ1RH7Vc1N5xDYVF/ArHFp8RMRx7C7wEQGYvFZLw
LpC6/vrsszf+ji/FTpv2PUZj9nLLsuXvDbLQt4vQI0qDJoeOEyqUmYwLR80HYUszfue2pUP2CmQu
AZ0DCw6rvttb/b/Wl4JL/g5yZ7m14vwOuStj6uAB2r3l+HEUrjuk7MIK6JWRhX2O8/dEKejCa/c8
n21jfZ8asSx3kqOSAivde7YApXzrWCuV4VWEa1YeKNozBo77BIVcXFUjDa4N2/F29PwN3xCEYWu/
HcJfMVhmTlqA4MQc/0t3b69nCovDtjDjpKW1AwbNYnXwdnnCKAqFnR/FNEgzXw/GnVV5EsuBSh7c
Syndeenrb2CVRoKWFiRtJ+glSRA0elrJLV9mBC2Hk/r+v1LQCAKdnUdhzD/nmNX2J/3t1qxBmudb
6qs00kYK5JH/Lc4TUHzIXlsgVBQpzbKZwfsX86SnhRvxzG+Q1CgIcdTgxtV1hUbuGZn13CQW0c5y
3foql2jcWzOMh5DPdLzauchWlTeiqrHUTND5CErWGvdNih5RvH9hl/5hMwfloKCk5T/r9605+OMn
O1GuX+aS5Okt9XjMetMu8Kw2RAbqEBpJOw3n1RceHJlVY3jCEKQ5aCnEUG2A+jKD+GGIajqQGNwk
A9vQdDzClV8dePvqh+4OdeHyMN9mZmHxHfvEnxqltE4Fcz91iUlpnqsKpg+tHfmGJzVFH1Gq9jG8
RN31SUFNp6ov2aU6bnLQYcaL/rghQFVjpIOEinyKB492JvApT5yKxZ6IBoYzRfoq2/izbl7PnzJK
E7E1U1BhKkqAOg2pB+l0rdsdGjdMwFR/q84KTooF7zJgndaiXZxh3OH9GLVeQ/CFHL4euVq/942U
p2JtvR3lPkadA6YaX0mr/cGc5SkKLLYNUximnV8LGLcMJ0xRVAehYTlBmK7RUP94DQd7ZoJkK/8O
uSrDZ6MTulJ5PZA1ObnCElMHOakl27LEGo8SChM7YjNewyy1i34pgmr4IcEpWhk8qVNpZK6FaGgS
sddnGjZB1QHaFgdf44KtZq7o3I0vhw5K7bqLv5bpoJySCwHw+uHkV2pKNzCjU6gIg5NOrjvNO2+6
wTNioIgW6kg6wqqkCo7p49DFH+cw3SyjSemr+pC73cKPdY6c5zBmVv+qfCkbfycoSmQ+y7PeAmuF
+u5U3UmCp7TJAls/E6SUYBh3yadOYfHffesk7C26MJr5GCJEXzm+nW9ran+7ZvHF0JrgrlxTIy8d
BAI7WL0pnjFi/fUc6kpPtHCZCn/9zVC+XgQ0kNep8aNmGKLjaMKJiaZqMw5L5ISMQr2gpW5XZ3a8
rQgztHu+nPQv9TfLFbJCRM60kZ4hCRTw5ZkTFcZ62NDXA8Asn9QV7nV3VibUHn6MkBd/qxVdCDvs
amXavwZsY49I5yc0/p8zB1upRzjiyrbUBdQ11clewXSPvFa5hy6fmwWcwgTS7P9zecfI+JpBsQGU
Ks2tU2oRqETmP0PJqtno4H0bNXb0/64hHZms3/MmvY/Tug1ONZSIsfEQzSFrvDEvN4FiD8ipPNeP
PNh+HRslxWcuFkejd9Gu7tQpt5Atxw7zmSXYgG6EtxD/3fdcc63JN3T3/whWY3LNU8LpYQLXP8IX
Not9qFshHUGcPx86D4HWxUC+jgjBhpvn8u6QleStgBcQpjHIgXjGNgQMWBNhpA5bSWJuRNjAbayq
Qk5aUo6/dNGYfid8Q4Rp/9VOyGctuJKN5Y8U18as0QN67ZshYVSL/QRrLsx+cruna6dVxqPj/eCv
dp63pbU3Sm/qlf0WmcwnFFpZbYv6JIM5BYEX6QNQV9vJwDa/mroxNSUcuGeqjijBy+4G2xBReDBd
n4a26LmswPLLeloFief8+OlTs8tA/FX/TYsQJ2vwb7nYmVZWNHWxZtMZiwy3j9iOqrZViL8Qev4z
xHzvD2WNBxdzL+2ewfMaxULk+MiL+pjRXey3AMbryFs+XXftbgPv9GyofolDwkmHip1VlLwbNoU4
ToXivaZcndPbTc2OqTn5L8LJ24fhZeIFMsRNu1KjeY8/DEOExr2f3F11BbBe7NTM8cFynarViNAn
GHszGpvpI1QjKagq+SXu9/kkZhZhSS6Wrv9U2+pT0rlhs8zmh+7+TVzbezeTDBIxPi7u+U1y4IVb
1C+NVh28PukN/AcTyUQrOxS9pU85sXJQp8QaS5gfY60ZyltGSLP+nC5fR/j4vtfJtLp62I7KCE7h
E58z3HPD/sacFkzZkSKI+a1aYvgBBYKK5AxZ3YDkfpDz53L365G+zQICLXRBWFSWq+wpNOXiqaJB
h2Jwnzjx71GjmFgNtDhOcVQ0kPUtB6yImjeQhbH9zmXUL9+SbB7rarBNqBg1no/M2S3MUQrBi1xl
RX4GxcOjKN7otrNzpU9D1QnxkxgST/P2BGLcLqZz5r4iRjzpieoULd3h4VSR8v1H8CVzHIzXZSlO
ssbZy23HoyDcLtBPQw8hV1x6gnh9DWbMSKF4T9NFfSTFPbrAjfLbC1NLrqIhHmFX017EpIg0jP4y
Sr0xk6tjuVLB14sw/x/hJjq28WXxGzMCeeRiGD7SW+G5dGLTXMWlXyg1YMFDfbU52ut33YYXIBSA
0IjN9uLOLntri/zNxdmXFunwXid2RRFLyOGEK9JAyNAzXKlbzab5elLzOX6sLqRi0Xh560cib4u0
XNzsHACqFfmOhmNwV+Ow0Fio20AqFEVzko4oyIU38/dPMm0NFEG0Q4bnzuLfsOvlvQBaziBQOqxF
9NIfTcXGci3v09L/+MJzBsZSrAlfjOnLWaioJk41JZXNxrtebjs6VgWBfIf+Zx6507tbIdiCRXlT
TULA06qlxh9LUVxc39K7MbzPLiIyrOpbEpajDtTOKvUbN/v/6QyiT/4cIVU3mlHH43BGx032cxYt
IWbDClT2hka1LD2wHs+xgMJfVQPtUSpmhGtzqs+1Kk9n+Fxs2eHI7CSZIQxBcEw+RiFRsAxet9yU
EZ9qZOzBMtJnDhmZs6SmX4PnwML41k4Metdi36HKKgiUMjUfrAzYZQZJmq+8AcdlZwTm2dAc1Vuc
igUMiRCnXbXEEhj/CApAV8DtOCmhlQsmfDkjO0qNAzSerykka5hAFcWAH+6P/PSxJu1xfxav9L9b
1XQgQZhWhbK1/kj+LBSR1E7/M2oVWYsIoTxjjRBlNGI+nmizQ/OcgRmBabjnq6qSYp/skjd3RRId
QMZhfaHcLsM5x0zNVHijUkXUSbhDC/HxHwSNmsg+EaeRABhqS8m2NgU6atsd5ADF2Gl2M051QmYj
EirJstNkBsUTWl9QzTdI/CTIHa9SCHYJxt6zVgkhSIdA9hMX/ZRYoqJcqRQS3QkhfThnE9U2pLq/
QFbSSKggEvxs4v3ir+zT+ht8b0TiDG6Y24yJHYxywvJXf4BKInEsUVcmTWj5OukkM9W3OtZBLB4E
izcRWVdZ62lXUlUd9WtOaf7jR0xXOS6In5TTTAasGLXjGNwDcrxqHezriYBTcokWT0dUkQmbA5l/
kmPZHLUQajOKCaDUHOba1tF1ocyPTJN7YGS8Ny0wCPxCaDOS9QiZ0u2uhcSBUoCKyOg0xvA8/FMc
sb7HH4ihIpc8WUoAUgVnHax6f5YV9twcPLV0fCkAB0r+o80TNDTesmIJNid6Y2AkdX9rEJxjZ2AI
/jk84Xa5qPMYYhWTFIoLTE9KHehdUeiMzrJzDf9Ypqs0o4ywq2417G+pP5wKPabeyCX7wi5mGfDT
/V9NyW6HbVxdxXY4hCAM5PGLrUZvMQDDZzXlQmzWR87Leeqd8m3dKOapIB1Y9eeMGTZd+amnmve3
Zlt9Yz7DtMcXiicx2TUjfCs7GzBwfrLbB07KeUKyWz76VoI0YW2/wwzmByIdcLru2ey1NEPSIoVh
HCm7sb7E5X47INMhN1uWuSMyuCwqkxo5G/Fe8mPnn/LE74udI2fEHZecwfifb6SbS8vzN8O7CU5/
4/X6CDL/9bpni/+39arPOp5EZZvQ+wBXv/MTtJYau+RinWazrId38xfpa4kvtEFKhQNkf/M4e2lO
vNFgDSd9NkOGIswUalU7gmlWK7IbZD499fXdu/sfWsqIz617yLXHO2jY+OdRc+KxIP8ho1AQrmsP
6JXmt9K94HSV6RuM9Tdeb+EG8IHAwnCAvUdkpV7cSsiNkqnEC9HkwPnCpEukojoUefIW05XpoEnD
BJwxNvhyeZCK06MjzMtun2i+KrV9cVXOnp4REANN3anNNKJKCScoVbEfY9iQOXyIMKwYLC9RpOcI
CKhb22sfAyf1AkvGx3iztsdjczN4cQMfmbpKMWhgZI1U7qBoFN1qITyA21gA/7h8MMAQlqnFhEZy
MzaZlsNiJ21bCJE22Rs2ZQy8xzF5wnVdZow96IYbkBaO1ITBmdx1ulwYvlg6KsmvPq11wIiWxJsf
B8WDuhlnKCsN/aB1jJB4JWJRl8TOoLHWZtTtvVR7ghciqcUONH40rUDfq2eDo6YfrDJZnOmWkw/6
Co2BGCXvfChWOHI+e1PC8NMJljCsRSLNXl6+khjnZPF8AQRxuzAWd18+JbphMtV2kPQ7QK1pOtHD
E6xyLo5ZDfaL0NDQTHVB145iSzDh0g+O5CJ7lyXBEPEMOKyuLjyOhUorTdlHtAvXZ0QXIW8w+jN/
XDb3PalNkJFsTedMusoj5ikwt24aP+dC4pMq+GgCZMQM9jf4+hOk6EOkkZHZDLLGD6Y6k8fS7BG4
bhL5Xi2qpdpeKZaeQK9i0rGIPt4+PxAxbWzJJEeWIJctmgJD5QtpfeEGl4QK1XYkx0LjE6BzlOvd
EeQDyXyPDsnzxko0lkYc6owFPbyBwtinmfgHg9e1iKp/J3+AJ6xR5ggOE3DpGq0bkI2NcF4lDdzg
mo7323iC85zlUwf1jiO772V/+ayhzoEax9YXD1z9fs3alDbnCHsyfqTmvBNqdIxuhfzlN/y8F7Dd
kohblEavq1tONTQ+xTcuCjzaZUWFxk4iDE2Ek4UTmGFFR1BsL15+eHGGWuJBU8UbLEil6zovG1Fe
0Zw+QSxFN58WFjreEONBNsP+tUHAF3XzDLgXMr3y1vISQFENrZU8KWl2xxqJL0D74kVtgT6ap+ni
/ErUFqwt6KaihHb9RgpiEd2omGzIQxkOAODLOBVbSN4wc2cVZXe3p6qpHpdxAZta7bQmb/OqyzWM
ZLtpyZfMY1mK5QWEr0atjDlpXNYsuMCi534+Ldf9/Jf9L+cAhLbWexhA9lcC6ncLIyPSRfswFCRn
0xQKKcLLwDVblBYR60FVCfFiBHTI8c1I6ev4Q1etgRapaD942yjtRPXtLlbAcA1cIeR6M+MWyEgb
5akZyIGzmdpkh/K7nUM76zfsvnZWS5SOxJth//e2/ji8kKlUawQ+WFrNJe2x4r5UzqX8Xq5hYEd8
gu9ySua02dg1bOXOdcQwIAbW1YaUhf24E2rydZnLS94AYZKFOvM4k+kRQRMY0SfOlXapB2sam0Pv
Lm93IBWueI6WCn6a48nX67eSFZ4yfEFLfVixjCP13Wj2+uRpBI/q/N0sIodB8T6b63wF8Oa3hcc+
pg20TnWoMtIcjk+UcIo9s85DwPOJyCRWTM34VcMPhSLtA79mxtgRZXjcb6GOXP0SM3d9KOtvHB4L
c4DIfGdXpjLtSxNMpmt+9Yj66/WFvTbAckCcD/NNgArD/5yB66U3BvC3d8asojfh+eDYkI7B4S6N
UClHjinud60Lq4bkJd1HEmcFAxvMmjIZf6tGTfV7rADQixcsqM9eOtIy3oXogIVXzuaaor1EEi/N
U2UzSGPM2LrT20J5p42wo8YB+rlM7XePJyFIh2aptvBnFwb8cy7D14YGSVPS27wu4kZzxW9pWi62
SdAqXTdIptqECrMqTM/3Z6tUSz5Nmupz556s+9MSicLemFHU1ZHEcBrQBAi8eCNRZ3yRJMRaj6BJ
EctUE1a7tqcvY6uBCezcQn1KzRxtmc447KUV74YxMA0ya36FbPnRj7QWrTb22k2RdtyZ8OVy6rgM
MWzNQQgJGfYyuJ94HgJiWJcxWZ0172EzPM2gQAQ4zlXndPVg8HR0iXCiFYECXG4RGKZsyxBnuoXP
7IkDXs24FhrFLYVS95fxXDPXcll19G9RTr6G0xb7s39SfszOQaMALfUJbaokkMoC2+m9RvyCMnds
41tN0yNMKjZwLm/D2uy9DeNNe6mOfcw90G0zngLjzINN0iL0oaR7jLlwvVtVL8CHWNhqEEn4GRMY
BSjEBBAMQjKv+JPSsxz20qI1l4CSOa4p29GybPRxFHeeqeIrBOzhKf4tcpb8fQGAhSEeYUe4iyrg
vJh6VxqTh86EPM8fhs5hD2uTQj0HrYWdTI3aqFaltKNOpH+NbBiduj/O9m/3A9m2Q1DwEqp8A0O5
Rd5a4J9vyUIf6f1hrA6uO5UcWxIIZSdHZ5jd6isUOPPiDUVyN3aYaYCce+KhLnkdhQYBZUD7B7l8
8EoRxE8bl3OOBlyXuW4EKus1D0gbySAmPfhpwEMLmrasAZoDR8vv69qxl0Fp89vE2rktr5OJbEaz
Vl1HV1SAq3qwhB40pkqHTGdCDDF4ZITaXIXg2S4pdCELaPfg8PLejH1uRSzyIwpzzQhEZe5MKQKd
f2buscyXZGfgn3IbAz/WHIh8YBRHQKn1isolzqnKsML8Yvq2NCbs00VlTSXUr1NnZ7MwbVgMpCGy
5QLg5q3/mOV0M185O2hvOoI6YfuPvYpLhFgNZNvZfPvM+5N/m5BcXzXQZJh91djgrBrh5vTDySvI
L4PXnF81KU+MOuBXCd/vb9lWwpFoUtLdwqp1Z4z/BW24ar5NECOlp7HW9qwbXTpYnnFAHFakI2qc
I+EyMmNKChH1dMXYVbI2o31qPDkf+kgoVahN1gOyj8RrTjo3pTfbKy4fLqmVojLIwvJtljP1rh2B
sT8m2vW32647acy/jii1z3NaehW0ooOzoB+wy9CefM4sxyfoNbIuIET2l29cC/mFKW0BVjN94YD1
vzl1jE/AOvRl3+sYqVpZvvSnTjw0HUAGepW7aFPnOvt7QXsKweavmtoUJtErw1P8p4W3TFhYI26u
140Y4sHcfRsXkETUNFrggELhMGzFkHAjZ6XpRtNv3vPP8sCFzwKKRvxg4OgcyJ19EMH//TIfxaj+
0CMCFmy3cIShvIUrUv2uH8ydbhMwTBQg0da1ystFh3acY3g0kCyN8B2aRhwVCv9DHtTbBepg7NKu
s81xQeHzAzDnPFn9V1jeHCHSoHZ7JClv+G9AO3Jzuyo5QcMepBXcTBfD5KiD0mpDqUfOCmeeawix
1JkfLTVEb+pxOiJXl2P3wcbPk1ffMDBx0IkbN022HHvRYB4WOlagy6V+AubMd0+t6dcj2Uxth/k3
Ewx0+hhEDvhSK1PlVlqjgMmzZM33jv26QYDv+4C4o+hQAbBWoFXMaY0P+qC+BrqURBhfFMTj1yPi
4T1aXqp5YcOBJ9SYoeISTOjFq1HtbzewHYRwtS98GzBagJLp/nGXEEyE34UQpQX3L/6Mzx8FKCR3
xXA91UAtMJarUqjWJGsdsjJp5E5aYyYgmVCz9ESLv5Np7SlLxBNKv/0chKdFzbvNPjpqMofkJovD
mRiUgAfjrsWacBM4O5l6LMy8KT6KXhzWCmAc5xuveuGY4RBnt4tHijv3HUKpvSq/Ev7m+KcqZYyx
7F0QkfL/xGBFkvjClDQ9YUMW8cuQ94lMXgyrQbuld1r+1c4WyutpqSGwATy4e3RTnDWQOktmYG6V
IKUrZUZHosxiUCkiCru3mbiKNV6mimMp9bUdP08MKFMYIDYAkLiYY7LdnMfZwqtpOHWbO63HizDr
+5Vftupd9Lhk/H5z8p8AFaLahLJwqzjtAqSyuJLBAIUxL/+hm6y8IJWVr6MPo+Yz66HHQ1t5ouoQ
XfV1fehXdDK5cG8BgZffviqkYHqiB3bNxjMn5kekKoq9t3XUQQf4PpjapBAjXfAiy5qwSyxuLDhL
XGDqxmwyQNen3INsC5sf3QURqzPefbuU0Gt+/lOTeJBedvPcs4VVgTdou2P7XS4TKWsKDppfRp68
pgxOxKRaNnbPfzT1hwhEjSRHBCZ4k88LCuLi8w36WQk16qA1pk01Ze5Cw84fkN51BTx/nbbx0tCq
t3jxFzwuRcy8vNSYQuG6KTZkWvQlC+mq56alSI6Ee7lTPWbD8R9kC75HMQBbrioNDg93gaLcNNeU
ADPmbyaROQ0H2YjjaQ+ppPZ3jhcmJzFbhrp5yQjBjsNFdprx//Z/jyyE6Mx73+4i+nBsoQx+ykkl
pPUucUMIRdCz2Wdz8LTQQXCVMcImFPj1m6GxAqY8v+faaE+xt5bgQDDsSCH8fx2o2Xr0gJ2eCIZm
pb6R+XFZVdwPvZioJbLsASLNM7mXdIqP5VFlWX+Ez5OHQssnTF4fcBZ4+eZizVuV0nDiU6w92xTE
UO6OakBgVXlNJDMRHsMsaMbjqRi4qy7X76HjgQ3DBQRyQ6NWK96qeAh2yXNT3W5uA/+wNrgALPrR
8bzwDaAkW6lysKG30OccRmHULYv1eUn4LmZAeRq46Uet0aGg/nn5RZhhr7tNLahHqcxwNW7Yw5Ic
8PeQEWGBJNGM1b3i//o1sHKwxJcusvLIjijYLfxIyHnF6AXyWPTFYrei/1hXrSPQhgnHo5HRzN0T
wMf3Z/BwikvDdS+31mv/wOuThzOry4njYgxzT0jp2UNz3zehMLFxuQgCQga6areMXJPkn27pyCg+
+2O5xVBZcrmiZgrf9lAaeGBz+f6KZZZysmJO6zZLfLBNHGZUSzsYSaQC0w9jW4yy5AkU+2vm8PGp
GWsSG6kamzasRmfR4n1xxt1ExJFut4P++ovIaDsBmluJfaHmN+/Umt7quzcbPr0vB9A0qZm1S+cN
/4AJTLL4SDUPoSkHgqTN5II8pzv1j892Oh0DGZ/vwKjobfh/nX4UazaEWW/CTCCvvEcZ/jrx9rbJ
sdEjX5ciCYhYMfRHejmbCkVSh2nDAfGyjG3lRwUMSnQNFA/x5nqtcu+NNu3gjt+b0wF/4McA4Ef1
aJNucWdVWIRECxXMynaUBJ/RalbrQ/P+x+eOihDnGaO+Z/xdSSK5v+54eD21R0zjZ8ayXfh/LUiQ
QKqjnrvS4/ZUJvZuNW7Ks5WNEBe5pSlHZEF0sh+AxNV2KYIlxjwfKFcPN4VIACAPVPH7WH1L7uX0
e5G/6yrnZ0a/+rrXNE5yX0ExEFdvz60aY6Ur3afglfx87fzplN5/2g7N2TqUkF+wzIe5lyqQXwYY
xmc04mxswEUBO4Z0Mv/c9aYTp7hKblJI5ZmMKUHyn1/UaXn+MlZcexIGSkntkSB3OsMFmq1Q4SWT
SFqpPkA8g7FZEcYOHYfZ2QzRY7sOGMMFZptjYCavKyVr/18J1uxHSMrS7AobXNwLi1liKCUf0iNy
lcwskY1U+okpXvCUMUh2R9gsOtCCZF8XAqFR/NGvvpJr396EiuBb71NCusoqwwALVhOjsScga/Jj
Fd/iG4255cifX3xltVVJhPtc5M0wKSQbdWLNZLtVDjQjypvPPGJleDe856k4RESjduAfoHpc4bq2
ndAVLeKb2dawTmtKwV6WDd461mFgLvQGlqgp/fnWPiE9DKqBq+2ZUl9++lNtPK9b3jNvMcmaxGNs
YntxkXpWAYIIKhnDoKjBInlKVcPvMjaAnoyYfXf3K0X6WwFHvxuGyHfSmFFI07p/E97w+1vF4EcO
Jc0drw5YwEv68sIotthwsH9LOxuwdDp3EfZIhytbIg1mUdNeErxsLEvMA1OM7QN2kMayoNs89qvJ
wrhCmvgG7/LYgPZTVLzrGYUWIw0JyoyIQnRHXYZanB10+lPvC8wu+FinWOzKZNlLICiua76TTyos
11leXSgjveM2Hp7cuHNGnbrToIaCD+pu6K2UkBfhkyJa51orIKtA8Hijuv0hvw+Znvu4CdCjMigC
bIih23vLbNU8bH82bnRW48/P0CGGzQZLF6f+RXWr3klpGkWRi7bxBjDrsHfG9+0XTUE09rKMGPYg
namkdOnw48LWjzKyqvFYqZ9OPLnrY77IfClPeLCbut0lxM30JvvRNwKC185XfyFgMbUibXKtNQ6F
YbVme7yahRslDro7hm6t3Gtg1lcQbr6KAVElAmwbwPUassPbygDYV3wH7Y8i8aV7wEsXjxOLdZIA
ELkOwsRIH1fRowoaeydnjfEJMXHHufnc/rRiDmxVwf+CB3/ydsUVMt8T1k9dznMUbTyK3P5oSbs/
ruQM90zdbprazlIvo6CdOt8c2srIZ9LxyKNoIdSDxHXpcFalrbZEOJ3BjyPG6GqnYrSDRzeCNTY4
Suy74+6Cl24rY8Zfdb0Q25+fs9zEFUuEDSKatcIbrDUOWDTA8U+4gnpe2aHWoEocX9nWW09kTXqY
/uLiXEIIfOYBCy23R9H1IKQImlklVKyJTIrp+saerfQK5kku9iomPhrmRxg7lveaK59lwyWX5Ll3
eVvzii9Qa5BxvQ56AKmCHERvoLp7e3+kULm97Qj9hxZb+r5tXWcp4T3nIh655IJOh7Ao9ji2M03I
VwtLBmqkRstFappGv+JwWG6LTFhe2+WPMYnYue9RENWhWZw6ltt0t5kG+hNPRTP9X3VBU24Ej4BP
a3Vbc89asTEU+CDKt7Gii1XheMGgV5i5lo+iD1PBv4ihgGdPQ5TlelbHmsl5UOsJ38xndNkZFFei
w9rGAUjUe+5evAFkKwMNPqMSCoeo0GQqZQ9ezGxxHtJ4xu4Enro3n7dqjDFsfDAwVW+UUmETQDvR
lL10V26IfaorJuRYohwWTMcrJdZmR2Of/ES4jtfx/i4NVo24HFuNmIhVTFDkqYcPBpS1YO4XcMVi
BVe7E7tNrchZdjLbg8E9drc00ntnYplE199HEYuLMqoC4DB8no9xGPIG6of+C6pKu7X+sXSAr8d6
kiCCxVGVkhGkqHDHYclP/jU/HkC+/9wTOt4+aQX/H1wtWICGE9odyfp7MzxW7i4s+6mAGmvxfKPx
+m4FflgyIdJUVI+hAO9DJI14XxephBfIkpCj+osd7NSVvXI5HiYW2QpbwVtzndMpbQR0pWD8OTpy
eNzS9HhRG0ZquTJj/g4mrcvpQzGIpzSvMF8krL7o97L0Fw9+S5+DZeBHeIzl8BHt5MeJwu1qZZKt
wLnn9o6TJkvqVHWh8ivr7EXGM1+bD5KvRUtBChFAOTmCNZQ77WOPtNy7kusdXBUdXr1rdIHMJASx
6RTGogs41PLfnyExvzq5o0119rYwvT85lGGJ7xhuOGzeOVvOA4fxS4hTcqquynCAsFz+uU+ynJif
m0dV79oeJV5e95PsgNa4HuAL6vKZdHPgVAHpzEyNs0VBUa2CTiDXfH8jmdVTBXM9uyW5LvwNWkzz
lWrpnVvuhp2A6lKfDNd9GAQG+o5E2mfEbVfFOGIPw4skAjFAYOsWKr/aW6GMdMp7E6YVsKFNO5Sc
fU6Wsvq2pGsX4g2TOV/FkkXGU6iRLeU80RNIpD/rCrYJJRMLlR0P/j3aWcPO7cEV96JQAoTZ/EGJ
e1K7waZhbfqotMS1UPj+Rnp9nbHy4D2DhWYgzPQgV7s5sqODlobDLdGw0H1J3f2kSW4iLfion101
w0b/DB3U6rTQdURV/4jTvl9LwmJmZ4ueo9EuWY6XMYkDbr1n9pVPW7gMhlSHyypdgK3wlcvwXlsQ
HzUSqp/GTqlL0pd6s7HNUIgl663dK55C1zVCrZlDpIePHZiM3VyAN2XFVfpoRvcDrBH/dz81+x8U
edcv5kFK5ioVXa76lKgNI7EqizjiSlGWmf5rl8tTfKULpneJqAdpqG301rqBtpEpaqQU/dFTqmKa
pHnZePkdeW+q26/DFji9C857B1uALV6uuLpqEYciQPcabh0KIX27yl5aKgrYVxVth1WM8zm5mGZf
oiYrOaviWt8P6olrzqcmkdPgRZdiccj2xnT3n56/SkgzJ36i2GLvwDZGlz/lPQTU6ojBWJuhrODY
VpDmwIQDWkBib8h6/2KgtJf9qN3DN1OUWqsGHG8EKVuR8PyQpIEZQzReW47ioCB5NRrzXgMAmDxR
EuIB5NNK7K91jO7HgKxBAHypZOJp29pQbw8ckLFUCOLUzBQowflYrD7W7YYZ9+wOuoCRwlIpTD37
8qwvUYmuSHkIjJ5fwIe0xHWvDfNyDgFpoyGpHId7cphcWaQZpZo1NjoWhkKTAABTY4lcnQVNUExS
09u9Gvf5O2+Blpj9tmxdwJqpo7pqRMHMjrR7H8BHcwLMHu3unl6mVTmCvwgK15EGo1JBB3jhs5V7
Oa8IJJyhokuPHD0PT9+gzAToc0XhRutm4m77hc76rINaPXa+4FbsXYYYgXALhIs5kz7j2FnF77vf
pA73MS65aP/mJgRtx9FuJr7wAvyKRSgAVDilOW4o2ss7uTaQc4K4WfJIxr4ymRJR39S/pZ8K9qOg
2LsiNakvs5s5rFdREEIHM3CACVxsFn9Mlx5fU1grmLqTQ+5OkMXJ1vIqGSdveU60F6pCGCUnQX1M
BDeLBX+9jmYLYDbulHEQuzpevw2hK5V+cbpiX8XRiHEMowc1o5w6x7DgXrU9IAy2GupF77o3FQk6
zkAmJwfbiQ695a/nJgPsiAghz2DKK3IKoCkgQ26//33QvDS2Al1aCCMnaty2Cq2ZGISaBhFdPaHf
0tkuouUIrc2pfWLWDqQn19YqmCEQNXPLPr3tS45RX0QZK9JrwJ0A4gmeQVLAXUx6PDQ6x/thiUEP
7VH39kwOZ9terTNklWOuYuAKA4cT0IiX15rSVByOCpwKUfpcNVouxqpAmMupxOyRi8Pa55rY1Jm7
XsILhexvnQuzmqZvjOjuLDYoRlNvhFqMK9AgbepJsrMcFE6zbiJOneUM0JTlaIExhM8RoCEVvCNj
BDADpQeCyl24GZ4kyazigKpWFC/eomXrzwnzefOGCqYegHUKnemnrnvng7bZf9rmA0gcn0ljaSK5
n/3LK8E0qsb45Rhf01XVEM0/iBrXHSFiGygbOuSW5w5ar7QU8e7R0mcZ5gLn57hW3nPpv2uuofBp
M60joM9IwnwV5P7SQWGW2f7RV+yu23uta3iVglMYXTjL4wHt6A7WYHJV0TMtw3yuzne1RhcV6GMg
QTZKGabiFtXQhuBIUmP1MT8yQPvh3/PA1XJwY5u2RLt56dDYhTvMiJrndHplLjn/w1NrAwIvX03Y
KIslQwiFqNX6U5x6RfApOuFeEYVuP/YD3LWmzCmuDmofySTRNv7WQp/H7mslqTemQQvlKSfPi2r7
T+Xj0R3/y5058fkDajo2PNMiMPN0wjtqarJ4FjRSWDbhQUGXZMMgEXvODdv6zmeTIOkn3SfpkFJB
OWHLDoy1trs6AftkY7sU/B/33Els2LHizq+hKL/mK9ldvuXONq4xGbHN8HosRByiqL6B9hePpx4W
DeME5ZSqgggC5vx44VAPrDBW6JoopNOz8gj2iC8doYVm0Jc28jifouLW6JMI3JiAbjUv+oR5QX7I
QrDnofMbIPi+KzoX946tmrlbd3d/XmMq1cwUTR9sQ7FYvLiyQv5EL7cQ0UnCHjR24C8U6b4cHgKs
+nvv0ozARcI0bDgsRp2eaQhBLPrzd8a8WppIG7U2xRMqk0VARevrNjm5rANxrc6Izpt4bAPk5Hv1
O6V53pa/3VlNWnmJlK1RdQS6RlZDo0jwaSWyqP/jsQZVGqJ1/TVm1CZ+6xQXCjnXO0qZiyeUemjl
qQSvdFkev6H+uVQVfg2k+4lhb4sbm/6oTnwWRr5Uw2O65dQXc2UZhvBJ3gDHyTnmuAIywMsL50Ou
HQavYoRFmS3sRNeU7ThMHrx4VyBkZF6G80+4+aKO/edUrSeki9tPdpmoGZdWO4nmX55lr1zVgxU4
3h84cLpf0D38nqXOpDQ9d3z9X8N1XIu9DQXbSPzcR+fO4rZZfpPt8uW+v3q6KxSIYDnBL0tHD8U/
OylRsOJ0Nq/tQaS47mil5FmfKwwT4qZx1VeG0IWbGxIDkpcCsMslQqUqZFxzNLnf6PF5wnKLbGda
r6P4gcY6Z1hZ7DTatdlW++2p0TCXVOB0QxOPXgd/pZD7S3rpCgp1g1rik081GAapZw67oKJdQuQx
3EZ95tsiHivmt1G3d6dseFB0FdAR4OZShJ3V1U97iQ8jQWsleuJXYx6QdHZzJltP5wo7WnZfl4+P
MB1O3w3h8qULClO/SwXLqs9q3LwKuYg2YdTKS/xbehfD0lp0ZzBuqkpFWpokE3lwjWEEyum20y3p
uCtuTlcl/r/H9cZjfEM8P322GjWK3Da9CNfPIQPyBWqF0lsIYcQm5pEb2rspDiu1SiGeaxpr9U8u
NCPYSlcYv4Wzc8G1aKeBry10m3JLo/5iigard91DEh6WQBg1CzPWJdm7X596r4OakeY6WF0Wc690
CnILui/tHrYIBoXgnP11rF77T1/JyCo0Q3XdzwzWQTARlOB+7kG4rQFJ/RXgox72SJaZWTVe9G4z
Psn6hzt/tc8BpUdnqqqNvl6cOaON3OSJlIy9DHV1c0yfVm6ikZgwvOKptC0lRGOUzekHDPeLdqZD
g8hT5UftP8+40MZWWh/s4R72WMR1a7ViEw6Ph7lW/pcUCwEHHhCmMSUIpvr8UaINeTMGKoFJ4RHP
uTuaS2Ojy2Y1vZ6Qbc53MWVm2ylFPp3CMT38f9NABdiDBfnmnjf3QGLMBh/3BhMiW2Phvh2m7FUN
5Zosqeius/GwU78iaXgQ5Ycj7CSxCLsOyJ3qzkA7/JUaPP2SFV0ebGzsKgvKEAlNyUgtz3Q3oXio
WyXIL5rLUEoai+LFmY/vt79yih5c4EK09RtH+awlsOEaVru3VTr5gi1mypxyUfL0ZliS0mJg0y+1
ULrHrRYgDkWvx/eoqljA52I3W4LvmAHegas61RJDqt+0gUSZJwR5f3REQE0s1MFukKhkAN6xUhoZ
QPEGc/88YZRILSOH7R+P6G/N6t35jRhzSqc3U7wT+QaT4+Tzt9LI3rO4W5MjTa2Uw7MaL6TOz8NV
DYbIlru0bzMkjGtGC3tSdKj0F1q95AW3B/e89Seq5ZTXCskyutK5kxzE6usEvMjcW6adC2FW9d8U
BaPsXlnjNgSDgBfvieEj88Vv2EoNlgodP35/jEHLsAAo0V98MUqexlEqXZ3Ue8oNXSEpEG5d7JI5
p6c/2zc19szI8VVE+M2djVDqoxCs2Sb2JVS5WDzhQqast2Q772R5wuLVn/Iz8zusHwzpKycYHPqY
75jI+VNxpIQdd9We8czeH0ZiPMuY3jM/4+5iiwon0qrjEih2PNH3dEiUQRUT5tjNTbybBF3Vb+aO
rNVmXhMexW0lKyLaxmtcrWESb9adtsefVuOeTxpx3KVLccGp4x87QzLPdphz4Jkklwgrw2rgeOW9
GeiGePHQ8G4IDMDzxKbBEZjcBFWQWw0ff8YB7j+AUIA3kjn6cs2u90EMDK6uOv6dC4ooOeXAPlbn
7+vHbpMb0vgYyLK4fypEQfm2ceB4zoOqeMrV0hmC5kn9Z5znFYdPX1otAOngNWXgBF7FRZZFIXqz
aUZU1alX7K5fNQhwCwN8ztkBEc2UtWoNJy14h/BZq+IoQJwJfKm01Q+4q7K1sXlT0VaM3Nz7jEoe
lRpQGkXU0amyoVEjLyEWVNHWsztOmG/qJSnTUneZC3L3Y5SDdmc2J36LKbdt0pZELbBTg1pC2Kye
FocaLz2fGM9+saaSmlDop87dg8/PxEWyR0xf9pNlfEGapLPrzTGig1qiMoGh4/olrwLF5fh8cZuH
kNVEiximG3XImeTnRu3UjGDTtwCO6hJ9WgtQ2/EcDzjfZ/7jwJ/p25KnKITHuNgXorVKfN3d/Yy2
GDH9cl5sVouzWwR5roBBzV57wqr8tjEi1JXzNcKxPRMuqt9UdqiRQpR1951/CODsByIPOjhc84Pl
yuny8BU/X0eCNnaBLWETmmyTJcYa21seL3B86PIgokoaYVgwwKNRv50r9NF+O1AEVDtBExCg1dPT
nEtswVWQSbJsrXTTEv/svjUmePvraupjwIwfZC9Mqf2TOOjn0mEXyW+XkLrtIqfJgFNaLmLioN7F
dxrMIBSWmec+SjZhUdQyHwP7eyjfs5g8UyT7mt67rDNOe1QS68YOryVoug9J5r96mvR4ClVj8EGf
weWKPxvFexl7QbvXtJHUy8FnKacIVYxMxIjKu9HjoCgignQYbWaIMnWYpR9KTB5ejqym6Z2s4d+W
hFs4B11jgwvBSH42iaevYz2dG0J/LXjb4ZjLPLwXn06e6C/pgCwHnVT99cGh6pGGMcLAOdJm8TBm
PHvdb8kpIVbcg1ER+DThLzX3dzQCFDf7KRy7+pjpUidywR0j0zmyc4SF2tBni6vQtMD0R1SbBezD
FZbO0Yreu6GIbTIKYwwjW654elJPPTW+SNazejeEN3SCidiYjxrwkOKQZyZvm9DiqdqYiwBpRQaq
GLQf3/aOh1PZIJC6YtAiootJ/1aazUSPcH60R/Le/QJAsQzMmgPowfWS+kHDGlxd7LcjbW8egIPu
B1dlwypYvdQHrbU3KPDZZvzIquJ5Q6aKlAost5LTj55QZfZKu7vQF4iw3o+rYM5mGhDzLjzfoS8r
wK8YW2oFRlqvXz+/4Y8KLOWRyT6b6LBQOL650r5IkwQXkykmWij875UNWEfd1wpaI0skY5aZ4Gyj
XO3VaJ+jGmk9tZyAX5XaXDDDjUYBKWWe4WFqXWu///LUjVH+yF45Qv1aL+R0LvOIgJkiU3DYYxJY
VVv7wwqWky5Rel0VY4ryLZUjG7IyjFLtH7qRVNvhec7ZmH4ShLHB3csvVqV4VrKAKE7V7egESa5N
BV8pUsl/scnMoqcpocI3uwYY87vfM31Wms70dPxrced0+/gczgcYjv7qZb3h0C/G0quxcKO4FCaa
5b7vqn2tZMykR9BUNqn/ywH2Zejh1F1dFHUMig0QAJhbmvOUp6I3/eZFhvfrUemU3KLZmUW1VVqV
1XwTYtW0taN2sJg6GD0weg3VnDtfKpH+e41ElwEULRaFCrK0JN/Ef0Q/y/8nYVeUJj1Ec1etMYyU
UrJ0cFEwzJC793NGMVMo0s/NHye9Gm1oM1aF3endDLVtJSrewwVmiQvVE1N91GDUvBTZSLjuF+Fl
9d69txdnWnFoGyjVjupukYFPtLsg/ffLhQ8XIbDm5MTDyXxjfhuvCAF9DmuuPaB0/qfnL8ajm4Dq
0qqocmOgO9E8Z9+frOvu6k6+DJocODl9W3cFvfIbiYPkIR+jzIuT8HZ5O4W6PVyyZltS+OXBfKlV
eRxbD+Zn7XEIiqJjg0FYnnlUgCZWkd3DePhkRMHU7AQleASOFLmE/cwwe1Z59MtolBLj740Xfj2e
duhs18VpQ9mtvtai5DTeVdpQcGWKzhxY2KLiWdap6S+GkrNLdcSjYDXaOHAefpuDoWOJVj5+DZ06
7Gf3yvgTwHU6LeYkwW6inKFQ81krvyoq10Dow/0JGsrpVb/x1imFZdFopzmv2IxMdfoxch6JgqIj
OX0xlQwoehyL8yTiCzdOteAmp2iVUebLQgYJGvB47oPJnR3akFR6Hknwq7D/MXHXRPiTK+oE78Ou
PZmwnKFOnPXjqoHepqcWgBRv6AnOPHKOLN17nqNGnEHlNn8ld8EAHnDI5U2eLAyNoxURD5Z5EAuI
udPHgm5tf6+BucP3zdA6cDe1osoG4bE/8jIYWYsu8O/iel/nBw7nA6yNR8jHR0kdSPR2TK/TDEvw
TRS5K8ef5KkMod7GobiLD8Fv8htfxxcA0ILAQfhi/DQsGFaTrhVsBd6dUD+K/MpR5HXTV6upnL7z
bgyRwN2HlAqO3sp95b9JJhQ2EkmaepF7bwvzYK5Ch7xsFlsv/GKClaD/IS84WizwXpbIYEiFJRxp
i8MkKHEu768SAcXe7cCAs/1kSkQj9GljxhlxuNtxBXwh9FfEZnAg+2S0mnqgu/mQTKh3/+88l0p3
F5/MiOemI2Z3SpyAdBzlKXsXO24sjnLTsWEC3Il+Z7eI3Brxi8Act05/u3VKeneDGSogRZdX8Tuc
uV1pT6nBvUBGc8k8z6OPolCP4E2jYS37zp2h0bWtyE71P5382LkjdrQdObMvmnTfyMi5MU0nfVd9
JUglHTo6rZ/T0gMIBTdJvREmWoLXaVc/BqUmWss97ZE1GhN4/VN1Y5VsWKhn5qddZ3uDx5E8lrNi
i4YVaCqyqn7qwxJ1SRHWq2I0Li+x1wmY+SULOSMs7iN7w5SxNfTcdydfjqX5h6Vm+mfZtTEsGL0Q
CBmed5G0wa2HELR4Wz6uhDdcQwoPGzGL4a1t6+hMwE1vi1ORLxfiCwxu3iHSnm833IpE36Ncq0vs
8EX5oLoE5pn+2wTniZKRS0aLHMceruSgJM/kAKqKdE0HzOmUc/F+jlFEEpmLQ+rbD+hOQNmcRyb3
fyZ0gsleIngxw7vO8TtOxqtKRRlRFfDyi11cUwNLUPPr7q5jbN6xuf+2zfikNaen77PSEYvQ8+hE
floEllI4JkFIMlB/N8qhuVFCrzIPaqUNGsPeP2gY0c8zhnuPLPXeAv+rGtIRn4K/o2HK9ynLgXT+
/bFk5ov3R+ARc1upKBUbQj3v2gCwKv7u6CgPIuPHMeinNXpVyZdpTgEod3Mp3gPlB8xv3zSGi+Kq
d95qiT0vkGdf2gISw6PodmL8YxUIW8Ml+bN1X666ufVc69d3n1fUIWKBe+1fdEbqCVQMvfDD9Atp
IKLrgkIENKyso7+6g+QVI6p7BUO7qcXoQ3RY5VIGNa0S4cx6E8luy7qL1tJG573BjsQiRcj6IX0V
EuD0+colxQSqKlMkvWmsRN3uzSrPJY5q/YVmWi+D8rl/MRnRb105OpJDEMPE8yvH0MBuowIc4VxT
/gKyu/f3ws5eJEcSgidwoeTP+tT9AF9VUg1oM1mCREJU5UEmV4Ok0Ptyqjmd7Y01QAaywQcrWFdO
vi5mv1ItO/f8G+XxRgQpbHqXilUFIMyxb7AJGQGbM9gj2Y61Bh9dGbjwhQX9W0o7qvZ9e8zBlWm9
fqs7foBXRRldot57+NEDME3Vxw9mbklinmFdWkoIVey8F2ho1nz6H3OZ+8ly1+YjCjtwjlzXdINS
5y4KZwo8UXCfVLpNpHxPZlf8oKxncEnGvx2InolG+Z1ceLVleiMiK2xFQNrPFJmlCQ15mkBmeQ3T
adDMisyywlV1Hai6ycqzwyfAukIhOYDoBIlL6NXsg6IhkdonvuahQpTWjiSh+i2/xwGnwB4Bb3/D
RX/HJ6XR2srqF04tbNe24JZsioSbBT2UWjG12qwHnuoUE5KIQ3+6BtWiu4OSrRkBF4azR/JIZR8R
fVu7EtzEgnKJCam0bykHx8u6334uPFCP+1IsbgZhDPFFPUXhM0JdAyGFJJ/c8ei1P4Ob5zmj0QRR
6BNtXf8CMlqAyzBuK2E8mS5IMcQQS8l+mt7fEc+J5ct7c4jAAkM4ivsDX2AuFonW7Pa63DqFok8s
jdK85dLD5TXmzJ1H446EfxB0XQVzOusOtJcytlXy8XXfQYn0zv4RIRqlVVSZD7LJTbypKOOU9SAg
9ztwnZjOcZAiHc6rRAr1P3IEmas6iIfMyJIa/gi+SeHZOKs5B8dYPszwtvQZPp2MBsptuhSJDZ5E
SKi0Ij/QL8D1xJJJ0Rw4Yae0JJGrqp8BxGYs+kpfbBPExoUEtI2Ik7bU2iqu2OPtEbt2blC6K1j0
yNjdNyDntKcF2zvKVhIh5DdoahiofbTfTS23dgcRPW+CFmR3zmJLXTs+UozJLA797wCyBEwiz5wU
i6uM7Z43P1QX0j//DO3TLlXXgkMk0yKLyOFc0UjqnMhjrnjeSsD0tPlNiSouI4WlGZ9UIphxnlvL
D+mIMRnbMEO61cUHQ/mMBtEeqdUOjsIAa9mIHgVSFIpbj3ZviA2A24ZYft6PQqa6RCG945tPxUk5
/lswdPhZIGJucO4ZyCvA6rqs6g40PYVdyCPhG09+WNRn+0+S6xprHhpw1mSJD2qGw+YXHIZrzTvg
3SJ8QGZq6y8HYCCLn9+ct0fjUNRFNhJ0egJBhQ/q32zvYTbqm6YN7efXnAJPsCgyTfmLmQagB/Mm
p8HLwoTWpHLYRwoUJ4M3cQ0yMtXkRJ7+G3wmO/2j2XOK4pQsyTL4nxCOq5RcqrrBv+LSt7RUDODs
Gh4kzjFIkLRyhafDfgYIQrjMsdrOVvfVin5JwzxfHa8Z3+KPz06ksluvq1W5rEWYXkw+dPsxkhtp
nlauvTs0R8lp6Vkrj2bj9G7qxaGfPzsGBORucFEmNRwo4pTBeu2VQg65GC5JKmCrFez279WG5oYE
tHqMfvTq9K+AhKyovbgpfRKGUO+ct/yrmrXELyW95yPTMmIVOhuY2ZAryS2WOTt19yg6bTJs69a1
j9w7Qb1K1C0fWPF/uDvZHYo/cRRVRlRJNIcXU4sEihoYHtDTQU2GqCPiTCzDkCvyJXutsMi6ntJk
CCPAePey/UUDFg1T9citt+YxdS87PEZRuK+4Dzb1hL8p+Qh4CsFJk/7UVZfQYLMOq+r7v5zimb80
VthRWLFfHDDaT8y10cTjT/uPFObuzRXLSCcvTRvRr8S/WCP4cI4GvGbTc8rJzNK0VwJSqcfNHgIR
SkkxcSwa3I1an74sxZPfKAGnGLeMrea1EdiwK7sGqg+bzNDUaTKfWWaNQPCE3B6v7n90vdfKB5Jf
1urxa6CnS0NvYB810PLAxwZJPBx9GreafGUYwAw1rAIEmWYMDsk0iC4ujlStAMdkBDGHdm/3BCBD
A5wz6lQoAfBfVgiUUutxZ1FqAxETU0QPPXFA2pn4m3JqbeFpsVpQyf6ypHx4jy90OHvaWUNPiuQC
lMEYOOh/5XfIW4jvaoSv40i4gmXKCoE1+zbCsi5TLgmyBagVmEIG0Ihxv1W80Qc7BhBsvO8LX/WV
vEVPX5gAJScvNjVYOOL7xjlYTdhRkHeoNDuXrLoJoSA9yAxXxbtdZzyEEIaCtOUDStEJH5+RKUvG
YvW/S2ggs9Hk346L28ZZS1fUfF5gfJ992VDKYIrr1dgK8N5y3zR18nYq39PXvYBJNNng00eBInoW
aqFxMcbzM9HAtJthl6DodLzQHaXu6LT2hMWvBl7g1v+7bTqU5NDAdt3eTNVdo9fTfm4jeCajtg7/
+yTvok8fZF1HIimTWbvHjnZtiuhlD52yX4+aJ3cJZqku3Bpva1YpceWEHzld3bzH1QPkS1x5azPw
05k1oPcndz0z2zRmajt4hmul+w/iuWZanKkXtq8U03qPNS8FmQJszZNcJae3yKfPeQ644+yneqlu
ZYs9Sp38FT3R8AOo4upYAHHCfqdyBScko3t8MsR2A+Xo+yrYCINRqq3VLD7a7Uo7rnDNcvzKHPar
kx2XuFAFTAv5iYCbVdYUYkUXSSim8oQMw0K81KT53/UtI2NIalyEUfkGHDxX5tvLl4nJPrV1GvH9
yO92RQoMT8vTk4O2lrPJhSOuahdnvUIHH5P+YwhaRjs02gwQ6cBWVHYkg4clOes014qI1ra7Bz3c
jHKUXmKJMvbbja9tvDlCWf0wBrm0qejGaUUddPmi4NXKAaiEOqrYy2vur4DVxF5ylMckRNr/GPBT
cHR9ny42ZaAKpbjbBgTmSqURNf354eQDvLG99GMqFm71O2aZcjCuaSzBZwNMva7EVsrr1bLw6fOJ
4PhaOyoGAp96WAbw8W8J51OaqJJ7A15UWaSNoS2XHEUOeH46tL7OFjlbcjo+l06yfOYA1DIY9JeN
hNCUe+9q2m00XA9aYDNAvcJaRdJJ9pqTIq6ryT2Wk61XlN5zQTnixf+xlX2xCbLkUNgIga9ej0r9
4SpwYV55T47DbyrUBi8nBdJh3ALZJcAsonJn1SWGKUqtx3S8mjQVNlgAR7psknXhD4byuoz7Oa5I
89KygQRXDYOncD4l1I7O4WqN1d+HBaePUuhXM3kPtap4oQ2soX2U2RvrsO/lahPzgfmPBL9YpbsE
rp+7x2654M2pURRGH8rLly0LXyE4bYDF8812FvLEmQlVKY+sFtdoGrEWCl3oYSw6KYJUQbI+5PmB
E8boPGpDjIQL0XEw0m6T+Y7sxh4VJU943+gGLp5ijRSHB6QocGODv8gK70efZUk9E8lynGc1D9sk
7aPDDR2t934y+D/d16XDYXJf7uL5f76k2QU1hR7S1h0m0awe82bgnf2c2PdHrIMhWj8TmhYMOEB8
QbeJ98c8RxFaErqUum4TrEFv8lI8A2abSaLBNHhMs4HB1za1AwkpU9vyBo8qFl/lJjSLnSIL0Zu3
PXVM4kVebTjXfPZmUL9rY53G2kErm7CfbTCYG6hp23ipghyinRE0KiIdTBmaYoq3yNVitwh1rRSd
Xeieq36wBttekQ015wCC+98GyUp4ZhlsfCArRvT7pja0ev2uG5d6xU1FBzHRWeJbA0gzBr6hzVQS
GcoAJOKG0BnHaPxh5/Sn8OySmjsyrhrxQEv9oF8+8Ywe2qy1/zReNGYzADVLY97cmaNi8E8qNLPR
lR/TSMhtLyeSghCglUcqnEUYMbD0q7FaWppQnVLlPNWlX5Az5Pe5je2z0d8ZEgh7e0OxUp088FRb
NIrvV0ZdbTzGQNO6OpL5iqqxUerfMqRt8R1e1FGURWK/oLEk38Lfpt6cIMaqCGdm1fAxW4+m35GM
u9YmkpmTN+0nk6kX/KGCBICPdr7/aSU+K6AjuJNRFVY7K5aofkRPvuRLRMeT2SBbom/Z5DgSZGQB
yzxxzgSPbQHhpICb/167jS4jLNPvZ4QwBoKaew5QV889gx7gD9aLEn7k+sQLq9oCGwCKsXP/NHHP
LS4RGP2yWvB1N23BjPmARjy3MMJ+fZ0Z+hHjW/aSrWS2mS4jeh1ItdvEwmWh6ssgjdb72TQUyMYl
GhMRgS6vR1PT5jZBrOR6Qr/u3FdstsVvQZRDWK59AcugAVEMPeEdq3FyYd2N2hVV4As1SHfnD0PE
nFX/ZSzQ8QEJs3bpQVpi2IYzKSrjGAGakkoxH8KMDb68qmYg3KWHSeIbiJZwZ1gIUUAgzAC9WnG9
nDPVGGBcC87vnd9Io0k/D+4Db7S6Rz6weZndeThMEjEvdUjODOlakKdpiTJ9RvMgL+1BiCyr5rtY
HzyNad/I+L8AKfvEoLuqpir6BOy306In40ZfJHNM4B3DJcNJK9u0pz15T05gRLFyoB3y9W17NjEE
9dFQm/viPsNq4RdPkRfYFi9EVw8nuCF5Dfxy0plkVK13uy+VHV9KZxWxFwFcxFkE082gCyWSTlFF
7aIkSXR7sDGnd1QyY3RajqpoGc5ASG2fPuB6PaXZ0pk6VFWHidfAvAO/ReyFjkMP3Z0Rknee9tjf
hw3scxc7URshXbm5FVVBOfPikbwIxbKhl196F3JgV1Ajv42GOBqiwTw/ftw0U4Y4IDHl1PZ7COs1
s3TcVOMY4ZG4zXHyGDTVeuKOwmCjJJ09nKUc6mcdsWZJ2roiaH93McPov/sBqkxoaDj+BCW7wTeD
LQFy71ruBe9OoPb/0pCb5j4lFq2oNMXwccErYsRRVSQ1vz/OkLjcx/eb2UqTPiFoJFHxJP/G6Enp
+qdusiOfyzMJ+1C4rS7NQVAoAsAY9yetWs2+S0rDBW6KbgVNf7n8jxyIfW/8Zsr2qmdbcjR7ayKX
0bimcHV439g3hWDH/J3DrliaDhhqDIi4KiGJlg2Vnky8D7lj7Jgyk2x4ic9I2+MCTs/DdzjDeJAE
qnK0EgFTg9aBwDTt0gEGyWDeqMVRzwCeO4jhEVTVi8MrJBq95IZsBlpNnH8BTgLQMn55sHu1U+Is
idU4NaKhTFCnnGzLRvnNRW7jOUzKzQ7haLZjyAnTLymUw7TFlei7NymPyWp5wMrLZa1dYpmgi2QF
Yhc0R0xOgtqIBY+sLYTxBsutIJbb17xM3GY2ex1o4jGX5pwD4gvKLLv/Eqnr1O9b1m7kf32HghVb
a8GQ220SuVqeIDgD6vGGVLoZqzjvVmku7vWCWmKrvGCu0UZOfUKPSz9tU7V2GHjdeal6pfzW86t1
RKrffwxeFeEvGIOEowMr4MYFgA6PPaYj5aMlG+bfOUYFqeR6tZgaokMfGQ7vtbrz5avkVD3/zh+2
hVfdDTmU33KN/w3oLWJlp97ungXhVLMprw0Ps3X3HcdlHlXIJ1NC638Y0zIA1cVSKLN5j5VQsnbD
YgxzjzbLRBKSYYhn3oqB5PIYOESdXr/QQvkki3oYqC2LeFmty8WXrrfil//lH/XqryEVHl6cl+db
8Mu9fLOdYkvBsNEtFI279Sej01qfFC2iSGfzWVyEdiviryOeqa9RkKWgpK84l46JqPGr7qDHR38q
n9HniZgc4J27ziGgX3CqPlZPvvuLGkqVJEARaNHvrJUlhCrksCgKdyFEw/6tpnrGvnfCm+H2EFWb
P1gSwzWfhQmNPArgPNX002QcTE6ZPlfMxz5Y0ZmdUspPXS5I9EOEISCzMnGCi3R7RUIELXAxxUpq
vcxX0COHUKKTNwZCBa3cNf5mI9kQzFnQSiCwoeXYebFNC+qI7CkHNC013dYvj5bTRn7stEcK1Uy3
RCv5KrJMsRQuo37o56yf41+J7hWRudYZW1Tm4+OeFU4beCno/j6hKiP356gZDjMS5bNsrRDfEB0M
zfIGHJS7KdBPf+XyaPBtPVV1ugrL7WJIGGF/7s4JMpyqsLFUUVj5C6x0zLPI/BlYmJdDNLn0qeaG
74XPvL7s83w6q1oVcsGgI81k86CWzJ/YTud2at8SDLiVxCQTteiZWnWkYfCB48Ry66XAUpvN04ec
vuXd3W//fdNdPUMxR+EX169BzI3DJOlf7/bTD379IqzflKdckWrqavRpDlN4dUYpP5NLBOvTobSV
/Cojmcyc7vEwgv0E+IybIrPFW/IjFps+nVQ0E8QL739QpcfEGB7+23d8XFeXag6r1tTi2J+Sil+6
KwX3ltjMcEhfrFG/BCBIyu8b0z+wqM88Fumr95WaAumgd2V3OSf7k/PvS0exeidIhiHm9WOufeLp
yXWbaixqoD//NHmRKO+nwBywn31QDf9l3GDjwshnutgZOQLfmFCkomuUTB7MEDWPsHX0GqNFha3n
hzKSOD/zjxe0R1CyINnsae/DKoikxKwF52P6Oprx5ZWIQlCfVqAKZdUl0Amo4ebU9GwCLuN4kCMA
BLVASBdsig2dxEAaXDANtAnaipHAl+DnB7TrtDXpfHmAQb4yx8qdCkJoC3Bsi21xpJXOGEl4P0y0
/tQ+JZsuCoVaDTZtOvWQzOZujxonecNrSeMMwDQaU66KL1Ar+B2Rk+he0QSRMwyHmWFaGWSqDPQw
/VVYb2m037cnYmUmXsn8/FhmOQprXBVJIWuKJZBDidwGkHuLyddYMsU4dELlxxD1SAxQgzWCdPaZ
Ko2nzagfNTicWACO4PCmSILl4CbLfE70mqL/s9yroKLD3ub57pd/ba8AdVXD0f6V+h/mEk2fz8es
4MkrTRAn4LQp7GO9K1xLmXEiYtZAjUVOXhAtiE40pTG4Jo+z0ICPdxwBmizqXoCrN1589qqUKWsH
Wn0Clg8fiBlj8fyz9CNdP2JMLjRxsLEbndy2TWOfHrDLlk+i6x3jsq9SWuGlEHW/8vLdPzXr1axy
TU5eNwyx88+W+nvX1yMfpnYDPLVmHXoRI0tc4ZaDhwfY22Y4lZuQGfNMtTYnOwI+0Qt7hAexlx59
kRrv92FQLelx0uSJYcHhwIdy6FN1a1AsiFRVA83NuoDwP53lAYfXM3PsSdRKakeNXmK81y1nhMhG
L6l+Hahz0EDAHX++zY89GkgY3uKiXOfg8Va36/dKqLtB4JnLzIA5kE7u3HtGcREqgMKZAQVlpdxC
BSqblqRqfS+bFKdYp1h5tDgIsyHqJ8vZtSFgNzwmjSJRKKkYIEo/jjI8pAMZSkoVVJvykfh/MHXs
ZOPvXmyLf7A4F+O78GqpS2kHO5pBciVfQTdRgPbbgD7GGMkEqmdRWJsTMEDvKP+UgLD1/IBrkRFp
TnoHS5HB+uORpAqb+T95LiDu3dUOocLwtMmai+Kunys5iUt8NfOgPzYj64X3nJsS+j3xjY0OHsdV
mu+vVx54h6konTwzwnFDFYK2hmt7AozrDjrXIAejPKCyJLVbynB9i4s5gT2C/+pQ5thma4hB+uhp
toPqkfK6R6uVsu8dabGEQillgYFgJaxCIwK18aquoJyXTPlDOt1xpt7xbaGZETzqhVvtcRIy2raf
n5w/Sbw/5K+ZjXdgJnWZSvSF71+85XHAOcGam5BOR9xzy6Syn/TE4ZyYlVd8Whhuj7krA3axNEL2
mVm6N4QPxJC+P22xTgr/PClbK8oGGTlTbLqJgl2zkLVB9RcbJZJqxPsJRLfrqnuDEldAYGZMp4xT
AOJ0Mtj02TSTRy4IGKV6T6mR6Ftd1bqYza4PLquqa71IKVsc5YTTslCZOfMNKjB0D33MrDr7voqM
ImPs/uGuiczJKNVoSTqaJKSaIWqLlNKmR66FlfH8DswhvwVpirMS4mWsC1wqwnz8N1X+sLWTpqnb
F66bjAH+CUtzYM4Hu+MLh2hJEtmqQmx8dD9qBYIsFIAMJwqCBfVDFyJY3bXt+DxcpMLvXX7+LeXf
S8WjO5SlUp0BztyQb11xCRahZobNcMdTm0PKaNAbEdVpZ8CXeZifVUgjilUk6wHikofDy0Y7pvsI
kwlcfNkMBxQzhJ5F4t9PGAU//gJXApkS+D+NM1G3FYA6umdrtaFgWYTnImNKSQ9tu+SVJO7AGeVV
fn5ZLSOsBfmsBRNgx5tH4cLUgSRHKQLWqNwkIy1dXvnunpEGtmZDKmMN2WAhSO4QRjqAJ21V1BA0
c86CLDoho41FAU6Ci+1YXWZpfCuKQ4/+DE+zKaEbq/F7pRL435+j2U/UosTUNKLUQi5Atf4nHAmZ
osiJEo2fghCCQ6zVNykDn9bomlHaB3RLqcGmy498USqNn1UU3jAcj+BywWe8bmQZnEaVkZdRJ48t
ZW57BAhOFxcE3OE/YfB51yn4mANZyIm/17T+qAhc+XAXuLZ/hRF3TPNrJaQ+sHCBFufCC5LTAoe6
qESycoaoXz/kPcSrHlRMS3WWwCX0PV1ynZX0w+bc5wJ+qh9lQp6qwn+z4rPZxEwnDdqJ4OsxtaO1
ZtwWJGcnPzitKOraxw+Mvc1yB3ohggok6mhpvnB3qVT3aQMMK3UUgNTKztcRbW6pI+rIpszrKaqW
fYX7BwDbmfrowBPw0cUEWbxNJo9Fhic9TClW+B7URSnIp6/l4YcsGTaKuIWRCn+k6qlgoRhWsGkJ
jy4Ot62Eev1yKzH7CPfi/WBeICmj9Cq3YNWI4V0Ax3ql3NIyYUQqdlxJZNWpEIufvSTRiThgYX4T
ld6XA523WBG3Skqnbi27op9kRt5UMKlpWGj0GaZaIir4TIaTDu3UC1DCKS+o9shmpWHzh29kjnJ7
4GGiR/V+vbvy8u86hZ5JFJnsEkvpWsFlNDqYBULO6KtXs297VDdln/ySjUlC0XHj+mRsmkaV3uLM
w/6Z/ouk+Km/W7f0Y9DwbXIKkvZMMIv1x2625m64FGu9sXCnujmsQuM3nZUTBgZPjXcoG3GEsLG2
U5P6Z5RvN16YWQD++i5Bl0YHxq0HtjMZVZZKosrZHuxaW29hYiUAxrxEEoP8ZN7hJEQLMBKONPnf
gBu+HZfVHyUHoaiIdldU2ntAZV8Jp3sKLnxCDH827SJUM86BVTHZsbc/8iHBNLwlbELbwVLl9+WL
wT56+p2abk8W5yM2Ujs5UipcSEMor+Wsf4lSy4NjbiRwSBgDBefFpuchuiveCsReLTS6EUtbB6oU
rOB355IhPg5bw+bYFSeFkXxpInbo1KXUEO2AFuy2doC367qj13Itb8fXxJ68szt51oa7k9bVi8/Q
eDMTRi1UgNRCDFyPlBrJ1BdSxr7KowkaJUhcvvfhwzRjEF2FccleaXXr9U/SUpSU1lpBhmSMEOge
Fb3LXNAxD2JWP6q/IjEnnNtIOjOscDieqYZ8Apkij9M0EVOMWKGX2Ck0rPr3C5FqgcG07dE6qyjz
d0WxHD50AYQc+P0Q266tZ52+sxeZDTmvYN+YjBMh16OqY8NtOKyKPZ8ZHo/RiN4mzweLCUvYnXON
8bGyXrBxtY118AyYK+e2RhYT9FGSFKyoDfubgiluJE1iTN+pz8FacZzsbhblmyL09+ttJPGsI+wI
HkY4a6ux5o02UiNzk3iT+lkvR4yRd2nmmyPNtzJ9HUWm2MDr9VYdN9YoVWcYtHp67FP1Y6nA24R2
/52eWESNwxdXpGZ7mV+WnhwYRSekv1ZzJcKHSzCthu+dzR4e+4QQTDx+BIswnN6BgXa7GL6mFezc
PsmKWy7TN3DuCtLeFACIsRVaPp2YEmR/dDGkYdFebNWKnOccayBwIJZ95YiJJ5HZr723O01JBAOM
M20rhJg82F30ywF6MpJSo3M0xL/llMDh9S0ICszNko2W4Vg3C7Q/sCgKMrBZJg2j6VJ9bspH+Gu8
FNIzlb0dqjqFhOqhjRSdMAZSKBqi5WWDvQmw3WNY6oQxIx8K3WL+jfNh/ORmg1A8bcO/k5w8+2Pj
SxywTaItj+SyA9Ib/muzfaaVR1ZYdGA8/Hb4CYnKup6qmHRQgh+lF1w0jKS1XYd6+ORF8xdr1J+c
e2cUas/p5KMGZjZmtBtQoKUk6IN5x7KNB5CUcveCxv1z/JZyACT+Ub2a8hjK1Mw0trGBBZgMGOhz
jVdDmBc4UzA+0rH/nYDiUzFarJY72p5+/UYgJ9yiL2M5cNuUZXTlIFZoIfFiZaQVg2QJV3MEaxYv
V7ThpLO+GKJSW6X+7QUDmf1DD9FMMpFbAxRwZdN+PQyJaYYoLvpiLcSDS28MtkxFnLOEwoSSvJw8
bR91jrclJcAO2nw0+aDQCOsxgPARDrhNrSvEwK8oOAX4mb52WGu0U6Wc4i+f8yHBICjXzLId+cXk
4GHs4P+HvrRjyMRShWsTrllo5+oARWaoPdECbeLLVLFLD+yvYT9CAQ4NGmOssaBhkYeOGQzgdIYl
fC32VFf2WaZFGudJ/qSBOj43SsmUKi33OWuWicADR0tTRmkoOxxwg2Zm7O0FalqQ1jIJeLumUpRp
7esjYqH6N/MPPjJMpvXVAQZz0xPwIXlTlN/u1b9MeQadvuaEdfSOHAXiusihqgCYsDrqo20mFUdE
YoW7sDQDPAqmSmqVwWiHve3Kg2VwANd+5FfnnkOcxRA4xjg3oYSbFCzpUkiANNDT3MXx/GLDINpy
HyvPFqyua1UMVmzHJaQ6KNYW+/8bDjzTt3+FeShQQ9zvvW3uB2AgFrTCUUotS32ucd4HT+4nAKHa
lGDVskH4dURuoHJH2MKNkMUJK5YL67rJODvL3nLWECA4Lu4e9ggK9aGzXAJL5Vr30k6g2FB0wITk
ZyNUaPD2pDFv8omdUxUutbCmTJrxtHfdrF6SGkfQ/8qMc+Do57xJ9w1q5iIPA5g7BYROOFNuj851
dnLWH5dLGJGXusjH+j6+KqIyXFXroMlca9xu2CF4DN1PBkjDyMWdp4E26JSHPMOtJ3b5PkPPDdGI
xIfLW67JXknPOroPfyKEu5RVn5IU+ePYPoS8LaclJYVbYW+rM1GHmEm1ssce/TtUK0OoT6sfDM+2
/PTTMkea1iDK+IChrJ/zjcw0H8DzPSXe1UOXXs9rOUG7siNFDvWiL+lGUkI810uPd9iwTEHZcde+
aFLSsXTwTP+pplVEJ8BRnRd5g2wtsukIOiEzMtziUK5MabTd6aH456D/czmSAi8T6sgu6A7BgyxL
cyooEm7Y70hGs21oNf/xm0taa9RBpI+FOQCL+UDg/2AgWno1IAJigfPV4olk+qf7voksdX+K3dGH
A/dE4Rm9bg7fLhuS6i5MLXZEjoACzuFHhQPbS6AB6p/P8gjW44Dvr5hxJd73FEUC8vqSFe8tPSgu
flEhlNySCO+YfikvzPTpcxQ/VSEJxBucAPE4w3j6NhFV3wNP40iwuOnlW1havN6lfb85Agl/Z6Xb
5FiI5u4If4q8w6EXcm/fVoIfkSpKfW0OAHjwKuZxE+h7zFp0L/FS3+mHek//eopCyGdDi5s0dFSK
DY64ENeqZRguSQWwgXyulk1b+Twqx0PALLkqfznkS4fAFk8uH6kLcFQ64B6pno80aS7tN5vW4gLb
c6xxliAYOGJQWXTEuYF3mgt2VuV/VpmAJ8zN0VM9XzRTENjN4RUHv/xuuZ7AfKhQ8h6VsRyO0FKp
zpUUpKnAxD8Hb4DGRAigwPnOz8JYvtnmg1vSVftSGvLpTh8HW+q6NwztAcbtl9nQpyrcxgX+xvQ8
CtdSJarMK97cje8yldFIc3tTJhn8fxFDnakfDucIQuLdc12w8LRLT/wCf0ussvIjO8VidSOwGyI/
oMIxnS5mR1traQn6VGzVXUArTywIAfDWODIDsKuQELNOo9wGqtPoC5D7VD3EyWdP320j04ruH5Lg
QcaMU5/1W/htJSOzcS5cgKNQ2EVkM4ywEJOi8TkJLhy3CaxW6hc3tRtSWYajoZLRKNG0X4atQvum
vJuBj/6EB00AUDN4eExN5PunInjhD/5OCodZMUyHk8MVyJ0QGy/Ny+NVCm8SfWYBOSiHPpUb6D8w
Zi3dz+yq1HZNEicPLe55XbT9+ZwBW+oEe8a2dlCL6NoDE6MBu7ccnC1QmLYj6vUR8P1GBwVrH7Js
a/DIP8QVEsOu9MJSlDKw9KG5wj0PRg7FgDgoiFRpWXYbIt5UxTIT8BavDvqjZAy0m/YHl5oNK9nn
pLkWZonX4HlXtyr0R/OAo08V1+Lgd0g8Dtn47D6AVzW06N82ARHo4D/rIKdpbg6i3NhpPIs5DwhY
69/2rrqhlUSU7XUET0X8Wf/zJN7Tf7bKgIv5FggoSOB+LSvUOOMba2TOe8beFHierwgmzqRcGOf0
IZYCv9dJQItfBXIGmEo+ybFEZ1y1RXxY1SdrhWpYUqhGa2om9+HLJlr8bzS/k3FpnkTGOnckrS8B
wkkqeTuQtcw/iMB3xUQQ+gCpiN/BQ0in5YwfXx0CmaBCFUtPyjjFXjam0xHfKIbqK/8zHIMWWTF/
CC2bUYxtZ9PJ2fD87j0fJuroLsl6tts1jsUzj4cJX9l5wQYm1RWPEm2eg8gABMvfIkmn7EpSMjBU
A4s1iZdRcNcUf4idCbupFB+K8GMaNBbxfNTeRvrBD4QRoqW20XWwfS414jd7p1f1coRCHnltzNwZ
fnJ8II3sUYs0x2QylFiFMeISHtxoUf1US4IPZvL/MMLKRUUWCCV50ka7vr8K+Fnhdoy00dG1sFiT
extyyb+3m525EDBs+WpCbncmXsmgAUvBsx7LyiCVsCHSzRzvItCMIhZPRaasMqrWiOD8NpbOYpCf
FFFYe+8uDEH6WWPSdkRwZAtuVdzTaKAQpY29KjLqqD3bPa1MQU6rKu9F659kIulomC7h7LXuU+Uq
IG1d9+KqvZY/H4bm5R8ZQQQbWD+uX47Wylab08GPQGAoVJIfPGevtWqb7gVtJriWwJfWgzpnQpbb
V3qgNgAxzScqRiONcg8Qzc0dPZDQEn8ZbZGXxQ/tNsdw+J3Am3wHOUI0UH4N10wQnpawoyDL2yy8
nVzpmJ3knBrOYgiRH5wp+eA6OWuxk9okr0Fi7LJFoGdp4O/8mN8eIvda1WAppU+HcjXS16OkuGbD
+6u4K2GhLhDgRlWkO+gK56qtlIDZFkV9UVFTaUm0nSo22OwQAsTzNo0foSILygf5H20m2tFxFHzj
nHTRRxiNBn9wH6vdeWxpWOCflSdNri14Qu1fFCVIopX7MSd4wDBJ/ZFh+ACxkHMfhlpk34HWW36z
bD1cA9ruIVvFsLqoBcpK9p9PBovN+GjXOryJilapydmW2cx8eW5QjxOjvrgsci5Y9FHCDhxew41d
r3p2ZwWQhOsARhBTMivM/rSeCZV6qKhSv2V7n//WrI3TERQWC+V+CRSZasH67llslzfMbQPja4HH
23ipfLY2/V6WRjFAKRIrDXrnEHvLt+kKwLgZ9pHtEhOt77bDtnn9Nslxwj6slgU0BUUZ8DXBF39w
TLutmL2SxjQVcSENQdniy63svEOi/EE36wqwzERN5zof7BJgMK5BSvlON0IqvGCOATYmy79TTxx1
xNsozH+PyNJgEShX2NPEt2UVO7/E+seoxHetoU75vwtGqFbcX9XY/W+ozOA//b5LveVDd7URfECN
lyh30Djxp4g9V068Vt1fF/izq4UMDs6JlqhARv5jVDOwIDtRlJ0K0pAn5tNzwUokyjXv7t9bMP0F
FPeYfOHQAV4NA/y+V1gceznJcpLWxEvRGFH/Zb4/7aDgfxEPVhAhHOq4HwFtHsn2p/svbElsw34I
N3Ptm6Vsep09OJP/sykJkVB9SyI34lDOESG1C/3fWmY/Ho7MCkxfafw1RwbtX8HXJ7kGI9uhJMcW
HQ8Fhv3//RCt4Y6vq3gCdaNrh+inkzeuc7iigrXkp+/Wc7kMOyjUJm1VOHKXp/1/wDZbFrLl6C+Y
XaS/Dolxp1KNLPXqoRDhDeG1aTJqxpIvhYlc13xuprlu4J2/uq9geRIx7ypaT76aNVZIpNjrbYFi
YwoGaJW6eEmZTD0sgdaI09+DnFZjWSI40jiOU2mU2RA69CgQICJBJIszFzVjV8kG3FBlP7vmqAO6
HtXFw5DnvaU5QgXacIMBACQSIDEahZ30U64dT1hiHIk0Z1+IJBHXXAzwUfLbQASAjANFQRYpoIcC
Y2pgubslE6xpw80qYyguQTE7AxjbxdLCSijl1LKA0DjOJSEsgzuWyQoI5XQ2VQPTuKXxry1u8OMy
hKhUCRSMA+moYJ3J7N/kKxt5K5+ie0dF1SMMXluklMkgv1+uG0MNOAual4y8cg8BH4ESPyvTcmdh
U6A4L22ZZzLOJ4uH2MffiIYDP2KVQ4cI78xlG6yl/3Lmbss5xRlsnqSYUiMI1AWGUVIqYmlZh6JI
UT0bOrt9HFDjbz0LTKd9zdaYxdf6AJ4u7jOzFsQcKT+vDxMcjx5Ulo6PviUgb+UE5g0euRpxYWQs
b+2qL07Gr7eavmteVkw2Ihk4ZAVrKfyh9FUbQCs+AlON+r7QJwTD+ex2P390g/29Dlpd5/Actxj/
SyPHqAAEGpRgJ8nKTis+euJhatm0UberVlOkSSFuRmAoYN/8nojvnM5uOlruN+WC127bHpU94hvE
L6mkhWp8OGgZQjaryxWUTs7Qbf1MLIl0IUxV3LkxmBIRvkxYLhRboKK8t3pvJ9QGer3c8Z8GUi1g
WZXC6UklZGTGKb7Qevl1CwqwflLfjj+mcnPxKR+dpf8RnGYEhtQecf4KADeJ5nofi4+nyijTlwJL
/JUP2PNh2epqLktxNfyYKwuG/6NMQ6jO1w0L0n8DmvTWeT0pFArjh/kJBiIw7TjAfIHp3NUxao4s
B7tiSzKD6GVyjDuBnIJAcKayHUAoF7w3O1OIt3oKeEg3XMq5y/si5FdTtM7XNyLfypcDmdi/GOLD
DhOaaPmVzgPxPGm3xRhzWWFpTCz+p5ob1/IO8NAJtRT+1l/8AQV5spZwapa3SgDQSmJ8WUWX6Zdz
87583PqvSdjNU/nXoUtf+bfAIb8BTbCAwyiJwzQwrNYNOnsXEvvuPJ/eIYfEJx1Qi7lIgeuuOwwA
iWQHLpGJ60pOpe8V/Qbv2LWyxsdK7rxPWad7PV9F3+JxkFnK0u+skK+ZMSVY03s/+s4ilTD5nby8
MZfUG4bxgCzRf0ev0vz2ocifJt+fuiridLOoXg+95hA2GtmM1nUbHvugTnJfG6eszKzkiJOenowN
F77uvzaHQWxlUd4U8rUlJeDur+HCmCk4LFNtgWnskuCN8JEiYBGPMTTp3eqGIESpFSSzkl1NDH4N
UrdJ5b97LvgraJiwD8zOmZR6l+NqvUO02KWF6r48RyHpMLg9SYt5Ef0uLvQmV4dk3wNF8I0xDsEi
MH09hC555Yuukks8nUrkJs4OihY7tsniQ7f4J08iWlqqhc0sYJHFl+LoitIJJ63sNrOVJxjNcC2f
dPSd5DNXlA+TcHMV6BFpMvS3puQwBf0s/SHpLGVYswsrg20odUeZG2tX8rkxosE4eSnABw2XBxdo
BpDtt3Y5PmEQZyn/6KCfEw5Ayy813q80Zf9Hd1Gp3UvaiiTUpha1QuDx2zqEGl1BYEkapPkTnTfo
flLswJTCO12K6QGqzJ7zjUNOejKBRUFqozN8vKrocwyYiVt+ucVFP3aWumRqC6borJkmH+ZAna74
1t0cO7vVDI2uXvvpeOowsdxc3TLtdwWn87+zCjkhspxczPIzwnSV2SAQE11FCLoI4ZLYXP+nVxMx
XhGU/qm81gc5fBUUb/mAp43dvwZRIltOcDeG6Db8NHfK3MNyc88PSXeWgn+MddwmZMJyUpdNuqIa
nWYFWguzsbdK2EyxEhTsPQm02+/hoI05aOTRLfqz8iVWjxco5T/1unz3jK9bkQs6L53f2GEZT0hg
/dvVPGQXDWOVPoVQrba3KyqyK0DNSnaYHqQ1FKv8qoKqpS1aj30hrLZbUPO/fUwcl/fIp31sgXbI
M96Ssp1HljG2iJBVOzpkY1UDukwFjwGXW9fS53/cV7rSQVtk7xY6G2RvAcYVVHOdO2K1Y4ygNXN7
PuP1almrGXakDsc43pXAtwoOU+zQmsIOoisoHSi3Y7z/Apoya4vRJz5ulKAXLUfqSIhadjrlIP+b
+jBivKrmZlnjxPNSK66eXEA1kwbryMLvsnrZpLKoceAG5lxfC56W133fZx/QCEZV2Y/AOMZRFNL0
BQX7EedG2KNtbv/YOjjkuV+zK2YKZlnPPnNw2F3PFMspeMuEK/cp4pNsHeoKYo+PffmQB6oZG6ZK
1Jvii4WuQ48NrYjZkgkpfYJmcCmpw1iIIrUBFHULVcbRLYywG+7IToqXxovk9zBw2wCiNscy7g+D
W3xnKRHDwYbWFNOoKypxECpnauRLUseuQtxve8FVJBjLvfU8znfrXBr2s188f7EiSrd+H6eZrWvq
YhSliKQ4puvmKCOMFS4t2J6IC8bZsNeSzoMW/0UT6Zdi8elEx77G9QNiFCI/oQvPOtmUuDqSWZ5G
skktg4DB+NS+15hYf7jKO+sGYwFBvhPPYm1KzD2vPrC6fauxMSMdrcYXEUCOFcZr0QHL1hUL6Omu
4exYkNmVjfUZJ25jNx2NArSSpyIssPSrsDkBoShxubqSMtXzRZdICN330OQ/649w6Llc8AnkiuGH
+M4h0KHR31yDbCunryKOI5haejxWJCowhiiVi4vgK6yIYmG0S8DtSpjx6SGCkD0yOL8MG5NwDQEq
zUa3QK3cbA4CVQP3gVwBvMbmNZoAcAAcrFtvpSEJCAuCcd898sMgbqw8DPtDx+Doatqu+OF7O72N
x86290NvfrOmXJJDZKX0mkn+Kj8gDzXqpnnskzub2O1+OvmeRspyPoZVUVFNRlY1sbnFyHXXoKLa
5EIVfZvcITXAbRJP0qdCuAkbK14+d1MLC7ircaVKToosrLyKUekPiVw/9QcSXoePFu2YCF8SvCQ+
jhY1fQPvpvZzdjXf2Hu9osv6+Kcyk3WPZTbYo+MpWOrKxCEWphyhjmp5c6dqDKaZjJLJmsbeqgBi
JXCr4/3nV0r/++YF5OAjAlu9GKM+pI+ELwNup+DbZZUy1uieCmHf/nI/v1ggH2PgpT00YDUa67eP
gOGvwKFhi5zqWUjBIq33oMq2SOkuZ16Ed6tQ+rh2fkqGGM1DLYFVvhmtb9HC7C/qa8kvIPoP8Qem
vAmxKoXGtqEkZx+zZneKemcGRlxiahYVnmyZNk6Q8FZCZmzfgKAB1ExO5CiyGbWbIy00c559lXoF
sQmPzTAeo0Kq03St7RaoX4PTGpmP+BupwlD3JWpTBYtyP1HAGaqB4zcK6Bp0tjG9H+099jXnfbRX
fnWxYqYh4fEcMgRdu65fz9yp+IXHBy0Q9X4S7cBpxLIV9qc5Z8GRkhEJZK7aGpR0NozvvoUc0giN
M0chjG+wpL/ej/8OAKGIPX+QRlfYM2vbk2PM4e9ots02vQLA/tQZTXRX0rLrZAk9aa+CmL3fPZkS
tJsscKnDTopfHdLdwsnVioBKMWY9DDR5+3JFfX1bS1PymuSIwaacpoil7eOqIPKEB7QUrvdtQi4M
YL39AvsR+i5dp+zYaXv2YFcxErKVwAFcXaSp+KDcVv5FGecuVBR/ubh9BzfpxToFVZhTe72SCdEy
l4eY9V+3Q6bUtTIGOh7F/cNqLxoxvEVA9BkH63S9RVurJpi3z0F34wyMvrlSTjDsZ2PhvnkubRWE
A3eN8KvThjJVa3zxu2tifzlxspzrvcCS3irIBOEgKNy9FLSwMZgqo5s8XAPitru6LmdFqP1E9Jy6
Kl+jsp56d/vn/8jzkziGquZVhOVcPXAjAiy3XO5klLkwwSy4nTGRz4lN3yeBw+D8s387mFBobG0s
nXFb0Hp0THF8ZFk4m59q9wi6O7cxFXatWsMDZCOe7dcsXNiH5WaLtyOR/5R3H6Wo8FYJgHiGPMJh
PqM1heutLllLQnEZDTV+Sxo1CjoQwm/Qb/11aLBjV9K5tLauQb5z2dBUuwVOMI/Erf+7h4vsDILp
k0r5O+4RC9+480HHepOXASlQp2fqvRsp9eQCS1iC1Sja8IhEvQxKfXPMAjB6okZTj84gAtqxeSxq
hMBM7i6Uw/+l0y1ZpJPDmFWREnvtdPj0xdHmzaiSRj1nkYKMbEW6i+KbnOfRJtf6R3k9RXRpv/+L
sJL/dpQ5tv7QiznxSiQfRZGl9DyeruQHInkROCpPk49FpwfQ2O5G7w35iYJHRFPPs4ju2zxkgRLp
zyJhvoQVIsPKR+Tvez3y9rGntEXFbwrPzQsYZukHEF0p5ers485abxNo6RuYFQY4DyoH97AutEy9
JApgBWgMxArPVk1t27f/HF5jCHlOwRCnEDGTWWTdxba2gUVD/4aQRLIQSME/W0QvwuT8jqVyXfIe
mto3ZFr9eYt3KhmJKCMnBVyqf+s3BitogtMFijmyK8qAcB62mZc4hOxJBKFVRPP3qowC378J7l2R
oiqi+wWf9V9dyLxJlysysv9Nq3hIVX1OEFqlCs0ZSDDcM7gAEJwl/2SCWz78A8fo94KbgS+IPwU+
+60hFowIHwH4KSvhewxGcjYSWpPSx87078vx4VlRNPTdANP0IdWfp4jKyQcFCqItP633ymTZg3UG
yBn2xQq/Zu70/dyMMcYWMbDphNFzANe2kzhrFt2arjDKZHvSr5oHwuU8ycDIOtx+3PbJIBZlH9TZ
2ScWMHJEsafqsuMy94OOCLpFs7ZEDDVKxxnipR6fOQYnElFoD9P/fdYJmlPwDkHFzbuULGNAHKG1
rX/7R4oK99jmETRh6HINt3+bqYwSFWbWctm95uFNDbPogH3sJfe2KVE0wtOuYDOpdWwvC8JEB3XX
R65tTXy5HczOR9H1i/bqYmDdjL35ETu6/kL3BHX/7x74jAbYmMFAaUbhbWwlDLVRMMs0DIfKOxTS
MdGY6MI5+xjqsa4/SgzXS6qgfbsfLm2fJzDZQYbPDW2pHncdxq0RfLyrrdNKmcZIQE4SxQnHnC2v
WQvhR5l12B1YXpVidBuOkbsmN6ACKjtVL94fKwUECXDpHIKL14MzHrfj81J7/sKmr7bauH5566nH
8+Mwoqa7fN30nXywta+8950etn6WKlhhKce+8hYI31sIB3V9zfhlUB8hSrLSIs/YT2x7ouoAYdLk
a0kOMyJwqaI14HqPjlkWE8inUPRAgSlWUDTD/2O5uyZ1BIp+JLYhWixrL/KowLFHrEgQOXmLhFct
4M9kasBBTfblcomHQqU+6ALDtl8QHMwMz7ZmJlG6mVUfnYenX9ipdcNGFFGXkwsnybQomexHkKox
9XYU4jLeD+f0ZiSK5umjO0Z7qBd3wK5rXTdMHOVPDmR20BP+sokkjYeAmLXWlHAn1EA+HvwttNFm
jOH3EOmaBz6YQ0Hjv5pyL1Y8fjqdZmg/2y2WAGjR2K0XybmkT4D5MnaeJ7gSLBjk+DFGWdvSHCwR
FPvxi4QJSHp8EA8b0FUBGAzFbP4rl6EOa0gspXAo5uAZYdC0Rwvy1iSSO3vpP9yb8wT/SiANS9Qq
H+rvQpUSkAPurjqZlcsfKVJGnIAU+oB70m3NaqTifun076n51B0LHqGJcHFgJlXMrqYm2A4qKVQV
Dz52uR9C6/zWBGFh8aQJmDzPM9VjQPLaEw6zrqzQwZstBtSH8cuRnc98Z1FxMvaZwpln/uUOolWa
23b2o9SpeXrDE64Ed/8nzeDWRNIPuVrYFS4N1KtaWi1VAJ8XzbeV2BG2j2uHhvOZNo1FSN3cgryz
9YSiKC+Y6iFjw5ScR21NjvoONFCs68Dvgdrh3/priQe1xqEljiXsA3kHEBwMA3O5xaV09T+2S2SR
2I9Rr5E2zaH27RZR0hgbG/4BWc3m31Z50rSVp5S0Eh2R1pN50bzDdFNZOt0Gi/rHaSQW5JP+DN46
QJAuj4sWEFIW7aoKtXIuycbavskhOgjhNLT7KmTdDyztWLMbBCSsozKsNu9nRUtpEEx+dp+s0GsI
RvDkuHGaLh9/xG3wcDqvEHKGbl5uZ3DVLnDoYwmGgqL5/k7Nzha5+jxL9La6e36wYHrYloqMoQM7
Zin3Cp+rlPXKUKXiBjtWoPyzrUg6BFR5uE17YP0BXPTReEX0tJpXlvWV05KmVjskZ6jN35WjL9OG
3vLI9lAO9oA2h1pl5x+EFhiU2zXkcUnXbo5mU6yXd44m2PGK33S3auWelsjrL8rdDGWQHAtmFHFZ
W73PBdtsP9XDTXo+X7yDmqzYnWM3VBVkXE6DzOTaZLtEK9HT7S2mNGFQb+cuFh6KjJn1kmX2+dIP
MuXj90QTa/I1dd6UvaE6yDKzeWkum6Gc9ARBOrY98xfkVLRzhIOYDNBGEZv8OLPO+gyY2dWmjJNq
nAs7RRLghSx2fDnF6+g1t9Ya4OyLq5nUQOXjA18hWWZ1zyHH4w6Ut2ThYW9EvEM1LcCstMe1iMc/
TPKxAMv9sFH2PrHg3eeJ5jIII/3fq/20lPgbK7NjbPZhcLSANb8Vz+cQRmyEMdZCb9sxVScF5S7I
XBfzGXKeNIWBcknffi+o7qmRxZJJVFhTFcmoPLmDFffNxQQK09LvCXNGQ+UbUyiIWentHlyN/dsR
xz5Ph27OBrjC5inEegJcHO/ecY2qo1gh7ixv76Q6iN0whpHihGod8G3QkPlncxGgSjhYNN8ANllc
dP5bdow/CD1hv712srbAeCR3GncAtNp9TkVucKJtH+CorBs3ixWyC1lYPxduuTolpaYSBr3WWYbR
W7Y68SPJFihCcvyTe4HowEmIfJG+bAroeHsmy5bDK98ojWfiSa3Gz9FgMeZadv5ly8rWSyUMW8HO
DENnuezW/7+0thnWethglHgQDQZ/w7/zHVb3RMN/PHV38IfHh+pr129BFnZG31zMoAi4y6r90zE4
2hs7Su1jkxcObUnFJOg5xFtm94pOIm/hBnAKsMPnOJ6s5XIjHgRiXmuP6S79Xf2gpEUSsmoCy6Xf
D8ypwGqmhqsF8a8ijtXXQhcGAZO/yYwmbzddPqGGwfwSF9UfhrVUjmFaNqOQRUEnQZnCNikAnjEW
Y5l2NPx3NI354364kT47NDZviAKvBdRaCHpHEfsJSAwQ5XcZGjp03Vi15z2MH6c/DggJ9fxeIlWC
3aPQkRbQ7B9OcYxW8nSfJtkGaEjohAHF0oad5Y4bbZlPcYRvI3BYLXAkMGvRdtpOqBbyAerV70Z6
8Yo7nlYJ6vdzpV5XaO4TBhB8YGSfrrE/dsV/LPl1S5GLPy63THaet914YH6ttDoKNDqu6AZCedIt
VaDPhmoExIwJZGr5egRyzSFefKPhIkz45j7oRp95jwHvm/hTZ/9Eb1tm3huhCuwVB3lMNZ1qdamJ
9Nxd5dtw6LdFyeol6JT6PxPKw9hDqT9aUZ6cbiLs/Qo4Tl8cY4D1zUMqP9k+DYGJ+QJQSRA/jC/9
Y3p6heQTsDp3zy9zOIJUMO7FD2A/CLEeEJV9VIv8DKxDio1GO95zz5MX9W+FB5pQ8I5TW2WoPkQr
kQCQzR2ZFSftxQo132Xq7Q9WfnDLiMb0oIdWbXZ7vuCmfF3+NDldiHmdZXlCeTukCO5Tyc1SAC5j
xDwDqjFHGhRsXNyuAFlDnPsl32qZhWRrN9xoMu85dI+viVJSxnSi0fgvTO/GL9eXqt0nvekPkqcO
kuqf3EE3aqAUNNlCPfd7jnbnUTmRutDqqS73TD1151mPjZkQpdMTqL1TK/MJ1Crg7uee275dxzIM
Oh36nNQSxRsuAlW6qJaMF2T1Vit6y8eZF4UHB0gzi19uiQpxMQ8ItzhZp3tOAI45SbBl3Xs/2pc9
DeRRRMlVe64q9Xe7JwJhH3BOrkXa12sOn5Ovl6WLA+258gdev7rmw9eL5vo6szqdihMqvims+EVI
MUbfbe6Q2UTVs0JFVt0u0K12YczH/KhmNjNT4FDLiQIpKNDRoDKDxXhdX3GppMp8Lq/SD7S5gNHY
yZhfYeX04gdWQFx8FeChyMnOgoOnEA76aBoWJy4cqQdd7WqCvoGxwIXWlLNxpQ9fLqJmwOZJkdiU
o4tTcn399iWTtMCvL+G9vLJSHBg+PHVqE5vdORUINTxsLjAd5vrUm/uviQ1kbRzyWDI05dzN0PUr
iMK/nttIQyUCNfGB03XHKkSQlxq1OHRdvx6roFbe3qu+VQILoPh9EqrkH82NJOGD0GqWEA+kzQwN
6CqlHt8/c8QndkKo4O/DRc56QuiJiCudS+Krzc+K9atIpmiIoqgv/7bqqayA+D4xSN8ev4jF0iNY
ClnQYbbzLV1WgBNM8lCIAS1umpIvmpuE4OFfmyyXUx5Ckv62DurO8sEDjTUvvOHYXIhROBNOWRXZ
XLmpWh/kM3259zU+434X4Qts1XaMSwCMU+07Id6u93F3EsqAxJOEX2NO/pCmWCXUQtPNxVfPIME7
hMpi90TEctCAnbWp6zjHj5/iMaSahsCXaH38USWswxHtKn2die8kvVjEq7ea+IlREa3RJm2G+xD+
Zt7IEQPWliKG508+mFjlLoxWTcAz8eQZllllIsJf43UQRHkTSxwU1a4TTZbROsY35eyljg7+Tsvf
UECtBZ6ICp/TFcaihvS5p0C8aZF2lNmDO/Heer+pTiLWecIiHniUzl/BhWsfIxlcSbSOm17GDXX7
oDiYuuyDueIE8ZwCLh+m6xU/bjysnUGOxo7hE8g7sTzxnaxJcSdCItGNDqIouXdzcx+Ad6KHxvP+
tD/ZO424jKFE1igifKSkDndaj4ZIMvf+TiwM4/WWQ+In2uHoMYxnRuCqFrJmwJoQ6QQiwqAPUoQV
zFAaDFMZ+UcP8xiwr3WNYrbeSRqUZLeRAXeuSxcXDb/DuqI9OpmkepDEAxhOwc4WfJckLLd5nWTp
VdGCSz4iuKbjluDyrFZcVvE5kGgtwaWxjUlgyUct9pvQ4Z5WHkMYcKjcG7UpugQr5xK9kPoJcibi
hLioz2Yu0QVzqVZO68mImdpSLod/2lO9M5nN7861ShIg5pme3pCEWFrczGp6QxIjrcQ6MS3DagRo
OIMhoWIXojHLV0PSSo45rtfPiOyosIw0IQBtoiNw11DCTR8QoqrLwlLIJ3Tum/oVBamxW6ee2+e+
WbxYNeL6Mo8h4WhXwffa6DNyfPFIzZLU6EDqzbo5il9UoQN6KUGMnZIgxHpbcAfwzsYKbGet8kCL
IoH+gwqusVS691wRts24pig0g/DjYuVjmi/l2xPfoDl3y2UtJwMQgDdLkM2CvpxkECVL15IJfEjc
CFHURfnxm3H2xsJXO2BR96RHfW01RtlzpcXqf/34s/orXbOdIgpl7sZj6A+CPtywoHbRR2xG3wVE
Aab4tOtDm61ziM5UZ9Bct7YM3qYHErzmYAnYAQKxd+BUwIab0LKvHRSUKRA2OYr3pUvat//npJjI
DbuD4BNakrp4tfyX0PaGXNFX21p5VQoDrtvDgC4AK36dMDyogu+wmO7KKUT6ypRSeLfsGdeaIYjG
X0Qt073UVL0G7uKbvVKHTPYN6sjJ29g/c+G85l56Mzhj1sPIYyl8wf6LOwuRzzQINVglWzITaSs7
LYhAQh6sZcxtDV8yENhnaRAGU92bbFxtyRbC0kctreVWfKN5erDknnNVXhqrWo9YXiZncl95dKRi
X0r1DmmKYk5naZWpxiAmDGPJk2RKF5vGb7xZ1ZP7WD10OJtJR89NEGpY5xZNg1gYN5PVyqPsg29U
wodJIeUNhUNaKzxqruSAYfgF6HOgjRVEIyRbTdYcUPfG93E23Wl/i1Jm3LPUUVsQH1xVhhFB+Kdh
A0AdTyMvsoV3JQCnwSnQZVdQ/KzvFmomAcp8uUPqkOXkUtnl3QPXgDCTDR6IkczyzU71oONJT9jY
RgBTh532D17EhnMtKbQZNRsO/cWxH3nQ0hqn5ylHfmG6+oO1Q+ZKbziHYgo038zUaq8RmsqV3kXs
Ob5HKCtvSRPliG8/o+ybrU2PbNi1+/9hBaEQcsRXQ78acrjc1+p5CfT2tPyQnEsl9noaJEu5xP95
idLpessHTPpjqZCE7w4EFK/NijwX8KtL18WcpsUKR3wOvPteClJDbZjbKy8nmM5KiO7xNB2X5kLD
OrpQ66XcZ9hfndX6bSQVWk1gy5KOjGjG5jQvavU7A5PqCGmfD9MmKJikLIPJR/KhBRDDMQaieuNy
6LmhDcRc9/ozC4/o/686V/NVNSmil7P51DOc7l+OLPk1hTs8ZeKqacsRR/jWNzhBKA/p7/7YLtr4
POiX3j0NtIHJvJRV3mxkCul7UwN+OqUZ3UyLayBf9bVlsSA/KFflwkfwG64+m1+3gAq3By6foxGK
Qb/8SX4sj55sSV0k6BeX4cCWiuov5eMojcvHGuZhW+pOd+Vouc4GHN2I9562dDpY551L+wV4o2IH
IykZaa06ln3tBoor6KiTsVv/yvj8Q9ijNAVn7Y8TJOJvgxQ8RqeTBJxzK0djiIVie1f5y2Gtrf5Y
+vcQjdjLF9mskF2BcB8lUHbi+Id1wCvOIBWrTyfxQru0n6ZrJf3XyUCeO94D3AweL/4vIn5a159R
AhfkC01LK3WUomZys3zG08jycyvGRJtpEpBi96O4d4YWmUAkH8OPMk0KN6ICnrhjQoaGZFqEz0Xr
InoeCnz5qCg46xCWecUslV6XSPkr9S2o9adZFXRg4Vg/d1QExWEroH+7Z2Jd7GE/zyaJbFiiSo9y
6YuAOKI8W5sazNtqqcurDCvJrrSHYk3I7yINtqCzUaixb0I74mNTrCninehU/UjBk8dpBuaVUmCK
HqKHK24PsNoBDTyqnbwAD7op8PX0btci5dm7VkF3sym0yC10J2BvakN9us09rHqCbEiEPZISnXuT
IXIp77vISqzMlpbwU+bk7XetrJysvy8zLjQJHA74xrCRDDwRmSXS8SlUUVKM3B9x3uiAwMstqtAD
qylQUW0v7fiyKMLSOQkSWehGwfWSDHbBUSbCjsYggXPbT5jhhkZInR4mdHhskzr5aBd1jPisdaKd
MBlr62b3pUenxLDVjbsXZmx2INcxCmxQ6b/OutHy9Ed6j+PzuU2rmrLw2+OWejG+jFmiKO3bXPiz
mgr7++F6Lixl5ZabwihozToiLrTWwI+IFn2s4iJd7DwSiA/6JgeRBERddShCAT497jh872kkY+hE
bjvoDDB4eufTrrxJDz2/pUdeDGbtE4q/BeDF7arxDNKYN3SmBivySRYZnNTBIKO/e90SHouhQGWH
+JYvSG0yxDoI4/yyI+rMpXz7ulUwcOtfErqy3w3oZguBCNFM4UMaDXfOhnfWJhFRN5XCdBvIVXhh
NpEIgolvwPyjP6hI/C6n1eK7DV5UrwZkv8P1PdSyy9iVpnoXNuhct6fVNox5nncgzVvVzaC0Flua
hucQJj7SRHrp9CiSWZM3HMp0YBxISXoWb5Opg7RUoiRkFqbfF5eoqW4OTUP8m4+x1Uk7c3CZGpRk
heRMeRW19NzoBIvIhN2uzD5eLQIZ2dLnaAl+f4N2Hya+yZ+Vwgki2qDMx6LpMPGbqht1rufxwzkR
G4EbwydHw9/JZuOCfYQZTn3ZdnooYseM9Xmpp+2uk2F9GZl+1YH5ju1NX1EJ0VUI95pNcFV7Z4Tm
iEm1HM+kUbo5og5nh8L0OKq0Ae6+YTb65UNxlqqkSJK+6IJhhSdnVXtKdQk/kOnUGTjQvUXw5z9J
QAAM7aZRPYluoLBC/JLs10q8M+uTBhqjHIROlKkFUYcc/uRkqe0MAnw03Fghit8BTCUpaqTtPazM
MhqM+6Qwfbg6cGuZr1oGcHGf1tYL8eHFFH+u9VjfoY9owzLQTlR1RyVpCzlGXV1ejsIPsZsCQB1M
8Da3kL7U+pXt0eFLR3qy437C6gegi4cqmEuJ2BT07gfPVQM3kMgRFmBSOoFMSIGEx76IhQcWjU7K
ZUZdSs/LDo0OD83Qda5da6HoAEfcZOXL0lDcCNNHYGhdqpHxmcJFrpFMLBG7QHneQFz56PykPSeX
fXxqNjhPg0SbP7V7bJAFjWRhmC2AiefWXDjqRx/oHy8/33ZbJZDWQ+LCl6zevg6DhqIBwK0FeRjs
rzSoAncVOzzJx31jcH73chgNi2SU+OThi6GFaLYYIdAWzSLUGSokHT+Wff1eVTO3p7sw+6YbXcrc
GrW34lYdGDqMXuV4heanFTCNpl29RsJ8J/Pi+oldy8tPNnKN/p/s2hEzM2K8dvkZIJusnaIw4A7w
0ryqr8UqN9ASsq/ANT/fQk1XQ71aO76N4gguX9nefAyXZmkZsO9zdD+Kvyy1VsPI0BQZgIOSOvrW
OgIQ4f4I5uAq1ZAohmODfCxuHpHcvW5Egh9xTFLrlywPSWk/W8TQCqDinjRPfUqtL2we4dp5rcbV
z0O13U5ExJPmQKzo3KIg6MlGJHMfmU28Fl3KRf6JhmOEHJSUjBh7ElKlArij7Z6Ei6obKCkzYHDd
SOIOrpoxCkgBeUYHPq2mntJYF2behyYkDNnM2GywbPP0L/7AHaae9Q+gLvA11IerpqXBDvsJ/8mP
9WnDiwdunBkwR1zDsOAjLrIzmyWuKdZAz8h2sJR1cDsOFt/b+SaSfwWaTzrbMgit7Jw7YG2FgkFD
SOU67AVQ20BZI+YtTKbEXwMLTmhLUeeEqBP0xpXnGyMI9OCy1x3RX8+G1+4kyMlBzojKJEljVcjW
ChHK03OBT8Aag+x0k6IeAx/Nrfm6fvgCkJut9hO2z9guTr1ikE41x0+E1kbHI+1y22FZkoPCGqBe
DKWjRnAqspQQkKqZ2SAyGuTk5W9Bw8TZ3qr23g/iQnBQw3rUDwSOKeE6S0N9Oo6FVwlqYUJYD4Si
me+7k538m6i0/oewj+s2N4dycPMTJT0rGCwJN5kHEW3ehaAC/jPN3p+RfoSd/NKQHhr22HODIKIm
GFnFR14+Jv8v7Usxii7nML3Q3O6MY8PkDbjl7glehJZ06SCsY+vn0qKPx+uu7S+iZC0lHdfYe1AI
FcariRTpVkuzIkir0V6fNeMczL3b6BWOIwMkc43eF4D9OYmdhu/t9MOw0p8ax9C4Ol41YKZ8kjRQ
0wXpaH6cNu/lUj8iZGZFqXFINN2Af+sCXSkSeVXw5vDuE6LCZ2lXkCjNvGghPfm0MDHsJBx/OlWo
/gYFKJX4RTOL7eXsM4Mgs+z+ofhWsVFovCpMVt0dfqlwXYvYW5UtHJEVfQoJ+v85Pq5QOXSEmsAB
FInFfGx7Uq8pZ8NdfVbO7q2aIhhGtumQLi/4jEjA5MZ/1OHX+CG74JMoreyw4v9AiaI0KAdUUauV
mccwsAMPEJ0itvPQVAh/vnXPntf24PMZtoxS0vn1w2JLUUmRkh0Lore9/Cude9vK18qfCEROlzsc
6ruEqWw7xXho3SKSFIiaIv9AdR0Q/XKs318SijY20MSEJPl8HR1U3AfU+hAky3mvvViSlCxhDUlK
7JaJ9cgJQt/bbA40YsCu65Ps+44Gej5WY9P+izxtbwfH4xQ690OZgQkT0auqTEH3Gq4hEUpYbs2G
rwYMT/u6GJCccbiyklrlZaWL5mXeAj3wgxlWvfrE1sJzzxehBStYQgDq7puErLvZKJDJGD008Tzw
0srBtb2iVLgv+caquFA+3kfyPOfEH+Nn4mVtUtLXBEWvuUL9l3faqYrOP1pdU77tdWe5WYjJ9AcZ
oH8CV34jwkAGasAwALf9nWGUMW7B/T2CDSqRRxbmzcpGejLj4Ba+/aIrokSUirs+brnyH260lHQh
/4jXa399C2s+rv5OkaDYC4zZrr3pKajqpGpKPtWlL7F9J4i/cxLDMAdK6rTA8W0zpLclOj/Goihh
gzViFOFvOAMjDZaSZ2qnlx3OkBraWr2QRVLsdxMNziFKGjZJ4byTAYF+Rfrn2kf8jsTJTfWcxqGk
f5IaOt8Er+hRwJGhBw3+1vJHgHr5drAkoxWtd7eA8F98VGkj3f1OMDOH1GKFlwjv5EjjfVdF3Jw2
YtRmP+zHz3OmTk7BbOr6g4bK8agelHv2VrPUY+OsUu4Ee3ZsKOS1sSCmVD1w9u5owMIQondYnK3v
w9I2KiyqW5c1TdbOdmxXBJv6EZQKeuhwx6WzenbVYzRxFXfJMiCRP1iPmshBd8yctIerIpN8oBDL
jCmftM9SvpLlcJHeA0gRTaoYU1Fj4gNmRv1jOl4LqCBrgq8xiPdc6TfYDGLKhLYyO1snfznhbXFo
dla4idGG+W5Cs5BHtVj71wMurMMmgwfJUt0BAcC+BplTKeeCTshh256GFrULtHcwoxZ3KEfWuR8o
gl10PMI8pBR87QVq8KGEw6XiCkVg9sFMmNI5dRAeUbclyuA+7NxCgybn+r851nLzoAxY811J+MNT
GkMkoy76ZNkM3290dVj9Sm0MHRJPEUYMEjbwmwz6uSlwBUI5atX8zS60oQlegyTCf/VNTUC/IlNn
YVg9GmdAc612uxAr4ugaEVyetdq/w2PHqYztnC28Eon6Wfjse9S6mEoVbfORk+/2sf7k9LlDDDuY
WpyJbzrm1oO5rejRu8onKcD0OEXmHHb9QFPf5eI8LQx97pwqk/LszJ2NR/AqUyi8rnNouAotgnH+
JvO6831tnlHIa/vlGSG8P8x8TBk4xHEj8uICSXOjJJ0RYcgE3L5l553210CvEb7DiBK49N/QQO81
n6BxPjtQ4e4SkQqsqJGI4tbwWA5yLL8Uzj4XY8NnQ/QilJ4fNtLbGGS3EbEXeGt/g+UEnDqiMGWx
/0IoizIr+QGJ3bXHUc8mkmLhYDUAxjbKNwz3a8Z3dw3GWGwepHwOuF6Y09WkNh3lOQzEEPbnCbxZ
/ojnhLzFMIc9d4dcVIF8NSr1O0LsXlBieMHQwLsJxccYOWWy6Se8ogHZOqx2/S+mPqjQnuCv7bEm
zr+BHCL0JJ+U3xvQYKt819GHSPiFSBfIdgfnTgHVkYzLLxjKvpnpJlKhlZOlhQ33CbaH365VWHM2
vMhBselt2/rXWI4VZ19XJRo0aMfNcHk78RX6xrMyD+lR3C2cNy1TccnpLnOsyRyjDfgIU+rtc8QX
rv2cmu33QbjrN/vNJYuOd83rT/Q4+fXRFaGoEv+TeRCpdmJWUHI/sO0iotgVk2II10Dxa+PTUy4i
WRy1wlA9d3he5fEgTko2Y/wI67yNw5vsokkPYF1nuL0YWAxQ9jQ5yBqJB57UkCfGp78L9lXjI7UD
qJEqYod0rZktwe0O5g8x/XsX/t5q9jcV8Qf3e5i5loYCQcfSa4obS3jVGZmXZ8erkhNOLh2/NhwL
1su3QPYmBFX4OJEur24jHAK+ruTnwJL5YwCYTlDojvGrNn1WFvS25hFO1FdsyjOCrAmXqvMljxsb
NI19c4mCyGaT8QsU3ul93wwGfY4izjnCUYv7IDIUzPgnJBVW93kSNJL1r1mEtGvJg7mDG5AmR7Xa
jqWIjgG/mR0ymCbIxbFa5o/I/zHMGSY3T+YI3kQy/N1nMVzUFh2zOO7+WRgp0l0IKrjf6E8wLR/B
gzWji0bS7vwdoyf/S1znZdUxidtw/v2bj3dPxRegevFt4oFPOoLyZnJhouX64PrFlWikTx36hNMA
pIkI+zCzQ978RR3KnjnfGJhwsKQUNWkTPQbRTz2IKvH964SDf6TjaiwVvRYtJ2/znCCDxH9z1Ej6
qZq2NTccFmqTWJw8Hb+tH77K02hZ6l4qZbosch64arli2ve3xiZVH4yO1U+siK6duUQ9+luuUnlW
YRRiBXedeuzkU3t85mVoAyj/pOJBFzUItndj6m2IWAo9r/M/CPHQBELEgQMlZrWLvH17/T+ewBpl
QN+zrenG3VygYTJ9WzmQRVSlmIRtgpJjqhwfvRgyBYuA3Tbp7R7x4z8+/YlsP9UR80YlgH9aGGub
mn6wWiK2BCenHW/3hIPgHjU6HE98WhTOzzY5lFQ/UrbYnLXHFUqNV3VsSA/3cNBf4l1WBP9ZO0fy
XYmuzke+8IbjuV/y2BtJH8SnkQPh1uKz3mwWXiGo10xJxW59dLTTm2xzYTJMxhUVXiJjeN2gya1V
LfpwcVtdlUYITZJWVe8xmk/5XVzj/CTwkghIohVwKIy2C5KVJNSVEhG8lQLl1Yi92hdhJysWydNb
AkcUyNpkMc9yCRJ2OiehBOxxQkRLtUcWiA1zwPpGEeZAkAZOpJPWu6P8ED7Idz0/gbmAAvLh2DFE
bEsqq8JWw148WUR5an4Pe1fkMfN7ZFQnrVfy0vQWM6o0NdNYqsmnB6xrXNVl6Hm/2sBr8dOvQ1np
SB1lkKkvvWAI54u6+rNf175UGQto5ud5sZPhoZi+Ad+AZ+ezXWG9xRPt0W2ib4AFqQNUW0eiQ1KU
QDKPYIN1LsG9FmhVeEBcTv5bm6J+XcwmRH2+mpyecmcmezPg5QUcqUhJ5p1ALUdzGza6EgRdHM0r
WqIxLD/8mu5Oy9PGuVN7TtOiuPPQYMrgG3TNunr6JN+2LNIkKrgB+v93ebCyfRhnrM3uv2P3/jvG
2cU7GZroBbuuvz1mBNDcfkzaDWOTg35Hn8jaFVuLv2qbO8qBMGDb4fDwsKzMPgYB2Fs9Ve+YRYKU
qgPNGfeIEwP7lsM9jgByll1qMkC7jkGwbggSZmWAvNozQXyMyOHFIUU3yhjGWukxTBjQ7IZ7eNSn
o/+1twGY7D70Fi90rlRTRhYJfp7XZIH5oPIQkzkUldtfIy9wrhzWoTtnVnuEFCLQYrx0ll6LzRU1
jla6iiaTNbPZRpZAXeR7Rfp86hijoh3kd31PxSIQ3tg4/HC/Z7n5N92tIvfEKIHB2UnySCZyxMFe
Nx06bP+/oGqMq/tT0ttLOIWNuGiG9oinYh9NPo9l8BHZxBgmMRa5DzHK8zCtbhPFTQExNP0qrQVQ
LlEf57eBAzU/yU/cWwkO8PPLxwS5a45SLNipjRFh35iucMulc4GzQip6tq3TitU3RVqN4nnJOuQ5
eYdFXOVvDlmiSXm7P+9kzaOuUy8cNPQWL7hN9Fizhz3DonJzTPMoDmdHO47gNK8PBIiwwWLhN828
lyhHw7+6on2hMFmbi+YU7Y5t6sQ9FZog33q0S8bkaDgWKd32qK3msZmQ3yLlrSNfO5ajFs5nHIa7
cdXj4cXjJr4zfPXPEsWBnwDJW+oNDoxAh1VW/wGQwWlx6BGsknzapd3CU1xJijmVmui74RANfXsc
F5hrv2CYJTWmUmzP9+Yby45tOQTFMGjf0yAa2gkxXkmN+CIBrA8DYQ20Art3C/2/1HnqhU15oK2H
5sWKcI0vbt33EAvagYnJgdLC6Z9KQ0tFSixlVKkf89Ul6NLuzwEQWWN8P8a4I74C8QN13VbrWFEj
FBkaKE5rpuE7+C9QA7heVDcicCkzkHS/L6zGcm0REDMX4Q/FjGBg1Uutj0JSB7+uHG9EFBi4wVH8
e4hj1Fk+3hzXA3JXAFnIKBV8lc5RkGsijmrMpz2FfIVo+dbXnZzBxfXrhpzcLkjbJ3VF2yvX2h67
SFb09oMKxs+/Kg1orU1pz8lrQ9jhKlfXwbaM5QAVgm9PRfiNh9IOWgz0pT/sSi4Fe+orlcGHjX8g
jVwoMMq9MvkyC2xaq/Uyic5oQfC528K+g64vJTywh4u1bMyVLjPuGyvtBwNO7bOyV1l7/NxED2d9
e7bxUOZbPtW6o2JXRSpAz2WfVOdv9DoQZ9gpmSOr7D4ISHkL4CvU0tUqOfkBIvVYxz59AOpTzA7q
x5Oi/rZrXk8OAb5kFWCnPMU/FdZT5sz0n+0xWu420jT2U0YfRRUEV1fBCYEo9nEOkbMl8gj3bhvC
v1wuEFvIxyoArXLdXz5TSNXCcY2ZMBeQTb6ZlDCkjCTdbfEyBjNO+/ot1JoZkvkmdbLQGql2BnOu
tZJz1HXWdevOIwaPkWp1Fmgoqaom9NnsAWDNiuO/D5wsoe+6Os81oItINewNOhnvjwKxLWttRJKe
Bx0qfxZzyEUJQBVpFNhsEkMxImORl5bURm1/ODdFmBzr+6+w4XIi/RYl6x7XtL4JqrMLTuRdYwVg
teU/brZBpbdtu1GvzxG1jb9cGfrNWJgtjLrj8+xKIbziESaH7dF6id4xSsRDpk8HVoT7d58KiFaJ
xvFSC054vhNrFDsl2kd6Sw2yuXYyzvpDiUl/uPHQ7aYW6y7d7mhqC6hDcuZjbedpf5YcMA5EhLUK
zQuff4bLwwYKWPpJa/oTE5E8X8CEWzdyRxK1rbnJYm9QhsHLpMqO9Qrfk8lGlbGe5CqN+fvOuuTj
cPQA8ruM0eOf4Jrq9lT8SzlsXP030/yzi8WUMvsZBHze3x8wIZDy9NSQ1V+X55U0fzhWJ9O+cvan
YpCia2hngRmDn8RSUcnD8SDzLgk0PHYLs+yvmN8klowJcecJY+ROsU1U7teCErW9No+7Rlwl1yNg
LAvC4azrRTJ7A4Q8xvbZvbpvk6jmMmzbwukNaWoqCkoc7blEeJ30My4u448pj/UsNrC0iV8cZnjQ
WyUpDSzCs6fp8sADVjNbfHyTaC61+urUxGMTLRmu+coQmu6T1TrCfYMUIruPXembACC9zVYuZc8a
NjEBMHJxmJNuWGFuFXyaxKdkdrAEsENtgf/XYaiTxiJxQ3I4GF+6ASSgK+g/iYr7COEu3Cdi2l89
eblAhXMf+OHjqDCA0EjWZJEYTLihysJ+uPZStd+5rN2d0dbRPe3byu/+xRKiyeLHBhSSbvPI66Bu
4PIfEDHjPKgxx+NRd0y8x3l+B0SeGAKsThBz0eB0nmVR7xkCFE8WSJZLuBuGPxr4AsyPtw9QbDnE
MNJuh99X+frObpo+z2h7OyJNH6xFX/Par6SDO9RPdNbwyKZWpWmTAparyZDO2bHu4ce7mWElj2ux
7T5U+2dW2/kBMN0kxOKcXU4orXktXZKT0NaDmeuXI0LHpOJWJu7z0e6YPw0HNRA5PX0mklSXXgxu
/8zCburtrYR8AgdepRNfNHRpd+0GxSuha5Jzn56y6syiyfwZsyADPn6eQtuEjxpd8LBWoz+kRgQX
ur7gbFlNsR0fs2G1s5/6wRLvMSvnxbeT3e7MzPU75yjzzZnE9X4H7v4x/2dN3TB0xQSuOjyOJ8HO
dnaIlx6zRrzi+RpizG/OwFAzP7Y7JSnbKfEJExPMnQe/PvXaWSCmfNw2cQaOcFR36ecm8me49Yn7
Wvkio0Y3gATOMSiU31lsCWU3bqbFq5wKuttdTAufZl7tjUwwTBUOexKSm+yt/7eK9HCSmLI3dcoz
qMd+U1A1buEXV7ML1sgQ1K76wL68FM11KjH30NjxUx6xUCSf3n8IxjBWmpY7q0goo/Ys+D1JOVP8
bdZ53p5gPS03oloqBX7u3xJL3BwTJAIlzXDr7HDlLLTt4y7If4+nS4/XTzQ72ihIGkXE42D7Ja9S
9dGCIjoanPkLc/8gKx1vFYA76IGeFV+y/xJVRgz7lXG8yo5HzO4Ly9KunHLbNLBqFe2cTN8brHhj
E6iljRxiuSwOnv4xDQX2PiEH4QCHhRgGGaIby0ZEhcA4oc0IB3QQzF1YI8ibdcWfdTNKXo44gx47
D0Q5tum1OscGckDavweCETQgGlzIGcDn1/0jbg2J1dcpUrRKGvPeNocLHE2io64VjzML7K6QEQKj
Btzt49HR2qhaGSAuIiaQrFKBzpTOoby3CXj5NiNTsAZ1Rsv1bG6R4OfZ9axoPnKelonxMgq2SEfX
fpP8+dlI9He0qks0BOtcYZ+WhZtACoo9R0rxSMjfviwogITf3ipfvEYDQcBF9IP/14OquonGGCWU
ckbCOO1TIZ/gQqNcF7GX7kk02egmQmU9ccnspfLsG0z1tdgqrZJUcL+Afbl/ikhZgMsCBG2CYVbm
SqOIW/EzDj0P0GaiqTlpki8V4zj38E7KkKfMQSY/iCAhAhmfMILTlfB4T2+q9ZTsMXHZyObCFLQx
XZWMYTwQoS8eUelHCGutlENT2DKmwWyz/RwTT/WyjPvP5T1vuU7UYDwm8DPVRMbPWOM3qk5zhR/Y
I5Mb9pwi7njg8kX7CScJkkBD1g4RAFyJFUlxqwxoY/xwXRKdJxg9CmJFtus6CmWr//xqFIZddXiV
U6fTtL6c+FbszTHRX3/Cp8Y1oNGbHW3UY2noXlcU/GHyeVPGdq0EXq9MWR7jvZTN5gK3aulORcaz
DWLm97lgCMAakPw12gZmccgH4LBTdUD6CBeBvdYg54GeWFeOdY4ca/Ld0FDwBHKaKdQog0rWDWMn
L8q3NJjQ59rPfLvonj3aTf7AxKvdIHfIt8eVFxzAizFtQESda6SpKBLSPb3PQReWGA8Gw3WxkCB5
jWzw9bdCa/qixxLfBasPmCmt2Zm/JbFe1gpU9cxWG2zeA18Shs2jpMSe3LwPeyp/Aw/I5yB8TB6t
d4bGAI+76PHzMxUNvB1QJjebmXoA8hqQrPYPMvKaOa+j1FDMWWv1Tcz1+D2ywsCEJcEXkla7AJ4z
25GCGBbXRL738BSB9aUGoyv9VbzUubt6CMUi28CCSOhlcAxxmHgdAHGXvF2AS34gjWNXS5GLcf30
I9jGK3SB7pSw4k3ikgK/QCVgnk/2uPaL98trMyuoK/1zWQO6tMgf9DyeGrCt5NjeDSK11W2MRV8p
mr+aNinBFrqr5Ptomm4QZoPVR9IFp81quoGR61uMVNBsDm1Pe5PDqRBTVlc+6c4idb/KcFBsxs1k
Wtw0YEuCXcpeJpp8JlCt0+yBY5sy4esANs1im0DGbNCO3YbBm3dYTB6VANyz9en742F+wjspU82K
KWmYGMVl+o9EIishH5/cdB9aEYSUK2qcN+C9IjOlWDk0YmVJsJc8yeGECXjSYslYvzPqu4wcW1Wc
8IAzaYm83yLxmKNad7XiFKzc20keV/Xoe42n0dEKznWGxS4KIKIe3CxCia+RjB81kTj0UCMDtShn
/NrOg8ZIuDwWQc+lRqyu88eJks6LalDS5bjaWVxQu5jjklaSUTlTR3bZfuIe6Vd+bD6IfBdwPRBr
78EzpEG3vyD/gptcb+0wKf8RtbCmsxeK3P00QDHI4UGM8ZKFCQreS/Scd5x6eWtazclYLUZheOkI
uBpVCL5RY+GR/cIFL/Q/h/FqTeDFuVP4fDSQ3Rn9DTUzEffITjaFLLwB8YnvAj7OIUdGl4cK7WFN
YDlLj0saRa+up3dhJzynFZOLd4Mb2+HWEImWtgMJ7HNIyX3JdBXUQZRX4pWrVKtzNARxBqhp/tLO
qo2/veXSiNOqixVxgbwmpfY0iKWmakagxtfJpIIo2/ra4xc1VnV4nkL41Ig4oNDhOm63S8P7j27T
Fq+r4hgmwoFjFU9Z3ybCMqxmkoBYOed8Tr/gjZsbVefpUgym49MMbePYoxNu7wgpcnfzzGbbfJYF
tmXfwc0a2/jSMvIwvACdagrtMBtTOcxLz9AW1adNHyPUNa01T1Pyh8PX05zMzuyswHR66kCZvzFW
a7JYSLjf628dUOYnlSZ1j9K3iilBZcFiJ9PTQWxBPOktWt3BR9NUVUIBNSh2H0uvW9Gp7BnPkTyZ
zwI53pbEFxp7y5Uzc1nZIzyf3ZxnqN2kgw78fsDjH7dOZZ6nzNGbGq5l1DDXKARYyrKhS/lIB0xV
wFFoLqMGjB5XANXTbo+JtUsbkL8t6VwCU00dUfWE9TLgz6mFSig0du+hRHyJ5pfSqIBTrUpwhwPZ
vrvaOwo1rP+QzGFnehbGr4gkbbMkZ+6IvoEQaNnVOddp/zuzhAXY/Zuhyjd0hU87gTBjXeO/LwjT
3oC/qZaLj4nUGNBtL4JVxiae+kUIgi1yRMs/cTNS2RU6MZJ6klTeryjvLQUfpJHj1WCLEZ6s3i56
aXhs/tHk4S4+Ce/vSSReGbddGmj5CZS7g4tcJRBYRMUzYO2YR1DIUGlwLIWN60T71vR8kkr0vJyq
X/gOZDDs+8ax9ERZG2oF1h1K6ytFy60DJ7DZ4wZBIwXeUPzUXm2z1GeVt/JcOg+YG7CMyhJmmSOg
Ra9ZxmLEeW02v76LVb7YoNzN8qUeFbuYp2qImc+v2bwlxaSbUvjaZF+GY6+NDRycsADwHSW719fH
Lq40pGgMK+Oen+eyjgSFOIfV/ks8/Pb9SHS5ZrHrCHt3DZJXGIQs66ciejmYC+M689BD0UeAGOp5
c7rjfIE4NfpnBeKifwHXypFH/Kn6OShOZ2UyUSXXOIxr/Up+P6/LlrVls366F5i945kTUG8mpBDK
w7wXOsgA6R4lURuJTkcsK04Kw3Dy5hwrdtVP2EAoMw2zme1AM9H5zQ4njfdZynopDud98JABLgUi
0w0qGqfWvB2El81SqJ0VOY/VI3w01IlEPCSLqZmOvp+GcKiUHM6Yg4Dj/zSvg470O+H6S1VaNdU2
goF5c+Z7gVUSE/FvMm45XBspyEcXrGoddp3GeKt6IPQIEthAlBt/j7Y+w9jyZyiVTgy3gFiSuwBw
J/51kIPSMbd7ZQizEHZpEQk1VJy96zpyF2Zc3sc70jHK7UMIZH/X/h+2ycX5cZr2hg0kHspaQqRH
I+T2iusFS+B6Nq5XcqLQo/A8PsximjrNZYfRocMSf8roDoGl47Ai5K4GiVs9pQ6G55G2+UHjS1vM
K/tnCKlV0SBFC4KOHcbKzojwk9fiS3Z99oinmWcQYM3WfaugO9rhRUo/iXuMBTnz4fAcr04mbmG7
zeVDjAVe+5LTFqHii9Otfm9efkDa/mPcbVXGLtFSgpCcCzBrSMYGZ9GNEzphn9K2ujmchq4QiKVM
8uhQA+MF3LkdHOOG3fgch4sDONcWRxa0bdMayOAnljztf91T1uuvDVeu9/+WsDFsi217OV0l+DmQ
mxe8mi4zXBFLA3T+hfyXk/VqhkDlh0mNeHLpHzeNTut14V7JuTulOC1qTjgKIEK77Wt8PaxudNn/
kalIMCd6fSoO9z2LPxiJzT2+aYJ90OnD+GbFQtFdR+kG3TlFWJ99jNcdf3AWgHgUuW/gaM2qxU0G
y9sDLfdNGfcaPu+v6PNinXqLF0u3FaOO1M5xEuE6IJ71m2emqu6+8d8Aj2f5WY4qEsDSrl2oD2tf
cv/7KI2xTzJ4n8R/vaCMIZVPh4RV+/TSQ1xmIHxZLIw/hTlP+5ugZkuCU0XhSBTCks98G/ryo2V0
MgPxfrs3jBS/awiv9SQpY8YJ0wqlTlNc5zsPkV+OCkQF2pi6Kfy3NXy09AL4U6ce5uhfnbWwRBQ2
64rh4XhVr8sdI4wuytWsfH6FuBY65+T2a5xVXs9+Lx4I4R5EOJGv04wOQ+70/z45CtvsiEAjFKsr
sRrrxeUsZCiUBywxleH22YjRL/yxOJ4usooX/49eNlrPv1mE1HoS0t49E8+kF9p9gcrKW19BtUL7
qBVbGCzJHecXZaUlSZ14dtvcz/C/uSfDEFy3omzitg6xIPxOcuIgpbiscBq10B50fjcPxzl8/W0k
Bcl/mGQralShlNN0YyvZ3OlTXq0F55UhKiEhPylkLU/1uGh7JV7Wv7kQ0+iUgAe+z+F+lq0ZvId5
p9NYJwlhC0l35par7Y8pBriDtySg9stGLqhgxrTN9wbrEzJM6fKiaNMB4qdIZMmunlg03kFPb3O5
TgjwpuJGdS6MHTI935uJ9W7wB5RenF0XiTGd8udWVbLP/4YSjvXBNL2sz6CZc5/qA9HhOxe353qp
2/K5qsrKJJkkRtx8JpBq6CDlB3HEBjCQTVOefKgCBs8bax15+VafMooOm0TfzI+7JR/mS2hSMV1R
1rFY/58OvV7uLw8G9Ac2cNJCn3645ugqJxQNBwu1R3WlEyk7K5y+O/PLnh4dROXlVI8ZC4F5Tgu4
2DZXhkHl5nvJkaLFGNNmYmPPx2xsGajRJUA6xS3fahgewk8kvAFgGyU3AUffYG6DM3+mD1bB96q0
OvHctNiH2lgcJRouBjdetM5Rhn/PuipQmz+S6GpSk8AdNvwDOcLVnqwRLdZaRA4N/0QPF+1feBN/
W5vKKPHrcSQC+jVNGjuAE7RCjQYLNziw+KWKcBjwhdqdP7tqw2YvK3FI5h3yOlYW2w4AiYznEiFY
XdjO/LamTq30qJ+jTDVNi7qVuc53NmofjDvDU9qwRhKagYgpHroh5yjoyJKanVvYq0CEYX3DZKGM
0QNuGrhqzsUJ07NnGWR3ZUGoUtBdzt9Bd21EWdXTto8tQJIIWofsgXRvJlk0tayhtNae+Z9c5JTR
9rzhABwhHybAD4gc9le4kxWkZNKBDe9c1f/o7u1UYO/fOJj0hI3N6cu0FTFetivn4Tm8Diac6m8e
LoqKIXxN/VxRs941KeWong7heU0Qn62+IdLjNZwilI4b7X9OfRGxVprqM60P+Y8MGjO/riijtxef
CxZu08oZQrZ5aGi9MCxG/M5mUwY51Lw0I+CgBjaO0I75MFrwTLXb9PgbCMu8xUSn1MBWpkNUQuhp
M90fetQCF3AcCIeVluOfK3WvXvORexV2s50z3XX6mP3g3Xyutk3t8V9Gh+Bs3dkLiMQmq3nlrhwU
w31/s6sCYvzNrzgb97cbaIatnJOT97ZHmn2ljoRDvx4WvIcYFs/7LyClT14FeZluMEfXil6s3MVi
GOvn4X/cwL3r1l7RYrGQmhY1/L8wo7L+mXi4MMntNae7eooUCOxDJAQk532nionwAPDDK1PRZ1ct
YXJDzsOyR6FpZ7LRfQ8qhJ9swa48iTBG7vyzdokF0vfWemn4FuUcAXPDkMMg7O/cgylOJaoPO2hO
TEw6EGgHDKi3qgwM9/W14wXBMIAMYlEPFnwD7+Ut49rQDYFGFK83bpmAxFiPZ6dr1U/y1FN6g1wA
Eb4h5CgW43WnI1MX/QbDRAKOuU+HD3ZpqrQ8Ekqwy+fDlrFUhlI7fe8+UlRI3CHNFGCMKYM2UNIa
PnGzH/WMqbQXKUoYlHt3Hb9pzBo/B6Zz5H7q1K+IL1pcdO+NS/zz3XdQ0Ds7ywQZM9Giju1dv5zH
mxyK76oTIV9lijLfkcp81a+oYOvBBT9EkKmfFVgABm8JyE4TjrWIqUexWyUeVrmXPjkYlEtjqO9Q
t2e2/VMicpoR2WhwGQ5Vm243PrwdUBpKk6C2/Nex3wgi+NvGJiSZPvF/lU/xW1TebhBL83vhlYHV
duqngVNL0dK18LZse59Ed5BS2FqJN6pssDpR5u+MSFHzd9NWKJjdureIhtm6/KUwm2r2bh+n4h2x
Havla2hqXH2+dsJQjJp2jWX+gRpQJsC566rsSECuxGy+wc+EG55DKE9Zir+YB2Hs8fZ4tjmhya50
F194dQdVSrVPt5q7MY2dpxUm4wF2NtwBPaLcR9fKpUI4KalFzQHoE/JMzF/UMFTtlRgrKbkIeZ0n
aJlMDxdKXxd4wcZl/7EZTZRvdegG2wdZZNEX7jz2MZvTYjUbFg9df6nLVEmdizOkADKqXgrXEs8a
7V75aD19GHg183EsZXasSERhaEL5Bs2U/0jP668S66VNSrXr5mhvXSzw+LlindF4pQCzZs4F4Q0I
o/vWQdHYKyYl+BIlUaLylm590FBYcrFN8CpgukPEeIa2K0+IsZ15I+Dvf9Zkmq29CmkQOwfT/cQJ
N64qUaf1vQbrWt6baCONS0qOpb8asJmEkBfa1HmXe+pBuBYNMAhpEpBUKCS8zBsPf+058xVGLac3
svmhuA1FeAtGzqsiqbDJFykVwT45H/AAgoSQCebyl0Tn9u8yl7LUGzWV/k6NsuRgfra3SIkezZAX
7yEEutGI+Plb7GQXCiKsX9aSD0IeELbeNvXtAP+b2WrRaT7YL8bv9hIVxrl05BLUiq4+uUlK1NOO
C5VnvUDNWfjSDw9sCIiplsiJUY1xkS+OGZTYbOhD2OS2aFvQJ2rBKBkmak21XY03FlZw09Q/im1Q
j3kZAjqj50mtMYf1NjSg+Jfe7RYl5CfHqlDXg3xdNZSkx/9La7kLKE5Db/nA1SCSk+BW+JRkFBDy
GJ1dxzx0oXiIHeO3ub29nss8+wNgUYSijHNe3KEiU346hCC86wpKpx076oIokwIY/xaZHUU6YVlX
TVOQfwLaKCUOIVx4KY9PEYsjcZHhH7wDvIDJiGNfkWJQbtdzohVqT3shwZZAzNY/IgRiRPg7s5RA
eNtaBuQkts9xOh4/gFRY3413jgCuGYO8bQ/6uEjalx9hL0oJ0TftOHYeMW1HK1Pw5+3/2rlzXTVD
BjM981cWjtHcOK0qCTVZZelx27kDZSLe+45OuywOgCyHcejKBLXtFywzYl5YH9XLR4M036IbrLzM
IsU0GWlLVTFb8W7ug3cv/p+o7I3/QUCEAlld65o2HOQBLxc8q5XL+dGjsspTwYWnBn5EFUa9iMNx
Zzzfn6wor0hECssyqkW3UFl/eoo0kZymSHSWruQVUwKvYXIbSEV3STBPv43TyXmbQuJOv7j8Fz/P
2mXCc7N6cPYFrSVYoCebTjGCH0UAA2XsZlVaqtu3tneqhq80i4THLD2T4mKOQ30n+4UTOP/+lVAc
W9qKd7IQJHbHW3zRbHrsLL7w1KclKjRqjtu958Y4zSb+mSiii3Ob2K+WhtS+m4kfsGVJBRbiKK5u
AQuegskRVM5VLWG8/UfZPcQ2lj3cBt2BLqAwbkGvxoFIrgqAyF6T2Cmh2x1eV7dxbDJJJjXZhNM9
Oj27A0mPZKC1ZEtD007BpTiBNt/LoUMEKAqZO2vfXa92v1PgAfbU0hBLIvsgikdhLzQnOrpV9sy/
UGMGgAevnt3NO9a4TEC7wIOJmCEOOgKH3Xd55JLSg7QdfqBoBxEyqudts/MauwxU4OiivUsf/srg
OIrqKX6zhFVkrY9TfepVmzDmq6iRaeGJjiLePKgQ8+dGXKU0JWtfy6uGg83sHA9LkLcSzNzoAwA1
tmKhl1VUoCkYZIKCtcXZ0DEM3tSS8gWP3uXDcqNx6RooIe11NNThnii6M//OajNYItpg7r2bR4l6
CTrXoEDtah1AbdBMCFKWUqW84GolnUThtMasM5/XWiXU3616yEr6XwBYpMSTW4S/2c+i99/Em0yu
8sBCS3yzGlyv4tJ1WAUPhBXYOW75p22CUA/izPgye/Azh0fEXkDR0iVk7RWDX+sM2LV8k4HnRS+E
ffzsVGNqHt+t48HinQlIpxF32X++HL1fOLfedhMXe0cmlM1cVoR1kx9uP+wZ0UV6OoOouRloVZ5h
mUTvuysaw9VywOWi68TjequrYBo50MbsbJFJHtTod1K+kNT5Ot6Y3ruqsUOokKU5SgHBNM2m3xmQ
bym7L8L+mcwYdc64Yno7iPtTXTC/IujvzEotFAAYM9KXnfNPjmjSq+vxeBvCYOh+5U6l98g7zLnU
winfL//KMvZ3gjRpA7pwIOCuwx4ZyuxEwWM0pFKIe03FngZCh+trk7ZgGIHMCvDAeNO3mbwX1nDa
mLjsnbrqMagY4knshxVgQ17DZxjkappwk+bm7AtQJSWkRIJcwt0/Wm0EoqdFwsgZpiUF59GhFOp6
xQgm5aP+7myU0TuG+gqY4s9zCBaHg5DN+O93DKAUyxj2jkBUIapZAWe5TRSKBAYAPwf954RDUdcs
fFkTR54/3v5dr8Z9pdcLCTifl1usHvGyZFZrbX/utmotsHBNmW/eyMO2wfX/s40RAvX8bOQRJ8GZ
/819Mc78/y+6w6bWpQakWSITXw0TcLQD9ByagEW82OE53ArhVTXqWrmZbVSFuKpEzYKide9OE7Mw
68hcGcvRMuHXm3slRg5WSGVR0Skkyjwdo+G2zf5f81kFNReHFIXjjKHIiBRC5nIeznZKV0Ln5o6B
wKP9uejtkDR3cGAcmGcDWYfzlMP8ClY82pDnulnfIgtg0vJzD4G5XXKpAWfdzJnW75NaEeElbDRH
XFtaoq0C8QQv1m9xWfk45M8Nt7tyMfZL66LIe13Hid8xFsF6/oxlLuRcqsChAR7VBja0fT8M0a0V
OUBuVKh1esVU/J/vu0KYftZYIdgBhsQU3SGlQDZ3X4EqW+TSK+zBc2bgg86kaZJ4GTBK2UtdvMkJ
FK3nK0yshKzvEMOlewTmRLO5iZHFeTMXDcKnuSxHP8MdIS3Ru71x3kiVBxBRR/oEpl16ZY/A3mY3
aG6L4ub+WDwk3ne+Aq+c0FYFQ8rf14yGLYBh1siFGztpgm3SqDWn1CAa5yQ8LIiB0eXt7SJw2IVm
As50pJ6cK4jrJlVmlGrG0pBxMjPqYJZtweYScBa4eXNu8uybl4yHoO+SRnVAjtVMdpCAVEUlkmPW
jdmv9++e6KFawtD/H+97+KqWNJLLAqy0y1+kOwMvN/zc7HkHBBNEYmLGPFY6v4uZxw5fpgR2Bd6J
2hJRFpHCnG/lzGxsuqtnFwVzCOHGqiyusEIpO3AMQoLU5COBbuE8pNRdg/3P1zeQMYOepQ85I5K2
0VjhkUOCXpDMqpGnJD2P92Ye03YE08L0TXEAxYgK4S6tceqIaYobqymr9sNOVx4he23adTlwsJue
6/J2YUAshDl4uSBL8FLi5xnJCu4i5TYA1GEBRcslulmNen7ATHuYfS4GVazcP2AN1EqI4PIZVCg5
imtuaoqX2JTjReAbDd4wiad1sGpySRbqRqWHCJHHecNqxlUr1v0th+MM8AziDrIrim489ja8cmPs
gbEPwGfAKW+yeoIfidwfTuxj61l0Gy9gUOrs5MLp6x3uC1iidT6CveUjaqtFR83aQQ4Y4IWABdZR
LoLMq+tJQkHlJnTTqqDTFow9t4H3KFDbzg/KjoQVZIqwcQUDVbSquKlqZc2BJS3khdwI+mBjJ7wm
QUr3gIGtULbbEmT3BuBRBjfRNT+kWu52x6A7A6FMBtAG9ghYdMrBUKIm8EB1WMuDXviB4uFzPQNH
ac1BaJarN7X75chG4NeZU7OlRAW+sfphkt37G6KTa4CdpeXL37tuQR4XPh4MKu3FTOac/ex2p/TW
dj6q+36H19KsjZSmLAEu8DR/l2D8pn9vi1l6O4ocRVP8cq+ONu3RPg10OsdtCWOCY2JfisQC9Pn1
FLlZGP0IBCC5yCD602g4UPicFhAbRHQG93I/SoFvimSdD4skt1xiN3e0cJ39sv/+deAJvV5tKA60
5+8sBNQAxaCt6feO3p76ZbDtmTVajBwb4ggpNMRjF2rsQVhg694ElfK53M9E7M8C3UCxE/edSVdf
dHjuVLzhw7gXumunDHKW9jPY0UTCKgeS4IhUsEDq0Fmlc44AXE9RotZgtLTUYQFmyHmkJAKCgmR6
w+xbpQE3rEufGElQbC3YdNO+ubTqcITtEf3FkwH1WDDXqBsBZBIU4qzakFkKsgpCVzTlvwf/En1a
V5BM314Oi9MhfcIg4sklYzVncqba73/5QmcL/+8QoVSgdYfo0XWrRoqfGgH2uUSeTFrCUCWOntFI
QW5ynsvaZrhgfpmlKqNtwvisst2CeZKUFQyECBY/oGNyRnsj0N5c3pGeaUqSzTf6lpZX6Y2xt+iK
UBywvr5J72ukbnHhfITLkAF9TiiDgsye7mwVLcUI/KiRje10fVt55fFToaZJyOLcqk1Zfy5o//ZK
5HT9XtiIYbaNdGX9mrnuqiGlIgvlg5pDJsqNK9LfePIhoHNFJCJk8yOqNU8Ie9tA1/1HXICmZSwd
RPlUyrWLjujQZRiy4xkVvE3KuvSzSF5zDhCCQxPY4uTmgp4S33qsJUwCNtXtVx2Hl7mTITnjRxuD
NLftl7ACpXXCNcaTPfMZuZ27Nf+BZV0vACW0MqefbAkMUglv0+pBW4e+Mkr3T7n63ypzLsZ5Mi5i
csZ6M46SbYIop9RNrXAoKd3XcCNj+CzxA10qs8PjjqBsS1WJfC5AQ71nguTQiZ8mp/Ak11qlFos3
umx7SddLbYZvFnpwU6cGhKvpAeoNuSmobWXkUlx4LDtXOza4ube6AJIpOnORs24EKRwQhZ3pQg/J
3OQiqI1Gq53h2NUrOZ01vIzgP3PPzvKQan0CYsfVjpVRY+BbQjL0Cmyrv3yFQj32o58L0EF2bTM/
FvqO1e+8UN+UyzJ/2TXWBYV/9Z2gWz4gopB3H/8gg4+UoMMlTTjAzxyjxXiLTAC7LpkxcoKndIrc
bpavdKgZ4qXDcagYeLez4u2D5fXEUD1wH8NaRO4bzJbljTjcjc1ogrp9UspLFLa7hhFdDVaAzzDV
KNaKMYCp+lawWj2VbLGCa/Fp+Y5K3i7SiXBU+KmixtHJ7MPqAj5NhnxpkfmsIgzEvPjgJumPxBXZ
+BVN2z3ThKHz8W8uKgdTSBZxvenchvDyITgFc8WHqLdFlembC5bd1PKoxa6nqA/GZX2flucckP3B
1vXd77OpeJHb92xRHIwPA5hnDDW8rD9aKDSraFqT19Ioc25jVEPYFCxiJRCE+D3swpv8sJOxag/L
beIK3T3i8hVdNGbS/tCxZhpxRe4+FEpcAsFYVxGd+Y5HTslOYVnaLrhpZU94f6hIGfk6/vpd3Pg+
k0dFBGAzukDIl7nGeNHsq8NzQLwO+WBad//rtNJ4faLmslwQlnRk95SyTIqcAOmVaT7oxDWrsO4b
lnrWheEYC7yxLsrOiT6SGuaw2UQ4CQnZ1A9eR40TzvvbhuAQRmggsqN2fUoU4cihpYsvkLNk8PiG
exLb2Um7SWIP4ho7E9L+GDAdAzlevid3fCFDe6o2XSLxBL4byr4M0/tu1SeskVh2/BDOJg65h9JS
RktickoHFjASFuVnF8rqXO+nfQkiJyATQROYZ4Q/8qUhTd8CCLOQ0QKuWpVbjdtmbboyHFDuSmOP
R1dZxWj0pQ3fQILyLwKY8Up0NWcDF/IwlXYQ9nw4qVxhBmo3X7ltGSOkxNmcKz+Jn3vCnRiWIfRw
QqyTUnFjiamgMxJJxc+vWJ+35ZspgVHpnpvroiT0eWGrvf/y+1ELk1jn8n6ADYW6i5qFx/hmEKPT
RDjdJrKHsp9Fv3/gODNlvJgKa4KQSPwgAEIYsFf+XuEMBSiWDIWJi4XmKYA2QI6cMZruviufUu+O
qO1F2vz2xRSYhTy6rmuXPZInKxTLsphLOFadzAzv6gfbNzRajEl+3jl8BDREgnm9Q4iyx2aLRf+7
/E9D5+EYOzJJnWFqqX7mRuf7mTXNr0+S9mWaHachVDUY0Zg9Zs/JZ3fiU/dibCFjZx7lFV1XOP3T
W4VV7tQWBYzbycHmYWm2XU0Md1fGVoEx6uE1DOyp1lBIU2goCBJ6QrYEa9mKN382d3X2GmV00eTr
5gLjiEsAdZ0IYYJeHpGFZIvIbS/3iEZg8YrZpVMLCiVvTVcN/PYenw5Op4ZQF+mfi+UGK0fOa6sS
CdgrEgrM53mGIwihv4P4LlCtwftllMt7laiFbugrVhI5tHy2P9V5Z6xXsxsp6YZxwnvWwtSincq4
j/LowNj84Tq3h26UgWBbQdG5uEBc3k+YkomC8CO59gvZ0yeQYkIG4ufXQp3G+YkIwxsOVdLykFbM
xkKjAYs4lryR44ZaPWiRIMJz6/g8ynTFnimTczaq9fZ/4k8zEG5d5eXySAw5kYk6yH3QoUUoFEOW
Xk7/UZrNhqXCM466w6TRl9rw72G5gaL9d/0P8IGkCEPqdJlz3I8V0aWGSqUskNaXgKJCr8K02Et3
V10ie8/WUaa99wu+t8+APMUSmMXM9UVCrIo0HSReG1A0HCWtefgjehWUxY2fQ3DojX7Gg92Xsg4Z
GfQObaAkQVqWBl7Ca9tY+F7wQJ2z86/sKNBHyc0x0U19JTk+IqSAM+BfAG7UXkE0VFvSpaelvTkB
PIqNTg55U0VNJ6PBhM4Y57ldwpMxxmu9q4JZFdNGst6uhTR4GSsBLKQXbZ2r01CUhQ9BbCC6sV88
O8W0BGTHYlo3PC1D2kKpw1QNPIIZio4r7+1AxmPphF+cKjCjP8xn2gK/nGLaVQcGZkdiloIqza/k
L655Pgz+NAdignbj18Qi7Pjq5xerfzcjI8KhDonqN8HfjUVCy3lssMulCuPBgCYSBydnKz9mcI9f
N6vrN9w0pL5676m5PMDG2MzVGngzSkoCpfiw5J8SSIgq5gMLbsbQSD5T4Y0phOFcCJ+sy9qvfSzb
WSjCUUVAjqqTo1D+JQR5bjiPyLOhHVcGgKUemCftU/g3YNU7JNHqP/zSK1wY4TUWXcU9q+jX6sZQ
KZfBZQsB3+2DP4C/N9aNnGeT6q3/5N0O5a5pTKP7nl6N5MavRvpHAFWpmSsguHYEXGk7HEVZS2jv
Rtr2zPWaWJ0EfjbMq12yF80zyIFvE7IP+htdJf+UTpLpjsFHLbq10sa8MTXEz/3OBxHtbD1VrpH2
vFr3/HjRE5lyXowbku8NfrcPeTPSlNGov9DkvsysLA1Sa2r1QBdhCwfMxDjI1C6/vDqou0TE1GUP
QwZ3+vQwQT4B05JVpM1/C+AxoIc9y71F5gKZFqxPGvol24AFlYP0Jmv3CHegJ/dfRR0/cKi7UY6t
Z10AZSKcp/W6FWHLTZfYGj+o0fHQe25mMEXeWCkDRuSUepFrhKMWaBaViBZk4nttl+M5rgZNwgzP
2YMpUCVwQPFAc8f3oxIsGJFKJuPzxlQFL6KkGTGlQYnFllTTiyyPcLcXKko5MRTjRq2TuO/ZTv96
JXK1Af4zyCHuBVRPh4tva9gBqWCMMWFmC7EnlfzR3F0V7L2QkM8UOz2aPvoURM8MR6fnxQywVPYg
NQRFk2leMsoc5jtsjL7/pyU2NvjxiMDe1OMctSdXu52ilLC00YlmNHDdIxPisGBOf4NldcDPQJ2P
yCQxo8H0DwEeipw8FfiAYxz7cOqBVIAVmcXqqB7vboxmh2b1Nt9CWDgfEb7Pa6OWLC5Z3OLVbfud
pwZ8au5I/4YNJQlPBpuS3pMEv+DKWzyd58si+oHqyMSrooCS8cNaIqphjqgjMf4P+JeBtgfydGdj
dEpHIVim7IxHDkIoXzd5GAL8Ms8kShVdQOyEzWhJkvr3RtGDqnqkjSwpvzOhxalO5mBLFu0T8ApZ
W2tA/H3qdoKiqI4kBxu2OfwSQDYPYxTmHLW3fG6xWxMks81IQzR54oCKibxSLZkJHUHpQEvrdJn9
Dd4Mh/0WzKlTLPKjuiDKYhv+OKdgy0XcM61+xNjNKlz2G8M3Rha8o6GBRq1rvXwRnRMwDeEXbQ6q
najrWKgGAPlw7NC5MUc490wbrMLdUid3rdlk2G+jWHvyhbg5NFNvDi+ChApu8NHHPsxXHno1vtzE
yIKOG9n7G5laUNNH3wT94RjWJyrVg77ROnOJcz9aAB9oaFeQJZC0XNSjPyqF+ttkd3VKpXzlcBGP
I+BFRA9Ol2wm7BsSmXPiU6WR7aYB2QPy21xbuCQmlXtvs7FXNwKP+/Fvh1xjx1hMbmkwOfHSMaTT
VKCh1gOajrUIdlPeRILvETa5nnaAYOJqWTXtc1gXlFtZQPlZAkJTWTWbvRjm+Mz3C6hHN8WDQYY4
gjqXzPP2qhEwKRnhmI7yCj0pPwAUzzKyYUS/pgeYGcaLmN0FTz+A2NlFXdlfb1oF/vPP1Ctc3GDn
uGW8HgSXADDBTf3XCaDjoqodfzbsmngATjnr608Yb0kBMyacK1/kZ5Y21pgUIGC5pyBNPg56K5Ka
eruK3LfxMO0mAdYBPlQmM8mwmJFJhiiuDUd8qBzxgykp1UPvJmwO5eJpgEn41E/psncjbqNydjw2
6DXz2NJ81MLL93wHmszryPGK2tlrYMpnex4t/lDtKDTUKMFuDK2fRia3N1g0LOrP9CI4VxOE4RX6
kAEyNA0aoXNnhXPwJIYy8z0z6SYaKzEoqYOr3HDUZqrTbjX82pknucnB+XNDoQpbYR7stIb+RT+O
WqumOZEOUXtZ0AnAYTRSncIyYOUgCgcGBB1tiFT3fbs3BkzBfFU/wa/zQ8MZVv/15TJPOA/RKXax
42jM8/zCm0P18/cQSvOTDLkGI87gjc3y4AutKN0YKnOTzJ6RMTy0clXn71uwHRxcXGGDhJFe28Bm
Yhf9T8K/ULt8IPWUZEvXlapmR94qMPE7x/+pTwirFjDyJCVfTtmLTqSOza1o2fwCESFA8/dM1pc/
YAwtnkfTe8T70gMPMb0XvSfqpJzAVN7aeT7NCi5rVL5Cd3vuMakQGzmcUTnxRdpclfEq4yLZJDdL
zr+OmgJbnPkkkBx1n+Kb17MgMPwFON1gIJlAkMcc0skXpV5+7FWbQHBiofyuU2O0Os1YICwUx5C/
0DLD5H5cbdlu/PboYLgloXNO6VBbdKGGNfJDVpJ0dD2ToNSS1l/cd9DZn4zxUBoR3eabwwZ+P4oa
p/hLTWvhqAQKRSJcpW49pJzDZcKD6d/mTF5PV6fMhpzIcDO0Ft32iOz4/8KH/ohzBUpOVdYNOMl8
W9gqLd/C3GVgWx1ekjUjoyV8n6d3jG7PS7Wh2zzd/AOCBthvcORLtsid+V5FcO9/9AUSwUC2Dewn
xcwJVj5nKQr/IFfPkijd2glK/3s7AxJfsZbF/k7jarKy2zpp7/pvbeU2gWKu8n4OE7mhuZ3wxm+Z
tfqwTciFwiu+AxUtqWcsJF8T54ydN+Jxg2aiV1vRjLsy8ZqPUSEuw3MgglH7NVrO1wXS3baGecZ4
jnimwvTdO5cQoP6wRlSS3CqnRqhHRN6HkxgkjVXG+mzMCWEH6kEiv3t1qgSC4yjRv/nIECE/BGYf
6kqijL502h72yxuz9bfzfdAGCsMKIwPUykVCxWQTD4ixNhJRyl32I0MJtS9mOIUsmRiHLie3C1D3
b6U/LUMkCPEprnK/GNNdtCJzqrpxL6BBykvHlnreegIn3IFt+4IjkOMTF01LVLcgzelE0D5FCGYM
74gI7/uVvO+CzSqT35SCR5t5GGe5kux4za5T51sOuY3lrebpb61neD6XNhRmY/YlWKY+Wv17tpZ7
EvkgZPTxcRFujfESLd/fshGEnh/tk/dlqhqkm0dSAe6E6DHBz+c70pIytApOba96vRJ21vzcsWXO
dHtnFa680xWsfSKWatnBtClvxePctTuT3K/tdRF19TczVHfgkSrP4nWhL2V/dhYNZmCUAYNZHnLl
LUYcv0rTPQF/oUv5N+KotDLFxDV8YvOwmdzeAvo5Y8HigTQKAbUjA5vf761dkN2PTaJVVdwHWcwX
HP9MTCcLAz/f+TnV2FylfzAKpwhzb/+/hkqlyCT+H2gUh41Qu4NuJPHrVm6XKSSEI4woZwQCQBTL
+1HBKrgnVEuEr1hQk0pLiqOOsXwMfRNmYzbJxtnPLvu+7gn8dG+uBh+iEjKe1F7g3fBiGZsy2etZ
sjSsOJK1TMn3iGl6mhyiqgKdcqjfNhQVJr5oWNXpPOXgOCEsIIP26mCDuxxuniKLMo2zHAP+iDjN
oM/JZz75pdKgdnbuNbNyL8KUpwoddAuWt8uHAJmQUkJke/34chiWcOEdrxdh3l8cROadDEQvnnDu
SZOMivzdRiCmRNXz95l5EgqkBpQaT+XrKVn6ZExzeApzhfPGfhSbJqXGHkVuphzgkdeoKLEbK+y7
+keAxhnWgMYDsLiML/K0rW//qc9caOELxEo8b2afKokIh4R0n07whMfllfiWCsb1Wf8sB+EHxsup
vsEAVH5fOuUuc7psvUTjoL0pcMY49KiNf6c/AyqNPzN2fhEkczasN2PmGDqnYDD1JAsEfvDcIQ/V
99HF8uId9JxNkULMI+MYeBr0P6E9dOWYFhaeCeOOuyKo19wlx62tKZBEAw2ueYwYSMlfaNUJFy12
K44+nTFWLX5lJjK3z4rhxK0H2NB12JqiFlHrV47KDovyw0ocvciOQxFey0tCPqIlUVYOvGOfNFzX
cU3/bOr9rdcDZo2o9hFih+i1AKS2Fg0eq9spE2+XcWyJJEqI7ajvZ5ZLj55U+FjPLJlXAEUWu1w7
vv/qlpirdf9rUCVlqsy6WPF9O9mT2SSE6HYZ2mUM2y8ItXUc82I2a3hW45XLq5L1mbpw01ua0KLU
CpEHjtw4+Bug/xtPcPEPhEFFpOvvnWIJQNrhk0m5QjUBpycajTtUaj5SrNVlv9YsKcQ8qVKRLMHZ
HkRaLZprjrby7l7bMB9C39UMv30dMHySSm/o45J3lPzPOZnpkUEKA5KBZT64mOK+CXBNFONhaKEQ
N/Mgee+VBB5jmjqN9R3umMrEFWJvW4P2y5/zAi78USstl3yg6gVO+X/RbnpnguMmniwZzq/D5W/o
f3X24Qavt0ulxAoMBwXU/SOT+7QZB07XulVjRqHdPHeWAlQ6bueseq8GPfK5bB6k6haD2eD6oKwB
IhID6hF0FnU34iBcAQhX+L4mSnSgwkGQb0vuuVZMJ4E0mFPYSOV61/x0ZCaJIBvpJooaU8H/Gmfg
uSis38vRB8s5uMsnBXlDi7uNSuPuVRHfup/nx01oe1lXRFgug63x/CzqPRPwxPwNMQtENzkDrHQm
NSBy7kzmQt9HnDAlCstdvxHvaB7IZg4KvHGTY8treoQ+T+reKDum5+IWSt51allApCs3RzZWI26/
G2VZnEeGDkWVMVVOZe+uXPDp9ev6vKoP/ywmYrcdiNthq5wMHOdtr3XvSwXJZOcfJnp4N712XXI7
ZQSqce7mgYqOcRgT8HpO0pF3+zhyWq84F/L5LDEj3ddocooJmChWZQw9eL5iwiSdE+RLFwpFMj2O
TvYzl1TPmFxa2QqB/nx8U8hRjQLBGK9z5f4OMmTikNklET5k73yx/tW1ROcDVtkIEailMhpNI2dq
lckFNWszHP2zGB+mMpQ0el2vlKjMSIvRpi8n0CEKYYUgIyh3e0JVrgv5PUevzQQSQ8zndfk6F0Rq
tiDKGjGKlocLe3yCH13LjGru1jBUs+F0/oDiJnuBIi8A+u/wZ9opWH+Y3KkR58Q3hJjiqkPxayZS
g19qqJRXRZtpgzV4wZQmG7g+AyCrr6rYRao+KDDYfcS/kBoSJjmn/eFl1gsdiTDZhAVpPs/+rVof
uu3yKrS1tLvmgPygv/KXv23VsCDfqTEGg1xgTEsG+F1KGh8kAFka972/xiA2kdBrooTbcArQ8QY7
0RCG65+IE1zv6WRJBzf87KNIQnQtOdSk9QLnCoPTAIMjpynZnA1F3L7rTsmKIbCCUVlmLemF5o/J
kyCkVDezXPBvRaHbxlORfNl8gshabC8eYfrcKuNJXpFZrQtD/PG1jPR2/Qqc0kh0kKtwt755aFJW
aSbbWOO9IhmbrhXpgmStOTE4I+yplIoIWfD/qa37i84ri3ELywE7K2J0N5iNWhYlmEeNk54MZVwm
vUbCBjNnBuhYHpxweRv/SBuh9Fez7Vnzn7pSd6QJKyFS3nVjIGMJ/qcY2Ot1x1x9mOdAuY73xgIB
/DTKl1/ZH5C61YAXTEBljc62eI9SuU4YUjOYw2eNNh4JFU6y8V6BSeAWWWmwINOxZdShXKkrz4+/
uPZPCvSpa9/t4I3WTvtb2JKeRgy20U+0F1F8EnHkj+0Zy5nzV/Lcluy7a1h8wo+3uUec44ULcWIv
uxg7lFbV+dHWBc3Dc5xpeeFKYr2EU+ZKd5nZV9QA3a+XmBBWnLXeX4zeiNPt1otmjqI14uGZOCcC
ar/VbLDQPzMs+jCEJASmMME6mtu/LPQY/YjcAATpe9apR3qXdall0OI4jfzUR+gys3JRJ7Ue50xf
bZgR7usMrgZJTzmzbdG91EjwlEIwmKSv2tbVR7slbgb2wJM/dfM26u/tJIaL67GyyNrdNjnqSDw8
+eP1Fln2QFD1ehQFASALSFgwrXGd4HEdEoHI/NxmbqCa8+k/NcTZnykXSEhfBTpQSbapl/4tc1S+
smSAfoaYqhGW9dzEctiGzMXPsSSvBiKCN67ZCNXU48Axa2t6CopurXeNShetHP8yMVrBJhWQvYug
ux1JJ5215eL9/rHg1e4DZC6G+vm3nGMxJzFmZExAgpu1vQ7iLoamIDHbZcvN/1S1tcH5E4gjxzKj
6g18riuM8MaSfvTK39C2W2M+pVLLtIXIXGVW6qMEFGTXWN0SfO8WWXS2hpsveF0Gw8Auj1tuUL50
QVbV+nk0/pVuIssYUcvSEVG/h/NGPjXFG4qSviOtXM1zaQCvvjUTKI+0xCF4l0NNnKhA4CBcY9Fr
v6+phbv9e3ECqXs414scHpRgnfLJmqjUdOchnu3OkAZZrz3hRQQ9Z0vIKBQUL6LC7+EAO75i7kSY
o50Trs0Gk7/Og3w2IXCEWkfqqhp4ozwW1Ar5P9lMnOSMpPecDSUoB0xDP4bhmVwZRCluH1Uii/5X
7gZsrtOEDHeqiHm7nSFnvGfUsDKUajLmSFa5LHKBYvFYr8+6HvbsLdI8S+i4Xhe0bBb1RDlFGL4K
M2KHGyKT3x+C9ZMGQyZmlBxoKJXGsnQGewlzvkSJnZy2qxOWRYJTbyMxMfO73b2fHnZYVaTb85W1
n9nxl/MONrya6ZA0J5vi7WOnTIYg7W5swT1gFpRZkTz0EB/y5bq/ygJ1bBxATDShhhNVtiDkUx3Q
0r/v1ck6C6s402Nja4QazPVEfg0o/olObIvHMteosQkmH+Ds994QJqCsSkOVR2TUuSepzYXwPc6p
R+JpboB9af/2e54RsIi8mQIRHDGTZyr8rdXGvvLwUpehursD+OXasuDhoaFX6jaDnol6CnTCnZW6
6HJQmbD1zBnL1PiRH2DEVdt1TijXjlspXsZhbUucAndyvUF4+/L2Ilvmby6JbvkXv6gAvqJDCyMX
ZUD+nYl6N+2078eTFSGBLECEaNefudQkUDZ1uctHlG/LMhnuWb96Dx9iQ3nS8/FA8f+HpQzQOY0L
mNsmsknoI1hFR3/91oxBZpYjqrLEgrsC1FocLpg85cTfuNPY/lTTqT6YH4PhJRfgESBYdnlvus3k
g2Nwy0IO9IthgX5vb/vdIoBWlHttFWjlnQ8BZIfbbBU4FNXNNpkRURPp0LUivv8EqDlSzcZt+6CW
OVNuByYcnX5SJ83AD7sneHnPK7i/4pITRwiHnAkdpbp063pM9Ke2JXyFe08YsvTZR5ky7/KsGnCp
UW/1uLOPt2TbXFPRVqZM5vUToW9BrIQpM3lwXJhfE68fm/FNYykLRrXUoRyIeqK22jOBDRyYKovV
Qr9xgdMpTwf6zKe1dSXqsf5oWgP4d637TBoA8DvaRdaGY8BxEF/np8i+poKRsxGrNW4hXxi7o2ym
F1Ya6ru3lKBW6ATwjNB+PJreTwcerLzmhe1i8O8XZqbTC4lIMaXjKFCntvKv8Jj7wdw01rVx3bPC
gp3OsrpAtdYz7OosbgUem1AH6ABkRhra9ZR4YoM6mSeFV71c2MQWWHbGDP2xpj0gIU2kBHU5HwWb
gCunJd0lujsxorBZV1CnM3L8j7etQ2fTEJHWYgp5ksfSAZlk/G1HtUSUZZuIRu6cCa71QpwKF6Ra
rQG6oWUJp1OTUwqNzQdZYYt7PWLW/nHjh/nlDRt/kVHPHfiRo4SRNMY/bq24BSz2adPZhLECElBP
EN82/DWOvmPWTsB3WDPrSO2Lj7Yd+U9NW9RztP1iDLM4JDliOa1j0LKddEjaTqh2Erzv364ySzwk
nsiat5ENPi4EX9swtO7uCXr6RH0kboTkdwWV7UB0ekwz5MlK5YCdCIhlSNLsVtLjGEo7fssstVLG
5HWsj60dqUahnmCEVSgtPQ0GvEG6PjLfmdvHiHVk/oapfZjSME+dw83oYr8Cr0hKM57tYj2VgYaQ
uyoEgr+2Pbd7qtqQNlKuEPrv0+ibnCJ+U9tRU8aR/JLqI8cQRiDvTYUr16CiH0VuYJUXcgGgX8ng
y00sIBqWi1GrKOQGWil/TPRr4wpLKUGnFZJaHJCHIvbnlsePt0YXfdw4BWe6/fQpqmSj9QdR4SGN
Q8WeLOoMK1alk3mfhLQuQnrOaIhH0/QMOkWOsZO07jQyDe/3BtrzD3asfT4zfL7I4bEzpSatTSbs
+9Qlp45RINXX6dMmMAULKnn6DUHoEpSxj/O8K4+HHah8miKG3Nis5qY1WKTl5lk+d7aXw0kXHA3y
jSR2Rnz/WU5fp2t6lkIGFPkG3nnW4jkB+lqF7jL75AiMYF1rsY3XhOt86dOTIIubLbzQiZ6egZIU
Am+vyH+SuQHxcqacu3SmB0zXsle7Xgarrr4gSbP+aQQBsF5SBu0X1QaTiym5WzYMDMAcJBHn3tml
G69oMVfKgY0LRbxLwABHQYAnQeb90s70oT1u2JNnJrfb3jyn7GOumRrOgPkmYx4mH2JBK9K198JT
TmXJ7ccKiXf0Lq2bx6AzgeJ9RaBRs+kzDxA5wXhzZJSQwc4fArCFuKoFvrPWjur/+6NMs+uOvAvz
DQ7g6Lr2hA0xhrm5+ym5gkQqUBMet11RJzdJOYERPLk0YDnTNOQAo5a/kWb/z0zotmFbXUHguYj8
ZOgI2e3kBRCRcCkidrtfE3KK50FdsrklWpItAb/3Gm/sRgT3ONjhjPR8AZBpZTDZCI3IkPeGOZ9J
vcItuGKt7f7S90sc+RItehgCsC5UPu5PDdh3YpjP2R5FO9lOumcqngHk9u1vwuztanEzDsgtDzQx
gA8dzkQIrqQ03NGQAvugpsl3JeKCCVhIxgacibWB9wBbi522DqHTyqG2/QgsmK6IpWFETJJ7rUZL
gVLG7Di997Q4V9kEEN1aBaYR+8ehDqgEqmyejNM08gf7Qv2pDgcbDjqDFAmL6w1AW6eoBKd5B4WS
TpDdDEali8Nq9ibsx+JEKI/gKS9QI1XOp3ZPd0Zt+Y5DhdklRazdY7nq/WSIHqwB+9Nh8AxZv8ln
3CxWMI/sggAQ8PKgft/HsjBKlVGPngpAv+7ZMJ8XbIU38CrbrKGralu27lMTl1tnZIAvIbF22mJj
9AsClwiD2LF7+PLYlIZbD6/G38T74zeLx9vs1MVEJRSvZo66k6NaP4+T8hsMUEAyggEDexm0bKbQ
DYsPX/MsX9+PWeg3b4GnI6OXQzz9eRNWC3fFj8gcgdBG8YOzuO+ZW3Y1M7PQk0w85a4p2oxYl9t9
hYttP3fiJLfwvP7sVS0hXelQlLajKr3LBjw/5DXjClxqqrkDb/3kbXiBZVuShlwlpo6kdbOx58ug
2lXb86Nb4H11NfsV+4o0ZWqSlmE7a8yKQjg82sRvDrQw53BcsEfOGk2HGVAKvwf4snjpE8TJJmdI
lCfTtR7Ywrua/lPyDdAHDQ9I4M0r55cgoK6p0nDOHsjee6q9exN1tqeN19NPH944sY92fzpNsA41
oCFV0yecicJtBldtbgsIBuaHPLbJ83ON9P0lTrGcneyerzcptuQs6DKQUrOyRwunpNWKLjagmXN9
myommZFnJbLGr1BAVXmCQ77zL0YiofDKu/rYYS4829yTsotdQ+46UWRhBuzLk0ZRg+R5W8h85zHh
f+qbLmWITOQ4L0ZIEye6jCBR6BHjMWfpHnsK7APajRDs3UheKwZ5EeGjs18bhgUJiXyk/IFCQxmZ
oiLJ7zZ13PvBSYVrvZ+HaEnweB5VxbHJUejf5tBYueKp/Tdltb7iCGANSmpXhvUocTkJ8WWq4jp8
RsWP7HI3ggrtTGISyap7vr4I3P+7qFWUzmnW+BzZ2bgm53JO5/NTbd0md/BrvEQ5E0aPh3DHeTR9
GZlKXN7tguysLA/nwWuM3TwfqQXfUNle7Y7YoE8Pl1hmj9pbBrK6V45Td2Z9KEXfg3jOQceZbsjb
NhD3h/HEBrJD1IrI/qUUtE93AMSThBm4O28eq3RzSYrmHcZ7d6G7yLwalzmLYad3oXzfSfwcBqtO
9ELY0UfqojHoXmRHrMRZAbVnxbCJgrNIuDJVNFnnUs4n9NUet9I+iNLkdrXhDdtUAnQbbc+ttwea
kKMdxwf4MBrxfRbkWVqwynqH52LewnCKY23vr1f23jfOt4CHPMPWXKmqPM3OJJEhNU1M7rNusruG
4zHqBg0L7eL0XiMpMJ3cK3xVwKK9Vf8MmqdWTKaZFUoOVDuasRwoqEzBZSlUfT9YvKZY5/AIU3Lt
W7akFXKtWCVTQruSAufRYsEzvDebe44jOLJBw3YlJgA9wJp/Ya94r/I7o+iU4cGVLk8z1vmVN24u
6LiWhcIoKOCTItxLD/4fjb5O5aPtjoaXWeYrhgrc0g6jZRM3oTdSKz6Iid/knbui8wj2CwJgeZDn
FwvCVcWKXpiqZd/DfRXCFC1s7Rj2ascKgD/La6iTzLbJhJOrUg0+LEbDPPB3Z2XUpPuwkS5JaOrL
YWwGUwYTCtZ0KXxNKumf3T3MPjqvS0Q2123fjV1bos3h3M/ueibSDH22Wwimm2H0cTUDBU10yzL9
WH4RLaZxRTV26vrCOTbgYuexdEiIuTtel2QfXbRxb2LaFpOUdzfVL/DYEkPy1Row0xlKLCapg+h4
vnS0S2UV5skDMIEgf5rvMuD9zTGgX/h5SAVXUun0Arc7cRXy3NUw+xkwE/cY5bQlrYjjyPfwsyIR
m5b9H6lOC+NRM0NhVsbT45OxUB65A2nqSYK6K75Vx9oBVg/kEOT6mgy18UtECUXnLDZtpjtAOpue
7SQEe6Dr2Q0vtz6qiZyW1OzzHb6T3QLA7xsl6D5GhU3etP/4b2Koxp0OCLz/J+FV6T7u4LsAG6RC
5pjVLnXlWhNfXzbnO671ZhYyVZBbUPZeHsmbQXD52R00sKneV5sv2qsAPHTYvKe3t4PVWVHBF5iM
cgWDZ9YkFR+yYTyB9l7Dh7zqlVZvDLH2d/dnmPDWyj1Ob0BLUD1wXNXofC/m9+6Cf32L35FS5dCo
YBGJNfinwOr/593JmlcjNxG4672NbzCbscIeVty/RNR6CSY04I4J9GKe3xk8cEv7hdDyesfgH4RQ
/eqH5iZS2cQ4zu3pIq6Of5QFMYHyT8ICcTJ7/p2/djdUn8eeDOkPR0VsMzthZA2/7qxjphNdoRFk
isTRsx2DuAJ/V1fso+iGHPAa1+1bmY/+PWKl58aiZ37nKv+bGoG5rvWlkVz8x9D9wQDRxVpWkkkW
V/hM1bfrO1g8Y3c6l2gkReTUGVj28gO2afzMy9byYXMPB0yWv+BJRwRo3qPiRGmtOa6jHgCc+4it
qRnR3WePnRQthtsu3pD2RouUIECiLKD1Meq31U5FxfFVam/9TFBBxzi6JmsxXkduSEXILqJj2m35
h63Ww+tnXpGDG4eceulkDxja0x2S+R9OgFKgWkgdsGdZNeiX3lMwoKPxlj8M9B5fyobfikYf3CQD
hDIkhkuGJb8LIUSnxYu/S6LTvwSSAHeietme+nyxc7IM96JrHGIuunOoRByxSoNZC0RFUZBtSuN1
BSxM+xNV/yx1J5ZgRdrEHvHxt8HH0mcXMTyK38D1mJr+xjVJpUwoEMbIBwSC1IdpZuoHjIrKpamM
uJ4RuRoqUsqIcDQrHFv0IAixNXUTGW5B5fGhPrMH/nCv2K1T57E0tqVfAc11hd5WW2p4aeeG7MMp
R83q8LOtDMoRh5S7TPmkiMEubS0xajou1IuZs5hYTekeN8i39IVqYlsjvSOc1q+KyyyLBBw1FgHS
4ziAfhhFOxJ4dhiQq2ZWx24pMGs/wa1UXalsicYhEeTsNk76FgCYZI0XzK4juVBbyNyQ9k8jSWoS
pGaeoPAnAZQuTf05kHyzmIbAjvu4OlhN9ZGx20G1pxJQTtcZdpT508bDKQbTBGdNlgxB6HiWvKfT
iQEakz9+6PspfyaWFp86DsY1qCKc4QLXHLZuQsHoN+F37LQNjbpghJbVJxdzxHUHGpFVOKzofuq3
XgCvMDxFImK2NwFlcfPc+CT0x+K0F5dBLmJ3xDTe3v/DFUQ34rHbkpHPFvTjkVLcbFdinY+rZZq/
G9mJvEeEMYWLA9H3dUYN26LFuLCcBItIk4z/gVnpZ3xI7QtTa+8LWOS7V7lqzOqHkFNHAZnbTIq2
sVSq53U5P76CDz3TAZtZ1d9VDnRGmcHq0EroBhz2DFwQTTMJwGuOpniR7OcXFyq8RfxkiJIe3Juz
7HueHuqClxaBxtRLZyP1+iUKW22Mz0rsxzSiP3GTJwmDIwN57GFv70GSCd3JWi/duZRTJlVaH55K
XNvGupEjQM4ImQ50SVjnXIIeiHzmzQ6oQHtuRWSQxX2oHo/mISS396QLI2NZxDAkoybyHuvLX1rU
4f14IHvHGguTPZTw2taWhX5e9JKmnROeAjf+F63CP0JK63ctqLPGchAhiX7Tx+54GK4ITDyX4LRm
g3PTEkHJ9L+9AkDWmcdGQ0muUX3u6XlhNk8jqQnnxPvP3bNUeDFe8HcOUEHgjTgjVnwDmm/qZhpR
KI9lf0k6a9x5U2/0sMdVAWlu2ZBMowOTB558qMI+R/sstR15T+CehCHSXoVqFF5FOipI5gI4zc87
3e6cKAdIKfFKCy1mp3OCHyu5oS23GMKGYh6LbUPLg0EJjqs8seLnCvoM98yJpUe0Ll63Hk53F/vP
yAE3nQd/a1kG2hYGWc6Iyf/em5YJMfVvaBjMf0sIAksDL9FLYEgGtDXt3kzYbtH5+UQhfSfDfs+C
AvZKZCz/LJhZhx2SiTFObgOSwY2MJnfNegR4BwshcreSDj2TKw84f4Vx2w6Z1iB1INKFybFKTQOb
dyW6IkBKo0NUma+QAi/4k375DR63TYEtxqNMrn3vgoVh+WTTnovaY0cRaVFPLSNlL7tcP+8T+a9R
jh6BlxVQmjd5azz2lz6yLFvQB0LTeVOgkKTfF13ThljPPUlZ0b7FaP5NaZa2c0hp3iZa7m1cPYgm
4tZovgT885ZTHIhKAEX1IlZHZuNIMfNH3n0xwo1VSnkGYmQCPQICWpsTTiguRK90/P4ZTdZhUBMo
6Iry/uSO1KsvhFCk7qXKoVNMeNKpZ/e66u6pIaTp7zubl4r+RHtMTdUOAkQ6D0IXRAu0Q+B36CfQ
J0MPWNvfZmGn7S3jxhIfZGmTQQPfh4bnwoy7iHlVhXq1u7LvS95Nhqzk/qJ2vL53MglaOA1GV1IV
7j45rOlLf1KBpKitegfhZR6Ppg3/qS3qgE3EqNXoJndd8uH6ywNAedIs2fst7wvgYx8Guvr7K6mU
1G8VGn2NvE0nREThln4XXdhHFb0fguLDPYk/NbIvrjUgqbfMQ/MWPRno5TtWevmGqCqt0fyIKglg
PaLpHBgmndf8IcayMMB+rgtJd3dD2H+avRN2UEjzsuTaRwMWenNHHdP75SWt7vtj1eybRDq/xY6d
H82PQbJtCq1hAw5uIbA4V+zBG12Yv+uekonoM5a3sZKkpS2xjqubJGmL0wXIdgq/Ujn1pxzq15/6
Ng/+ZbTrVvs5a0DI3vImRVuiQdf7gv/CDgAOKcowWn+f8xu2Q/YfexzS6lDu4tSvWSm6gdSzkWrT
bI4RQfXDGrVkxgCMV46lq53Ojc25FRFt8lUNoT0J95v+uGk8QkQy+m5sqoHTk2BnY56iQ/6QzXdA
JF/cfel12sfN6gk/Nh/24iSnZXaLdZYP6T7oJu9eQ7segEwQ58r0P8Zqk3Q5QdN4YeSzycZTEYIE
DkugABi61kU/8t0oeWd7wfmr6mhl4P6iRkA3favVIydTD15HBQxFSfvhfRfXh/3uK7sEz4UcRNk6
kML8Ey2xCXoTMvqNkPU64VKc1soSPi01V66fZHd6/Dp5GJOjzV7wJy78gjO5tzHeMSfiq4/s+PXa
d4eRSSZPvuv85UFKCvB3iNVP/GO4+0I2s7FjIgWOA9lfndcL4GWrMPY+U4KcF5yCNL7p4WzOWMVY
jS3Un8jG/dVLdFnScKCOft773Most8rZKmCQnl4YtusKpI7DWgmZ4GLxus0XcNxE1K3nZNbCrQ7k
VIiCWpiY5c1NWNdcEq6gmlMaQTg+dOzh/UdgFhQOWOHP+C6nwmv2QuVlAJqzegVj7Skuhnu4SoaR
vwq9BSfEswqSVSlZNG/F6tJlT96eBhL/YZjASE2VU4qME3DQkONZRBJrFomxykOzJ2jdtm981LoP
o85N6lswn/3DM6f5HWqr1Nuw5pFSSLYPLoGRvIkk/KY/PuqHdxOeo9E78dsXxvGVtzd/jYAGC017
BnlZBxZnSJDrzVArFTTWe//KjUxKrqX7la2l6p3Vu5Z/XcRQO/pyjF/IwiepF5x/p+eY1o92roWt
7p4jlPK50KY5aG6mTVJ4GRRtuS16EUClywM+mZwaP13l8vA1vmVAqLhLQ2K9Sh9tpUztaGG+V9t9
bR83deqFUvpfDIPAaToHFHhqOvR0/6jLK8o7coy+uudSgOv6O4/vxFCE5lff+HMdG/FEuVe4E7pj
jhd7QLNzWD9Mjwcj9ddhvI/U+ZOOrmqtZ2qj0yudeSK+55+vmW41V+oq8ItYT+Hb5PT0+biLIq3v
//Km9ZUFTxtHv05JTHjW/8dE/SD0GriQmOQEQH2jWCsdNHEkpRPB2l1OKxU6ANIIrfpLjJ0BeOp4
0/7qg59G8hDvj3TlEfimssOJK3Psxn5UfM3WQifG3+n9rJyGEB3Mlh7FERkbSpEo0AP6ZLcA8e0q
IUJdWr1v6bHnGQIMDg3nIIvO+l7Z6qhk899LRqiRxuOyQgOE7JkeVty6fxC7liSp65qnVNaA0CA5
WyOvvBXfK8I3a2WHsTQzyuDfIUx3VQ/G1T7N8z1TWx/eQFzXsS8nrsB+XibsoB4tv5Fe2L/CMJsC
Ro12fVdlnXtwNmeXrQvlkQb7yF9V0PZ+dThVhLtP+Ylq69VVbGwLKPG72wAW860j/hx0q5EV2syt
EGt+kYcblrQFvHRwxWgQc1hsj/evlpO72PlKY4UHSNGNORlKfeJgZ5jl9S+nNlWyPKkJDib70wtz
Vzjttf54WScyKXCWRFpDoSiniKyONE5lQP9r/oCPF9TDk/nzW15A6GqIhGMUXwlHmC5rbQ1CPujL
3VspOWHIvbXKmOcqZRbSIeoH9XxtHMmLwqhaam2iiSWY3wiJSx8aNJbx7GCBxtqtRj77r0Kyh7PQ
cGTvt0nN6cqiC2OybHYzBrM7tYm+nBfyEXJVs6oeoXyLYSplxm8TNAJ+Vpull5a+nlca8lS0lQvb
dSwb6Km0qhdsg/oDoh5XvRd7cg/CrZCEhHRV+2ZP/0wm7pw7JOFVoxdtr/h8M9+6gOza2NiROyI1
zCcIBiPTGlEbssgKmNpSDqQEJUEdOF/5mTtYcZDOD7dhggG0t58NTjuh+aiBgVz6fSdbNLdjP6q/
8MQ4Mrxu8Y/xjEqPOAVynKuQnOBDz1AAs4W4m7uGtERwnpnwcbRKiV9rflPf+A4T8jr/B8siDKIr
9EzDzg1sMWw5+S7GmB7U40SB3JQd+raPsF3hZImpUhb3ugnpxttBu+wqIAckZ8l+Uvl/DHW8A1Ay
N1aFqqdqvovetgyXMYaA+Zsx+mRyGGTLStFTo9zhFX546CLfxLvrCev7QOO/tg/Hv+vt/7Bx8yAL
128kLxULBXO8VLRq+GqBUHozxunI0KMMEYhJRzwTvAiCqSwDL0Xznrr/S7b2Rr/1XfuVM1naAuvN
GBXvZXr5nlGgILPlo1lfMq46/drnfBhRbg3Jnk+dxIUvOBAdHUklad2R+Doeyk5mpZbwh6P4yqj4
YzHS/lRy7KsTX+2gybtraz6MariHhkmchU2rh6h5eIt+OhPxtMyrU4EjkxYlFRMLxsRGBHowlHNb
sRGKeQvdKCFieNpx2CL5zNvKC2HyTanDxeadZhec7N6aYBgkVKSZeSieMRdO8BS0KjAZdfN9a7pZ
ig6bRGVMdeQzpLYbUoP0cA1YCir1GoAx4h01T9DRPygH1ebwDNsnfTzBpKr0giQFzMWIwYHs+S+v
eAvM+MzsI4pKASaRuOEtKZlwW+jsMy0GrE2OVFusTjbpFBZkH4Z9gQU7f3x960Zh/xSepmC6Setw
2w/c+T9AoqbCj1akIsMZjvuR/0f5kbrgrXI8pR4s6kwJDIfOBmpFlI1geQO63/zkR685rwY4c4q9
zhbnfl0ETS77DVrjFHB4mVuiFEUuvQhu3rGAbCROyzCNDIMG4VwesMCR1VOnBAVowKQpYGWZCZtL
sI3+USZZJU1CL7v221V7i6y+vqOJfRoQcXL0zjTC8xKz1cywlU3Kj7GRG8mURlB/OXmZJL5lBSeq
+6myXLzFlKsMBGHUt6HMcScqwBWaP05hw7bGC9BVIOOxtN+z0ngL5QMCGrLZnDdEauw2oxFJ+Qij
Aciww+gcCL3U6hVF84HZmXnBLCSkd7wUVCnAmVUkJ8+JRiVO94EMo7TGuPbmcq07mbKoo5g/2xGL
A3LfrLQfP5twCEW9+E2MUIg296VrHW+xUkHCHxQgmMWujIWZQVJ7po7xevjwsAhYnv9VgQXiQrP3
xMtdJP12tZ12/oz9ePcb6zR1F63JgtDPk63GnKYbDelFfVqBbnL+KsjT/3Ha1GyiPWxIvA9n5kcv
NJKBuya4Ubh+jVDEPPWKHmiXdYl1ZL8/lsz0cjmf+vMzH2LzphuP820wrMKB4hgeQUoIN1BtG+Sb
J/g7N4vnv1sNmafN3a3mzKYtNVjwrTC0ZGiXZEM8rZjQ001wQnqsUKoVOU1E23oYkVgLnReBLZLr
g2u1sdcn4HAAfN2Hss3VnCodDfpcT6UNUIVno9kXJCaoHQfNVInBdunFx+gQr40Iv2jujp3eW+2d
hyoue0WmXMLd/QeZWjZiP9rJMMNNfAfET/+LYeHDekjjPhpVTjkm5ghrScozcznW5xCOmX+43UaY
w9Ty0nnZCVQuwIfkPY2WnRKO4WcB/AwYBRNDInh3SK2THglr7dNIrorWcute3xHe4onIhokhRTy8
nf4L9kF6v2ZKK0TmUFs0nvrXDhK/E8pHBux9Cop0Y8lNiko66xtxRaSi2UCsYhExB3I+Yiu6gZYw
AWkp0kCSy7GjsDv7FUtdGqr1JrnjdyD9b1wGjPCrtFolfAKS245OydVAt7HLzOA6VZP+K0sbyaWU
i31f4sHXjGu6rsgNSAll7ks1lwaqDg8ECKkVnxaj7qaXWhzJh9EOvF7eKRg6QLAd/YzjL6/8vJjC
rtF5fm3+t2042fo5gtFzyXIKEhg+t1LwIO6IJxNE6KHvdBbhVgyCA/pnA8EsRnQQMe7da01jENj/
qmmXOS5QurFV/rdJdHv1uOkM0FC/hAgIq+facIEgRHBAmj//6IcMLDjKqnchPP8keRYaxzTSpdqq
l6ngW4Mb4kv10DRiB+gZ93KsU2x9MbgnpCJpaoIDU97LMWjwdf6QukONzprzO1KxIhaaAC0hGwHa
7kCSLlpV/YrsndyyeOA7lyI5olm2u0pjCxaepTPkfvzgBEEEgB+nvvBMJ1K87RcwHZzIx/x/N/gZ
g2pRreaJVhPuwuvUqP4VS+GRCxZzwxCEGVZRfzWHQIYfsPG/BObnxtrE4crTYxzwi6MekNF5CuW4
syIa/CfS4SmCpxO16twPWpoA0j4E4FZ+NSmM42j3GtAOgFCDZD3+sA/WMsYD889eNqbU8bAnfRtG
VuswZM/UtdorKjukhjKvIGPs6Dxv9KdZ+dU7rakPv9BhXV6l8lPEbq0rcsU95lL38vw99Go3y1Wr
2CeEtfNF4Thylai4C/QSYdIWiHDMrBmJNnonKSsUoGay79/2DgaZgRtaQpDOQlcIsCrVpMyaNFX2
8v4UkL6xo6wcm3Q+qb5FXHtnrGd9fFL+Eu+Gl44vGk4ptl+hXvj6CkcCYFVmFIgEPTxZuPGLDWsF
B5iEuaBkSVwywxKWEaBol/p3joSKpH0NIO839aU4t8QEYx/x5Jn4G1oH7xkbbBFwY0XMaTlWYDJX
bXxHj9/xrFSz8nmDiV/TXqu1LfngEQlXh+c71d7hrFonAyWWaAc/Iler0hlr1Bg7QGb5v/H11OJQ
l/e6Uof10koJ0HBL+uWWsSMDWBSm5JwOwESVzSHyoP7YIXKzEGnYx6Q/RUZRowHvswSFNI/GUI86
/7oRa4c6m8IxQVfK7awkZyxDIB8vYO4V6U+y7Xm+/sgJdYtNAi3es2A5YSHtAxV391sIlzeUXIMp
Pyw1F7F1GbU98+OVwL2jKJxHC6B0gRtQ9I0/sc7LP81dpDS+jMG8+WolpAoupyoTuG/F06B72zdy
k1b0fNsEHpi9ChbvjySl1vCK+nBhfCe4ANgv9c/97JaViPBObVTpkGuJ/whnzUiiLoCRSMa/GxW+
qRYAu/da1UnQJochTD2QJr70l83gNR9QCKrQhS/gW5bWJX5By+kQ/5MMcWnkbYzW6aq3JMguAG8g
YCGdmqMjmHwqqzC+/5jjYeU2t2mmqnM9vF8tM1/gR74C3TOHBvK0+/VBRh02GgJGUBM/SAwTAxGD
SidQlUm5HDjwnVy1VzlTsf5CjoWzPslWoL0rOoZxcDIurfPdCVL695LNUkHaP/feHreIVtVBJpUt
lcsoXtcsig0EEj21D/g2Xt2N++NGtcJkk8h50SKkBYp4xMa3sBFJuO2vmpY9/abdRRl4VzpLN9WY
yCNsN9XNOCZe00ExIoYGgUoA9TO0xugm9dOZMbApoOr6v8FKMdm9wQGG4br9T+lTR1ipbFHIvy0u
P0nkIkQXuE10jiJXmgvt2n7YJDyhKnd82oLlPRaiJ4ei1LGjcE2GkWYiyLXB/OYNimyjOue0fCpl
q5gEJCDtD0MtVkj6J3eREKo/Uovy4+u3CeU8uW/MmI/GKLxCBtzt87T82zridervyzuUFMbZDcIW
VMBOhJUukq5Fg49JP+Sa5FJr56A/cecjohUTZbtYmJr4aDKFY7fa6mn2U0nnFfTit3cGpqEx0suM
L524b8D3jATpbnKYYI+KVJ9O3SijJhRRYgmKktgVWYiJ8Jaan5MmioBD5y0yLtw3UDuGsSAnYqmK
7EL+PFvI+1Sx20Cv7/aUKQpk/erVp5vLx1npeohzQBZ4TiKGoLao2fzNjilj3GxA6nrGUnNILk78
0ghyJumyC+IrHjjkDLvr46zimVIn99naU1bRvUW8/BV4CCp0G8fy0fQ8f48p9oBcqwg1ehVnYzQH
YzEtDlS1E35b8FB1GrtnUsAIKY48bA+DqsWim8m3DzH0KUheu2PvHbfHgICUXSa6A0AbCPuGq2ni
hWYwlS/1/2cks/N69sujogvC2lskFv2r9tnrGoHlQixeVkpu0OywwQBeHZzb9kDUfqkJXsXL0RjM
yCOYn7m+hdPWkrOiN66RqbmtLVwbpKDLZBWoKHGisaa5lkoZ72BIDVysCGK2V0/Dm/2w8nyh78DU
hFsYEGvUbOXRA5nrNlYGlG7QZ6/Wwet/TjWWYSBwsj2vZ8IvioyP097eiv+281Ss9lQ/yPUvMh8m
HI/BleABJUsN7MmjY70WsmZwyWD7E/KBb9eKy0Sgg2Xpq9lh9WHRuPEJkHlc7G9MVrM9iib2U6TU
eqzLWoTQtPuyb65MGwy/2ljBPMHbAyrtLQyXdyQKAmTUyaAT+U5bqC0sdAVlUIxlCan99f2RMeyh
v2mxFZW5NNh8AgBi3gM4m8x7VNSvSE5dAOpk+5U3o+75in/03bJNwrf+JDnh/vuHM6AfR8+VXKmh
Xiv9UWuY3mIDK+RkjEV85oQFiYIPNCNnKzuOHwGQtAQM5XSJWhT8/Tc0YGqFDfl+9cjhVDpKhge6
9YKJEv4GJxsgaAK9PVAniBV7i7r3H04IwreoXmp0HhKmXLYYPXk92/9KdtqLgOwBDDAgfpAJd0Af
7XBvmvY+kzGzD80gzzWMigOhSsK7p8Jn+YFfJeRdl5SAN72hK8MrrQ93DLMukUhXXeZqeoKcn3Jp
7zOIwxNRAnHO2i//l3uunA/YuVNF5qC+oUzr9MmXcAUV2d4Lrh4523udqQHBVmwLyHa9ujxoNixo
j1xtXRIcqApCtSkLjOwMPwCdJbL0ftE77dMC+3xCVNfH0204J1PXbSFig0rKoohIewtS2S6A/dB4
9Zmh5hu81x2Zufkb4w+LEkwvv/jOQ7kNQHFG5SwEpuSfMORnqVLdt8+cr8zAhJElfwykEqgo4x/v
c3bwznLp+87iBUuAcp6lfJCFsjgfGBaGhXAzLZhriq3G1rAkphuJ1UBh8CfzkIOfiTBBDO21dh0g
Q5OkiPpk8JZnG34LFT5cZmtDjF94I7iCjEqOdnFBHylxnAg9fFhbum0T4M085mj3197I/WXdRXPQ
S5JoRzx7BCcrZF2J8vIzJ3beQ1qroN/lahlCmV2OtIojeYGc5loCvGWNvVCily/Q5DbIeahFxAjc
Nq2p7sWC+HuHERMo0jnhjEkwix8LwSBV12FTMlmIEkCYzaGZApgnfv8vKFdlZbM2hYKYvSUQ1bnK
ig0GOxGlr08Sed+KVboGshFfNdB+NnIJc12jTOEmb+v5Ets6LaXZznk9dKJ2g9fOLwA99wsVzkxp
8UtPBvs+GfA3mcb2SOz7egIfU1wcOap7hzaI+U1ro0MG0UCtMvMmlxccTq6AT9NAQrHNo0He5sPv
Cd2PmcC0ey4W0p9Ovd2KuvOTT45GU59VwqGxV+vm/YusaWjFDsMR4TJmWqvsIO6xCBdoNXJxQfGm
cThbtDhaxalCQFrEoV+IxGF5UMVFyftF4hnglFjgFnARsb77Z5SwVyOoFJMRtFvIlOxWAv7osFCO
QbNMoptOosMudYbalAAw5uoICvQd/qACFjb0txmdQr+6+jrTGexR2mxnxQwmPNUqlWBfpVfuz2L7
f2m3U+8KlphhZ2qsj1dTU690o3UO1YAWEgcKYAF1gL7DAQmeJIPcWMTHFYia7dQxEgpOdvnhw6wC
jsx7Ca89W5z25A6oH0s5Rr1XGNCPkQdqgLy8yibV/7uyWdiXA3lxlWEYieY+N6ISCmpO9LMDR+c7
prQKSDHelw4FuGeJ8+oPC+4TwzttGsmCpTqIr300ZOLURdjWBDRhbMKU1k0lgvfAPUh0Z58g+Hb9
m/Mu8+v4P2vdXFA6/3V61E2T9Eo+Hg3W0BJ6TpJMEK9MYQJjjfV/HO7gpxEo+OhEfcD1nwg6+9+O
8PIH9uU/BtZa00vGkMpH71FwPYorUxg4dLo+hTZ+wlZVkelElHFsUsDJSuuVPV/ztzAL3azKNyyq
6gCDzheppm2OUkgzBH91uYRN9BsQ9mrV4VUZAvNQAGg2J1KoVLOedGrkg3wnybX4T5oEXPvQcCZw
ykfW+4rXQAY40wyTFK0sF/aHHk2Bs+q2cvyjKLX2kiNcuetYkJ19AQ201ebHG+YPBfsLOIBOOAb1
ZMDTGxfFuWqky26Y+alC59tAy22Gl/nUm0i+ZfInaVOSHs97/ryvY0UJWYabrOKFxxglocyWcwDI
Z3htoWXvawDD4+vjxcZ0nyRdiqb3Age8XxLuGeU/9DfeILaape1fSBPBx6v5wI2NMhJ/Qc38Y7lm
hvZedn9+hZu6x4eAu2qBa4G9nR4z4954Q3MCN2MiB6O6BG9xB3PjIauM2N/pI/E9GSIFqyb/16fV
Y4J4EkZR8fg4PAp9cBbgs4iXiKYji/jKrTsSpx+K2iz8obDHjxUsSgNds7B1cu4OOHbbCl4ybqbG
88qA70HDcTjk0N7J6HquGkNvIi1Y+LFsI6ErB85u9Ao2L4D+KibIlGNIAxTP3+9f43AcuGIYGgEj
dA3nMMMSCOOLM0RKozInjmHqXFhcRR65hUn2wXwG7OJ3TmNTDvW95MLSu8uPY1haSyxvKGyL4MqQ
IVsuhsR8x57UlnA/QrNS4ynkHWkXyJyBA7Fx8Vzi5mAc7MxEUAPjHK1Z/GVTjsl+ya93Itsnm3/4
hDIp0WYj/bWSCoKcy/2BVa4wHaF60gi4kVRNuSMaXXtvh/0kriGJuID5K3YkQShZW9N6FzYsras3
84TJ3NHXUCnjWUy9SSDN87j01hAVlwpBn52TspGLA/unmLFM4rFOtL43lXJxe7PJ9dr+wUyG2DTf
jlE158zg2G4I7iaIisDNjckCrFB+j5tihtehU/t5cNHYwCQ/ixOfpEo5zQLREVSCWPjgas4JyUSB
aMnw/dMUgHWrUPCm7btgLVbfQo+0Io9oWrE1VJ2ut/o9UJ4QPTp05Zmn1QAwj8rUKs+k3HMyQLCp
ygc66RyfgJrz9DOllZFVHi0LwIdvinjSbZW+Eo8jLk9EaD/JABNcab4qQ8hWjCs8bkXHUjMl+ab8
yT+26t3W3REBIxvKxscvOYDXIIhjx+p2MrzUCTxk06O5tE5Q/VuCAzQmTjdQfsHeSk3bfNAWznHj
4UZ4cCPFNAH093YXAciIeWHkA07MWteTS3aV1uWk3IORQzUl4AsUxMWfnRNsOqKP5l2Lj7/6XVkh
A8kobCdFVgrboDrX7cp6oAXIWiF2fkRy9i4euxQGRAt6lAcT2L2hqrybAdoUbDZeMpdqFkkfUo8O
cTZxTllT/SMYFEmIsKDRKKltP5EsyDjdJHkTQiUBqNkdmtHJJ2ElpL1fdTYCO5sI4FqPGzBBwnyM
SD11qBHDDwEXVerkso5PE8nVPE1MpEahkdedbynnJAs0rIVdfZsUcMHskGn78bRIllAo1y5FFi1G
oQXrch2L4tS/aOZCGh+gBHBjlojLAG+hVM+mmpQImt6e1dZVDX/Ab2d16WEs8YPceAt5kgmTUQDs
RU0YAV6kB2Vf6XqPwggXInfENynqCIR9/Mvqalvsc8HmynXdUz6gidbkbOhJUoVNv8EQ5o7MAxn0
y13t01ERIi+SluNqR7xSorxRskAXccWZTfvk4bu6dPfP26vKQ8x1H82+RM9aO7M7S/RYmpN0TcUB
QRabwYFI3wqKda8zRHiHvBhUcTrjc6PxODGJ++0IlMTNVYnZCUVvJOgWwcfnTyj1Nmft3+EoEwrb
ofhPBTXTt9PS5iibKVtJaoFk89Wnm+zDZb/cRcIpJ4YPw3Ocsg0bo0Plg5snKJ+0zaOMPQzvXjy7
7/mJn19g0ams0VvGzi7hQGyVsn8oqMK0aq8zkG+ZrVqetZfv288HO78SM124lErf2aQsYClKvBuQ
egHLU2EzbB8731dC0BN51lDkwk5a/QkVE3+fb9tMrtPX1kJayx2YqgTq9D1YmkY6a1cRlhV5OBzs
3pq1RztO8w++DWSemO/eBR6ox817H2/DQMLZXgX9h8UkPNHbWvD33EFXCP3B+evObu+BhyFupnop
tbo3+KrgeOlxdqfKqTTCeG3U4H94EGXBscWRpmH35wY0c0I1XxkITKNQpO2GWT9vsagRWa3ZWcbX
KLSe9LZ1qIf9W+KrpbIQN4OuwvpabiEFO6pt1bB7ilzbvlVlSkbSUR+1SARp1BCOW3Ja3GXI4Yhh
TCwnqYOlUWkkrRyjJZHWR4OdRl468PkpCSYkB0AL5IDAJLvEI5rzsPLtlS8tXPphLeQwESCmA98r
GJWedpaUVn/0l0nwkAMRw/GNY5D4OLMhUGBprtsImehLeOF4wQ7QePJR03JpgQnj5j6AJE3BJjTp
xZPOYt+Y4Mn6PzPQY+Ta/aH1w+wIUhsXGnJk+temCGklA7+8Bc/k6HQ0iDPtRiBw/8OwffmwZxQD
c6NzSbCjFcr2QBZMr9CchjpZbBcQvbKuWai2DkL3vJPXOpSJdJphwT4Nmp4kGZHJjsxTD12o9uU6
VZyFq81UfqaSyN1GH9Wfh67vdsBrO5jt8V4igV7zvOlFcwmSwJlBRNkR8d3Ip27pYEio+jVpQM12
8JGPEo3Ry32GMlQaz3r0c3fySAxMPI73FLX/sNx4KIUXYOdlTEKec5zsq0F9ucxogzBavCjiUBLS
Xypo42YfcK9oIngDS2i/5osAPt2HeTTzn4ldl8+g8uqPhCkhyQCe5iqjhkbCS1whvgg7egwdFYDT
ac7B7ackKCIEBTLBeD1UaeOKHds8vWiM3jjTSLd6qWmn3RcKzYMltbzJ41eGdrJW3yI8lYi8qVXg
Rtd1QBBHf0rweh7w+znEJmsDv8WEN4uR+NZIMkkhKvSxcoHzh4e+S8tUtfm1AQfAyb7yYp/4UVcv
3VjFmjFSVj3mQXu7zhFeoQtRrC2r02zQhmTWg11zbs7kRiug71+O4k+XhxBqvQ4invgti+Ysr9sh
DFOV0EOom7NA+HcrwcbT7FjP9wS2//jm0tDmM9HY3Nat/MKtCSQ4f/i48M5L20G3l2PglR8utD0Z
juFG09dLpIm+T0uOa8TDjqMmYI0tXVMVqxe16tCiYiyD0Q/HVadsVLsrdk5VdKl3f/5e5dNindQX
QqkNqKu6dLOZjsR0Y+uhvG5UPlteKF18FRSHXMF/BBQK9or88CtjBAF9A7o0Om9JpOI4HhCC+gJ8
3lFmL9krowUtxhTI26jwGdFlmvwEfcc+EqhEsBJDjGnTt/QbxAXu8wBvKpljrlhNfF94mQfP4Mgn
v5GAHmzbmOEE0xaFk7Ok1FXjDwrAMN44OwLDoE+9BJGU6DLLtt0Y7MRg522vJc9M1QO8tQWm3tIr
w7c5SpBcOfQyLb09F2aVQHtrBZJ1nx1wg10DHhUodeAwDzT1ooMbZFWYtaDfYCGTLefFWXRxYcYn
Nldl8dFFvl/x1UQJ1mfdYV+IPE4wWAbhU/ktAik0s/Dv/SjdcyAiGb9Ri3Kyb5AijcJtRUVCAFbO
WEdoXF8xF+JWLBI+Xe0Mcmml0mzfI1/LeL/81AcI9LGoFHQXRRQbFqjiBzlVBfvsJZj/3+CpP3Au
Up39CG3XpZ9tFnd7zNm4HFlJ100FKCxDKy4+FtZ66xyEdowJWxSQVR/D38cHj7+j7oYXp0r5M7yA
eLrVgkaAdLfde2v7h3z/xw4G0rwc/hMTEYwcWtt/M0ZHEWFryQrDgelx+YIwB2eLILrCX2tuOUrs
dJH9JCi/1jSMeqYHEjH4rJ+OpMMzEedToiEVXMEthMfR14dMKqmYBbBeJLPJ3l7aN7q4ZU8nQF7j
7f+e2eO6qmPuBASWr/f0DEFwWnyI5x74ijRmVfaTU2mOyC8uoKO19VZvhuZXDZKQJ+gpl4Cp7XN3
q1luaT4FSX92sQXkT6xGs5fphn/ZdpiGW4SlisfLJw9JnCpmjbH2HXsjTyvytnK+ccIeET3wzt07
pDd1cygNr5H81eY93snH68jt0/tIpoWc11/eniPAuGiIgRVpPJCWXQc/2h2JwbQNosMjo2PiRvt2
yXagTXcnjra2OnF1EYBId+ZadMd2Kfw0Pm8bo4EGsFsqbIQKWmwKh686ZeXutH/7EWiCSLuFtGdC
3QRtvQiDSoevtF5fe+I3htuGsOd1MLUfU/JZvQJhUuCB6RImE3yRvKoU6yVQHkPuCiX99Y1Yrs1L
Hr3q5ZxdO/f19KwJRHrYFF/36ddlrSKDVUYfdgB8Wbl8rQMjeRHLQssnnUdEHahX6Sbz0gC4+wnD
YA7KYwMPuvkRXe9RDcfafzEkivvGGbbXEfdxuShs+wVCQ53rdKUhRcWVQxUkv0dJfPIh5ZYd0pKh
qNfcASIy3Xv3CX4iSLCRQyD94hYFSeRBZi8pyvMV9JEjdEdZjtf37rS493SmNAChngfqKF6AbIeN
9rcrfVkxoqCoID93pcmOmxuxz3gsoCBZnq+D/ErK2LiRcJwc5k3Sq943yBL5PJdCRDozqMlvo8H9
MuV4aq8yLc0jncQSYpI4DvtMq7J8rJ6ZKWOdejEBn+K5ECF0+peVy+zW9GQcp083F3agZhpSTiiB
2jAtClonoPbbbt9hAQHPcb8r23Uuv6bc6fPWkof3PBD8jdHMEY3yhjIIRtanalI08tbpDKHehURQ
gR+WOn5RkVnxDBFvkfyYBiu15Djc9qVug3ILRrCFvy5kfh8ODJJSpxbzci1A0mDtKKPL+75/cfpb
6c03quH0GdoHZCMFHMkypBQgFVyesnAYrpEKG5Ixa2RXeohXVLi0qZtcJr2uz9l6xlHzrJHqYqEy
q0S2WlUMKqK7sD2aVdJffEAPT01AaMIUuloGKupTRtIHYicMx1CYzxkTNJep6MJ9JtIaxq9Fo2o7
kf0x67fbTBO7saAnjhqHT6oUDQ4hMfoqzP8WlmLwW7Qgc7pRF9m6NQJF58XHBmOZVK7XJDpjRA7z
wdDBy1htGAjyJT7rppmfIFvXKQWU6wzvppVIqWLplI5SzJbLv2VNmWTW2jEmb472GyVCe6//tLn3
I40vv5E3nj9nmfFskPbwavctcumhPHtGUgJUo0Ks8R+4BvAune6+aD46fsFXPqPdUVrHkRwdIba+
0eDWRKJEogH0bUOgQQLZhzr2+hQFsygQEJyQQFJkCDkTBvSvIj+dUhcazPXp9w1PIrh1q6aaAGCb
PuSTEu2ENdo2cxdJSx0vF4Oha/oNIgKXNwpGItcoTV1w4XRAad6jjTRCsVJfMzrCyR0jsPTqh4xE
TLA9/xl8AGlTU8nfz1n4iIUFjvZP0lxS9TpB+TdckLG0IH8+dmEauHiyec1GqrF8Txy7NV6BAP6p
gCF7huaMTfHMIvrF4GUu9lW6jf17hGnCmMuw46Qk84Zjqpvz9mJasi5IrLyLCecKVApYGjaV3AWS
9C/e8eLfol9sd1+v5j22tyxZppsuUrCfziziRVou862rdF2URc5XkqB4DKySD/pbdKoHwO5FE25P
vyAcge1UxGWCxEcSq0BzipfXYriWGSW05nLykrCyxV5S7bNdVPY28bMkI2qg5A5tc8PfVwMUD2sG
/Taaw4Ap+WgcUHOW1YyV0pz/NuliG/4P3juoWzqYTEZqqN2DU37HXFq1eYn3wHHqShLaOEO41GWm
3vq32YVe8PLR0ar4uFqBkn/A57Pq88svxOOxfscglUdXvvRXNB1WJ60KGVBzdMK3eMLPkjJDUg59
c9dYDlvJVhZBElaD6d6md5jJ1pkc+2HIKwxtXY9LNqnqszVLETnYK9EbmdK4YEOb/lAVjdiKABos
2YnJGwfQv8OXUk+zZ05unOGc/vYIDFvlZOV78kAWrS+LFXA+JDjJQmyNConcLhzwFD3+tcXaQqcn
rXO8aVFR/ykeOmPMT8FjTpXmjJTGgR1MJ+nJP7fJxNeYsuG1myO0p25wczPBB8qQ55/H+KATT3Ck
n1VhOIx5oBFeYAmwluKAALwHXmemRlzhQRgEL9d7D81zouu3WNTohVswVBkbJpo0vmPyK8TTj4WX
0u0gqqbiLZNyM4ZGlvcrdhTmPN8wUCmOOvEeXAmfn+Z5xbBB12I8oTExK8oBqmmd6ZJkul8QRWfU
JwpdBjeiKOelzXpztrx8Vg8QfV+SChc9c2LKcnd0JHfTi50lq9XUHD1SmadnoEb2CSDdECUoI/Jt
9fym79bK0me5P0/8LZwpKwQIR6fSVL+Do4sITWTy5yzMEDiNJ6rIXw9FXbXfeOnSCwqZOZK8KYBs
zhVF7xcLc4sIQoBqkIaKR8WPah/RZcTXx/tNbjOCAQfGo8jmoaCnb1pXrZCl/tdd79VBiGLv+gSh
MpDG9+z8fETsiBwji8eIfgsmIIdAQwb4DBlzRfgpAqs9TLcvWi2jwnhG2ve63rvKZ8dCJ+nsRj7L
kaB9KmK2mS2WVXO5kobG5/c5ItObXavQU9/o9QcbDjdVpkfk1TjRs/wHGiVUrJM2DrNtbTqvZGNT
vcrnLJtNiZMpQ4vjqjmjI3dT4/ScIN2XDyeZm7bb7bEIGN+T5YYPfWpc+6xuFG4AphsfMCozVMPm
oz85lg2YwZRGlR+QQLHrskrukwaps7QpQ8wp7h5NRWTyhdQIweRT9Q/0gaa1JZGitRPTtdH1U0mV
WotNmRWKej96LdA8kOrBa77lR4E7rb/7OFDDws5k0//MqHFYprJR1UqfTz/vyX/tnjv1vpq34K57
7KKgq7w+8xR9Za+2fxMYV8VEp9350U5q4x1VxF/xVsuuGGBgWC41H7C7jRM2bjvtE60PbzfonRZ0
0pRV3g80p2JsLCw6E+tNrca2lj+J74i+4MjETpakww98KmUMwBU2GywYTSPDIG646Yy1vSqQ+Wec
yUKpaQSxUWbdrTK9tsoWzLB6b3u4PL5PZlZ4XtxlfeKDJu/CBRasQFlq0aFnrJx4aN/fH9meJdVO
5rqW9Yf5/tw7FzDbflCxxTz+RCdeVWZSTNgbV2pPfIwW7EBPPuweFsTq4ytk9e6YySXGnH+vSWjF
dzis26fTM2Y+CaCt4ObqC+rLS3KNIKZ/f+VDBkaNriU9D0OdUlOts5kZTRqQKb9U4s6PmFxxFarV
UV/uat83iqL2/S2iTYB+O+/1SZYqKINrfomy2xQqmjfwz5k/+V2xXS9cFFsSWf08NZOsLUahtPWB
JQ4FsOzAji+WS6Jn9K5yrQZJv4hAheFPwhZHU96NjbJ18jjD9FVCU6IwkfinxxfMDe0Kkyar2G2C
EIPAsEzSj/FO/Hz21vhtReSwmNJXDBQVuxvKV0D1SKYOZ0HrFDfzWcwxSUcQV3crCrXcJiJ7NtV6
ZT/R0cgGmj2TXceDBwUtQCrzwoq3duluonFJTWHZe5Mn0egVRPkkUj/SzubrrCzUMqWEh9/0ULAg
SlzD9Vqo23GZ1Ddmg2wbLTmBIz0o4a+xaodnw8t7ZfbUo3Yhdc7ODAxYw07tEDaWC2a8T258+HLs
j+i0VOfIi1ZUWqhTVV8PweBxsiTb5lrKDs+ax3Gi/tUkjdz6TTjP2VC1q10x4ddVkCpyC+WaaD7K
YJEkE0Q3Qm00IANEgv5UgD0BaYEQisKWNIaRQASYmYt4rVrZUvnRrf3e7GAwjVjVP6fSbsvF0HiS
ehDehum5FDVlzxHR7eUhp4d67VXkmuEJJkUovjEtvgkHegFjWdarHDRjQHy6FL93b8TotZZ0WfMB
+rv3w3sj4iYoO/LA4mt0HYgBAkdVDRr/ENfylC7xbNK6GtCxs136gGwA60KAdW6do6xbHooXOpBS
DMiOloYzbUhtVf3kl7UNe+XmgcqM0s4hJF5XLfBL+K+KkeKnxy5OQrTA4qmpb/98Ts/LePhBlS8N
tGG43weXxC2I2zcJdbPCuSXTbd18rcggts+6F0qFIKjatQIdbv411M4W6XBkEeQxiSwWGxgckJtR
cViZyZ8DaLyUGn6Rgm4jWZTWWfoBPhheOHFEkZkigCp4k758+CopYFcwM7U+tk2PK1ZaqD3VmeBp
DDXQOUMBqH23gjoD52+MrOzhazYDpVupEbwegYH+IVO+eemDClSae+fUlj6VPvNOD/ajOJQX2J8G
I9RgWTU6WeoIB/qHHJ9GETwgBW504rrgEmg13IGGj6jhVALmWF/KryaW2EL6lal5ie4RwPnch1Hh
GwEuRWJnfNmcODxPth+gCuIPuBJPfx6Rr9VRpZ+08Rz9nDR3mWdh/3O3QXfAVsolObLqHdiFePgM
VxHZSicajxV9oYXXWhu/QZPDNLGdytAVv690y9eWxs0lQzeLQXB0yA/w41tqXsKl4rYV/yZud6D2
xq9Us7BxH3ZvJd9QDeEobv7z6FRXWxEAjjfF7MvgXNennnkHTxDlMEr+FR0LCl3e75e3359EXWw8
ws9+OzF0h0GCkUe9JlhityQDUzzOHCRvovOdi+3jm7CcdLsfBSzsIU5BDILAHBJbi6sxODGT+g1b
SpvvDBT5JslWAzH+QwJ3AIMRl0WWA58kw+OcRuOCt/oRqUACuQv36etPZUuqQfSLBqG3nV2YWEXa
5fG5Bi8MSJpxRcgeACMDepntidGz5CE3icI0MJb6VLzbMnQ2QcwA+cHFvLBqrv572pvyawaciKED
GlSrOOc6dUlu46GgC1ImRZO2KQ6lAtb+DAJfiwetIu/FXnWstWdfmfkbv3KJAyQj0rJAMKS8touO
0hp9jj+jpycT7bohZUZ5dN3dd5qZondhcjZ6v2x6qiSHFLQuPx9pLFDx6D+HSeQLJDgItA/cYTA9
Uu51kq8SEls3A1+7gkM7Jihh962vEeri8hRiwWzidh7DZOxMgULoWNc4usD+i1+G2TPw1HIAX8su
x/zwZDq67JJTXnSGashrx9e1Fb2S0qxkvRjQzJqkb2axywoDSOfIWddJeYOoP/E+4biMZedQi2v4
QI98WzqCQfMv274iykzSyyABwC8tKLgrJuV08LpvlTcTzp2spWcYyWaaOJI0SnQztfTwkuBxwp6q
QvSwsDOuEQXDL2t+30RekCLbnYjiJ8SNEvjghRlFX2qROvWabafZ5+W5nCKRDx/BSMsZ7PDvqsQn
im48xT8FotVj9s35X4yao671oZtjRZyCSD1+F0Pt19j1fDkycGUyM9jXWPeIGHezVBoCv19DS3C0
itPl3tKR7Mqo5E1462YPGWPA/gdINTmPMRRUT0dAsz0+SZjiFERbgOUnB6sKeXk0JsVsA0/5aNcu
guSRqiCz7wafH+nB/x5a75lrtNRtaq9S2R4WUPH1Az5kPd9n10CKfB8aRW4uny6WXEFPjWC+VdIn
WksSAkte7MK9JpSaJPBJW7gOKH8zzBQrDWvA+mPHdVt94QnIMtl8kq8cBcN5siX8m7aqI2wV1f4C
/6863WAc3FhGYNDOWKH7ghVtnux7MVDURzQpCMlvvpsL2DSK5Jchb3OV+AO45MBphOwCIcg0QxZg
VZs1YY9zk6hh48JRQempkdIvNKs838lq0O/E00+AjqXGoGah3ISGfimI02Cqsm1IX36PaU3j2r1m
r0J+Wx9nw8Esg5fOEw5q1cjR+PiGz+IyHwGnRrdRC+ZxcXLzEH16ysmMbw5jwd28U66AG7Dwh2s7
QBCAUT/I/jHNe7n1aBfGxApGwdytb88maxwYV0C/x2n+PwWVJQQosMEEv4/bG4ClB7HdFiCNhikU
mJVJa2HTnmbITIJIzrd6fZmWJTEbEVERCWYo06G1kzBrKYegsmI40aY301XWBDpBYqVXlFr2iHJM
5FnYaL6uLJ9q6VsEotgC8S2+4Afc7MLintJsbRs3KzBRIubtdTZNaNzqwJlEatMAcj5FZscOg9I7
lHnfXgvwb+SfJsL6We6KERRo8ppqQ/dh9VSMcLyUGBbeJTXgS95AtkDpJapxlhxoIsRQBkl+Z3nQ
M4foQ7Q0bPQTPg/BbXHKAYif3zH4bI+X6jR8RBQ8D+8+LRkSUcnbmIemSfikos7aBfMdT3CqFhAI
QSDqkSPUDJK8n95mkkyN9OV878W7fVFc2lkFhf1El3Mxvtbbkgh5j20n2a5emPt6rCX2aLVD3LvN
3LZWVyta9ic7gYNRf3spU73FrvHQpqe+v5Qa6D9q/BhtM7/rmowhwTDiXgCX1IH2jVzS6PaQRvjG
7SllBDnJBdZE3aVRWrBVkik9iIVYaEyAVTlO8g/gLCPVEdPO75NnuNUy/03DWbOmcEXgc72ONkZ8
05rICRIqQLKokuB6ZUvUYXbiaiPZZFqMA0pycicY7fp+QIaZHpE6n8BUXBZjp0uxcWxIdeIEn9PT
jAnDpbb4ZcbdG6rSNox98EZSf8DoCzRZWpHC9n6hGSSBKwmTh9zh59A15X4c0g7p+e5IedWo/WZJ
IewayNMf6w71ANM1u1i92reJJV5grVLhh25c+4YFBEGmMgwctoi/Upg5hcdecPStm158rszxmTaL
A/WpiaBfzCnD27M7j71p8K6IVAucZvYOBQhsoQfBqQYRsnNMUOUboLQ0dD3xGLrhmDhztzy9X0XO
yOiFWqGC1DCyy10FtW1eTAdYcuwDNpNwwBV5vgiZta9zwxyIlbvWzKym5j01UkEQaNJv0Qahg08U
mF6TKcaf4slrQOwZEHYEG1zyYvTPlXJ1JDXBwS7lzbJZcsYY2VplVU7e/vMMPG5DHCs3xwvf0mBW
U7WXfi5vz6hNXJVjK4wNHJHnuyQL1RqP4z8kgVN75WaoTRIPmRDg7Z5xPARcZJI6q9i8UdA8E9FU
aL79HHX5UhS/UyPvdkShYhYEqyhgk4M6XXHvVxEom94ide9gZ/z1L9RKQS4qBc0JPx1FmfTssdlv
s0LXnaXbFYjsEFnlYB9EmI5A0o2/aNqiKLQwuTdv0ra+IOfZfHPMgnO92RUbs8g8MyxpIZ6wwVEo
1NuOLyNXvaG3uEiytgVil8sZJZg3oNiy0COb6A+GZtQiJlJER6HZhV8ZRbhKEiyJm7nihW76UWz0
C/oG51kAdZYIbRNeHl4gIRIL4xDo8kIHN4fQmeFzFNCPQ7wYi0l11h7MpxGUUS0XioysEM9vNELa
erY8J+O/lbzhGeBn0HHBdN6ci5MawFAxx8wo4l4RLjvROIJsTiDRj5APy+mGKYdMkInCvPayhUNd
kA9BYJCX1saNvsCuRgjJei/sSNvquBFzmqGPT31cXltdVISzduOpsJ3eko8tN4GbegsY92hpDVtM
ffyhSqnTrpZ7n62UEuNSwjS3A6rre7KCnM+gS7naGjDIZgm4YE3UENHdVBjADPFCvZSWSFg8f6VM
3ITw18oweE1/dZ8Ma2/SLtrkvderYCD3EYbCcTmPwJQ/gpHe9SRghivDMigAggbWm1y0BjT6qhs6
VXFBW3l6x9d1y8fr66QBku9TZJ65TQLJkZT7/wA8GGaEp3Tfxc37FdnOzqEY8tEULgi2EtJJjIRr
EWJ4Lr2uCzB+tWEH+KRO7pbpiUzlzW4cop5tCAQUC9zgKBzm0dFdrJN5aGtlF0LCIXIjWAElbYD+
ms6b3fdSTmpKjzpVfILVFEDLZjoaiOlhxbRoSea6d8siQFp4/Cqg1J7zXWxKI7WlM/x1AtvwsH8x
rdJfIs+Fk61XT/zK5n7DEMDWhQhWftkNAZnB0vMrwXDutOLSenxtV/a9rowELvDLka79iflD34/u
LRQ7M45FIGyigflFtQMhuI+PmL8x9EjltxxazqRyLfNrr2igFLWg9rBOkoLEUOqlN9Pv6olc+Oul
LVqgSTAKFnv66x/4kR6lvfdA9P7gW+eTFmUppjbII4dIHu2iXw41Q1fUhPUwftlqSFgy+0yF6Qne
JfU2KnSn0xTAUlB+aR+6J//+B2uH5qoQx127oA1ejQgMSD6Rpv292o0Zdrnf+1+KpC6vZ7iL4JGD
n8q2f99judi1ltGT2C0M4/e5mxgJXX2DhPU+wuQPtlboA297jxQNutIo1/1k0SFPodcbzCBpG+tn
sXXKuUBdqMdWJnM42cfVYoHROkXZUe8p7MaMhAk/e+KPdoOMiLu5fd4ANr1jcSDi50RK7rp0FvuH
+pU6FfT0Y2DmFCVdHGN4tALVK6i7t79Ej4cWHRlzO27ZouC5n3UqDgYhUsz8CIEP08xg0io4M/TX
g82p3O2dURGhGyCTI57K4XWK3pMXVKGC49NOVOPAveyUQzbjeK28ViQ4ZXz0SrYyxYUbEBpz7zH3
uAy0JqO934bl0HBp5ORJ5gIyh1/TEuexuDsX6eYbjeDvdwZFDxYcXKFopBuBRgMp7ZWeLxtAIMuW
7JTkJXMWQzCO/M6SLs32svoNSu/drBvqpGkrF9IQzXRVv/LLJtNMBFFlOzuyzuR3QK5RKjOEH6KU
J5IUeBPTtObAFjitVrBclAcC26FGpWzcElEYl/1LWJmvdP9ZilEAJN4+Nr2nBStpem61s5z5urnE
U4dPbldoBKsZaa4+/UXN0G/xPifbjIbx7Nc/tAM/f2NDGyrWIBoz+LZoCSnHLHkJEyPrhR+IKEOq
lpBstZHaHc5hdSHPZhut3UfwF8s0/zB5SIg+R1eBm4NCptSvRHIBA3O4dQfj5eG4oFUgosqRzgou
XjS7nx635BhEbFfrlwov728zYYpadtxB9b3pHjQzZzKExnkyE9wJTjU8b9v1PohxIr+wKW7QK2jv
8SUd1v5L8mJjgU6RxY677ODAFlJyC7n2yhRrl8VKHAyN7qjm3UfuCVRk84ebYGvjamMlGcaZp2/Y
MzDELpKjN91TuVXKFQDzJBe6LQ3tuyW35UjuKHlqAlLl6SQ+wv38WCEVuBhsgbSPvQ72Cza6PxO5
TFImTvDNasnB9Ey6Rnb4vULYxmv5EEYfOrL2P9b96Gjw99SoHqcscy2267FToYxeo1/6WKvPwF0b
+vrs4zyAY8D3tNBv6346HJX4tF1H27fNXdEI60jVpHev6D3YB/JZBCxJYhPvuLEdGS0HEftVIL25
d9qBVXbr+MCkX+dp48f/48X+xEAdZnwLVxHeYfdRt7TWb65v688fVgofpQaXPPxdcVfsRxyG3DzW
caEUbySRbCwGA9By+AIBR9NTP3xW0FTTy+n3CsyuaML5MPnoLhpBzIwBV0+DwJcaDuTPqMGAzVqy
gZOXI3TSy2HYqPFkLA4rR835IeN8QZ4kIzsXj8YSWfzGRRlvfQJGzcKAtEoklGdBfqt9Y/CHoLAJ
YwzkM9YVMDx7WqoDRY8+kBqVuKJokVdzWIG41eSjw0i1B8HVvRAeCtu+us1FljAWg66h4ud7yJLx
+rNhBpNHLo3kZXroNxCr1YAtxKElT7SsKohYRpaO7MgJ3oALyok4GVaT8qaKZvZGP5vEhZycX05x
wwppVeQwmQtDeXtQwyp9Urgqrh9173hr2fOVM7/03dmUadaXHRaCFB5kGkEYmkiqGMm2pjB53cqi
Q9myXtGOljMQoj20Mn8eh1Gi1DyxrjMaBtJN4f3SYamkDZPcF4G8MSXh8APxH4fZJA6asPB+j9Q0
ybmH5z+N+E9JLKEuyFktJeR8rYnsLyQI08ChmWSb/f3OxutzOLy0DcwHDxN7QA8URUgUodOSgz5d
uxSn7PSE/KwpBw+8XaSm1Jd4cyShPKqdaAv/riYzNtvusTryBYd64JHb0KcsaCZhu902hOwTZHuJ
rYEG+Rz+vL/5gOvhFSlksr9jLEbMx9lnsDf9ky1KNnloGc6nNKMiFMk3Zo+otZRq1m3QnI4heIPL
BcYxfJd2Ql8hA4tUAKaCGM/EpWzNbB49uA+IBjxgYTWZ2MUOjqi73H3+UVAl7L8p/aJ7C7WEwcY7
3qQQihn6cr+Zj47olo7uh6aDkw2aoq7HWFv6lOSxMU0RQm9S3do4ULTY8imzwyIYY44/521OPuWo
3BkuwP+k/eR7wU2kSj8BZPCsDoeZbuPtj+AtLvtLIpX0gtEF3/x7x4AznMsF59AJOK5jwkI0TPEv
ek9M8pEJCwQfytl61+j2Va4a0iA8MP0kdk1e969U/mKYQGLF58Mo880eDP4vc/xIsUZO6fAHDPjD
UBK+CRkd7AUKbkbpFUwrP7EPiApJQdaoN4wDquqLV6FYBoYZczaeDVwnEPyexFzA1zlHNHuMFWea
JvRbEuFIqZ/ygSeumjdZ/Ib4QXg6LprIskmHbZbsuPxYzM0vUBFcLQXfCwRKRF9WGwfEgVXbzkpM
z/qxNB7R4vIjkvYm9cUnYApZhc49lFhLLUJiLWqr5rslqerwi9mBEABLzt110XdIS+Pj2KSU38K3
sYlje7F+fH1+glUl6npfRcwse6OwzaW+jorMRhIObUEm81wwD48f/xgnxa323J0lg+8afBTEI9Tr
lwhenvYIBZ82LNLyZRRcKJU5As7lMMiAkyGueaXmdz1+t27E4iR+xTMlDIR072CA0pSNJKcntHdd
EwR3tIrPb1I7F+M1Colrhv/KnpoDsFDSVzE6s8r5pmZiWIBOn/qUOF5x6cipJICtoVXQhMCBsBxP
3w/TVg7XbKnT+tYnLEWh607XsXa2lMu4yBQ58CAa1hmJr4ipO0QCSQQJZCJhbfAtj2BnKjaisJhI
y3RLPZeOgLjqXlcEX7flnQXVV2fO2SQkLPvQSeOuP3x6xtEwo31qcruAikfLybcZSB9fY08nlWQM
/lIEI0dljRqh7lOWIuoQtjg7zv6rXJ9Pbms/mcKFBLss/BcnFFDhMjhfgvhNJVnT4GmoMRRuCJVi
K27DXiVpsbcyNX9wcvAgy2beRqCVyBl17B0Uy23qBbucWRMpGdZ7tATQdA5TqqUGMgWaX8yPLgi3
0tBjdxPm950i+YT+vQq9ZhxdUcYTYYRw2QK2VlAQb2Ipm2DqR9xXzfYVg02GxwUJl2oQy18K2VhE
CXo9pwoy1PAeQXR6+J5q8iGg6+NzcKwV3JDjjbrS7XUQcsRvXZ9ST2xj2MNlOEt7KkTMmm8Kfvdj
3wQLIHZ3aJwXSm16DssJ8vb7TXKzE9/vSnymRxZiya2gVvFZQa92izjaKzf0hHQKZqtFMOlIgPTg
tbSXNZXHcg1Wve+NKy4DphnrbtLg5wPV4L0JukmO0dw+Og0zXdxHUeI/oZdprCnnSuvP/3viQXgv
fh8W2DxBmyx3gRdNZ6HV/RkyyT4k9X7qcB5RS5v4Q0NwdPcTUQsoQVKBjdpYs3TkYVWWFDWzEMHO
4uXiqjjswV8A96phPFVI2m8ra09eLkA7yHDe71YI6kXT82FpdwpUD65BQJNzsc5gwSqDNbDLw/HB
kxM8upgL1ILHdwjjY4dwjOZNA6oZW3dn7F2NI8TNQclV9JTqoj5uU9li+o8nbiqI5k7yg0WPuVuh
tydrIqf3gZMdqq4a8um7X31Eh7wjcHU+AyWMq9nksixUkh34N9QbKqzsaWzD1B6/NbBNw6j9JJra
hnKY9HJ81VnIC+GqP8OYLMauev63/B8p7xGQ2ZQ7QRbUCZmUNUotB+yTXsuQDdHUD776iCoa3dEJ
45ijjLU5Bfoiu36oC4D8i7mCsiISA33C5CXYJQ8INDWcJuqOBIpsPPBPOIqRa5Tghn9fO8AqLg+T
qq5rQkIBMsvNlQHWsSb6doI5oCOJkchBNcIiY0CX9AdlrS6FcNRWj64dcNSWG+5eFI8lJRJyvQoh
Ti7XGCxdZpY0HrUdAfejQgkM8NxQ0vx8qR0MQqVup3pipOtTwE7RWTTPYqyo5gYGpa014vhaEpkb
l7vixb5mMdxPBAuglKvAk7ocTF7sEEy3S+FyBxkPAuh9WxK8bkqAQJfb6ZNvsz9245a6lx/O9dIb
TYUYzlEcusgaw3dagUEWjhg9ncZf7cIhajMMSgGd4iD526swnQpbXtYYEXRt39iEZ8VhxbNXmjFD
siLxSDgfPMJoUAsV6q9BU9KrN83siSlnFQLXMwMEyP8Nt8dfRy5MZz/3PR7oscWOub7CmxqLZukY
Ttd5x0xjpw7nMTtLgSfkASo9r/0sGeg3ISBVYFtYLdoT8ozzY1V29VdkzdDRWTsth3DLgh9FgWmE
SAZVA9+yYIvD8fUH1rEoDfDI2Zmv3IHz5VpyzxrubuUsvkEF2GTtmn7dtbO9YNQTQ9X0SdLa08uj
DFVMvnZkkkVJd01xtGV+DvGKfJBWK8G2UxXkaB+5TN6aCITDPB0VYit+2zFsPYUniRZ9iFT+C5/f
tnyHPUPZ3DObhjnSjjBH6YF+3k/6AR4kEAfvTFvhGqy4OgQdYRKQCP1VSFl36GTNLM65If2EbKWF
ZF5njVECQ2GTZrX8NJA5UPgxs9pAMx8huYzSliXf7Jbb1CN4gt44Ud4gXLbDNk9SauNvBIsSKsvH
xVEnp/5fGhPMAm/TDJZIbH8K+a3lg1zecCRzGT8Qjc36enh6XdqnLJZyuc3praPqtqL3yZGQuZmK
neH8t8ijlsLy8JTfNjgF59iFPZ+8MBoPwBwifol0vCbgxiLNTg3GYD3LFCuz9sizWMftAaqM5GsA
WU+2NnN81PAUlDpD/SAX2OC+MBHafnDWiDDGmier/2yev5iFtPRLwOFahSBtOpZ/uHE2n20rdSb8
SuYd4unm3UucXDpAsfkpBeMSXawaUdO0KfdRxREcPjWW+io3cnce80PkD177apGt4H4CdgsZWPJ/
B0WClUm4CdxamLIKTdmN4/PVwrzXcut7na4wAs8CQSIep18MlHUT7L3zcb1cQL6zDVj4rfvsLu/x
C9iWvXmBwAcAPc55cJDY4c4Rb1JJCy4TEpjqv57dUgl5yz/B9KNNddQf5VVzXRU6zaLI2VU0S0pq
B/7SigFqAfBhnCAEOHjQBzMB5cOKAt9bI1IMxton4adk60nBjiN18JiBsWguhoMi5COy38jw4x7e
zpFqXWXwTpZulMUWJ/v+r0319KXm5T0ZQ4G7qxlLTUGQvyHp5Of2s0iPZs+zlK6RsXnxqRFMp65E
fnQK5u7C63aB+Z9a4uzerFwt10rRNACnCbn30tFJp7M9kw8MDDWNFC2YN3NiIX5YaJCgOCXSUcqd
u5S6drEsA3QpnyzJrYGFFCm3TMeRuKlycLVfX/r6NjlQmXiF+wFwhOHNn0vdqhNSPcFqdk/q7Iit
Hun348abcUu4Bg/lLmh0uQXKc+SOdubXn91pnXNUiwVhhhVSod1RDfl04lHuR31MQWFMku56sPtO
seN0o3PUkbQa6X76yJn7+jxYhE6A7C83t2yTHjUYWwNG3Ar8MAMLtwba97BA42v2l8fGpwyns/F+
Eusg7SQJTR6hSmWDHB5OS/YzTbMA7aPnJ13crGAjbei6/loc1H5IPHpTv3JOr6aG7mAoCHWiFNmZ
fsRCyx/2gEevF5ZIHOaFdLR1Ie2Lj2EZsNeu9q93nfa3R7yvFlC9okDwaxUcjM08Zcf1QLve7a1D
4DiZpv1ORrdigxFGX4f9AOEzonbLP6HskG2j5ufAe6+2anuBEqm8Aw3vVyVhAwSolitf1TxvDuUb
tCMJ19dPph2sFvv4WfPr4A46Vm09HkIx+32OSZyNFtCqtSHHHfzqEbeEx2d1nEpjqVMjQ3Fk26bQ
aGkErXmXQiNiOf9g/qfVecAKwtFeJw+VmIUpt0EJmZy9WAlGsyb4JRVf91z0rHNSqHhBSuW2kZO+
DrtG0II3ntbKjjDI1Ru8TjAmJTQ+yyNmtG0EfzudxE4rAxifdpkInzO7m34BoiHrMZ8bKW5IKND3
z+MMnKajU7AwqODjRvVvsebLKiaTr1jEyqTQJJDBxel1DWNvXm9pnGpysdV5fNr3ExTtrGjRsfZy
egRaU4yAe89Uvwdyqvvs9GqdLe68ek02KqeMNqdj/T1WCsMIizvDe7plmk09vPFB5soUSet2N1WU
hqho0D5E/N9BI9G7edRYMMfTwlE0zPSkAHb7D0W065vQPMl1F40jWTp9JR82fFEELQvDcwA00L+1
fPzrieFBUt7fyFi1wef8G936AO5En6DdJu5TzEET6ayb28/yfqy+oYgTFCC985oRXISYTweSsvMp
rMXYh334pa034tsRoNrI5/eJOk7uMBD60wfke+OayUbOuiSrKQjtphBs6PbJ5UnIAZk4A99TI5An
HlYPI9f/cAgnnJdOy3hs4m02bu4sHwZ5YSRUysp3c7DgDp7ny+hvf+rf9MNNzfMG2/e54YvjSV7I
gO1jB1Ov+fqSEkWScDdILp/uJPct2IzLVXYoI1EZmz1mxv7dQR4ATOBHDQifLR66BPXr0wGV5GqK
+Z5EwMRct/XdGzc/nCTLc736Iyzq8WpIcX+YSpgSyXV5BhNJYCy35NyMQs5VJW6d5vbloPaqI94Z
284lQdoDdwv/+VLdn5m8lJGMncnSN7JWdNX+WaQOGMBclbrrR3kWPSOf6uw2vMeGejcUTcwKJydR
j+eh7HY5CAvYCNeJSi1q6lfC0ApgGaIVwZd4uDU0x3BJ5JcWMdQbYRWu6vXCj1zm0SxwIcTYzYSc
/dhwE64edHhHIujUBa4GArqUBpljAUwKe5XvU5vZg6/RweZmcekQ8M5kFV8hwcOarwTF32N33tic
zzw9lb5tgfsiIGewZJgcoSvY9GWIhNPD4dYOlpFte9NXRcvzmCrzDIbccQHNtgjsqMpee98NVm0X
6Rm5fN29k5c8FAPFEabwYOx7TrADlPnjmNmKJ+CdTvBagc0vxhZADKugBC1VHbXSVvHdd5Je2pN2
a7AeCscv9WnS7TrXWhu2W0JDuFBfL2pDhvjzq/tFahHJtWqJntx46XhhjKcVMboMoHuofCZaOda0
bqE4ts3oflAxqVbso/wiaTnLx8oBQZ49i0StX93iDZbFK9AUtG8PsYJ/m1/RWhjZ/1KGr90I3H/p
ulSwNVJQU3zTdKfzE3ddLEog97q/gTb5Vu+RXKfA5BgVloV5GdvCpqI59WMPZXlcpPn12EkgO4mb
beLtsE/aUmh13zUC7nBHitqLATMmiQ30UAZydfsibO0rFnPM4I1vOh37dTLkw4h/k3ME9nG9rMLG
bfO5dYkhT1/8sUApcXJXRnSFDA81n/6NSIjpbACvozUBcy7qvXzhLrwddU3NqPK9Ap9V7880Mm/e
Tqy4knIgj0Bcgo172PInn5uyavrcuK7w776L3FnYq2PKPrfsE5NPQUxeMZ4wYW+mSqaLlHOjfZyd
NEQWwtm4EKIgBuVxmGFeRA8aXz3NpPWRwgFWSR7yBhmCiiu/0QSThERFJ84rQqWn9b2JQl3fmqHt
Ejq2PYx9WYdDrXCpQqsCzaALckwKHM1FV9+H9w/sEPemMBh7RIglGvSOFArPT4zgqkKxsK+G7CPo
PYhzf0MTOQQZ5jZvrYnDzdCxnJ9eduROJvZqhrk231MZrymfULUuwkIByFa+brRL2bemyI+OEvOv
r64Aj/5VJe9lx6OgyVq4cKjTnqUJfN8KZ1SnTFqDjiDHrLpEtWrMoCZ0x00mkwa+/dkMQaD0Y2fz
2w72WzFC45gvN+0EfcIf154HsujPsDQIiQ0IsNVyiVdVd74+KIermHwsFUTTKB5LgOU7JOfOW1vm
OJULtYkvizIL1JbhqGeJk9BWyE3gurcKCovkKR8dWmNPz8N9Ow1c53wI6Tagg8Q0oA3o+S3raaHR
YnZF33TqkS9ChEatiRwarAFO0+BOfMFxYdPLcpMxE+wMl9Spxl/ARP47JOhRfY3KGGZRU0gwM3PB
QlV/5RnAcm+o1qBzCvq8PhsxoE8VEGtcIqvn3/rUJyD/MpnFgUJxuyvKGtDf4jBc5vjEqf+H3BXB
2o70H2nbR7lV7yPNzL4ngkY3zNunyL+3tkc1aCqE0n2c102PjsXVx8cimLFLan14n8d/lDGLnr76
4mNhIr2tEMmypMZY1kJgOxSvW4io5L2vfTpkxbx8hLLh+vvjvB7tHiY1qpYXOcLj9wP5YdtICtKn
KjMElKI86ZWYhqBYDP1hNmFpfyWRuyuW86t3TUygRTQlwztvJZdLXpk/u0/ZP6iTOSCRoR0UMlYM
xsjNUJyPFQZq7aFw5LmZrMhPrC3wjppFMQNGHpza6lqe+Jx9aDrFe8aQCFxyKx7RvUNq2wgScLmH
6aVRRCUb4XkMNhnBejEO9wB8TLCk0GD8RIyQafrkQG1oHWhQwX2Za3WB5k36KITIGFPdHgkGUTIY
ZzzkxKIx3x/AfsdpiwPrYVvD+7ElkQ2ymaipJCDytGzwHz+ycyHabVjj5e/tzxiV1VfYH3OGihKU
MKS6o3w4Npgf/8/mgJ8k7x5tFQBpif1lPyqhhUxst01W8OiomRphAetyaN/JVQ0jrnAkoUJ7R08l
KkdAYhiWCljvKYvOtdnb9XX5KnQMKoRimPndCDbO81vPwCGEnRW/a5TTiPsGH+sxApZz3/7odBUL
cgTsM4VgM5Kkje3n4ZJWcjakbqBWTvp0HUSsJ2wZMgTVIPgKLlBZDcFxsHEUrPqqZ6p2xSRCCR2x
LLAOTgRQZMEzBfYBAFcDGlR1u//Dc2rptAqC+NmNkIUsrRXDg2LM9RQenEK4CfiNyMmyUAumIHNH
9mUwPkAofFB5//oamMkOFsi1Y+vMWuE7XkAos+fBUOxdZgwxQSAvOzJhZ2w5CY1pFfZNPyl0UtsR
qeV+l/HwN05KGp+vikpWT7Ojpk9YlCY29NF+qC3HvdTBPnyVwNLEdrdGE74LHrN5vuytve2+vRH1
x2PIH4MFn0EI8hifxkE4QfYHJV7rF/ATLj1zbaZ8E0fDjom28wK4jjd62qGdEUtpVmObzGqa4Och
gr9J7JeBg//8kDx4DkfbG0cMcnnq+ERXZuVZWnerqQkwrOlta61psZHqZK0+1XbSZK4vv4VW8tUA
YBlW0JhaZPN9AScApBsdHwz0qETXbyzV4Uvi34GcYZDrp3edHSbFr7Y92yl6nAKzpNYnFsJyTXEf
3Y3ZhUIEofZDnXh/1cxlzQV2dG1d5jfv5RPQWGHO/6/jRRdX/iDWwTwwjLCVv1H/fZabM7GF6D7m
VUsxDuJeJ7R7La2gq3bWmRYe0v3Wmz8mUTqQO+pDETCmiJw+r97yO7iafNWCq0YGkN5/mHMKcrx9
JfiDLKL3nSo1AIsb6qpYgHTQMBzCayLb6i9+pL1hr8xTjiWOf9WwD4GZKr2rjWLiJEzSYO4FwwKG
v4NEOvJvSHhr8VXB8xbaSXMfBZy1mgl2Q2J3DYZJpxRUsTn1hndHUvW1arn44nkzoMO1E9pcgpTw
ViyziRmTdOTHiRiskdjlUiPsKnKkccO8tFeBmxi+J3eQcHXRn0YFUsDV5Z6c2s3GJwe7YIH93WYo
M616zRnk7ycleNLDKfLtJQ8ejwCrPZWG2ZaCn3REPYvcP9xzaYYwXNYATy3/ItrkWOpdm/rIIjv4
8dVFFOR4bsOYfQb+etzrSybXmjP7kaaSmolkoMTbagXn59GuDL/ZgC3NBgiENrn7PE4XR77ir7yl
1Gr6dev5CB/7Z94ED0Iv4UD84s9b52BMipH6xIPfcrVdD0ILFCQW197+36gSZCgeCh8zJPgfN5yv
864TuKazCr2Af2UEsPYPZhNfnC++tGlFzgewI20SUMpS7F0oAz57MW3czMFraolt8wfFFHtnMwRu
CtzVmNQU/I66tMKrWYvf6LM/3vkmBmvrxlNAjEgefhLDRjbVxmrINJFueHw9LXD+dtqssU9D/V0+
LPSsS2P6/7Ss48BIfkWa/g6VDj+LncBvefT9Nd533s0bGul7hqO3XQh+rQ66d1KTlCGvNQaIme35
gzUSJ1jUmrSBhhLs/X2fctxv7mFrmAmaQfC2nXO5HC6xtpvCeSkXNoXhqDPO9DAyNbkLCMB1sZSo
zzwkfiPH34saK3hLql5/Pb5NKqYUK/JUwdYtrEzK4alignm6NrayhEZAaCulblZJ0LmRHV2l8epV
T8rX8qPe3wIbaK+GYe6RiRAY05asXQ6zDrjPgY2Btn03OGPvKXyeBHiLj82Vg1fMphMshwRRdaHj
CF5VhPG9br8dY7WPHv8kr9ERNZMg4epgL30Tt/TDkaPrbf/O7LVD3K3spNWmL45a2mBiG1bJ1LBA
yW1XggOj2v2oMm/pOoJMS2o6UkFTASOdSWzFEEEWuw64D4iHN8wG8cTyxbIl2yKz98KgTgQR+7cx
2si4tGAEhcFa1seVvZH/4CQBPYJM7yYCzHzr5qKMidU8iEFmLOApiyfpWGcpa1aCr1KIjNJxp1Za
FrKnc5IOEpqtxMAkm8k0nDJ7iZf7vb9UcVmlddbbu8Bw4pIx5kuNhak000NYh8vHkyqJvmoONi4v
faYPBY0kd/qIQocD1MNoOdaoEhxXVPnQrsgjlMC5HSNjYGnw7oorJLc+eCaspBAKIlNoqgLpPth5
Q9AK9X9JYUfgmMx2upP4wVVq+oLIENeMM6DxqBPrZ16gfjTwdMO15sSYhSCVfD0YbndfVauXJYO/
is+JNAQtgdvp7Q8NwlofE0jVbg8zRp7TVrzeRP0I/QHFdwfo8gbWJEy+DPbDd2rH4DSnvAyhlbNz
+BVfd91M/R75IHHUS8afxf7pc1K6bj1qLlSMGRBlT2nE5q6KSpsDWTePT0X+ml2iRK40BwHc8+2y
W+Ujp2UsOxCWWexSAEQogLvj2GUldeeDqoVVHNoPYc6d48A1AsyA3+b2VwW30FFJBTn6/Gh/JQgz
YjYXsVcjFww4pnEchB6YtRYvnVk8hXrkraqmcF8A8gHA0Y7fZocZAZn0Lb16gpQtdU1giMfsLCIg
8zRqN9jXLKQym03RmKZujAJADjPbwqC92bPJAnYHiU2mn9GPt+RyJP9IJeOShmZcAKKuERrrsxkf
Yu1HAa5z3WDVS8HzXS6FGyr3jEchMyR7aTXaO43lwkA/BaBQ+jGtVWpiZPgHw1by85Ime0/9dssF
zu1CldqlNgWVRMgWXoxN3zFJ/FZbD1kejnbYEuyCDjvsOxLeVg5FGX/sKwFVylXZFfxwWENKPdsV
TvxOKBtUIM5fdRP1sCrBoyC86p9D2V7tMrLaXzfh5OJfgHoOmPSp9EkDAVOsGEeWUaLMZaWpLOWW
EjkNIsOH3rXP3p7wQAsBcyIGsuRZRSkbsqq4QlFRm3/6MVFUoSDmWiX80YUpB/sZUlLRaKrKvAUv
pAeUIYrkEEk26aPmDgDBH/A/wNK/nkXbHUzuI4RSs0zhl8V6VyaK1Mz5QupdmjaR4NddnZjBMyki
CqAVwFS1G3m/VvY3UpOqf9tBWvPNLa0Uyg1CpaNI3XbJOxxRjpDzZYe3Hdbq9TcWfsY+ZcjIewDZ
3RoHdHSgLuxTgYTnOAMfw7ubRUmzA6/UrAAMx8GJI1NYVj1kydC5wpJamaa2tImJmZ5A3nemKv/Q
OrndKAMT74ms9JJRjKVKAPsR9McZSuK94b9EdmsTRTCJSR8Y59CveAO6OvY8DMtkjIWyH7+w54Oo
nF0C+tnIbJk7KtXA0/LQNI58gvJRW5mZR496cNo441K0CgFRI2WE/Is0mVgL56vzqpcf3VtbpT84
Gc5geU5ZJ1O3OsBhRjDKxljXPnPJmIB1iSCb3SnCvKbjsBWRvZHl5l/qXTZ1vFIUh+tkJY6tC73t
0CrGQUBpCRI2dpT/8OPqqewRO2AqOY3WEPqaRHWQGG6aSKJ025mFaxmW7yZGXMLlF0CVEDUtYWv8
fHLPonhJ2FvuayrSpcxiGMskBUwEnM5wR2mPDTferSo2hcF2M+AQE6VodJLlzbzdU7DSwhOU2t1b
ocNfHW3rThmAV9tXgSk1jkD886x0O0H5iFdPlpPhxju+qgXp0hAEHC15wSp2/ug+xy1IIddSVGBq
F7eRIyz+VYnkjTO0zP42viQFj+i1/7fRggpeKz7OU+Sj0HpT90q7z7k54Bxj87SQZrAkCSSRkna3
3CYj9LmAtrIpODO0OMVCkndKa+uKX1QBIFW82eWCO3KCXiC4FaLC/hI6QolYuNscIIYbq/cE2VFo
cWInE0V9SNr5RBjCVvB3iYhD41J9oVuZwjxWBCuGjTz8VpR6puI6CmdmegRr3TTSdbmj8TJGHR8d
4ru6I38fErYjMHHqIApuZwj2Tdu4LIJ9BpPPFCOVeHGTZrMZ6Bx/MnG8/5NyEn8ocOSnnj5rxLSZ
8bGv2xDbyoXp4zB9f3FgyFbJPmUkyw24cDVdbnYKi2WnJYRRI1GqeP9rI3VeZHU/l/5jmEZ/N7rW
8Rgk9QbW9tk3RrphR12smYSj2Uhq8DLh/YBeKKQVBao+33UFx5FaYKnf5MNhdOYkoM5WOcty5fGs
wF02qDlQmlcY7d4kuq9dL/ltkcdV8GX60AgAFOOqAendj5eJSrqB8RwJdz9uGDKJ7rXhK79V2NOF
inLlT2M1iF9SqgIHBDQ+BUhkf5KRB3331HTz0ODRZm7rsUek4uFQqiMarlciAKbB5N32tP2Z6gMV
N6zIBjatJTJo0zLTPb6oWgZwmPtb7mv6itD4Gu33CZRlFo2QYClwsLCGOoIkavolWUTEGsKJrAMO
fR5Xagrg8YNDLXm1Dpr8CyrkYu9LiB+/E8blrvBGCvvjIA+NJr2hJmfQ8neTF72DpCRjFMxKZI+n
uKTbEZGRRhn7f0aOs1tBjbU0hHmQqM8YwpboOKZL1NAYJc4WwLDSLW2dlbWtmbfcx0v7qeeOdl03
5Y28z64P16hxC91+bfwLzN7P7g4JR9kSjnKjBjoIInxrHzqLoXcCYGFNyfH1O4ih4SIEt4Q1YZG2
aA27NS0zFyMWYm+8r/D5LqipAdszFiybZfiC7PKlVt6VW5AGLvilzzptBtFICkL1PZf8hyNHRpql
ivnWPZm+ncjMo/IT7wa22WG1a6CGEOqf4IWwdW+oKKJSRDVDAR4oQmEYV/n6SxPRg9lX5cJbfZCE
0UVBU35V8t0tGtkaNfURgeHl8PvTlnaWNhwrTnYRxqvS5uUpsf429jGkKaIMwExO4cJTCaY+/XjZ
xW+ikcAx3z1FpP1VMW4+ARSkECcU0G2Wl7MrtwLTtmSyXNVvLMo4HQbGyaGWkiO+Y1iC7AyuiB1V
ClhZhQSsfH0maSwVcC9MTHYzDGxw8DFBJzjN7IBIlY4a8wni6h+kj1jyRZQ41fIS3ApAoT5wyN/p
unCImcLMW89GA3EqfsgQZENniZ08hJx0cr1V7oB9sWfLKl1lmWB8cG9n/IWA9ioB6/4tvGEAYIHF
Xgx3bY2XWKXL4yWFjJquB6XiUv8F9jYYUZvOYLGTDG8YdgwfQ2E4BvhyS9Uqy3UIlJwN7c+AIYku
RLiE3QimNTb0H4FYYnuY3fOk+Re3c4kt1+YIJCCX0X8xviEGrFT/UFDVtdE6YE5fvSAj5692FEDA
VY15cnXi64e8XGy5jyFmcQHSklvOLoDqpP0xDXqSiLogNGri1shfGsq+LpSsNDVm7Eoms+6oJ+JW
aAqaSeDUIJgTps/oPjhjiHMJ1K98ltKSjxmbQ89rPuVFIso7N1+DTI37kV3YZ+eOhHIWUwlCFbTX
zwXidhwIJi3SbsNFT8w8aD7+oes/RS1/SuutYAN1Vfd75pCahY22WnegQp7MWT45JSTYEYjvmfZM
xFk18C6Vyhj9DwCp4dLX04qAqk+Wg3Df0WfCTEq+qxoz+KxQv+gcfnIDh3MFF8NQD2SoextIxKfS
T0wN8m9S5q3Etdnkz/aAMG6Rr8aZtm18nnKfzJEAy0o4v4mSqUJCVFO9XqgJbANnc1QWECDJAztr
hK/B2tFaao/ysTQjqK3CPBejatrfTXFP/zmwIT/LAFCGNwzGk3MwebwsmFRW7tGHyClbeJVUU0/A
S3oPLJ5/OM0zvKvhjwIdbtkL/AkaRQPpmFlSBpuD5BptWvtYYIGBbOEfzArAv6dGFEiqRRjgEMFt
4baZpm5dFjFLvb639pIGyzIfoipPE5z3y+t4QBjUF0awhRH6Qi985ovcDLj4dxGSA/V96hDrgFri
mhMNNzvjB7yIbU/lDCktEoGivQbAjrE/wlFgoV89vHsevsxOp+gSCyilQwUPpHXkqoEWNGS3WKC8
9/SE3jcBXjjID3JTKXCk+t80qAPrluIsl50AepFh5lFSwBznDozFjf09Xv4rmIC+2iipX2XXcITn
N2xY0xF1wn2XM8zqZoU1uC3HjSHh4tGJak755eE61w9G35zKesb25RIooU6M5BhdncCZU+b4H8a0
IgEp1oHj+OhHWbxJqLz/hOTUF5gr+T7/JguDwNaqJ1UrUjM1w4FQvcedQ8VNdI9RRwv20JqV7OUF
gj3fk5Qq77nhbxazmnwDFnMDd87SjGZtG3WFELqrml4LP7zzSYaTw8QxaEbluNtc0n8/ZqXDnTH3
X9WAx1Swc9pS/A6+1Gb+7z+sAwp03btCvf6ejfKc7r01p+DArerVrygwM17lz9Ap19zrL7YozB4E
LADKdd//0BQKvu6ODSFDjWLxu19zrOYkINA6U5Eq+sG2x1qlQ54tqlkUUmuREN+7qgPvilYwSSY6
YLAi9CEvU+a/T9J4bt2c89ZqhNDk+yVwV3nnv8oNAGUOF3cgMnjRGGjLR5CyQhosTCHJ4iSgiD7m
l+MUSJd/RormdiI2Y4b9Zmdv7rwC6YgcIjF9yHBC6S11dGthdX4REY+594rFYhDtpITg+/0icN3f
K2zmk0ARjEBnbl6HIZdljiVo/JwWu++7sJbJRKN24MvRiBza4eJo15NITVAjWR6b8Xfb3bV9sd88
ZWUV7wB0SDmt/t8z4J09x1a7iCC9oeCJ8XDgIymo7DhdKVs/Q/XjajCZoCADfAFy4oBaWtEV7jJ6
S4CvRwQVMTVPJn6WCU411WGvySyXjHsK50W9oO2kRLpP/8FeSfdftirYwV7MKX2GzgbKoi25B6TU
Kbep4pcxAJzwwe91strWG7jQZgOHTL0CICH4mdKojJrHqzqpTs7a1wGyPO6aKcNs5qDNIQpZSsrB
VoLx/HwpfPbMH7QFGPdyL5PvsUfEVtcmkiO8yJxW4F7B1/UWg3yh6Wqv2ps1INWc5r3PRlblG9Q7
CjiQXTxzKHPGuEPF28gH6XwipJZ3eQANCUFwNRe9gDE/Vm077xVUreXovPJ29XHJNG8lvTZPlQ+o
oV5vtDO+mhzsU5QqxsWeIrspuCmFWUQ4KzgmnTcmwc1b6zVwEOMI1mGR/JAB5aX4DidjCwxewCPg
ugjmlu8+3euIaYMkf748nglRiBqR9LDaAdu/AIylkt4A0VJMuquc4fIGqA0umAyyZnxUFPfKTp0d
BRyeSM7ZhTot9lSP7L7a+Hp1wbhNMSPUd/bVCvElfinejy1WloOc1QY13tSEYJItN4rUUJOl8djV
IHU31uC8ssgo9kymZ14BUoR9PupCtTROlmaNT2oTakxQQ26stRwI4Tb7ZllrUtU3pY/BRsif/Xaz
rVqNMXMEbu68U67yZNVU8kjmNAPPYscCmIITLo9H2C2VQNQ1mjq1KzI3dhCShkRXWLJW0Let/6v1
zQQn7vvRRbiEa2RNBSBRsvahEnyrEARl6Y804RD0KjgLZ0e2pjycUJw695Ub2+E4CUhamuoGWZsq
POrpE3/00bK90ztpiT2XVDIq4sP1TQwQoUEULA7ly55RRzdAAtL9qLc4VQBcIjMjGwxduW14oscL
DNQTpnsseQNo3mdtvqvGydXIsSUvgLdeVSfKa7zmTCnosKgyH63Ix3xRh/K0EJCUGEyvtASgqe3W
Y5SkVRdrF5wei/c/xGyRzJedZwZG10MNOq5l+hlyVqgcMA0NjxpxeEM5NDGD1lqi2RUS0+Gkt0M0
l47YFK0VQu35XscnFYiLY44HBV/x7lJ+E2Wrzh2B8QZxUcKNCqie1B3sztIAhHl6uElneyJDko9D
tyK77SqjXi2nKE46gzSkc68cOQ1tOkFMtbpGndAZXEufBtcA5LL4sJS7nFroxVjSfoaEZn5WLeGu
0GuKYgzzvuzEVYyLu6Dv/y3qSlycLu1dNV+vOgGb0fU5wqQIp7l4anIXKcZjVNLrqjejnk5BQsDu
hQoF3fP0r9UbDF2ifJUsrWuXN8vLx+eYK+RUpz/GHVpbLoN/URswkA7XTyiQ9/f5r+SPEnfgDp4s
lOU2AScYelMYXX9VXPztV357e0LZm46YZkB4tZdhUu4V/QqC8aZPyRPyK3RdhGl/jv9O55qSFESc
jdWDTY1yEweWTKvw4ysxLZ4F3NVpXS3Wi3C47VB3vSK87kngz8yvaWjV0VMANXkCg7R0g7XmzP7c
macmnrUktNPeR9Q2/4rQ5/iYLOGOW31WwS3eaW0hcCDJH0crFq2ljUR3jZiQIjqqqzuoLO6YwMYK
VSx5m4uQN04aA6u1I5jYTZwUs4QDIlEXM5zkeRvRsOKqCg60NKn3cTQLZqN2+ExlV3o+V57/xfN3
oz5MlicRTiRwXXSGwSpeRHjH8kVo+YykNC0UHMHVnoM7wjNo03yaK84PArr0+F19PBOy3RO7QdOo
pcy7ImIKV1RnAsKZSZIX1S9X/r3BzZZhyBSilklu8yqr5nyJQuvR7Z50ktXA0SmWXsMK7Q3/Uw/v
i6ZCp6aXxtL5DbVhL/+iwWc3EJSp7vj6wFfGtC26rNCeM9IJuq7in/XhrARB4Y7Q058Lz0Q18dWz
zaDkOGCLx6pgGk5hkZSxAYPdHXnObn2XIMh/aU7Q5WYQFLG36Yb3EbLk8AwMclTHwzi/2CelnhQC
fztJAAuZvufBGrF6ShCmo19T4aD+c1sS3h5zahTm2yXGILzc+OfqrOC8G2FYsZyWb9/8PIIRuDZG
RJTcJ42fZxSnVCsodVe83ikPmxzj95vyyPurTr+Uvty7SKdFVV4R1Bc8ACv1baYdGdquAyiYOeXA
ZkPPDCAbe7pknDaANtXny7ONJIrkxLd36HxC2yE4uPC8JV+Bf915tFvNXeGhY+CreTRaBSZJj3WS
S2yWmTOKsRfueq8JaGJ5igAPEnCWaKS8oZ3ha2GK49CYK0W7OV+fZ2RYJJIPpvjQA6cJMPzp2M7n
gFVjC+JA2ISx4C6Wfk0iPvoqHiE3j+6ip0ffA5S/qZoP1US/2FSJf41S+6qukuQp9GfqqVVwzOoW
imce5nl8o0JK5NAvdfInX/3iuLUX4BFYUiI5MLXmSfZyiugJEIXQkg/E9aRRmUTAVlv4FQSLYqDr
oJOayWkmSwO07ztrHIX+LPzQJ9fGAQwgiPc13bAh/xi+Wih7F1lcD6sdbDPplG7nuAK4z6k3uBG+
8j8sVIOm92eIys3sQjNAU8rknkm/BxgnCu1frOkzNvd3Jt2PTzQ02rroPb0Cv+/9rWlG7RFjpX9D
gbIyPDTmDDQSBm5c6mW4Q3iSsI9SYhS3WjsUSWpKtojXsuv4l/hLtvAtBzpdGECaAQCUJFttVMiw
ozi2ycmaq3tKy6AND0db5m5861ldAzJBt06k1A863W3GmSmuX0vWh2wiDOj64VcWS69ggAnTrX4a
PDMc+Y7fsZp4w3DTAhF0ea+gXKWOW/w7dE3pxXgCmVgSp7pGrKlXi75AtmYT2k2sayhDw9HOK/G2
My36JS+tTFDbjnXShWUBpGCMLS0HbD1eeqraSbviJpUNVNLdfKivJN2fTVYchEVsGwzydQ7ObxyJ
Y5ejMPP/xVyvC85hi1zOpQbdGHKl8WJS9opTV4g+rXtzi+e5vIGAINRt2/kE3dOadR2ClUnCK22B
SXGShvO7OzMne4AyzClLCT27ICsQqZyyzZ9mNhCkBGIa4YYPHxIR2GdLrr+CJ2JTEl6N7H7mqWBW
x9jRb8kmH3ZF48lqMiMusFD9gggz8Hl3HHjEJzE24CwNCeP3Bx8U85J/BDihaHcGtawzEiqK+xRa
2Q4gsfrS4X/WMkJO7je5u84CHR66D3dgSJ4TTlMggVZjSJi8oSZ6vKCq9NAHDV42QeUyYNLTkwVv
i+VASWAtQlQkvEXCYH2aex4c4mtQrnYtuGJTSf8AQir1c07D3vko/u//2dEAw4DN2xCX1kwkP3SH
xdt8fiY0IzCCnLZkedh/0p7SVnFe6Q4DWpD1RKsnZcGe80pUrARk5Urh6uOYEabTozJDYj1MASET
eopszL2iYVQ7Na/PDOWSs5kPJtYzBLaClw283KZx07c8rkX1tpgwmfuaLxAryTELDsH52Uf+PLrd
paL9BPquIveUAAgGAgRLG2lh4+kijxv8fuvM9tIuBC2tW9GReM268TnPsNHykoG8pux3/pRyNrM8
kFSz6F1F5gULIzpOosZ1C+7ZqSEh0qST5so36pPQmk+VlFJ7F8nsrOGilkHaQfpjPCDz4FThbPMm
7Fyr0j8uCrmoeYqCdnJaGQ/pyLIwTtnZPbmrtUxTuXSptF1tDo7AAu9d64G2wZ0gUX/Ms5ANPPBm
tAPPeMkV2Fvp+nqLySzeZxnRQkGJtMEsS/NQTl4hnC4LnzsQOX6L/9POeWsJVSiUtI2LKH9Oza1b
iiTWJ06QooCOOGAokfz+xZhTO+Rc0aqHMktltCSSOdh9ku705gUvnQiWri8SFDvfqqgXA7SFSi93
TUnokJylCziSrEjy65x9uzI2NTW3wPT/S3fN2e/Gw4Azisl4WHLoPPJ6bB8tlii3MoluWPGQdI6K
TlanrRqzh8J2urQKw9FVkp+IG/xFBLMpIsu1YBHzQ1AKlMABOvK8MnzqdTQVskaBm4Z/iW5xCNJY
peMIqz+FyDzziHatw06Gt91aZgzLX3d0gnJ7MxsaF2qg7ukT8MX0x0o6nPsCbr4caxheNpNncpnm
enREm6l7hcB78XErl365u9j7udXNay/Q4ae0UGZxY9ZYKBgzfVpVpODXpujo5JHWE4UWiPLOZMZk
RoQaTIpVl35j2PNyPOS6FTez/IRIHOwm/BzEjRmLWRrY+oe+KVj0X/uioi3Q0POrKwcVJT9lmpKT
Ptu/jDd0eIh/Y2tllRcXmwLV8Ov2lGIjwoDnu5xlMvenC6CDXaQ70vC82fBG7liCENFPaxsG54GA
d/ZqNoOJKvaszbqz4/o18a2Iw9Y2D8adQSTd3D0MFLFu/rb56NsTSvFetxRgXfL23sK0DuTCz9LD
j9ziGd7fFbfuujzj+bOPG+qR39NzcanEX7CwnZCwkAHXoV3n8sfnn1cm2HLRI2kS/JPTGPqvDXQU
K/yAgHS5CTijLZL/Ob1CpvXZ63Q4uXviNkIodZ57w+a4Dy7XsDora0l3RXJgDrantRl3lwr1v5X/
GqXKpbYsRyJdGCZMuqU4FBoXCQ+eNPewV9BayIJ6YwBG68O0trvXK5tULbF/6yvPdskNQhPslhHi
akCNX+xr+s04bv82w24IVoJYV17IbYf86djzc4MofnXqSHPm+kihMMB9iZBWU7VtXhQ47lgWl6EC
WREOfRTO/6U7ejPmSgb/qIcpHhFUjDZUCxBPf4qwoA1nMruBKV2mEnFbAEE2vAAhLmV/oS7/25PD
i8qaNjXgjEKFANSsiEyHF2FgWmohgTocgl28J6TciOte3Jf13kgIXyDJiMdlqN1LPmJe8zD5IJbS
AxmTvHBkJ4LPAW+EvYbZ7mpBKWGHsY9lvnzVv4D33jvX3G8C76GZFA5ugrvPHboHSOOVNuEhPVr8
IrRsQrrnU736JHyAxX0aPIQiJf8uUy9owRQA2UEcBQloXRhsU87U5ThWyxlWSKEiFVau8bXLYS/0
B9+P3k9wDFipQ7tgkDOq6wCtShIicrQ8bMhguTU+rEGpFtEsmrTrqE5IGD5RAwoFTtjOP7Y9PZuq
L4bC4g7uSfZPwyFd8o+MYnJnG9QoVjFhvl0tVrKx+0lbPr73LjXQkNi8QmsUZwGowROieH/TAweI
D7qxLdVyJfOPZFydG9qQkp5I4tyVHM1ylNcOBFTGIwVdlRB17Z91ZWwI0IWaWMOOWtyZTkU+M1I4
PtjbHXOq4rAYQK+aBjNnEu/MwMHvulZ9bDnONQnylDtNxPL4W0w4voP1Fw2ZKZqbkEXAZq0dfQt7
U2BEoEH9BaMrlfnBnAZgwNAHFIP+2QjOS7/OrI3BNa69n3yLKQX4KqZsBMY0mrQDQla2w0n1FXoM
ivpYKCk0IY684yBW7z1F7fTWXJTQd3NkEC4g8JrXAvNSLs1a2F8PDKnHmnelticS49yF7KzBvJfA
lTc9rl8LoVLSaRLtij//TGNW6h9QgtK1Ou0JlhwCONl/875Hx0JEReTZUghv+TVboHNV9ucYcIdf
1kF6Jnu0v0rVYCb3E2jIYrRhbR865+HTu5BwGijVlmeJstZ0wuSRqQa00A3X0ES6CimRgEQUA0Be
eadBrT9pSYyl2gAfTlt5AY3M6uIMWoB8yDS3sMeMjkKmyN8PQTIx86YjHrlJT07Qq+NrDQM10akU
U5FgzOG1r41rlDcf18ZpmPjxxYpkXeoNnebnCWN7k4i24EDbyAFrO/paINdGEJ8M7I9z1LeL9Ty8
Ua3aTqYzBJN2s3lPWAT+Dd3ooucQhVdLdJ/phjUtF8WP1bhfkOYcHpvR+NC3UDl+fmXI0BycNT7i
zF4PneBDx5P8OMBAhkuJsm4CSF67oIuZ+SDcnr3TReCXSrLJFfXASiYJBRNh2p7VXzOpUiBRIdOJ
HDvrQS2QqGM0Z/19WivrYF3N27dwTRE5AuuixBz9eccubZJp8DGxGnvx0fYVxiWchj3qfIK035at
FhgSkuwZPETH3PNlBhHD9uJRsQ53ZglGnOj2Ig1FWoohAcj92TowaPQ9c5oarfhvXWdkxLHoXo7Y
rbIPYir5m/cJl29poDfPQxrgYm23SOMTu4X802VIuT411L5S4BLSYTUQUaHf8agohMxFfAqTsNk7
AO/ywssy7SLDviMR0jY78eRahjyblTSqpXtxh9Dj24yNSdfWq+F+oE2KcE11onpQKXqLoxuLODa7
8mfyTwlrfiYqnjUSRblt8MQOMqRjMi4n1BFCad1vsqUmd/XFhWofTxrRT8n7THkN36JlasC/WSoO
vSrfozcZizCdfm08EBUHy8cD1BmrpbGbwYiLT8S+QFpMs99v8vtsI2MXhGv/jOSZ+r8p/HLqsLu5
MvfM642aY2Ay7DfCB7i2GSM31BYHXdAUb3Uo/jSifTQ58bsN//0iAeLSrSYWOX7wA/9v/oKZRmtG
nhIyR4cUZ/l6NbbCI3AOKqtnhMJuyJf5zXtgPcdg1jxjDYarA/2jIis98KpDgXKohJdViPq1/GQY
2L4Lw6MDV38Nsxtxst6z1Icesa0XL/dygfqhUgccusgARSiYIXMXyvFLh/busyd62ZZZ+ruXg8Cn
pxvXkAtFyxxYmcV/At3MsMHOKwEMcU7tOOqV1Kd428hJPw1Fr1wij9YOILtB65tm5pcO4OuWOJ+X
iItPtqrnzmDFr3j47PwjAfUyR+XfLhShDpyjC+pFlf4fVwJ9Puvc53TfcRYL7ItX7W8B9a74fbkO
7qhgFy1Ye389zRGxBylPMiCDGJiVW78XpPrdNMo+rDrDst/DdtR5/mVvZa1X/a9zsBHx5JeQRSml
mmsgTeo3h9b4PC2EIQraLv9kuhbgFrzst1DkTl94HvUJLjE4B5g8vPjkgaTV7iBBh+7eI7u+0pAr
HQ8rOwvN23WugHPUVho8LIcbfSWFSlp7AlAbg8Qy7XR0YzPXs8wj4r+xnC1bkPzXddw5UqHcN3/T
e2qiixdPSxL0M6HF7xDDOJmCKY/nUEL81DTa1Q0T1t8iSI1mdAmbca6Y/KW/WU1hv5AcMkYZtg6+
n11ECWTBykyLb63PVqF73mTMARhw/EjL25pge8HSv9Hv4sF026ffwZfGXCl5Cm3hovltnK7rXpGM
Eh0tgd877QTyerJt2qrZaDd7GuHcdGAhxqbX/dPDjTPCLtELlo98ltuyH0dlCCFY/SCYwZUtfxbw
CCYZsZzJKmfwJEEM7r1+hLh00vFWmPkCZlWsi4nbGjgBptF5igSchhSFRde8M/ZfjtbD2sKoCr4M
KUEa4KjmdvFf3WmtK+GeNb5k1h0c/CoDMEUWu4s7iOYNLkTZNtS68ul5TKYJFKS39C0EEktMhn48
srDPSgzC9xSQU9vll8G0wq/XVC1rSCFv9i8fON0oMKIeWp/eyRBtZyFg5cQ3PxrKC4GKYNDAjMb1
sgvmtr/owy3Z16vlvtvi0LwmXNdSic5q2cHs9AJFsYk8891Sp2uEZSEBEFby7ysl2alH8RVTMimu
h0/jKWeKQY2Xcd9RKt0JaHziQbwBeTtsgGX4xI7q2cONsl28ZPIFPMw93CHgugswZVu+WfsHX+2d
4MgdPLMd/PIFR1lrTqHMH9DbfWzWEdUEFmxKIagz975baHXYDLXjeMTCTwvzqaSQcPy1wHdoonqz
itBOcfZuU/YCcY+gG4nh9zfLSNDWOd5zMidsNDwraBjhjbNyJwTZaGKR6X1cYTNFXjLbp79Dh3Mx
y0NF0RvbO6nIG9dndj1dWTYQLpkpSruBWFOPhZlXi3S155nexmtbhxN1q+jIZXTPRDUZ+cWRYgGu
sxj4M+MGp44bZHmxB9je2zaln+psaseMXRzbXhWFc+99gPaSE4znkvZZkW1TJhUBze3l/6ZdMKGU
0kL0teD9Rz9Hfqx4M8HdjPDAoWxiv538HQpwDA6KkW1IsZxJLyrQEE6BEm+74jBgBrZh6JzfVNDh
NqWwnryOLaPPPj3Z+QsbXnfPFZuCwJOMTzgpPDGV4z6G4Fi3fapcrMtgH9u1SySsYTPoQuHwP2/y
PDR5IvskHqROnZ2FKSc5WvX6oaTH5zZs0Ida6p0dZ32ia/wWnOQXbcxBm4eWPPgnawHoJZnbpuSO
DyiQxDYNb9B+R3uG0O89K8SaUKdGXwDyTjLFWhbL9Gd7pYNUJnwS+LCggXLxENWEdnXZmCZ69FTe
nRrOQs1u9b9oxbRHQsijhIQAKzRKF3+vzLrWif/nhRw0IL49tR1bvU+tYABP2q+bxPfwqAUaTWnv
0bqW1V/bBXALBZs319CWx4Ss8Vf6TGESdsD5oYUmmt62GM/z/dwjzO+L/g7rIgx0ZdAiC9NUE94Y
VkUJ4aVRxXdQ1M6baUCaNzYpZHKDpWjqRgKHPijlY++Nz6l2gsnswUt1pplXWHDVHrmn22sGiimD
78DgOA1Vz8oYAoRIwrUZrec/g+zF85RyYCfeLysjsyXR1NiChR4pl2V/Rou6OLlzz29KjZ51kU8L
H3uzGSoJPEy2OMDkbBIAJZBR7myEURhXzyT+Gkz8m5EfedadZXpCgNm0GCF/UfCwzvNQNnPg7v2X
yUFGXVGRXyP1/ws3wlv86ziMKB24TVF7vxy+zEsledHynNHPm3tuQLMbssMuA/2TgCnmIoWht1vS
Ghi8fXc1jcBKtarP1I3HBjYA1ZF1WO8XTZipE5DWFNU8IQvhvTI8+Bhl+FZxP/y7XYFzsSBMRRPZ
D7vlDajQVBKg6xhzgvHJ3cu2w97AK4hkLZR40rFLFixqxTANCBRN0lF6gH3mlCxHWxUwyY8axCfI
3yGPjwDGsc+mdR37E5pedmAiErIiEOyyO9xsgpQ/Bko7tDyDBrjdNU8FqkNr2UuSqU+jrh6hppL1
FxKb85FF6JM0DZrrmco8FhJ6zvMdAL/1zzk4ym7Ly5pKehbHXgpMYwnJBBjsRGjawD0UvHOO3Dzp
favL3RKrsG3bCEU6Kkdb1w8o6J444Lc/4PciYJQAdgry2sv9V8zea5amvo/U+3QFcJtqAxp3+6d8
lG55FsuRpDSIFjYpyKVQLuazkHT5LRCqMLSA+o3r1ltyA9+ie3Jg6yhYO5LQa8H1fG19wE68MD+6
hY4RUOCQ6+IbzRYQFzhjcloa2lRuXKVZIs6CvbqJLXSdDfXfVvOypiIW8+A2kxPuzJjK3Euc3Pqj
/wwba7W93iOPJJPSOmsQiTeqsCGEuu2nLFLM150oVQWr+QrMO8ahNPO5Vstq8NIdEIiEP4rudqEr
fDhXgngTtGLvxhWfJhFJwLivKHUbNpENjAPCE5kBhdrAbfk1ey7MlOGVZwgPAt9xEIZaBYV8o9O7
KMYACTzWFsO8EL7Bv0T+lE1azCEJjLq9Omncjx0UVfHaQ0CM4kgsBZkJjBl3woAt7/iM2D9dURuu
aQvLm0ta2BItfvOE5W51phijmrGy0syGpwOFzyaQhwo4xpfm0oSCOQvy1mi2hRZJ0m2RkzJ6rkYF
0UbgMpb0SWWqmfqXYzkDpJQxbIakLiZ7p7CF8LXTKC9NtratkXOy0LG8Q5rrSZ7FuEKLL8+wcDEg
Ja9/BZ2eeLUNX5/AjGemPtJHBWE7CVjz8aLRMbb961/u5yVGARwJc5vx8PGhnLLm+207bDGbAz7M
Fm5MgU9FcvkgUoOhG01h3SNahBKY78wg6nFZWxrIue+tAn3WWX2hRXfivUZbCLebLfPiv90BsA/3
q5Tby3I4RUoIeapJAvjurz4tLIsT2HFSy9v66lzzVhWU1fDXS9F1BMJu2LpCHpYlYt722McjxVBs
LwTe4FxiqpZc6mMBocyzFKF7Ek0NnUx6Lqkl9hEkGvBc+0CtrYiCrlmBYTPySOX/t6deBd5uuiQX
2OaKfCLL2xy1Wuy9CkuVP7eElC1sVsv58oOs3xZn/DikHh/rcH6RUfQkg2IpEZEeqPuSNqrjYFLB
g1MiqKoOjvUcLb25NgLPwiE3C3MpV7BTDg4g1tuhhtUyoOOYwNMnH5M0/6clwmtwn1NqMkmz+Erv
sudOI65IXnXtuFWdjXAhZbTHlxg3fSk0SDYQLQK7iKYmyMkVLCfUwClP0qsRnUHqGbwk/8Og/cEX
Kc/nV/qa8SK563pDvkXxbC9Pb05SwYe3POAXGu8CI/Ycbqr7zahoYZ4A9GAOE5q81DT1X2O1uhWD
jQFn1QepZLbdeL3IdCXhgmckkz9dgJ4JiKlY3OHb+MKyKF8Ep24scZbzXsito9ZLrWxWHNjkyVIY
KlTb9y5pvtUY2gsDd0bu+0Alm093W/h1j6yrhp/H4nn8kJS0e93/iPLJEtmtLm2Dd1sKGT2N9qGS
BL1bzeN5AWhVoI5dXjgZlyfpfUmii1H4F9aDJTOPLakl4xB6aIk0Lf/GDmR2lEj7xI6AJfMVPYUi
XyNpFCSETVqiYmzSMd3LzaznJ9WTRLpekKKdoblcX2hSEljouqaydw/ukJNghLxL6chBJU12V1oA
ZiesIo50KzIfPavjsKaw71ACsgoeKp1MVV+tXaGVEnk0aWYR7HhihHPg8l0t6U6tRbinUn0yNl0e
nW5G6N+fblrBmDXBsHhMDFbbJ79oA0XY4V+yadSQraapn5etkkrP19fXtbhyWw51a2kZS3swkSko
7t+CdMjefyc0PPspH9f9jCmLvOo+9/BdRNA+RIeWOuDwcKhYh5EnGay8IcYehWNcZpCMO8UM2F6S
uOG9WXhC3KR+6VLSRLZikm/o01xtrXgCF6XeTKBBV0xjuw/lv9KZSo9+DYYiC0BQznECEQ2aKPnj
IY3sshgDA4KIzHefHt/7Ayhd/+QXODHoXC18ZHCUbqesXpGYJpBRZ2jH/W+EUVMMoBsaKnzpelKL
sKYaefDcdYGDBG/AACR5i96jx1c11fYRPOsLu6beP788SFDhaiVXLTc9p3vm8k8IVG+eaYzPpuap
C0KdDCAO02RJHaOgH71qbVMEDKWlNopgTYBcQKfB80zu4x7PZRNUU9fwc6HazcBdZNITpOYVuvsc
1nDjYWZeFQmaxrMc73CIeBdH0KEGVPNm+XXY3sXKyEUewM1M1xY9XwxXGnp/OAjQxyYWian/xbiU
D4EKP3dgU0xterkjd0smHnIqSqe854AyYTfNshpoLKeiHWAoqRUnylhl9zdasMQRyjXKosWnckWp
lCtOtZiR7U2pKsdgLeQk5/SQY66JWWeINRFEBjEfMhK92G7c89zMi51U1Vvl5R69XwDS8QG4JY+6
tj2xS4BrzGzGvItrbTwCAq6HoHv5gPD81U5tXfQdwlydZnwmazQfmTbmoImzLn2P5vSdvQ9q39Tj
7hl7/I/uSKn5rSTzsmqo3iVqi0OQHbgBaSc5uWJmTpx6sCbI1w713WPrHGzcwmg4PDLMzAhRVjF6
UjEqcjtLDplz3aw1HoZMUso2S3HLF1eOajXPgY9Gea8v7B+K3IM9PD3YkwDNMdsbH1aCpXh637fY
1tKdaYXWgkMJA14tBiQo/0lbCL38bEAOELQRBR2+yKAbCJ3golHdOfjcYjKc01BvBFRJeBjiTzec
7neXoys93NJ3eqZFX4fR/C2nv+DqasX2c+4jHZqPUmSErqo3JwMCo9ZefTYVw0hAqXiBM1GD7Blo
zffStE1MIxXwvJV9Bf+iBjxUiDa4MSyad0i5LJD5+wVHAQ2U+RKkEPJWaaaS39L2K/M2ePhAKTdL
qs1A8rG62MzyUUasXAjcqCACmqf+nkm1GZDEe2jI+Xjo3lZktsmJxws13jb6BPxvVyGheoE7qSn2
00Bd3bNSujfXOt+OgYZDy5TbRCl5MY40E2dm2wDUVDIK/xbKa5RQWbeUBNsmaNkqYYDBAjIVVqeI
hg3TBZr/efbFywjPUyMmhgQkfqZykEX7hf4Grg3P64MzVRKpTlsVoApqM9f+U2XL4kw1G66vyfh/
+o9nk7VmBI1G14OvzjCgcVDZlLHRw5HwknurCN5KBODYAWhPpJB4qkm+FbPAoDpf+GpEt+jwrQ+k
IXaMk/DlvnmQQLHS8IJF7WLC0rIdR9J6CQlZqWMq9QJy2iaV0MG9FyLqogDkH5TxqSe86CVC84bc
Y39erDmnubaTyEpS6hkzM2A4TeeiX2LMExHniQcV/N/c/ybE3iTrAKMRRx8YGx1xrnxmP7UcZGDK
2R8U/QGUnErAxKiG69lggJelInGbDuokbNqoPxFBIlyC2xu/WGOkemRFTP03bi0ENqKj1MmBsMwN
scdibdG0VPMO606e8NITW3HPrCj7FlkV2jgVsUdTZ4DASImPPvIk83aHr6y3q0HUzjWf+cQHKTpG
EGjBYZFN6HnJYHCltcBvXu5xVuO5wopVAkE6EBm5K3hxqMsXZwkb7gzWT8WoOILtnQPr09syERY8
AYYssGX1+Wl3guwkClLq4fygxRozxjWIrFyVhEbHDh8zFaTi5sZLTpf5yppisX/+kze3xrGy4b5r
A3g1wIL0ekLz6LOr8tchQMM9m/CHNvz8SbYPFRDYEnB2ONojo00poAONeXGUGtJuSjmcvGEJxTOq
ILVCBxf8tX6mux7CaUk7Hfj+FidttwrpS7JnAOEtTCx4x312rmX+VH9RfPscajo2n7SYWFrHp0q5
ebbpCZn5OXo2y0SR1CKH8HnXwZ1IHMHRCCNzCOwrnrE9n2c6FmK/X3YjwPvDrsF1Wv/W+McmP/fn
Qzl48sDNMm+Zo2HliroXEoClVntdKhCTU4mso9BLCOhbyyyOcwzhCi6UV5pS+aCiRVn1YNItGbK7
wjaO64zdw3Tr0/1cXJMHX6VrW1YRgxxF+0ev80nHgagn2SP38wItC388Eyi6SQexig1RH/Z4JcyA
OB9gucbrG7UPHp5sjOwp9MiGWEgjKIrQGcgfo0oc0zGPdbv4PZkJ3lMFC6I8J9sD9mAps0G2FelT
YW4eA6Idn3MPgbiAnQ0HrKc1LadBMuP5E2ae5icD+6ZY9Ak+1Sko0bdjTRL3A0qZeJBvK7r96MTC
qUE3KR8ZHjxYuarrD9ZlvDY3EqUuZGYp21/oGc/X29cHuofy12meB42A5mgySeLp+Q2WDHiZs3Nn
K9dNHuGj4wTfX9qvgc2hLrqzP5tY68D4PkzFXkCabFinSDFtev8vryUtNwDlEorTJenm7mSUfJQN
nyDb0tGPHaPEBSoBzuy4dmb3KHVRUI9SwkjH5FAXQYQwS25uWT1r9Q2GsKBQj1thJ42RF9ipZVjj
d6mcIzwwD9m9UWYo7woHgYaG2YYkG341u91sUTThUtUusCPCY8cbVPLHF8RGS2jexXau7F/eOwJk
2QEjyhfCZJ1VLJ5x12EfCQ1rUrzbGhG0cDyc7TdKPzN1fG7FQcMH9jbHni9W4uy2O/iEdTXixGf+
nQ7sUxO0iTYH6XuIFTgMt1IvEOFHtBNjDWEmi/7cgsq4De5136vE9cKPDOkQwDnazA0vvjrJE41R
cWCLjCySQO6SeOuuaAfDeMkeENiMXvWjoTexrFkxl0lnNig9E0CjxVBgl4Ij/MnxATsCk+I2INt+
4rn5l4UKaIV1u66Y74dNqHCkJ7B5B2XRDJVWDRAq3KI+n6gSWHsTG2PKVJwyKbA4qH2G0G89PfSf
WyQxdtZJrOq3Oqrf6z9RMoAlvPGGTuesxjf+UwRoOV/Wf3UonZa3/hfCnji3ODC+CjzhcO3C1f/P
6h33aLSMnZzSlelR7vhxtlkhobKRWD2Fythey3M/QfGeKhNa7Ab01XF2anh+o0YWt/kZ2YaTmKsf
AqHQ5AjkyV6XP7Vq16XM9uBLTjzI3MsPWko561vBy1cijlqYsz7kUQzbf4rlVM1zfsejAJD1kX18
67kTRDeiYMSfo2uYJ2rzJkbpI398aziu2MJmzO3Eplym6j301KVPUE8wqHubNxXZe4HxpJf6sWrI
NcbFM2T9y8gFwwCpPOEHa2y3+XlHF7eRCGxZqk2/fg0G6lj7vHa6zApm9GaSWxN/wVEih4Q1Gx84
QXc7rxuj2RGAbj9XzOXrb5Pj6GGZW5WpZSZBMVkB/gth0lNud7v91Gyz8hR4oV13XPqiTK4ow2UE
HypYxZqdEcezW5HG91OvI7G+RJbpW8ZhAY7q6vtYnFZwbio3KIwP8Vma/4fXNLAp3tZWTyKIhIvf
Kug25bkf5UoIZIYYhEEeEkNYk7gy7VVXZIxrNKU1grWOe9m2/FGPeVUYo++Qvr0cC1eOrEe6D1Ga
OI0k3jtycCpIrLBQHfSFaeP3B5mkFegnjuth9rnQcL40Kg4DuBGT7TevmHH94lg5JDtf97BDDFAM
/1KVCaBVWT40LBC0LmdXC0YGCp4V5Mphgk8qBmO+VW5nZiTI+JVy/DLI8ehfinjk5oMZf0X2Qjvh
kGkZF1Gulx/EtoCyO7H1XGFapH+LjDJYmOlYT2Tx3tAKz8KyaO+O2vY7Inia4oJj+oycZBZltHEG
dOQ159TxGBzXG7xjvbNGo+TJykEN1gC7RyBS50Rr3wu7NDL7dH5Nnm98uFS/nFTdKG/UCWMRwWBs
FEExBYA95Sv0oQIOsljlr3DN6uD8Yn46sSmPPzJdJ4B+YEb+lud3up4G5raKlBprHaMEiONiBB4S
h+A2dd5ruroN83WHDjtJzPufDF0w72nOTGcJsb2XI6iFo42wvIZ9znSJSfUuC4nwJaF5R3O6aF9N
xvRqK04V/LKsP2zT06ufNJv2DFX42RZKzy0NEzUkHNLPC4YD/7ldxD0ALtewTfgUbKcv61rFJ5jG
87NtPpKi/Xy1N1BB6yhnAyYMNNyHRLGYEckKKd8b0t5dk+nC31sVW3ZHRU4XlZgWAxwkCnFha6/1
WLjyZNntUivedbCNM3ptao6wjQne4wVFSXt65DWqyKmXyqdeqx3d8PahQMR3YPmFyrs9CIsajNUA
46+fvwE8unE+HwwSmSZEkbLCIqpACVvgcKY2hdCdG5pgM0hToWw9aHVGK3CaTLpUO29nPOdlunSC
MMFE225Yo7dToqVNisd37Sa7Et2zoSA7Q1UF2/nqK+8QIi29q95oimjkjaRbEkkp0NT6eIKxc5sW
e4NdDRDCAWFKWYC6PSXDiYBqvjCgpSN7EvyE8mLLT2FSbhmRrM+c3SA34DwEVMjBfEU9IMwvPwMQ
9kXqSY18Zelv5y8f/BndhttmqmHohVHu6P8WDe/Lx2H5mFtt+7TuPbZ79HhuRg2K2UYx5GYjWfZ7
MOtcLmCfyekDGdy5Xmv3fZea0OYR9IZB02Rl2tgcJGd0r1kUVyM+eBQNKoyA7lygBjCNIgo+4966
ROqlOsHeCSJ/1ML6nA5bncZYcoW0GgBBL7DW5JIGKwBXFTT9ztt6Dqpz1oDqN0Gb5sPvTwgBItvN
YPhOLeyJU/URywvrdOiQu9bElRssP8WtyF4gvAdEC3vCRQjwCAuepgL5eZ47jxLDZhbsH1KKIwQ1
XkSCy/Q3RlmtMFSY0P0PM4DhR8PsbZsGR9slFHhffpGdU022ZfSRGIfsVHSpKVJSYSQCmLmTW+/f
Sz+5wT8pZ9OrTXvR5xdXU45DvUZ1MggVLZh+H/MOu2HUj36MxPEzZBqCvYWZMBtdCD1U0HqnSBA5
HAKcqSDTr7LIy15kyoYPI4GKoXzsUf5hcpPEQV1Z1XzfCq3nWkvTLMH1Cu6Jr8StBep2EcKjANF/
FIVVTQi800CrR/UB4uwfB5+kmnzT8CPdVV3sbzlD4lWJJZZ7O1HSKEEN9Vg1OYMsqHyiqFYnvlsW
Ndmu3rJ7avvM0xrFzH3alZBVB8Fe3ox204bGEhLnBcdtfaRVtf4y8OG2CPXk4aX4yku8mKjMZQQY
yxmijK0Qq2zO6I9SbDkuAws5UL1xysBFaTb7LSvYfmHCnPx4ehb8n9jn3l2OKu/R5L7eI4JraSlh
Fpr0QqhE3RG3xunbC0t89VTrgBD8BfpnVfLPXv0WifyiJ0msdTctU7kjQFIYiKeDAB2RPAfsI5Jp
wvhiwN0BIotnfx4PvdyD12uCQks3CTpXvvjlzIhwhHC9/eBKjhtitzjh1rsTnyGNYD/i0IyoW2WK
yj9doXfL800WvOFC9T+/NmoOWu0Z5/35PmeozXaOFBF0jOfQJ6qNoAGzFMGjlXFLnflOahTiG6ua
tJOd+D40osghLDN6xmhDYAmiXdSk9ta/5yimqc+KX6Cf4skTDjtnT9IE+adRNHbMuZtbscKA3dgO
ybyvNauZRuhKF/XvGxzNAqT521z2rSjUOPHx82Dfl5gBC+e1EhevMAC0wtZELAiOn6D5VVs+uZ8z
NFJZ8QbnLyO0PdwTUXrDrn0OrZ6tboCMRKXyJiwMm7BygqrTycHe9ED8iZG7q/sw1GkxsmIPDs2I
OhY8C90SOkFN8x11VdHpj2uXjBpSxyMU2E/TwdMlJ2xVJcaWAGjJ1WQqo+NPQyZtEDOOVCUiXkWc
VsQj7iaGpeqy7CUvUTuckk/i5qgoosuOopUVVsHUEwqhRptFTGepas36laRBKuJ2HiI1ra/yvZsF
uXb5ZSwLhlArJU7n/mDC9RuEm6rYSHrvoRmnMzDX4oVZXEv9uhEJcRmzTjv5H5F6c2TMbPdR9v6W
nNOg+C3dWRldAwWR0FLnJoGQoT3ceYKsfm2S5JI8Sa/DwN3fiAuBN/+ZsKVFihk04gT+FKlEzpLb
mIrhMsMdm0Ug/rcBA5R2dL8DErOJYu2rjwshJMSQ6y37B1m3ykrxv8OCF5wUW7xgcOhdBYhq8euR
DiLkU79OUjWuxQkenzdYJHBiwUaBf0UKNOxFaHkOyr8HwNH4Xk9AzN3MWeJ9LniwvwefLlHq2pMo
1A9ppvCfSu64allNH550EMRHLZ23bb3w80S3u/Vxc92mEUHrq6ZAT0yttQqaZQ7Bt9MZ3m2QHA1v
MElMzBAFg4HX66b88/383UhdYiKkm9vPf4YKPVUWg00uPnGpU6LDjWHZUUoCSvHPr7VE9p1FrrPR
JYTUb4ZNn4vfAzTzVaiGQ9tTQ9uOjKu5nkr6R5qgLhnrNcTwwWdQP//Lyo7r/1RvVqxoPGlnAJ6F
DUD+8X4yFQZjkXDPn8CMI7KIcjIr6BAmf3cH+WH60cKlBA5D1lA2JOxZn9ghqHrU2qp83aS0b6hm
fYdrB3/xruhp4EmHNeJ+a/lGI3i4zR2qOreBZqEc/RoOk1TW8vO6OqFWug9KB2Ge/CGoDDhBX9o2
yC3x3uSwkvVsRJE5zKdDHBEuFcBH0r5s6N8YyZIpYYildxi+DHZXr7ymF+fuKw0A+Qeh6cMJkgCy
2dwG9X4iHWLKtad+LwOBHb5BixJT50mKjyKe6fjdW0dZ/u6smXiYYqNKjUDyBQ08nA6LOBnzBZk3
ul1RyOlvVMSZ5c5k5Q/cpyH5037JF5rMxGxp2g3stqJ7kuKPOboYo3CtZwgL0RtqXDInRQ6qJQ9y
of4VeLk+1ROI195M3S8ah4cLVrCk0yMScqK65o3nH6bFKByxKp0K5E6L4skCEgSeq5Mdr0X8Wcsf
Wi0hP2xEQQ09wptEsU2wf3JDKBqPYqPfRuPiNp4rvTBLUVNs/22gEJ5HDwP2ZISOggceKmpcLXX/
w/Rbx8eAPIK3EjFyHZ0ZZGxcfEN+tlyxFU7OeFlLHZQ98yXGDzjXN8ZG9c2nP8T52TW6uf8qY4BK
W1vAdfDcpgtWaeTDvwZGPhJh3e7hzN1IcsNWlUrcszzMZJwkyYSn/GrVWxcR2oHxa3Z/zKpD55WL
2UMWuF+1EIVP0JDgcRTOlurK37NAYfKyRBgp771uuxgoNZmzFolxPII3TbHWcyVlKc3HrnL5Pn9k
M5fBkF53yOzvwMl+9sO4NOxebuUHdTdFwmbXOP5G94Qb3fAiDUraKOjhRvBn6F9qbP4mTuG5PxoV
pxOLpuHBclvxXYA+6q04Bn93w+g1hqtn5D58oXTl6noK7uGQFP23px0l3YWzyjWuc0lMivsn28QW
AJwrcWVcVqi9qGwkUvL/skmAsCTcZpSQri/duUnYhCenmILk5qIMEtx9cfVulNNsWjIqun5Jaz73
SIlDbcGi5OqzntWUh2TjaJI8EsYvcxz+ffBJlUrheNJPHJdqNXs8Rf1Ik+0FXgmbrt772IHmEqvs
qTcXkvxFj/SJRPoDkIa83E0osCO7LzjIcxbFf6n9sJ2xLU4dpqq35dJoW8OskSLaggZa54JhJ8cH
ITCpFV2+koyAbAYH/IVjTc7s/raQR6aPPobabDCn8bh2ftXWGtlKBBKpormpbtW5zE3lDRmsTdjG
BQIUMpAzbL73dzlz/3V/UYW7cZBYS8Y56PYfE3w3rNivY/PJJrG4rF1lxHB+B23YWxG2+NyWwNps
NwVqcIi8dtZr/4MB31en2AArj6JajZd7x3WaMIKzMT6KkebmTcCvIDDyUb+c5Ln5761u37p0ChsE
W111ZK4byxPRmnwZXdd/qe8xegufeEPNDqh88gsBurxh0aGph8qqMExvIW3VCkXCOHWwYHB+m8LV
ITCJulg3935XYHxsGOvkRVW/8wSxodpU5ZS02QaAkEjBGQEQ1NLZqGJLj/pb734nym+JD4U8RKjS
h3Petmyat6CbO3spWN0ad8N/59yvRA9aWVqyYQnBRsfy876WefUI/prRFK2pESk/IfREInH/1yHo
aXe8f/Hpz1gG3SjUvvrZ3LNYfYypsiyD93Bw1UajBfKfocY09MqUUYAF3a7S85p979R4sNcIy84l
guvicXA/Uwpjng4X9/sCtbujNa+5/EbMrrk/YEPP4DEbk+oq3+TWXwOmaudWjamTJEkO0lQQteSA
tSRRj3N8JL6SNQEXmxJQXxNTKfbFjbHxohbtoMYhH85GiErAPWHaUrDG/JtcGbhOum31GQmcJB4/
gFU1njccSxwiiqOafNHdeWLH2f4sbyAV6z5E312Yry1hx4oV/S5qckhoxxfaYQcuZ04oMaI5Sr7d
Xi2ZZor5mE8fv/nf8hypl0/KQ32G/f8GWfvI61pQ6hy8Fe/pbvBV7DV4ByKgTG8aqgL/Vufw14eR
bNSssriqmTm81PnZxdLEuGwuGeYqDr/+BsqC08Aa9c0q/N5eE28OJbL+pM2X4wiv04v2r99yo7d6
68ujTsJyH0pz1DfWRp1LvULy68JmKwT2LfUcR3HJIaHOiO+4xGU+EAlLLyaiX2kp8og1lm+89bgW
QJxA86MEr75rIPmXSRwTJNVjteWx1/57Gy65e0bmBuJWcWeH4hasz9Ciup2O8Bntc0BB3avoJDRH
RSa2GpcsMGSjBXzl4fsboKvCstpD2WE1/flS3Afx3ryPq4d5BaSs82SxmdPxa76z3rXkOuTPTHed
XIJhsFyR9KXFwKl/KIaz+Rat7yU0aI2OK/tzWdTVLf4Ov3XDcxOFlR0l0mgMDXgvzc4bCrF8386c
VObReh2h4ul5/Zg6gtvufonercoW9hy5DUBUo7iDv67F9Ubg+F4tiaktUJ1BCAf4K+R4aELzoO8U
0ovMcD7Xjbi2v8OkBNK4UrF5/hAsESnnlc8bTm32naLGzjr/JZOkKQ9bnZ6qP/gF3Bkw2MeeSGDU
qJMKi2JCFRYC9g/RiWXUfK1WfLh9GpC1JimSfJ10HbONZuvp8j1ZYfSUxSXJ00MmYKb/icYjyUmQ
8ajIRvKmjN11yMPBiI2m9xELO5edMEJ+n2fSNYx2Q1su+zoCxUnZhYGg3lZPhf3uJme878H0YkNi
IxI8BLEaRj56Wtt1M4b/m4NPikUXSLzW3ppJ683ygPP5TKZ5dCHMNpk6J4tsH/rvWqo4HMOuZEul
CbYDCnyS6J83+ZQ6fK3QxFwrG2B3E7QKozC3OA4OjWcbHAgZojNj5BN1dUzE+mOVqnS5SD2Q19aQ
E0a3NckrtfOZXyJKZ8Tc8X6tUiIILWLjdNK5OQ1TZyzX2qDPOSG81qclMPma13G9vwoBR5omnJ5Y
uTk8bd+09wHT+UFK77AtZxS1ZIfkuJNgq5UlLPauwxpDA+Nlmo+A1J0NUKxyjwTjCBlSJ2cZV4Qp
Mj+MV5d3HDCTlEQK9sD4CiYFqyP7LVnvod0ZNJxoN0b55kW6QInCUL5O81SLqRby9tgZMELr9Ad9
wAVybt4srqZTevVcjMIoD8eUwNfqP+tSUWuRkOv4V5QmseT5yxdPvfyK1aOb2xMIAW14yBTASVv4
zG/1QMCLLgJBxhjFmKAuhgJdx/dVeWdAlo3s4APj5XWaIEbyub6rvZ9mgJO0MBsx6nnfI6o+5Kpj
iMtvh0aTj34s/OXRMFM2MXBnfEST1JCqDw6fw/abXpVn+m7z/CfsXFbIdZV+Lc/qwN1ZLxIL6qwE
iN4av2s0XwMRC4TKrcio7bIGXL5d+oI93gEFA8i62WZbKkrRMN82NZvDtwkiJ9wTdMscBEK1cHSy
vtg82PDK6bw3qmxVeAUvpI+AorD10MGDTeUqZBsJtjGXjEDkzbw29trTGflMQoVToVC+TSU9TWyb
18TD6q1HLhypQhG8IKiUQAEYOlEMijBt3NxJh/v/ENZrlByLVyGSG8+L0Fglw++2ZwpDGHeMx084
l0DDL+hVo+bbzTOVlcKO11WzLuArEul0GTt1EpO+6BkT0xkm4LWDpLtI2ecZVvn6OHZVde6KIWZI
+qJquk82LltsaKIo4pwif4dvVp2nOOPXyOK6uDMJwNk6akmD3nKazl6cE1g5B/JfqMuIMmyx1NXE
kKs3lRzRGSu+Mb+BNR5IuK9wJmwZTpHq0sUstSlz9TWFVRTIfemdD1M/QwNzc8eVQz/E4VZWa6lw
p1uyW/a/BSUWKbcH/D4/nhOxTaqvFIvVyrqoNe6DXETcCz5mLf4vc98mlNDXBO8fFXCBbg3ii48U
l7nsZMhzACcu1Y0bNQsbIU/jLFaJH6iF6QxMDU9a3p+LdV2axFy9WFgpMS1oo3l4Up48Ci2B2HWJ
Tu8Ux+qOyARAsfrtCT7likXQDzSVZBlPz1ZUiKWZKrqhZmEwyUY3Fo0sVO7Yd+l/YF5NLIo0o1pM
Shd+3EeV8VUuwFcA8WiX5mMXLYvqIuOn8GVD2zVdutuFpP5eYeZgC86j8NNxRy87pqLdNIVwsnT3
SzVs/3XA+QKAaQfxF9FE5Cm7Q1B4bGu3qF37hNCeiVTXvYfrR3zwPjWe2NI3IV6wEwJCW886TOOz
NN4obdigLcEYgiZxZhXAHnuNzkL1/SKZGn5MWOJmHrCV7Fs4sf7zFqjaQ1Cg/Nzul658VflJj1x5
2LFuXex0tU2xeA8z1sksQWLgt6inyq2u/PO/yb7r4ou8KZ5RISTbK7OhCc28SWUu55HApR8osz2w
AAFTWgWo/QzrJ5HONjrBISmfhAx+iictD8HcVHfINKODNJDxFWqD3Gd4nELqCd+rwKs4RuFCc6SD
avH8vzos74XRLRcWtrHMgtleThM7Zn9yQKE9mYQh+2eOrRbVm0MrXM9AvLBUfBX9OHBszD1W8UYk
0U9G4RWXpmnJ5lKTmWyVvOdo74HDtndNiB6SZlM9UiXMHjLl00hCsVIZJPyD1r2wmbQF2ulbx90V
DuQsXqLx5bEoKHYTQgxohPlCgYbYqJsIwJLJXZpcAxD8CuiTevXtSufArCQ3nWa9HTpz8E5x4f1h
Cp98NHo4w224MpwKd7bHGZy2rwg33kuttlGqFtVSXh7BqkClmyVZ7Lehzj45Ca5Y8P8auSkGs4RJ
mpbZjR/2mFTF7oNc/7QB1r9Qn8E4HFgBJrK8R3NphgIduvECWt73juYUnCx7O66Rvwn0uUL7r0iv
dorcM5PyziHl+ML3zBc4Da/tkzHPRc0A4QFGJIs/5O+5rKb1RSgo1dumZs/CXM+tOxlHKSRcEWdK
6WXoMhK1Uh3BXokVOBLS3Ab88E+s6MsrcfKRSA8GIXckG7AHeQLs2H/DyFEw3NUD+xUty7A2Upfr
WeAdZUgfsrW/8bsC4Dl2qVP7SnofViL0EAeUWAgeHpi7ypx4nu2N6etbLtiMauDF/dNmdWfZXpBY
qVVmc16SZ/6kODqfGhOeIhYECm82hWWnYKJXcNeNyzpchWbn3dQ5u3IsK5/X6XYr465usuWmtSwf
KRZEI55fjugSfgfdOzgbN0NQ3dnm54bAJ8B7JPQ6+pmTFL7RgCjYL+HJVGeKxbN9TGtd+jOX2a0+
kGXiQJtPNELJc2GUkNzK8jmOw/HLajqjCJDENPTL09OgeWaobowq5pBwSqjtf43NiAnsFQSLUfSO
M3QydCNlKj8I9kE3pZ4GJE7SAgBQ/RD0M3MxSxLsOctPOKEUwgK67Y8zS8X4ONj/Tj3600jEWPhQ
gw4UkozpJvjG7Z5Z5WO3dvnGaUnM3Qnzt+WdIYggBAHjq93zoOOlNu7Of8Aag4CiSkkTE5qO5Z2r
wZfpC8Q6tAeq2US2XGqaXiUiiHIpoK9JeKPYzpMvlQA9X2tHJjvVMJkndocRposIwLDtPUP8o/Xl
tNE1QA5IFAIlHz6VARIMuJKAF/LNSAHJVF79CNlU4DxdPkEFr5w8rvQM7k6nLtPND4b1z7Hy0Cd5
qk40AZwNGgr1NGm780MEOEeC3jsFrjK/uMsHSIBa9EMVlDW4/2kZPOjrYvQLFPK2LGfodirzWWKb
sOGtmnjOlPeUie+9DAL7d7oKqg+5knwwjEet6GK8dFBBohvvLg6HuKr2TogoVrMTM5n39aitf2VF
THkDbZeu8/B69XuZI1KxDDbVibqjPb9P5WGMLyIwmZlqWtvr1mqFXjT4nH8LOKSnRQlfCagKKpan
P5p68estrtGx3+LPGzbzWcSwCN0+v4etLTAHz3FkgJMykCLAid8hi8q8qYdwdGst6f1chvCza0bj
04MevKqfrQw7U46RqjHSXsYkV6wiDwcRZlXfkZnNM/eWfparrPudc2ixHCb69jAj7F9tssKgL0Rd
kQbFYVIhNVcaJzlkkJmdY6a89KmJZNDlThhRPPztIH6BZ/QSf08c5UVgedGjaMim3Ezr1d9ToUpY
9k2FOStwKiLF6MZF7mNyw0vacC1Y1vsoq40pi5JNV2Tq/5hGf1L7OxPNq6VevWQfQ4qPeZmkVgWX
vjzEHDku1iKdEFo2DVlJvqvwAPy3vp0/o6CKKunPk7KKn2YruBsSeeAh65NYlSll8w7ssr8+HMfS
H20zcxMsJRGUd2hA+Dmz9YN7AE+mrvYy5do4ZgcRNzlO+oGFFqk91s4PA61YFWzkOxCCsMyGVlY5
RDBQJxPgXBMvwUYSzHAApozXnh4NKMRmEM3hFZBLEMvy1jfLkYv1y1q+Z6rnhDHztYCCOnq3LuM0
BdozrXSOHfdFi79ggm0HqAU9273dnwuCgk2gwe9JylYRzB2WzS/2O0ii3Jb+P1usFBIl8WxHFdc1
7hXLKaUdySMxunp8ltCvr3ijMqFb4EgX0jSxUfwOpo/G8wr5pkISSDp0DUhFn2+yCuHzaQ03r3zf
tnoqHXXI6Eq8e74A+nrdAAx9OJUuLFFt9u735UPwdJjFxZRWwmWiDpYqBF+gzp2dgPFiYcq+jnWh
tql6iGFlP2c7JZdhiy46nptlJVK0u1kWdCuanz4Mz7POJODsw4HXGdAk3IUSYST/oZgxGINaN/vw
XF449dKMlAn0JxnIoXPNlSt7bQc21YV4C89dgPKO6KS5Zsy1ffmx5Hn1IWdCGMiqe6p3Xx+VnCaw
n75zGeixg3iT2QFtSkWqdiFhH/MaTK2T7g/tvN3TEcMFg7OxPqMxtLy0jLO7rZ2O+t1UpKyr0R+k
+bRWc4zPn9sGObmtkWu7q6FYFuHpj6zulX1iJwMZuSQ7+RsIrrxMNv1IdgNiTQDAjq5grbORWuSj
BtqJbp7qshdihd9tr6guzcnP3MBdRuXDPBG59AMeH2XftnooVuvJp45LTMKvGKHkiQT7ML4dabRK
d4yjbRD2Ro2+0NjdoWwp/bbA5g0JlKFpvbLiQSGxbhB1sR6hIM0poAcak19O3rUTv9k338OFxmmH
RYKsofRS3KSIHeAOO+Ke+9q+/pqzR/Gx7luLahGyvkqe9xhoZJc0Q/UVAUy54saAqiW/um94rsuE
0SgEPvJDQzgqJxrTuwbFVyZV/X4iMID60FIevt91SEvh+Bx74LKaD2duA1T2vgaBNZz3mhNi0YJK
TLIZDtlEUvJrM7D38av5pof4tVqVHHluc6m69FEHeU12wethr7Ibm8WlyEQbJOWZ6tPk8UZUVOze
XxlHMg0YxOuzOcrO9+gZ9VwP5nUqm0Jiw3c1L3spcPaFqEosmvaihRhpmZ1Y/Ys9C6vv/1Jl6qP3
TgZAJbZNidTstr30BJDh7eyBkhuPmdnAJvvo/u75AKF1+x8TZ+i249bCpyFUj+Q08z6s41Xt4RUS
9O2xqF5MENrIamqkIALOzbeqYJXWSwFQdufe5gsHDI0kzXf2zU480qzEQWKGSxKyL3Bs3S05538S
DdaJC+PrSLczgOqbByE7AcOAJ0/8dTSeIyHDRz955RsuPwkTEQJl1EZ63Ceh+ERfEsahmfVRqz0K
dtnY8JomtEVlGlvH6TrWEnO/WghMfdp1XsqmaUbFKH81tKXmrI7i2eVEcW3DSZ0tjx/LE4L0zR/C
mIWORF6QtGYUBkxw1HQDl4dYa07dG4KrrC1KEiiuLeVhCyHxahQ5OpqQ2q3+xqTZ+SPkoKRsOd8C
q94PCfwQ3nZLBlh6D1YSBrNgydtC0Ciupfof1lpNqqnJTROPk1g1GV3DrLS+WYkdLEUTQrHKSImC
db0vL6JuYbivfm+o30TPKfHZvPsEZzcXHRtczJZrdQ1CAx/9DjOIBYbvRkn8UyJP1SutA7W8tNHg
ZM88zKnvyzRvdl9Cc3uqy+rF3QaW6nBGbmM+8MaqB2KCER5SSMbnCS9nOqd0+Uxy44/sIY1PV40O
GRj/8rZXjOesqHCSgOscUKjjCGbeSDS7v/SduumqzrExLtHgV9JWbXmhuXkef1o7oJeLsDodD+cz
Q6fxQxy1zxjv8mIBcKMdDxPKCkLnKQc1XC9GE9Yn/zJEyt2dWNjqFUw8Qhy9nblnq2Keok3hjvtq
u/JS8K0Tbs/X+3QXFkdgJuOsgLtiG0PH6qgk4xog7WqDP6kkKMKEmCSnWhzjtteXajDuLp30gGJq
ZXV/N62Emoaq4zuoxP7Z1LeMVDriaXNksNdWENjppd9jv8cQLWIE/9VUlOForeN+qU53P5u5PSPd
Ss2D3M58f0Q2aH2EPPvtREIDDhrNhOO+ez0iH6W4ZHZ3aSZ2bBuWUWXac2q2Uu1TslryPOvRYfdq
AwSDGNCxoIZs59m7EAO2t9qi2yF2rynAPWKVrKTUDPl4xm/O1/IyTu+xZFt1ZhwWhZJn7zopcmRu
JCYgNxe7GMym2lrtI6zkvcr01MwYi7G3ZYfK4WoypX7M78z4SKsEN6nwhHb1dODn1z/WwYsMsXOI
nXiBlmfn4Ml+cxMjESvDi34DlTIEAKTj9HM0oyXLuq5r0Y8jWJ8FsIS38yEjlRB0pSZhkSxF663e
tSVSGpBqBIXY+iz3DoAAzzf2bZabTXY5EKat+MH3BzL8vGBIzdIg1Nc5ca8zWRxSIT8PQYTyiyZh
psoL6AKyHzswdgsnUe1+18F6UXYLEjb2tOtxgy+aDrJ0NkIw9czEgCrBSpkzO6Df/kTsUVOIbS+s
eU8JRvm5WIzRW8osEkha1us1Q/BxTyOmbz2VG0QvhpZuMCpZ7IZvZgBNhhO/hTfjp9bOfax6FqWB
nIVG2JaugtxaAC5Q9ELuf/+7QSkqSLtK7QlRc/fYqra6gYRWRm0keqyA2nildAXCMzAp+krO5VLO
pujzq6uZqJNaVpHUqMgEOQvDbqguqO4u/0dYuhmkSbmU2AizgquXTKm3kFi0wcEkwJwy7YUawxMy
F3cZ9VEQaQwGFF2QtObq53zB4yCrE8eO5Nv7EMuurVn94mMeA6EAMHs+GNCVHZuDqZMUCxILYH6X
4V6yvfSw3JNoMiTPCzkA1a4v2Vgd0paSrO/KhglMGrJq/k0BwFY0Ucr+saKWbxnz+qsSfyCaO8Nv
FnSskwzP1dEtrwuiGHCClHyZ8YpbYcEr4zM/29Jm+hODK2btkEO4FqU7zwQcIDknLqmgXXOiWVAY
XHtCI+DlW5bKQ2On5dVKRKl2XRuCWkRyaA5c/76VffPlO+rjpzgtLJZ2kSlQeYBFX1y9yreRPAJ0
tvlxrvtemoImuE90BRaIs35o77yc6nNZP5r5Zm6MSVeGqc7W+2bIyNsdmJ5oodPgJ5qOWYUSi23w
e/g6lNfXKqGvm3waNg+7blPNiQ1hUvlYCR5s5/izcf/oliuZ/oeqaSd/yS1s9wh+ue+WvXWSmczb
FgMqzWuEcUKzqwkvFvlwn3CRXI0YBJMQkHP3d30IZ0n1oSZj7BCkw7wd4zySTANWOaBUNUAwXhkZ
8cWrfUozA3Tb3/lvclRtWMjsvNGGpniAAdjQykWRED+WY3L3BClRE48LiHFZGa8yv2LcX/txAoxr
KGy44NZ3NxlMw/U74RXd1v9OmdQE35jRyiHT+Pwc7lZJAHSvOVOsad6jEsTP8xTri86nkJiAEfdE
IY4eZP30vTZij68llydjpGMjdwISD9bhvqxVLxaHgt/LWZTw36PYn42ueGyVlui6B7crHdmtTRTq
zBFdCWMKPJuiLzK19km2vtsh2+3Xlm4QZCviq7KAK4FdC+YuI9CbMPJqfx20gRX4fqIogspu39eC
3PzgMmKv4MWgaCmXZ51ATZbLL1X9avG8sJyJoUnRLB4231rTCayd5uYJc+Jnn6m5vZRQ2j/P/jlR
Rio4FYe4KSOAdxvdnbCPMVvCL9U71Cv/PLUPGbOruDcL38bvELT/ptIINyhfZBL7OIEunSWWomVA
1JM5JCfNDNrhE0CJTeNY5ssZhQ7/9NB8DBDBZkCyHkpBnAMYqBtPNnzzXKQ9MJ/T67Ua3WCdMAzc
R8h0fWxj/VWU2pPYChJx/+zyDvWTZm9EyLXgWLuFgZe9EnxkJqHU5f9plZAsiuiSW73K9rPT5AUY
W6qKOAnIojexOdK8pmSloUn0C30QaLeOUVTNRjNlBnlw3z0Wqz4x1l9FkMITwauMDq1RuCgB0WUG
MenR/BWYMpFZyAr1/ujQ2LQdRo9p8VbL2xdPHxBILEUc2y8fP4rqorsFS3106dgVhgbRYY3NYAPV
zq/JUlALSKLP0PK9Pb01vG2i0dF1bhO8NNyVpE7QwtVVVakQuhWQmfOazzoap7tZZozOuuhFQ9A2
EzvYgcyJpQWk/V7X0Dl4/g7Gie05eJ/PcRrmJMLXEcpivzG925QrK9m9rIvYPrKKfcB0aDkBk4HM
HvnyJVWeP3vz2A1QLS7ULlaFjiLWduYKnX8vVoXl8AKvvKoTrLitsEhhEBuvsDDLj+1e9Ftk2VLB
j4ZXayONkcjc2i3EiYXV+zfUXFUVNa6ykDQb762O9OOkYinfPyhEFAjfvAJc/Qvd84MFdGzcLWlK
8Pyc+zm8jMgEjlCKvk45iMaLzs7cUGnwXoqoHVY0ZkXQdAsYZppktgGkhGMQeBJfmuRNlZuQAF7H
7NH4B3T7mPJeoaJO3+/Kblu90qNE2q5zw55xGX1ndZGRgnhQ2vmMYwz4Xu3wWvnOWA5wWgkYcqBD
u5pFVHJaSHPukJIifiKftz5qUDiqCVO3QjCWCcYAXNGjt1GbY8kMVqZrDC633mCy1RenvyXzBXm5
IFfilCS8ykRb2aKrZDqNyHtCKHsPTYUkLfsgIp9YETh12WHwQggU9E2wnGyom7Ps2kEbyidqvmS8
J9jgqikccq/+dx7qzi1MbOIxZCn6nWhWPREKUTgau7brWolkYmWY4Jh1TcRY2tJRPabE9EAR/IIJ
vWFbcivwZQOBoqwMUJ5xkTrIDtDgAd9IS7ILPUHVf2pyVEsq+QyviSa7khchpZ9wNuJFVoAx06OG
Qq2zp2S12YNbo+gi8sBTmm8BjJLB/EQtK2phLAaJOtDYJSOgfIp4ks1gd4wSzZDw0D06JZqvG50j
O6F+N4eUtu2MqeLBTXModkldkriWMrrO7+e6W5eBQke3qgEGQhcYkvmiS825x+0KboCgel1nf/Jl
0z/Sf8hSaecnkx3762p7p9sIFrM88IvJMPgK7Y+/JwjUwMR5DenaBeD1GjTz7AMCGyJiQYlgi7iu
NKaOTgOD7RRQWu0HZWa3Q80haKjGpKt1U0E+qIgDeaf8gk+OgD2wUkuG9XPILx+3Q6+e6aPzyhsk
06djWoG0yhSe0v4IyZGgCwjXv3DU44UjLfTP493kA/T/Oa0aWwXKxAJzTcpEC+xJQkdGJnm3FUlv
XvcnR4pUrVHqYZan9flLVFYxQLDxVWHk8zDNqWRXl309o0XmGcugxUR1P9n+1t6yTgxdMEHmXCa4
r/PuUL8Y68M6Jh5ZxgYHRmSxKUqF10UZfywPh0rckyLuVgKka1a6WgVf68ttNp7Qpu6PpNWlFb+5
lasEkw4ZfFoTqUB9urY+mvWgRVts69ezOPRK0YazYbyOtdIp4sA0R24T6yijKVBidlf2xu9gQGyk
2lp671uvfFHfOXOG63C91rdRF82gtg3I1ZdN3VuG3+NHryhkZ0+qgmZnDubxEai9u0oRyDRVkeaG
U7CWVmWww7SzLJ86NQRSM54a7W43ho6cp5CU+5iGxYqxatL2BiuDG4cnmXwRCS/hVdnDYZwnKHu7
sCqlk8D7XCcjdZ1WN5Rh63gSjn6eO7wEuA93nviCUtP2GHDrScWHLS9LhxdtIo5cH7vBXzJpBqfp
5jaUerCNrq2kCZyrtWyc55x8ZupC82queBVQyVGagLOUwotOfg5x2CJIfAemXdB/UWBZGS4QM/xv
NxYNqkqY7t4Snmp4/qyiVBlE2PZ7CuZGnEl9tgsFhZ8tq+kjop+UTYwv36lpbpDFz9K9GKEG6pae
S84fRjYKAo3qdENdymAV0SUT61yC/JfRwXc3aGWReO5XoCdp59BPrZJGMKwF9jPPAcugCXF4o7+g
lg7AlARk27xiKOjGl9uEqJfYGc8ZmcqYF9I61kkEZu5XevtlVvK70oprRSRHQoA5X0o3HFpucamd
BOeX/+0rBoP/QkMdlJYoXsbRoz+SxcnTG+jVJMc/3pefEvjva+SA9kyC6Dvvk83wpkaprKEaGnCe
zeckskKD/NljWPixID5g7JowALFDakVf0A4nRt1ALeHmJ02s+wr5V7GjO5tfGFnAt+YQMxLcAgnC
UAQd+seuMfEn5XSjQmOEif51xajCx2DEPwl+xHlB2vauwbKzXGWupXpmc0vIw91+f0dIMbCC08M7
revcyboSC3d7E3XM6jbma8sUl7jDxJMcFZ8dyZXTsn+brx5g2nTAXR4wSX9E0JBNINY6ssVbGBKM
/d6EbOqwsUFNOCGLasq4ndL3cfuQXhpiH/xCLrAlZW+74uKH5Acu+CGWNwVymADoCGkwLt02ryGL
kHgH60nbXbpAyUIa63lgjrk++fbTlHh9ccKvdA+X8JMvcpY4jQGR5OEVfYMm4Y2GS8JL0SgVYr5N
KGpOUZwhgB3kmxdAdbd+xC0VB/hpYcEtmTA4wJUXfue6XWlpjV79e2tXiOB1MIs7OgeFbHgPtmej
5TmtFNx4uqntoSYJOgJXtn49RBevMk0cp2iARFgvPRh+2L65QSBlfC4rG0E+RbHzNokIF1h77Mto
ZnQGDcDN7gPrd7YOQ1AhKjVOg9OcMOBSCduhCrsMkUH1pw39AbYnK2pwutQm2d8U/ADQdkOj40nB
zGC8wHqRYmOu8VkF2niQnJgh2omRW2O4KswAoXD9t8NGyPFE6Jx+pJw1Sz2uOeEUvsQZDoHrwgb5
t8MioPRg0ADb62b7dE71JgGtjYsAbjK63cEZEACuVXosXcqEBHdL0mHQPBks+74rkwbkMxWTj+JF
50hQ22wElCUxM0JpLu6gFQ4npJ4XpHoULe+HvTBPJYf0YlNxx21bYMDV17rCeoXIjmHLlKjdHk9Z
ZQMBbHCXz7nGdTe+g2nJIMKTzZolOw6shXjznlrzEsHzQI+t7xm0wqziBZDdZYNKLCqcwBS6mie6
UBgRY+NmEIOr2a5VvdQz1hIAbWHSOHOpF9XcaVJZZzOObWLKZQMc7O0AkZ/UmoqZvvLCUIN1yvzT
HFPNmuL2jhAPbyIy+fFpze0IRjcU5963naf1NmfIUBmerZMkiGuD0AdSUTPYBCckVCKnLDZMf0R9
Ks+T/WGWwa57ERx7fA5lYuST/yAnOgvTs65WQgSrMaUKuUaZvSrhTrzi+pcctV9hdEAS6RU3cKQx
LlI+5FUUDDP5vYDxTsvXmsFDoRpzrCoVtqGyIwI8ouglkWfvfqwVY1TUUFDnOyHMlNpNDOToVgHr
4QCF6mnqucJTCXY2DM+v7Qi9kxhYtR+cphyQ4TqqUxZfHHmfFOLNHJR21d0zBBBkVQAnArmJdUiy
fROGwAm1pGcEoUGNjsYr+qNMOfIMdCCFtwKrlJOtM/PCph3DJVuAN3EK+Zeelu8V82k6GN0N0Ju8
HGBTEt9G6fxOAlw4TTia8hW9/4zGZ1YKMoIbtVa4rY9VtXQ/mbgYcduK1Cwp9IKXcOfTQN13UlBV
gQi1Zi77jodVvQb9IIO/nd7Xim8VElMd3u1rf3kFtFMqbgJG1aDJ4TH7YRvOTbasLlbqrOrfDR/A
BUP8ilQX2W9uuPffIruYwhekzmO5XEKM6rk3an76vgDSoULvwc45aGEFl5QsPdIxvoBugeSBeymw
rw13sorwcZy6UKXFTqtt7IWg/oW5PtC2cCtOX3Sn+7ohmAAYrtLdw22gKgzurAyaAwahJR3U/PWo
YEh0fB5PnpsCQD4sPwYgyZ4RQ0k2fyZuO/iblOyxNfT/kd/bOFC+AdlcKjTCojqlVnTWJ1ICOcS/
yNo4iAHm3Y+i53nzcApg4x8sN3RSEhd6rhJJlikGs8gX9y+nERAahlT+27RQHuCUFrsbHYckGiq1
fSaf+m4lE/Cb5Tus4iGIWBQuGmkQRwmfzQ4UEh+GqDDOqsHnedxm2010A8RFCy67VCNrWon75huv
fYZQJcKHeopYQbvACjCEPtSiHM3qIR7UkjAU6DONwn23Rce87EgNcWhuQkkggV477UWPN15NZj8o
86iulKAg1A81tEi70sXc76ajngCJcDUL2Aan8DajddjcRAPcBTSyN2v5rOmRcLmd7mDI50YlfYq4
6ShJfN3lVAckOWqsJC18QsH21PV4Bf6YyFLzAdutm1aygDIB3cgR+S4h/wSSpNkkNElvlfTM4O59
V5b40iWgu4ipoiMCJRyzz72gtOqpWMfOOId1vz7UwW/C5yfsSkvHbn/2usLxdYYJc1KAqqPBm4PE
CKbwu6oSfuRk+uS7/FOIFlFb0KqSxRCrVn21Meg7E5WbrNBFQjIktmXQfMXs5Jpj3zHor6HQqo+8
ZeFjecLZZ+9Au211K4flnjhcRaMoK0NNVtHLNqO3Th3tEJy8t7/6D4foEWh8S6HdodEpUB1F/VA7
bEK7p8wCnM8jk2KKPBrpLBt/3P5W640TNS4P9qQXz+BTBVkkDcBPJQWMyAkhbrrCMW/f9inV9Gde
n6le6sr19EOpUr6EROcJZRlZRUvB9ChrqAb0nIvoQWPKQeaQgrQxlNJ78IF4kD3WuKJPQqfiOYaT
Uv1uZx/rA6YRy9q/kd4RvezXILFLgXLT1J2AfUN5RMZZs5w32bF7q4JDgrp24P6UnB81cAmDoKcC
mSbpj8bVRcGgIL0wo2mZlH8vVFMunUuRi8u7zoc1CB6Ntue/fru92RkdDG7dxaWJBHGmhLEx1QcQ
bjaZyHMzWLbQHAkbhsUXLvpjhFmlUmNEreCblbwlHM5JmR4MXBxgq91BJ5Ih25g1PCwWxYlgVxDY
rb7Cna8bFUvQrjI5dabGWLdJ5xhUSCwT4mQ40J9tRfPl7Tn1DIMHahCT5ACHQKdV447GjvxbgsMS
F601Z3y71QzfsQECGLT9d+LyBGkQo5ZR2EUQOxDpTZcaTncQuowJi2znb8dh0AFGDoWbxNHlN/Dx
GYcbewPgC9xde2FXE3qnqZrQKssTPK9rVqWW0ID3IO5KOTbn3RIv2rLs6nqTPo3NqvLLuDbctowO
I5+1kj4pFvIU0m0l99dOZoNDaLFHW32f3ntwMvCkndnRM4MQ/Yh4KuJ2oi73nCVGXwyPormO1I7u
lsIgsjNBdU3fNE/rmI/qht2113Pg4kFn47DzsXz4LSfYleR1A4c3JtWvmeI28bInpNdm2JiaowNi
ZpPse4C2pOzW9ThghkLWKTPeqz5THPUDFM/ZGHy4q7I4NnlgZkSE4cUTRN1G8OZo1AXf3jM6guKs
VhSxPgB+MaL6ExMvjQwO0/Ri+0XNMO6U6l6m9rDI1lUYX0GgibSuKSsyc8ueFteaCXh/JSFX+jwB
9Sr0H2kAOOBlVnV0p6i1GWdRksnHxbNDrZk7z6o90KNWhpMj9AIxPhKh2SIfToCdlpr6ancj/JGC
ofH/IMtJwp70HL2ltenGu0IYtZGjtNg2TTRJp6daq9IHhjyD3vy98nqYoqY6VKcuegGGIIiKctqN
kaSKmmbECimh+tWsza/g+wHFPPPcd8a71FcCmfX7WdaVr70kbXHDYiobAGA8hUdGDYKXfGVzLmDC
Es+rB2wJxepd4hDaOYpDGy87vPhQSx2gEbyQ4S8wV/R0p1MX5DtCePK8KFsqBFOJv4f9ArZ/4A16
XQWJK9q+CKdMzusr7sQuGG18ELO5bVER3OvLh1Wk1qnH5neEuLWAylfTiy1yDtewXUTQLS6Xv///
KDKW/nPnXDQcCqrNsDMRo0Mnzuq2gEwEDzAaho8wCgKnB9GGGJzUux2lnlZ5THZlupxUbv9pwe8K
BgyP0IVjCHsdnX+WVA8xjutDmM4GbDWOTb5O8/fRt0Qs+LiB/s3EyvaJ3Kw35lRuOTdBBZ7YtKtS
uoWtWo+wsRLwbCaIMeSOrJsKeWlK+XX/7CYvXivRWAT9xALiPx6QI3n6pL+kJugDVZpCf/5RmCqv
FT9VVXHlXAOI0JC/SbWsEx7MJyVq246MDkVjOtEt4dXxSwvj5//MtQwEFIDtIwwY7h/ZqP/Jng7e
QsB5S8kaHmKUflk4BV0jZhnw64pZrQvJOHApJzYX4YR8ZmvoLr9COdJyH+X4gd9JarHi4IUB3//g
mJbj2SGlUGcr7QzPcw1gKeqinFfzKY4DX4yrvRi/Gg6+rvL64WIaICFwQx7MrspfIjdEzKi6h8ZS
ATbrS0iUJrzl1GvL4TZZiLENEBBB8LqfverLuszDZ+capphLkmXXhL99lCE8U8FjqQD4sALFrie/
N93P4ZC/pkREHZM0r667LO967kN2CIftxOnU/rIadN0uRBqlKtRxABLOBV2yWmZGGHmXnBRIyQeD
UvUgSY9KFz93aXIDDTfgxYLBUG5Du1eYSE7jEfZoVczw1x8Je3sjiByRipm40ezwuf/qTq/AWIMm
xgjIGGaUt1Hr74m5g5LDiPz6P/qwb2xP/4CvGJ1ZQ1qC4Z0AGvhLHOo8QInvwVq558wMuBsnu8vd
OfnH6bz+CzshrUaljYYLNjnY4kzOELPbqyA8SewdOCl7whRh4qqpgmn2sahK6Hrss2rjXvxzTa0g
mHNTVgdDErBHirejce+kuC6VbCLLxhbwcs5+zbN4H7GYtb57cVTGMF4ZlUlwv0Je9bJ4Mcgy3LjS
pQ5EZ2/9PoNzdk508MDmlEqsRIDM+0JdjTtgzKF6STlRMKRW+rngh/HpYyC1m1kXoAcQMt/oGUMv
kZOpuJOxlXFpnZeuOkwC5o8AdBw6ksZIWCHDoTSO/8tVOj1UNNxs4rpAS9VFuNQicnh+loO8Bq9Q
sIO+5+DaNm6BV8PkyygKxwscL1nijDnQXPtwfT188EQ7mbnycMZf97+iniJ6bwkP2VO4mq+Ur1AO
Yybz5Wn0Pz5cGXiCCF+YM7wS+lrh1wCsj1D1PkA7N9IFylOS0wcaSpypwsjRXkrhiU1J3EFAJ9Ez
6QnEw8fQ+tfTPWVJDYhOkMKAsRMI2ixsGSNsHuf2YHXEVDc7f6dos6R1j4a6LdXYNP/q2TOgkLqu
GxuNaGuAt6AvZXcJ3HjDARp6z1yRHnG1DSL04uncd3W93Shn7Koo/msBq08X+DSW3eMmcf+bdhR4
p7+rm2htENYR5109RABrFVdk3qzytC+c6rQQIilOB6I5wC7jc4MjGRaRQJyGw2lD/xAOaRE/YeZ9
I2QfoBE1uEz9C4WT9XMsSBs1PC0c5/OvwJnCCYJa9KWjB8Zmk3zCODzal3B/XTql5N35wptLOuUU
oDVLxkrR4mZkgfWGA6K9+GRI7YjWJr24pu7fdCyo1JvKkc+gvI6/jSCH66KvlzDJH5LmobLQw/nC
EtTIBzHTh7336sBAM5mR5yR/EEvBCS8HIBDh6nMUM/0kOkfEYnWfK/FwE5/ZulD55H6XLhIFIfFy
SiXgEfOpLaYpZUjth8nnAdPoXZezWFltn2CnWEON0gafWRtRTQkLm+5wv39tMyiLt5uXZdU4swQ3
uoPo4fVKWXY9QKn3NfVUVrJkatsobSTpYemXFd/f2bjE3R5mgdEpZFS86RBCVB4G9d5ZquUfCPXB
fG6D+d6MD0XXAWxs3+lh7TRvOBCbJeaywJ6YkDruwvw+Lv2q4Ol1t7gSfvR8GyYONuCSBbhS9z5z
tIqWC+bAHqUKRDB236r1fI1gXBpNWAtfIf0W0hxs3RoNvuqC/6dEb5wxQenIm2AzhrWHm9Fl8H/1
kgUyNxAr87h8XvUh53s95o8hgSCmriXLIYEylSxZAn3FYM9OahmlGkrUidohNmwQLah7LPvsVpa3
5vEjnOU6WShjjq7MHLiWKOj4nRAZkmcAIhSV/0WKSiP3sjLZ6W0dT82EYw+RElnjwXCRPxxnWbgB
iK6eKps9Cu7OurmN4+GSFGy/IrKcElGKs22ggS0Cx+CrQJsjpHf276ynsUrqXUBqs71buCdbIAHS
sMPnNJMZS+of0eiGlqFE2TM0Buk25KZeHXuu63Curi4eF9AYUkvcdOyqBxOcmr3dFp1kjJUOV6i8
NnPqDSGmKVxk3ibxzK4Rp8ymIW4LjDo5YfYId0mZanzIyvilDqcXcUXJ8J0cvltWevZyg8KqD7GL
Yup3krDjYSIkPioddOOu3rFIv5gQbl21rt5pLg5qsu5sulT2UlVvd+c40Xak8FsARUDszyqt1vlS
ffoSkNQXv7AjwFd+huM88Rmrpnppir7WxCVtByVVcLiV9E1SUNNcLLqeYjQS6KWvEm6s8GQQpily
wkJDxKVxpKGUpnNRCNuindkgkMC7mZsoW0DZWlug6ntrjzn/aJWshWurAVquTNr9WOTlxu/edBq/
5RYfVQSW8dkVMW0IoXNk6Fn/5iyvOt9+ABQg7G2j7x3kB/9q4p9DUOsOdIzO6LP+JeaxuobH+7e7
EHfj93sxZVoXng+UDptyAJrhkbarCReZL5+vQfWaV31fP1YM6jTC9mtwEJksqkGN90i0j8U1oWm4
i8/HVKFc+0qpjCKNyktRgnTHWfmDy2xuiht4x9hoSszLxdP5bgzmZ1aaqKNDjAfJdNF4/xZXH0TR
rRbsjFtbvpuezana2orYwishyMeR1Hqn2QdhiaTmwBoF5OS2NvGoJaCBwhuzfQwSBz9wDyzFoDAM
/dFs+3J3T6ms7DguV3ZhqTxKHcFFYsTafPzBjq5Nj5A0wt3MUvtX3FxZ4JW6e9oSmwgGEijHeLoV
eZ8YfDfhcB+ME9d29vQyKkdjqyUU3fYM3ijCtPjEJkvJszXMP6qeZ7hQOc6UAWU1K2vRAljkK5u0
1ESXaF869xtcx6qnDMe7u0HOzL619ZFT1JuMargXve7n1CZYY9pQbpHYCx/GiJO9verlWTtPylSt
rtE3E6lNBw837NN5xOy55i1YVp3DAJmRs6dJMhMdZhEeLEyvfKdJrXy1ceoWiC9YAU8Qh/JBFuI8
wtC3+OcXE+6HWunbsd43FAFj0YOB6XoS2BneeodqQw66kiODoFahzAtYKL6Um2nO+voe8Oa361tN
OKUgcd9PdOIDbyX3b7uPHdbxdyWHcXmdYwWcfkdEMRcRP94Hg7kRHE9ber9z8aNFqPHdChMx4Z3Y
tWL9bBwhYOxW3A+oYpXz8fEPdKpWB69CZKserN55LRilTfZ5zLDvZfHeDTrp2JPc5LmDuTXechh1
qteL8QTAoDnUOkgHqN5P8KlB3LSt1d9nUhcL0J1Hl2wBmAVeVDMDqFNL355nTv0nmDhWMz3JDIP/
57njMWxBXDqN7zsM3E0Oy3EbDRalpcOiyaIr0r2PaxSnPYvXtHC068sbPvhlnaGVYuzFK9maBucQ
URwxOly9v0C5uKdo5WsQFePm8QWGEm+UvaDVPHwbXUhND4gQxGYGD+KU0QEKndvqqdLuHlgYGsKI
Ud+BI4WO1Yd2++2PBrk/gYhESqNf31aHpDvIBrDWkhZW+9rZOm9fPDaXFCD2Prei42V50r3DPDUz
dd47a3/FoIDt7aDiu0n0cM4+d8RV8tRKEqlmCWkfvGKrrBKHYLeQTjy0ttelLqh0zEwNUWo1aucx
Pw+bZQcEpEuf1nO2SV6BIPvHVcNYiwnU8/04N7yxNsc0BSUjOf59a2V4rXrNXxVhVW/8oSRbnGNJ
8XbhYy3bWkUJPVACgWnNKhw6OUEXMI8Oqx2RW8Ao0MkSzDw1gyqIP9L5cbpQbfuuKn6YWjOzgHNg
MiNMh2rXHuHMySQeCO7SnkEXWKW8w5tuBWqLFTWwlF5fDFoK8dEWjByxN7STQl/Y58irbDRZeGm3
AO+80nbs6JoY40vj+/rDK0hl8F5rIsV4B4ThUv0dN3Ml33BSOYhYCbN3O0AN2y197CL6jNd06z/+
DksFvkYUgC8+a8rIxcBnK3Rue1RrD5jIqO7OVPCDoKBZLT8zmMmOgASUKJ0oMtxVugLwGRQS68U+
bGNtOMDRWqvHbvCHomqAH0fcvOnI0HwjEzNuJNlnJzZtP35kwpNz792qdZjSdAb0ZQ5oc3trQI8j
kV3n6h3MDvuMsUGGar8oSOcqyrGVy0I4pzhsCGqP63NyoSF5MZ7OdBc50gZS9CsDfdzLvWdMha//
9sK9ZVgf6+UDdP43qQU/ffAmPHY7vlUxR0UVMEwChNHPJIxO+ZPfCmUcBkPkO1ujAoeJ3HeZ5/Vk
Yhdfr5qcyzC4EuEycjay6vnU0AtiKv18H+c2gl8+DJxcbO8ipYmOLoCAe9Q3H8scv5bE+wahQ+xW
9X4wZPBA8crhX7MrEmAf94HUW4EjhBb00ZZowAiAR/nyipCLPTNyfAAfyyipQt6OPjBfjZ5JkM0f
02saDY1oXozjh1ioAfMD42QOPKh4l6tZm1xeDpMIOQSBwR2vzBg2u7DZS8PH28efVr1VSqQ4pYkj
6ov97cZaSco1RBjIR25VPd7faXvAmbcxquhH6hD/XtPd7FIe24+XGOwaW1lAhS4Bv74Qrl8l0Ebe
vogJSi0GCmJX9m+en6OTDhZWiyH50oRZh769eje1Zg8YxDw8oesTZ0Otjs9CmGHYgn533NcAJf/N
mtwgK7TXoaYSWV1KWscdC1nWn/me+Ag9vf7urHZ88yaRtMhIhLFw3tp2dwDs91grGbZjxXi6fyX2
Nk0UllftDeBg7xKeEjHqZROPCd2+b9siKZMFEisBOx2bPkkedqE0qaJjtXh0JEOfaFkP17hmpdHC
CzDB2AQeH5YU1e3vKN5grcvh+TUAJ+nhJBG+TbRnoRhAvYC5bhBkaLmH9EWknbCVylIBvzvGLot0
boEQfue09qs/ASaAxj3/Pvjc+ByupriQXkcVmg1ulUKli/Vhoz9JM9oqg9dhhSJhgsn1P55DllKB
mPjlpaQJNiH+ipGOYoBmFayh3QOQdClHTwWL9SwCP5XBMwyqXZ4WNfaUSfW5tBCDUGyCTYGCje50
mYaHPkUxAvWUEVXSIi7QUWQWy9v9MR20u0SZXQxt5FYO9VUOc7CTtAR5ofSPl6uBOQvmtjMXrpMw
k4gdXv6SkTTPMhT0xN+1vLE2vyVGUQNW4UC8fn4IWiWCk1hCaHhEkBCgP+1SENTIdyI3mdAPiBss
iYOdV8nt5cOYoLXDQiGwH5d8zyvrEA+1Cl53ksAia5OBfV6FCC0VSVxK8FSHFBB8QElrka7szF+S
kSxLqPEEIZRsRUvZJBkHpwRpeViMni+xPp86R2PBbM4OZoViRhbxKtcoxGwGQpMw6MHjQSkBCiFG
9PCE1RTVUyaaTDB33ELeZd1tC2PiJtqCZjcIdnavOA4tBTOT0OAE9zniMF+/SzRjBK69/TW2yuGp
OWBSOgjQTY4kDaKZTzmzzNnK3vyx2k3PR+e3eq/6Pmu6TSFnEfHXmeZM+f4ONv7n9XYiuZi6tzfz
ejB3OOkdcsyL2o2KwHpqOg02mvySdARx3Dnzd4A8S/gDPAdAbxsxPVlpFFnFmudpWEl1RpyoExsI
Iek29BH8xAyas7tHccFm0Pux6Mkfak9uu25fj1viZzkX5qLFQ14Qr2c0A0GkTQxRUOlzgzb2g5BF
1zP9R9y+2kyphdbJhf7GfEgU9Gjfp/l4eQud9fU8ojjGlRdMS5lRRo8BqJvhCJdQJSl3D2Aom3P9
adU0vusrMOuvcoaPlVxOyGXEz9JFydrmy77fm6OFCglRJMGtBsBzYwiMpyIvVtRbjVbUbTQoBnAa
t9oZnvHaf/fPA5dsvGSZXM0hffo5C5dFkem0bxXxL/v6qyPC38D8qPKipDHUNYV0ue5IeSHncfqV
jE55YdNzHcyuXMRuOphuO6T4jlu646y6UHEPQVnnn2+eMnsb7fR/nTq4HI4hySuKaEDIj0Ezc7W9
yCmlHRwj0JZE9bQVs3dNz5vbn5AH8AxN/UoDOwutDRq8dGAUBxK5UdWnm3C5R5swy3h5/+UFGPfV
I8zJJeRTDv0Luo4r+efRImQKAboY5t0Lml3Pp/s4dvsnMKXZossiAv0qBhsmdZ05N5yy8wMiz0MD
OrSievG3QZIVOrx9LlWF4rLhvT6SgowIVkrImZ/r7XbXfvw7ZSHoHGxxg/NvGcWF3IKq5rroct6C
syafTYliXGIOKrE9NZjbDrgMiuhcl/vsLcQAbTdVNnph41d4gtwPzjvC7XIIzgDIZxU9nNcCHhNl
4l+7DsmcPrflOZ0IS8JqdwWVxQDccj6Dain1sZyouk7zOqY6Cs3CfG/OQ7tiLYumDnO185aFNkHY
yMWhjKaLjeBNm23R11EyUBdR00L9gekewwYXU5qEmb90qsmx62LXGKWIQtJqaqRDQd5o1S9X8MDt
9RfTG2Wj9fJ6SccJLN0Sm6TOSnEsep37hlZFx3m8i2+OmNva5zzU9U3ZuprqYRzZSYrzMfypunRF
BA5JRFkwoTfYfFdM4MPyCoBQHk4IeLFp+DsNitgCeM1xx/JohlhbG30xmg9adbcXy7Zmff/J+Vdq
aCtSv1FSpXhjz8u0LWjdFTCZTiu5WCvs2KsGeBsE18pi8oqvcZqPeleIpV552sMM5Bph73EyZS5k
Wpp6Uu6JBsPuyX+biCwLnnTtmFFpaRqYdNGrbZzU0dkzQEfeqfuMjJiIq4V+ikn83ZrnlJsKduDs
T+d9gVeAyQM0GrPlW9Wi4A4npBE03ymOzhQx5TYnA2e7nFuuTDZxsgPCo3Fc1lzu/d1FtD7a7gao
Vc8ft3YDli8rYDtaT6VKiMDZXMkvbygROfMDxHwuCG2gFHwC5xzie+h5cisea9Q+tSzszHcw39lf
aw2A09QPuiTznw/MTD3a7TGJ3RGrCyVQA/wxjz/BmCLzI0jv1PBPtoCWMeqpkmPbqKKXCyHP9QVe
nuf+VWl7dmnb6v5a6H5v7mEcGP/iJmJONmWKas9x3+8AwhVdfKeWtk62yR0x9CBpXuU3YPIPmhzz
jHGk2yUhCI10IEWVj8wlZqbsPmD5XrJG8k56e6XFuEiGEKLkVLbk0vdq57EAo5hznaejlGL8dj+Z
U8/VZa2eZ6jmQWlyzKBD/7HxSLuuct6OFs6dwgT5XWAPZUpkXzhM04DXry7uVzubhoQS/T8Eb+cd
Yc8JkyxUNymUnxh0q67+/teHSjUW56UK5WcrDeev5gLSB44cdkp0brXC5TcDIm3nhPeajHXy7Aob
HMYqA2CXuVz2VdLLEXvl/fzejSn7P78OGFUatY1c708TtLZC9N7xkFYXr0Qa5TzExpbyRYt1NJwg
z9VIjDac3fmZmrMRlezVh54DBuMgfR224csyjBsF4WIZ9bZHokCQ9BgBTqutlUTIQAKmKHqv7Gow
xUShpZqnSmyRwdM+h9KLUJ2DnCTH+MmxTgco6XKxz4rukDgpzbdSW15aou3kDjGsE6Sn0r08dxq2
E5EM3pCJTrfdRORmuBIiocnxex9xrAw7OzT0gbU+hnrYAYpppeBkgzyaQc/ExMrQt/rAy7i3Bsar
0N5Teemyf2iBKI46yi6Bd8PmnLHZrV+xgnTKpdTwxwRsVw7ihJLyOMYRzzc6qCXYV/OzlJMEAze/
SvYhIrE+vJXtf6a9+XT2c/HnG2XIhu53oCZPVMKeMghhfb0o/Lm0w+LpACNtd0hKX4m8nQ7izY0I
qMBu1NbsCOAi4CJ2iaJuuQGF2CVGkz+lErsnOAQZs2mOH8EU1Ocn7WeGk4Jvl8eSDHLlda4lGGoC
I3mp6FmLXxVLzAUix+W24ebL4X/jibypdB5D4zItPKRovO2JpRN2XG7wdxmNcAl4fqi5irvU+d6i
w3vQN08mZKhwSyQrQyeMTV5MpBZ9ghhmZSwD3YbLjZqMr6nuL1YPhkMW4WZcGWG47JCpO720Iaa/
9l9uGYTsaKMEOOSaMUO0e8n6e2W9S/jOmLegEL8lWXeJelEig5W+tF6u8Kx15/h/Kqu7swdheUix
4MgFgI1x5yPq6Huq+VgHPiVgqKPttin/2mrDWJGVVm2dPzWfqhsNN1csS4WtxCTi4evCAeyovf1s
nueY0aOLiB5sGjdRCsgklU8nn9WU9kN1e5kVCvvHjRyfM8DDHDC/yxGPVYx7eOHmW7RgAxqfs5Io
Fl1MlySZ2ypFF21S+NZnqNWE4gTKeZzzBlQeELDepP4U8/P6pUdRBMdN2ukL+H14amj1TYFnHgNB
ruUSAK9g3xkzk0Mw1rgPbrVJiYkwppGN8xRh/TYeMXwwbBsugFTZGQnNGpa+52Cl1zE2uhE2UDGb
QZnX8tJIdS0hpa86oUiMAzr65GwVni1TGvwsfelu0wm71wyDQyRKCzLx6AR1fLoIX2j8ujQKbo7m
3Y0s5f8JrGEymSQTNJUzAVY6ux7BNEWwWEsPxnFXVOCKgQwSDjHeEoqHL5PzffZhPjBuvzn36dKN
ochuBrz2eXwKU9X0z04c+KeVj0PUCDwxpG8qiLBw7mU0XWNGaKMJ2CQiZ7xualUSAbhkL5F0XzBk
RxT9JWluI2jvcSp+CVJn2bRhVmMqxUQVTvFqk9lU6uU7CzIb7UdAThAqVGnstl4IhWIExEd0eOAy
t0SFhtsYV6HIcny23T7glb/2THZsa1fvYooIdtip83ZKdoWR398tXAZiBikXIeoJHVfxpyYsog2x
ssMKFzstURnDVD6RrScpyJyVc5UEqaJTxoA78/d2iOyMCvh1OP7V6O+aofuLhApvaEC1tnQRGOD8
KG/M+ZCKWTnN3m/KFRr6exdc9gVG7091cL/SIiBs4VQ6BO/F3t8bb4WadbQyYOmpqNb2JFyrpF5H
OhU37geIbVOVnZcxNAAzg5Fwgu8S00wDrjLnBuo3TbhuMHBNU9fh6gzF9zfDnmR/T8Bwqgvltgzd
VwV/oc1wx+xcpg92UWQ9fxwsp93suto+Azap79Eknkc+NN9aHtGSfpJC8dgdat4TjbEsC0zaiAZ0
tzXAbxttp9dWbhbEZitSEF3DtbYzEjGdaPIoADXpWikemfcn6BQkPfKbtGlGaqAYYRpxc/Nzfdsg
d6M1/DeZ2dHamElPv5ELk+Wwtp1aJa3P4/mc2uzlqfz+rWnVKwD+3ntdfh2gb1qBaVaVsTPwiYU0
D9/vpeV5s7/4kGJrUZU4YQ+cKugNgdKdszIv6RdrAyNzvE/vNlU7pZq1gMFwh9E32smh+gmQmR8W
N5xXktaW18ufNQsoKs4aoLgldYhXeB+/sUc8EcCc3h8aGFC6Qa1rpXMklrxekw8hEFSxtB5H+xVy
WrNzBmwrGHlGo3QrQEGqnR1Z+PXJLqo9VKt14s6lWnWABhyMosQhh/EyqV9fVZGZ9PtiychHULt1
/zLmDNOtJrpQgAtj0Vv21r73P5AhwJ3/zD7HETIJzCyzoejOAi7KfsS9YoQi9YhWAMegJs27G6Yo
XVzTPYVLAJtbWQJ2TRGELgbezDZu2zk9o3kQSQoM0KpX+EfLRrc8LXbFBt7Ts5QmuVPr0ZcF88MZ
ycoseI4yzpzaxwxpDJ+CvWvvdb7Ps5LJ42eoCfhq7SUx9BLZGyVMD8pNtTVlFin/kba0SbI460DE
HX4htY2MWmIZwQO9EtQBWcY/gz1lSg7AZbyD/9atKUTfJPZDkoUuOysRmf/9Zetgc51G/6x+h5cS
tBwFmOdeU8QWRi9Cv7cVNdiM9rpLJBurLrmHXyXfKtR1r5yHdmNzppevEX8poG2otUfjGR7GFL1H
DUNcOHBuDK5ukWBUVz1rH7bI87NHE8DLR17wd+Oh68q9mAeYNHuWmBNyO3OJEl24UH76O9KD2/NR
HWhoCDmQ4JyaDGCti8NxayYes1vF3+yV3lfHhFQzfw0BKxdS7TEanMdG3b42lZPtdlXxY5O/+0wQ
mASjM+eBaF0G18+n+rg9z2VWVc/UUuZbu3xTOeFMsdtNlDUFa0roRZpqG4AuqkHDhVbZ7Gybq5cS
h2xgelyotH/MTz8D5lUeSHkZOQ/K4f2t28R2E20gnUUJrfeurQvqaU37fBRqlV9aIm7dIuwrOePz
W52eAbJpadxS3njC8DCAkWSUu/E6+aQSyT/xYbJAheDFLKmAqQUHJOXN1bP7dPLldcFNxQOSJw8M
/G088TwPuv3T/ixg5OnSro7DBMWve16U08s040C9NrKfW/inRpnSp0xGwefMmigI960kWypSBwhs
NzdFsZAyjCGrCUYNB0Qo6dAJrDNPM56Q+GQGquPaplhefXRtfULRxJHwgjFCinVz1Xh3WpEXcULh
fTIOqPbtlxiHBGpZh/oz0ZzPjMj4kM7aLfHCYb8jV2x7v1G7ZB4jVE93ZzLPN2U//+kW92j+nGa9
Z+sUvW2yxPsmmVaiK8kyPMlnd47E9G2CkVyzFhCYHKRt5xufIPYOO5omT/MbrNtxIj0VUSul4xp0
fS4ggAKAQDOjhcIV/90ucPur2Ldeb0NaOe0KxykznrPAQVudPIIc38eNtiLU4MFfqegkK8zbD/gC
Ib/EEAEdt3HjMcK4MY0oZ62233mTkmq6M1DuVQ0MLvjntgjLJ1d8anB7dcyD4t3BTBTbu2ZoO00k
WhgHvGw10ZPVrFIgrJm+2F9lEHOIJzOyaDduO36cmOXEWjwq4YsbCxN8ttNgmJyXkXN8JUlLLkip
aWxLO1npDTZhsAiOrBiO/3rPUo47vTSOXC7WbjOHYUcrpxBAHRPCBftIn3JOafD4F7hI1peVzQsG
enqRW2zfpy5qS0xnKIdFEi7av6bmP6q1gBZNxC7YTBSYZxJzzonISE+86LPnLuSotMqtMX1FYjJP
Ck+tHcc5CWlZFIB8rCFXJbufi0B5D3bxMmEanzk88wuUu7lzGcwVThCe0hbrmvsomYKlUBGC7GIx
KT7Cj5J3UlY7m0rcZNy5mfPD5g5cqq4T43h9ACfoHxxnAfoOnxFp2S/DWOz7k/tY4JY+6ybrmj7y
jm7V+UnXdLFQUn+33pP0L4dfziV5u3XD753JHo1S3zkvFQdKKCLxeQVnAmOcV3PEXCKDollfYjvS
+1w1AInk19OBkcvgmHZ+97q8nWW80T8i72CILcPGuFd9Lpo3/lkasxBrp4rv7tNp2NklFCiXluFA
UaO6nQGrf95bA7AszMSZGQeDhSVewdULsM56ca7nahOZ4nCXb5ndHwvedithnzV1suRSIzPoXZyu
SByTItESD7Af2MZPMWMT6ccUWXaT8wxe5g2DdBqrmHX/0APxMte4saJWW/BD4lyXfAWuHD9PZwKJ
R3BAV5DtnkkpO9e7vpY+z5fjhh7uvUkH85QnKiirP1B3yhEPbUGjGBVLXiioFmhrtYJd1slt2hcq
itAFTXzgatxmN04vmYSFhe1reGzkfebRhL6ux+kP9gbLgQoz0uZsuC/5ytg+HA78/4XSWrupCN09
WP+kIilRzJYhh847GzUDadz4Rg8WuR+yOU0gWW2D/+sfloyFdKrjPCei065V3LscO6BT02tThyDi
XDtXygQAbWmIgZcwMnexKCCrdeZmiV0WbJJMBlCzHnpr6qlAJpDN9GQo+mThCiCKrA5hH3At0wF6
ToyxtLV4kE1m6J1b2BRIbREdJabkatk802qGGirk6lxI5F8PkYdVghslYQBRx5+mxerjkG2sUGhF
QgY7G+7QFWU8eFmoGN/++Ry4dEXcT//9FR33v3datLKkVeaiFs7fx08pe/fk/TGS5FSip2MI+sO5
hEdgKeYczq5uV1aa10Td8XEbMzGMQiDTnECLh8zCpAG63Gwr4o7sbArENt1Sg6iY1JP6UNxo6XkG
Hm+H/TVsJneF58njYdVowEOPRLNHM+FKqjtT2pQzDXuPl5H9ChNTg9NccBTUWurcuMAl8T2yArJX
TTcJbC53RgtOoMOfe3pZMgEfpQXqGfs837QS9OfutzSnABccNV+vhQ1rqzg6vEJ+zFpUYzLc9Adp
kdak8g+ne5SwPmqoDU3pTVx72VZkE7MAc2PwJ2+/bOq2Iovp3Z02i/89czCEaaHcpbEItAQkfeyq
d3P4y+neDIUQIKqTkHZYvHyl8Enl2rDx6ZKG/XfIlcOS4rqplX8ssA2C7sxu0IWLh7E56ShEx7xT
IYgKVgbSPb0Xh10F8Jw0cuG/E7Np/MQptrAy3zgT1oyTeY4tK3cjaBv6/nce31Ec4PKrjkNmRo6I
c1RWiVzG/OMjmxXy8rqgEusOkYayLSOtCmHj/7B9Z346Quez0JtBYAXQxGMVKBHE4FnN8U30L7dM
HaSr8ZMgqNC9WfOwfNeC9dGJsluPhDZVPl4L5IUmEA3ImiRp6Fx4CC9vvAWN6p6g9OrUKYiUt/++
9brLkM/VcJFkREtEVCYeyXEOtMiysG0yor9+Wgju55xC9lFEtIuAI0Qd1FjnMt7G4uDfAm1p5PYl
gAiV2cLOzaRJTAKCk9ObZMqSxCIZ3tCDPGmYrxubQtQ5u4d/nzJUnIrmhV8yawG7ochwScfaw9cY
fP3Q3Qy+0h/8aldQ7bHqsu6/5924EuKJ89Y5b0RVuKiHqmdHbhUIY9fz/eqYGufH+pBJjdDxh2aU
G5Hxk86TIGOhFNbXqEH7CWTOPDNNlPU/S2E86iZ1IgAlq/ISFxH0inL/zP9v+6KxrzR2F+WyRabc
3OvtVUzuPzS9LxxT1yIrNsED0HVVqKO75NleBpmTjByvbdiFWCLAYTsnJGfO4ttNutzo/oEuRmOS
C3w9TjpmiHWOqxpP2QYjfbA75/0JMgG8K7ur0OzJ6tBknFw306aHzO8Z9+q+HnaP3slwSo+C1Qo/
fRlrxmLBKKhunCPd6K1/1kJFL2nDObShmpDDY8xnlPvhvNdO2tFt7mhILRecei9oSnQugzCDOvR7
ifskT3YqeUmNlBC4NuarvhfrRVDvdo/c2sqI/mK42QDw31zyYIXeF0GiqxInDc7Ay3bnQ2SyMgbX
ZN3ivBL0IFsOk4Qn8NOAZUdUi3fb5V3WoXw3fNAseU5dIe5Q2zjASc7Z6qNEBzNsuaK7HqY7/i6C
GBghCdv4AkQ5+fYp11U8AczAnwQaxWd5yq/djgXIxTTfXHKbioFLCT7GJSn4dP2KPoTTt35hSthr
igSaYlumclpnMiHjcxvpFSNIfJVFUg6t9HmAKHd/j80o8KEZODiQWGS6O+xtov6H1lllQP3OQQUn
Tr5pQeay0ZCU+18WPesriG7ltLfnOnbXtUxgGMwi/m1EJNQIseCx1xwe8jrZ/lv/jrB/zRdyp5bh
eT6tJsvI9onggLnBn5rq+WpMX6zw+xU1N+pz3Vmse+YpEiDVYpeLEG36RLELb0QhOwoCH+pYrgi8
MiXpf8AjyfAYFZC0yxgFiWK59pbrrrENCVVrisSLQkuYaWwwfTHvZxOWyL7tQBIbVadRdtwQuFxN
kgB+Mj/UP3ypZJK/BJ3PVkrsDTpkDco/iA+cM6xHLXDYo3sR2rFLUmrDpma2Ag/WGtnt6bNlDfcJ
DfyoGpD/u2HsOws8nQVMMtXROZG4LjvLdHGNZ0TiTcLPqSIF5G8/Z5HMsRCBLDHCPco/qlYZNe55
a5l5KuSoKnaqvUTNZHzoOn6/j+WW5GFSwctnVON/3p1HgKleUgHMszKEBEN0EYGLuA3qPLVvgpuX
21PaefG4k7ip7B4ubb19fPw/cISTueBeOIggF6wEf7qYxbx6up/S1HuwCIZ6NmGjAySZNkUPaFIf
y1sYjnWXNYBU0e0SFWxAjGntuz8VFSGZFHi0WyiJeiNRDQCOjSt6TbNrE+zRG5P3Yiy+FLunSmDg
kVSzgz0gOhl3wdtTPMlPxqDvBrFl0uAEEhFMqQjZKIWJiu+ZFtg+hrcVSS5yAosA058MA7jz89TX
fStgnmTapdyrT7zs/dXBK39ireNAFpqmmFj2eAL8VcfJzvW6+lkap54sxYN1TlR3bd2KOyx5gpcb
LJFjc5H0T6hiDoGVxXtuEiu5BIK7h5yq0xKEASpNnzlJ9EgXXznatB4O5g08UO9FU28tLhXuv1bY
CWGl6KPa993wHah9wmoARwHiYR8fInvA8on95V6LY7OiACHFtBVQZQwbsfryNltOryhFAM+vimUi
IC0qjMznNK19rHwXnZmxC7hNeS7YI8Lcrp0gAX+ag+VKKjLRfIM/UiuaKz/sKBUWFxz5MIk8KbJN
T21qCtkrtOKWDZ2A8TTwQ8qPZ63XDfchy+0a+Q/azMLCuSJbgZ5ZOZlQl9t+4nGCHU+MaDhDkMHj
mwqhQTqhYCWCN5ELms3jNiKDj6jEaJtQnW+I7y0nRYysUbInE7EGXJv7wnFvl5mYrC7vTCSmVvyX
aBxfJ5pg08Ld8Qm21+s8Bha/wS+EM4a4q59KbMbrs0zerKZWqxMH0hh0UldDkgL06G6tHQHasg4m
ZW1Pj1AVZp0fNaCnZud28bQiwSD6kW4IXINcoQTkHNuBCJRD72VbpTkLeDiULMurm65WgXwI+mnX
PGu3NNwgoF802gR0rgyO4ZQAGnbgO4rF1oV1z936y3TtzK44pb/mpVrc4AOSk/vSPXGvgNNjcwe/
lQEDlFRZtUo6wH4XgG38ko2EBiNwXaVJhKnY0UjkvSEQSt7cxaxk67D9SovOKOafgaWKg6NoUhmt
U71j4Vk51m6oqt+lYsPIsuLC4bRf1c4k8YrqXL4VtyIcmcorIqrCRv+Dzu3D7e7cuCYD7mcWss/5
Kbc3wM+tcSFQWn/1ycfz4yPJ5TRvHDnpcCCWES3o1q+3yzlct7LHBeKAshj/Udl/3m8rbBnmcYRv
y8e0sWrPDmi4lvfxhLo7a1DNhVRW38PNoBP2qBsCn48cAloSB2tJqtbnTlLt98iBjsTQb5qZ9SCO
M/zR2wE8C7edylDGCIgq3I9PXcDEVKK+CtV83ciUtjEEKo51fxl75g4qGbSj/HqHNvXXwUt3J2YB
RfpxhzmzaFgOqmg0iztQrCtbE10vllGwuW/S1eUVXRzKYDdvQ12ab9DSHeAJ1Oxq+yD5ioWqqf4o
riVz043+iIB6Y3DevCj+t30hg5lCD+xv9H7ULcIBp2s0aEzeO5rk0VPbs4V9T9gSkbbnOy6aIbAj
dkkqFMtUvzoSdJyHUtzjdu8DUxtFJLeglE7mKJmTzog0ovnImIPwgEZmFfsbL78TAMd/p9zV8VpE
suDUm4rUZzPpAekNmmQKGCNF3qVRYxwaQb6yMc+JutiznrmCeQ2K8b9+yuLo7S1EQdXbA0vtCkYn
XzasErGU4OVMAs0Js/l8k6dJb2KX2YPjnGC7J0x1svc50xupL7/JXxlH9ycBkhVptmlgn8hVwvhU
L/+32loDXhFqmDzqKgnIcl8uoQH/KLBv84x3KUgKY5+cL/mt/m+02EbpxKRcSY8+16z9wKerEJEO
iMotjVf7qFmgPZ+nd/l5dikJOxDHJ2wI+1voof4/1937a3f3qbII8IEENchSq1ktpCn/oUXJvZFO
U5/QW9vOiw5DbJtV6Z9fkmYmHQ9aBDHpa0uVjhnWyAbpZBEzi5c0cp9i1CvcDEpV9sHLWGzte56l
NHef3RrxlQhIyup30wF3C6fABqVWx2nDTiuMKG6cPrvT1BlteTvVYNK5fjVPpJyJV+n0b6yjQ6O3
ycqroxlKOq6mZHuN8SLxYh3ZHy/KYIhK0XHrdDdXehiW7+ZsFt/cwrzkxCbiuEv/uNVfkr1OWWSr
sgOe1Z/te54glOtOjwLcHgtW6iQimrkg+Yv8KrxrOnYo6ZjGN6mU0M4UfT+g3fK3JpdlWd1bMX+D
4aU9eHsHYETmmd0XoXtydru1UIE7iS7Y0uElxY7Kf1JlRfIJkpyLVth7bjCFjbj3bTyc4RgNYm7E
+WMKyAby0doY5j2pBVax7nPTmWhcWy0Mv0kPO6EeU7uhA4XPy3mjTBbu6pAl4UbGhXeo4upv3w+K
rE95OvyvIyG8vJY7ANdhmNJMHUYEpa+0wKRe7UWB8e5rAuqgAQA7u+tEBetxzhklAV8dBUUrK2Oh
hQTZni7Do7HkRRcRR86+Gr5m19EHT+pKWVFQ9+bUuIyMzy64fSubJ8coS/0+cNg9EgGxfvHHFJhs
Ooj1A/yuwuabNt6rN9zbK9VBDm3juSQHnXxFj3b1L3THRveX0V5GprthGJV5AdFmYBjJ2hkD2Zto
RILT6Sqv+E73fZ3OdGXSiAhSX6wLG7x13Wd92GMF/TlYtVjPva1LKZZ0yyZh0Ekxw8pCF2LIIxH2
jtPL2C00lAVBoZdwGIvsVOPoubP143iR36oAjcTV5Jsiia2Trzh5Z3rq5tha10U+ADZx+xJQCiyo
b4N9vB+SiKtwcSz4rrwH/sIXInOJQCEvcvYXT9Im3q9PnqBRIdJsEL9JO6WahOmjTKoYUU+FfROp
qSA0Ok6q0nhuywPjDv17iBzJEufAPg9cT+AMiKwMHj28XE2ZtlzlDGGMVUUwVY/D9alOab/9SVil
5WodZVoamlOytpbnsxtIE4/MY8DzthaZSAxtQz9mUFCgGiZzd/nkKZU9D2nWw467EgJ07042vj8g
F0PT/w8frrMF6VGwYVfvqwU3GxMKIrOggaxfSy1KkNlrVGRqQuSUKzzTrR58oOhB7itTqePM5LTo
iecfitlmRjSMxVOI+rzwBEzadRjrPQSdSqE2KDrlx5WxKDKpDmUVZSylMlCUDJlzBRDetP9PiRfF
CPq7+2sftmIotC7OXLd9DT1F679VdfWbf9DN8SSULdYVKc6/lGIEKXqb/N7PveXS30zSigaRo1TY
fcK4sRbInwShZMs82rphdJlQFPFKrc9cE2Rd0eWInw2YIw8nR+BRK110z1MXlqvcczdyg87muGh6
SvJ/BpaqFs/OWk3rTPwO34qbtkxljDQeRuy0pF0O22WWkDzBbyC5CrEeFbO7D5zuoPkzWPa6UwYV
0WovCNag8gFHVf3DS6Enl8wYpYWb0H1emje8ziKSybSiQbMsMYcLxgChTb3W24rbgOtAiRrOtRvX
fQseGY+aZuZe/M5nhINXdEwBpdLMeoB6c8owG+FqnAVAi+8EVu/XW1T/PVqNtIJ+LnkPk3xRbg82
XzhYtIc2DgcOR1YbMze1GuQeTZ7i0gEo/xZhJVJSqoT0m2/HpdsA6/rs60pagR79FlII21CwSRbJ
arcsWn5Th2CCk7ZFRIwQpyuXEfbTpFN6ZrFyFGeWTSRlRwBruCxbcjkxsE0zw5lRPHfFKo+1Ha95
ezdX8el3LgmobzIykaazqEhCfmNOtR3fsxg+WSEbukLRrsyJoggiiMnPCttjHgpS7YlBGd2C0CJm
bIIGUwRbgq3525BSsXyYo5cDW6s33YxB/41obu7MTVomwZoiOJf1GNPppUQCmDfo2wu+qd8an3d7
9DN/tL/8KRPNWo9AizNLG1VJCiuPQMK16yT0P0OzLOBVd8rCP87xImkOSurbgFlmCZ4suv4W/yWr
UOfKPA/EYdF0+5sU8Q2QFB0QUcqGq/pZ+hGUs/uM1HQ+WK/fWLF5FQUpKKfDid3Diq6LyoDjHAF8
hpoRwllpzrc5HRiXj0HLeJgHOCgZo7sHtQJfL8dBtg/Y2EMwAJAaqOfRRec5SLGnRrCP0SiI+6I9
y0ft+sjR0XK0UFS/MH017B+JYf9wkePgfR0MZvBN0jUl66MPVUVTaALphVyH7Sx1lRMWWoAeN1tO
/NBQOEVXq9oSgjOMjFACLujMA6B8BLAbvShL7ry3H+/Feau/2uFmTkmPqiVsaWntLraHBNzIYzcN
3UR8BwHEwTdNdMU+X410+cgRTY4IkZ954+zh1XWOGV2wYD31DG+/cw80hhoJeWryu811rKRbFmq8
oBCXsB1wx0T+OMnJf1OXcz/tW2uaXcrKa+SB5Db8W0XfwwgfONXjHFwMjaOtuBaxPbWwHsiPd+sz
4kl3ePG7Y6agw/v7UjvJb8az6kkyG53kAc36HW3yG692ee3J8rtIIFrsgSWYEApFhuGzWVXGeATC
5sWfsvJ4n6LH8oyQ9opZ0TUPSmDVmd2oFCt8BigapYcyPYbeBXqWCuMD4V43wh+BSOY+/HGccLQB
BBXARjuJk0MiBlNux9Jzl08ojyA+ePVJYS0tFnN36XKUnCxQonQJIead9qotR5xUY0FSHFeYbakr
3fGNcn/GU5mTek6cJiaKipFnDER3IxClgDC50sjCi4zli8Ggp1hobMZkexJcYeBOx140gSoEwCFA
qNonVJ+eJ4VhNHU8H6kYUI0ISmjFmmRDHwNYFekqZssXevgKI1IfoDJmjrUaGKfENBmmT8/vDsdg
5z3a020l7lInufU3JTBbO96qCnXXpqEkfWmLIfH5Mi/J9xh4L/UlnOlR2BUNFrWXtZ9rGiqcGItD
B/RVOuHHq9v+gnrf4HmQB3EofcPIas2mKdsgqfxMwZuwTEBTt1evZe+dNk4ZMApFW4M3xXrvVUdK
ozpH8GQD+tqVeo2YqeEtXZC49IpKUxqDRzSI733tSA5duAPXB42H8gefa+lNO12j2JN8hqsxYI3D
yAkDaYLrsDHvMAKfj+4oTtv2RhIHtsJPyMoUJO6h8znyoTeu20QUBJq7Z9IrAR8BL38ekVVHS/4J
l2Xkh/UdfQ77u/g/c9W1iC1Uz2xiWdw4fT5B8UzcNP/V4EiGrxNNK9xG2iiieorAe/rb8NQuj3GQ
bnUmiPHSI0+Lpr7xkZlvkiylkcnJidWO9dg1jLxLEbooFLQa6qkdi1UBHkn574ox4GGDWS9EUXPS
AVCIhiAx4NCtXYW7S4hqO0vI0U4wz/geQOLVfquyn2TCzT5FXgTc7DlvUsIOfV3hGpdRuTOxIMSM
AgvJsYHplMShxUZOeSc9psklXs5aqjfnl0ur0cn0Mei9Yhtkuun912FMUnoKL2kI8IsKj3yjznrq
U2KNjW7FbPonsTyy1DhzJ7paOXPFuTTiLK0oY7vIJAHOGt2og57o7izhEOP/peKs3hGHkDoYj7tt
4LPhKc4iy+vGn06ZIgVlltDW7uZsVjWbEWM+vnpagCwiayHD4u2OyJPv51y9ZofVWsBTBIEvV/a0
FFgB5akKseX14EBYIeSPuFrNOnA8UMRbrVEppJqKpo/7JUFL6YGb39jFH3lvmERL3YUPlUXoOGaG
M2wBgLgVML+WF8VLqoOr7hu7bBwnEVme69J1H0gPXasoYQxadUFZEOGFGo1zGK+s5ir+nZf5/sOv
rtAz69oLx62bcJM+ecgYSDHBwT1AuRvfZ+IxCQJVCITcFXv1zcZp6lGc2biv5udhXHu4N27W5vdX
QrkdZzlwlK+K74ffThuuz2+tOxMYg3l5buhvWP1/rA9pavwSFatpVjvWaLY4UpLBInPLuHQBxYv5
2Yh6UWpjLvz9x8aeUEN1R8vMklKvq7eAbf6wPPp6DM5L1VmcFFi12f39q1n7FGQoEJFLsGGJr2mx
oCT/54Ihh/iwnbvPyCPqEp186iYymdUCQgPnu+Po2e9m+CCVK7ASsEyD0GX4BeerP2l7qW6EXqli
cUMK1vmlh2yaIWUuuAYD1n+7NugxaX63rqgh7cwPOf2WSwziaNW3jDkzlzywll4znK/q88+iEh/6
UECISQU6InvYw0IgrfiX5SwweFIfxbAGhSYmPl/i5rzW2cOj1+Mq1GDzF5h/4JZvs5oWcpZemPr7
XJDk2IY/+FW33/3tRJ6bCM0K6I+XcN+MoiH2CeIpJCzSvEhVYfkhUnrc65kxSj8KPdLOHPyJlqVr
WwYnRTuojE0a2PwgRfSi6TDNoKojzUv1n/no1e4JLUCtxeriCmvvmsZu6u4gxj9jNiR2dJIEq/oL
uZ1rM2AqMoYTSWjkHRCKXb578hGD7nJDXa8octUmCKoTDPxoluNPJtiQsZB4D0XmsmTuhVAaE64d
/g+wQd2c+AviHxJz6zxLUjkcCxMd88Fd0YXVZ5LgXxLxGynwp+xJzNkmuqF9kGieSzXAtYipf0II
S58NXa3zBjbQS7rVQNm6X0O2SuzWl2I+z8VZCbJf1OD83C60qE2spnaEbq32CrzybYxo14RaGNXZ
0otymJLOOIFfzFLmMV/VfAohrEtc6Eg855eRpPHMM4lhVps0RzAl1fdWhqb1oSZaINQGIbA6i2bY
CVzbocMrpowelF1cN2VEO2M08keYBDozmaknlK8I5xzvsTmzhvwYCZTgi5Jp49RsnWvFevISb7lB
pBovVFAqx8U+oBDyvTk4dTcJ2Y0bdO7Uy8izpbnyP9DV202dxaqZg9bhUteYnrDPompYb78n3bGI
6p0rShwuLcimMvCqdk5eNrm+sLlrWFsK+NbZbrhDVjq3hBtf/B6AHbYfDuVr3rSFJ6Aytt9UFZyM
Ovm7eDZGsWpVikQeZjx1Sro3b493hnGtIid8md0+SwhONNu5wQEyuRZcagvs6CFSoOaDeuLbcj7y
VVYlU9VsLxdJwOec+7taGC08gikzB3Ci+UKRU+zhuwNI3QGHwfJlMxdChshHww5gJKEa0AkbPbX0
VXKSzxcaD8hTevL/FnQw0qRC/R1BVc+gBxfbeEOJ0YH7a+q5AuMyqpxWpLsb9TuKsPXisjFNZRrx
IS6GF2SZ/UyfCc6iEqyico1rqaczj6UgmYCnutrGT91MJJz7lJBbVBvkJvAUyJfpDxdT8kKEDMeh
ALuzN1vgidooHsPGTrdvB4WSl9PDBMPyawB+N6pRccsUrXcMwa39g1NQLwzSATt4gTKqzAC+oiqK
vAM6UAWZjpdfSp2a9JzvYwrCsKPxyCjLE4ZxyOfEx+NILWijGZqfiPCgZeHBzvlXakPS/eMzW3No
Q2bqZafbn2bl3TLxN+5slsb1IByWfr1jpsXyTGg+MIE/YGxnNuyLFS/jicMd+cxEm1xuRBgL3Wn/
6ZYYP+59O+uDZjnY17w9ps2blOFIARMJ5GPaTwNXXDVNknaHvKUpcHPfxxqr/flka1HLSXKMeQ2h
QJCIUHnfov9vIJLBO2BQbI0YPy2sl1d6f5yYMPc0vHo8U+PSt3bsNJlafP3VzHXUssLwXehradVC
w2OhWt9WaE0Rt2evQOSmwQ+kIXRrVqIxui9JMFVDwHWWXaLhd1VWJyAXDTo8y0H6XT+ufPxYKZ+p
lc4Summ4a38U+jNIu9lEBHolmACUsgnuO1nQ3lKS49lRcVhbHw23bKpa2/O/xhbHQ16zlGq7mu07
TdnrcnkoRpUvrOh0Ld0v5dda5NnMZf9NJ/ChbWLhJfkl81eGWTN9E8DQMJ9Ma8No3KfTgTOEGdlV
s/JaIrU+GG8qALR5k2Kvby8GgUzvg+8QITLk1ZlizubIAyktR0RaztrchkRZ5b/c7H1qkiPKwqCb
p79i9rqLvya3Mici9bOsVkH2vAx+je4MADEnM9kl2LPGfdEzMs9Tx6MGsUUkhNubYTm4L7Jz3Uyc
q8wo9jXVqFRvJ2ynvJSLt9giEVhllVvFx+8jTQRJffKYs9oahRhPbNi7pX7UP2Zesed0MHQg9Fnt
4PNRvOMvFi6BgAmP8EUecZBLCzcVbdAeAbJAeCyzbSHqKjd38JGn+fuUcFtdVul8UjO3ABCnzk4b
kfawQTVJErTeGoHFj6BWJfopW64e6uXUk6s8IOSxBYln3IOLWQ1FDO4Rpd59WFnGFaoHACOKGTu2
3k/0mxSBzNlOE1NSjenCwGjJnDDq4pbfXDmabxAe8Vv+fKVLS+DyGI8K89N+mQ9L5Lna5YgLu9g1
UKd4JlHDft2oyBNvJrLY/1ydMWlUf0LrVttcz+75R8HuzrvdzE96WcNbVRrDngwQMq+KNNVIX4re
VmVvrPv7YrP2CISmpPrOsBqNhG0FMCRU0Yo9DxzD4zFNzf0PJznkJdjBj68o9XDZY6g0DMjgWIvY
8XJQ+MhEcKAlQjM++h7Klv4pG3wf+A1CxhLqADq11GCOnEpbG3ktSFjqmt5swytO699m58w8wegC
QEaZ2jp6KiBMfuXjhrpgACnLY0ZLDpRYhH9pz1OR+QAck2ovRut7jGhhdK4qumpBdfHfBfLpftpA
lPQlvQGxSBAZBCaxdPu6aMjS/16nIZoTwGeYiZxZydp5KLaKgOfVotmNO3h7vtRZEnFKrfzNcUB6
DarytQm8x8zKVQ/rGSJThJgc3SlRAcaAMmAaDPQQ81GkTK53MQkFcKrmNJm9YBtI07TNficOr90C
eHBHObVmtUSPFWluy81r310tZ1424cQrkIjEGTbGhdeI84TLgYMc6oIyxGsuWhEUErmewJnDnX/V
HF/UhagRRrLonS2tXOBkxmyMewy4X5OVZbGF4hDHX6XW9IksI9Hn5O0+WxT8YaivyPVCQfVy1Awx
jn/M9ZpAWI4cPoJpiMTxnyZnfvGTwRobUHl5e00igwAqb5aBi1i/ro6b09lSF7+9k5dBDwZW2nYx
rA86kDKO6YfDOP75IQsUpJquvcCFLhfai8JWTzBGIw75XKaepFPW6XhmALzwTamjeK4s2IfwxHND
Pg+gS8JaspqK3rtjjfUZ+eQJBJQF7eTS0VKEoz9WaEF4r62DtsT2/9Jk/veiCIt3bjEsUQ7psuGW
sb488uRckhHQ3TxDjrIJ7JdKMxh8XYdyhLPiuP7SnwBe7oFFc1AP0J8Qw8XzAPpDDKyyyyXx6pO3
ig/mHMUpopx1BMKHaVSzytEoCBM2fo85EvJA3irXFC5rPTF8kB1rITYgKGGFrVrUjVXddRdv9y2l
tZ1u7sa76aULTZk1toBTJLlUD0uQ0TBIYyy+PnTmYbvW4qaK4Dg6yQrgglByy4HTNvV/bqKpjIpt
ICdoztUBhS5UVeHsWptUNQ0Dn1tmLGFCv8w5J5e2VGlYTYIMgMYZ3ASM3igwoEqESGjMGjwDcHPs
QhBr1+/5ICihVBFFOxwRIcXKf7ynr+F8ocYKiXsRAdJ8iLUtOzf/OwpzxESq4FS2oFiY6Ec3ghw6
BATcHZGSRyhYUd5Xc5aDoTmTvvvMQsbu4EGpiZL1080ZeZCb6OkVHsuISiZKDK9UO+9Y6Nxqgf2j
OfJTGBUbAiKgfwQassf0OYxfazMN5/9u/a1BngQ6RiBIwZJbcBRSZPBhFGmkMrVn8dHmunziv846
ZWQbl2Kc4O506LbRBhHnc8ElKqPgLFvXVm+xWegCNqtDln/x7e6qfS63RJdQWJWY9Q94mPp1Mi49
n6owz7jY9Gl1ED3K6MfyqfttfpCT5kDt/z1CBCN0cf6/8j1JaN4e0xHsJGAm58G9K1tJwIPYJ4+3
uBVFtqKLKR7/WHG8RrkYw61rK9a97hjZ7zkPNXy/TlxywfaXb0ICZA26vQUKZHxA6b5q6XXUhCYS
FallEfieQaVq7CgYgXNEdxUprW80niLDff3/P7xQThv+bNpbincikFO/GY0dVeiaeiecsKDDhSNm
b/f8ulkl0uUHUHzTBR5KKMZYxKGgLnmggBoeKblbyFXMP74dIDQ3eWTIvVVJ09xIPAxK6CDJumma
tN0vpMrAanq2hM+9j9v85nVJV73GmEc9n+nZYtRANp0QTPjTdkvXii+N+SOHL/FLOxK6YhAS8Kmr
VGBQqU0Y8dnSQUuCOGF4DLnF9dZ1cuVrSrJdK1KIBY3S+Dv/fe2MG/JLWYDmToYK8DuvnY4e5C6O
+rj4kXGMojEX+p5XSJUUnBX2e06NCYR2FZ5aoU/UkU2IyzLpM3ILAQ9Z5uk2kTWOMtG+w2mFV8b7
nsjG+05rWlieHulCorgAjKHXD/DFkVO5RN1QxtUbZodpmc4L0OjtH2w4RgxjLRdMor4Ks/uMoLSJ
98EhuZoP1oKQhADAHIN+5de8MEWZmUC0PIlxzVB+XFUkyrsO/tCcFjSK77X3UNEWh5xJRQWccu7H
tkTdg85/N8S7+vDd3SIzaDYgFzwUza/34htNKZPPpiDayjaS0MNo6IAJ8j1QUC1EstDxmsYruwn/
dT7cu31hAyae1GgaQlQp5C4MnrFkOPBpxh6kTq6paADopHmyWzrwOQCdoFzFQmBG59g1ixbKRs6W
WcPcwziDVChV0YmmW50EzLwbvKQJNo6v3vi6KCzDc0EVZd+WkhwEaKehpQ4ocZQyDvQBqQOBvfJf
TVs2LTdxRZ/VgByw13cgQJAJOvptGD6i1d/t65FE/nTQg4+SnNiP8hoNE9/+KM708EtpGRTeCF/B
HYZR6hXvagBb5fPurlmDmClftYau1Yz2BPxtSE/J9Y+kNveAx6OBwY2PEr2MJLajNCxML68r/cZY
/YAXGPWzDcRtFGngd4HolW7u+9FzlzebzjZWhlU4Cj3Z7GT7xJ0D3gihaUirEWJDqm6tpbTx8yQ5
hD7eRHBbz8pa/DeFfrwxQN7T8otwULm2S5UAt2vt8vjgnPYqMzYe7hLzPNUH9BTJ0iZ2zQbvXB/N
f070wYS8rZDb+506VLIVHvmyfz1eIp6OmuU+cFo9OdfyQd2AFdv/pLwOQe+ALVoVpRIa2nsx6Jjw
d46jTR/8UQUcPbyrqtZnm8TY8fSj1+Syrk8WaEJ+6c8mGdFz66sc4GwtIi0T0JQsC0U8N6+qhmI1
4Ip9vgxvTonAtA7xeTGaBGAZrY2YI1bBc0vVS+6DMNFGx9nYZHsAsOHsfTVcJING3Uo9uXLFRnLa
MxY3nczHqgBRvea4Y2ODrPsH4JFKB/M8Ubh59hjIPx5BCYbktieYzL918tC+/27eDNK0eKypuMLM
DdGhG+neEgNUo2QEBF6Azg7KB3EoVWB7zQ5kDzmIcxpBSPljkC3dGT8qsF4W2Di6WDkM89a9v105
o6h4Y38Ab5Vyvr7Xh88j0bfOCrASkYGXytEuqeY0uEVW+r2TDAhkXzfbLKRVHGRlUhT7/J6mMwOY
3GPpQCBEN5LSZ4yYTY/wP48lPiMd31m15Jj4pmQEMav4Ul2z98IS/yaQHALOeybQm39Z+x4KqpRx
VWY8Y84mjcQDi2lupe9eCC0Zib4tqWJa2Lz9e3zSW/LODk8KtQuSQLFrLIb6++S65xZdji9Rdb1v
4nYujg7ilYhVex+WScy99O9JI9iZyeVY8ecfCafANvw6/UH3Cgw2FKWjL9y0bJKDKPrhWtECicJe
087kw5LttSWh+jkNHz9yT28SwWA06/EOpdYMa/wjkyQiKEbUHT2uWx/G6SsIm2rsqzZtdZHy1tlt
ZTuBBV/ROI4fkBvn87li9RLqw9O7VFP1pyZYkiydaA4FssscD/tj7wWyjFnebqyCgIf/BMPJjvZD
9drMLuPQnbi5K0ZrKexN6iKD8ZF76qAbHah3bHqwmKhueLNdLaPYxB8epEq6wtlHWj651Mk7pn7s
HKhOCkqll5p9k2JrzqQE5Q/L7aRmqwXKS9lsNKmM3UPnaBYlk8QAa0N6cv6E5IsGDQLTUQqG3a/X
LMnGXkSP2gdI7GU/KWvUG2kF3upvik8PUJDzR00Wx6s9zzwrMeFMg+ghPUhhYqqioXNZNyZHvY0M
6wzJoGX+VtPx5lGN7sn8+47SQSYkC3iuWHaa+UQjJgvtB2Ngi8PrCPo2UtHX4idsHCNTxl5NMXds
YbOPr0d0MTsMqHMb0M/JoHZmq0MDLhTGi8kNqB/cUmgLFiXwAtiLMl8R0YQd44iL0eQAFRoCqmrm
W+rLtefCx/JYWbQW8X74eR91lUVeHbgnVWv/7Zzo19AlJVgPiIijYw9UUVJmsMg3NG5GgLIJ9e6d
dFSLv/ghB80Xxo8zj3SLKyUwDeB1XBvBoXVVxQ7crJXweeGB0JPRJdXH0Ddf5JPGY6n6kLt2pe9O
m6ukrcauQlcB+Wt06dyMlhBw5QjJVkDrrtupa+lhXib4YJubFl0KBXCKZEeC9j5DCHSxDQ+BkuRL
NQXZLeuP6jEdCWKCDxjKBYW+l/AWECAGeK01a1q7kqJo9ydJzebcagGtrAiB7JR7Q3/4Uy70lVAn
nhYxnsXAIluOh0Evt81vpYFE+8QQDKRAM6lG6U+Xhy7o2aE74AL3olexFnrU9Ocpkeee9Nb4rkYy
q1e4RgJhQ/1IF3oPTMrUwTaXB765gPwCrP3aU9tIl2YlJeCJRvCmYKH/U0MUh5ov4VM16oAsl+P2
VhRMwx+/vTbNYqWBsv+YZOvP//4jlu9B0QnK9lj4cVDAtpOa7TpSeFSQdGUoNHTBo1RkKM/PjnNo
b8/Rm8nddhi+seqKRQwRYkTXOrc+AChMVboLBV/QluFlQ47eHoXimC2JAu4nL8tJiAZPy78IL57A
lGeCjRmAsSj+Meyi8c7D1CeUNLD2pgGpHlnJprPtkWUJQeJt+x0UWWgqRCODO9TYHT2/4yev4xs+
yKjLkhceD2UArv3bqBPVqzuBS+gLrirAhA+sJt3/wagC8b1SBwttZG9S1srZT7bNqPQ3FSgrv1am
2rgwQRMVsSOrosNW1GB0eqB/TehvWH5wTXohR0tDLtjrUXE6RAMSGYa7CK9PbhTbtv8q4zB8FsgV
7fyRjIcSfqALk6PRh+b7TFKTcowCzhskOZWx77nV5xKcRmHCRDOM+AN2OeDsowhTbZFmoaRsH1fI
NgRLM7KbxInYdrW13wg9V9/Q5FenzhU74bjC1yym+EcC+8d2CYmbytVm6toJDSvTnONyyUCtfD+d
oqTqj8+Axk7KINakGWwyVF/SY/bNJ6Ssp4ZkErwFtzBxay286pkbAEQ/1sm+ZFd3X2fqnCPasAYH
5cUz1a0X4lf0juy6Kzj+cQFnZ0AbBNzx/m/3uLXv9osh9g7g2uwfhVfQ+dxYS63QBxRkWIFja+Dy
VwRoF1viNiCxCmx3+FN1WmCOOwC9/AjBUkP0GhZEIhVv1iln23tl0J9G61/hGgmdpPYypvLe2emR
7sV7JboORSoJOHRwinXQgCT1nAcebhYzoNiuCL6vmy2O/vNJRRcusPKMSaC/aeomarQnjFn60Oil
ZYNoE0blL4JtOyhoUoYWtB1FKXQfl1PIlVLl2kPFhTXgzbuFQQ+D1TZTBlbStrkp74AysPaQ8H5U
hJS6LmaehrbVpuxfZocqiyhNbj27Cb9v81loVgvpoWB0FLvpX+FIRHVeBLAGwbTIc4UcbBEfxb4V
dnT2S56l/lG56x/LI9X2lQ8EyBvIU9ME8gBCM7SeBWInK2vnej0NBBDfZYx+3nnOuQ+BFbbNOTU8
HIKIlc+JxU2jGIZdpMx7XW1IZOUNk4w3u/WPTgkJFIjB6gjjuy9koEiCYB7TSCW8tAyp3AXoMBJe
ZrxVPjapBnu+CoVwICayrjCD+jL4L7hncqxGhE7pnj319FsuspItkR3h8uQEo2NX14VgR9iwriKj
SzpfJexRX7LVdZquvii9/3ycO3+0pblCQQs9XC2BPaKRE4FT6svhKM9y9NYAPQhca1yhBaoARQ1+
UnUJOh6INIfVByYiA7brYbkJn6Y7iD52hKHdiED8t6HjbI1Pk/YJpZg47YEB4NotX5BXQxu59TYi
rwTgvenLuYkdIuVGc2pBNdeLmqBn1dvkzDlp0rm5VBiCdp5CaVwkWpzIlmk4ynxkd/A0Stgtr6fY
FmWp0FgvYenDXq/xnTg9LaEQSI6c+fSkpXfOKsUdoOMws2wHAsFIh0OiSmCGHJG39Kw+PTwZkabA
kVnwdq9Nv3cajPU7rTGO5t6gMpMkMtpgOj56nOa7WbvMlOl68I7rl2BiqNnbFyuy01F+1hMQ3WnW
u8ggvnRmNls2zsyrEeShy8Kp0PJYuFS9Ac0Z4SYQ1zw/g5oYAZQdC5x2j4rvT/MDiztDd3mw99oD
Bg1qacxjYfA0ZctNlkUO1tSEFodZ7kWQD/QhpmusPlW49nlDHHU8Go+HmE4AOFff+DfnProVqbnL
KPk+SOlK/cspufbujVYZDMxKQwvLc/sIzjWhqU8psh0EgHMLxfNjUcsHbixd/k++BwOiAP4yrNJv
AJJCspmrMHZTukrLnbm9lgnamskHH1jSn10Z5bBVxceyvgrEiXcPlX0uUufyx6ZvcyHgAxY66k9P
rHDipMLRgbfRbToPPpc/daZ4HzCFWM+Drl9w5woMqVTN0ZGc1IBnryxovy9fegnD1mlhMGIaRigg
VsAUaEdrPmQx1VzvcQuRoy2YEQ/JXoMXMa5jkJMB6l5l+i9gQs4GC32HYReXAwdUJ0Tz7Iz//qsj
kiPuGXblSTCZ/TN/tGBWKAfYGsAZXU1iSxn53RJOznm+SGX7tc5WinW+CN2In+ws0K2nePvN9Sta
blXeyS8jXHOfsW3BUhO7AhJpYm/li4dukrxQHic7IdhB0/Mlh3NluCJ1U40lueydVUqcQZRF9+5e
wp2rZySlbQ2Tz2a0c/a0XB+7nnYAsI33WRb5AnLPRCtZ3CUEZTvhWPKjj1ismKwq5PLo1PEgLTBT
xb9TVipdy1kJ/yK4R9/5qULAlqPyytu2r/EwmCaZnqagpL58zBdNozwMczPCtc1dqqnkQMJh3tiJ
zGc7UuG+zbPWXc3rQGZXx78O5ZPyMTSruNjLX5elyrZNU4r1I07T3CPdVYqJhptrGVbFQsz0RAJN
ck0yULzQCHPuTQ/zOR7hCSAwsOnkwUKSzct9IZz9pXMx5/qJlAVTnI7vlDGajCEJX62awW8Fml3v
YlXnsVhYpZLMq+3HHxvpj1KWmOLKkP3H+yGSzxXB6y92PzupU0h1PKljzrmAhEIrENQvKfKv2SAc
7uv/YHLdIXpuP7HlS6GfK7COND2M0vmUAvt1jL30nVxvFFcaI24yM5RaPiQMZ/6H8nf5ztX3aTAN
tfywk0cpxSiiT01UUAPeZ3uJXrdhRlcBZposNeK6BAKjpU5h3fVliiifTPlDwuJvqtBxcIoWd17g
UquJwOesXL2elqK5rjNAJZi7R1TvaBGAmAj6HHGrg3+UkG32pI7eRnXT/Vs0qb0iIMamsuveAhgm
I3YMmmbb9thBb2iT3KD6bDuRai0GeTIZ+KNkyXFliVY8/UQ1IZNigPPBm6uLEFUzjA53zam0Au8I
06xUdK9pn1GffWbRnrZQnvW9GrMI9zWAkVcauRbE7xTpz8ukIe4JWUxNBRs1jh7pA25mnQJ69gsj
RnpFaroOEwDHYcYLIxj3YeKKww5wuVT6GVsg05m/FaQIHNnUg20ufsGS9e2RIW8m7a2EAamHReJg
aONx+svlVvrVqg/C/mW7+DvcrxS4uhYHY1egFw9XwrLzy1mykRlg/MbyGNU1PQvra7tXu8XkBXhf
EfCBLRZRi/IxtfLdSn2Cq4vCaEi/O7gGHP6huXGEb6YZkBOzqLvjNPh7q7b8Q3RI6vPjL6GWoTxw
tbceTVP5BaQtNrfeiTVFfIXoezs3arWs7C91Gzr3eDcmvC7hr0eBsBn4mw4DTGSrUUGbSTnx9HNx
PN0f+2CEYf3pEZDksn/Vw00OSBh/mFL2Q8Dsvef7y8DBeUocz8S+fil/iE0zWgXJZ14gTvgjDiXj
rHv68C+KrjtMv2U3wBYRV7e5TjArphtF5Z6zS1OgvL54fu0A+tLJjQcYaLXuG4+wGVGp0hwuqW8J
p6NVyuqzCFT9qnUPqqdy+ibMkzzyHsc9v/Va0ag/beV2KjR2gPat+fIWfVxWTm1H28kKurdNJG2l
IE9lBzV4hWrcc4mDpph+BmhLCSENt7qEnwMiggERH4fgtgK/XqTf3HW8LvtnQMBLuHvR7CI+4WrA
L9l5m4Tyy1Vk9ALiPYb9pkFMJKKpKXTq1fzVm+UXW/ciD278dIkphHGRm5OV8MZajqGm344MkCPV
loO9FklpNbdTu46uv170VI7DnH78izgTpdFajS+f8/xRr7bT4m0j07CDlfZSjfLo1X9QeaRhipKp
Z2TPMXEBnEh483CcJnmUoG8ZqqnTc4VhlwB9Ska1kKdIwQzJVpqm159BF1fl64zudRvUTbxjXllM
DqLK2u/JO72HtppM5wW0Et5058FeK5Rg5QrBPv19r502EIvCvwCWucdR9uhfG/Cy2DgO+B8/N8et
TGpEENVxkohifkzjuOeN8X91ioMavFZUFntM/XGPeme5tlM+9RQf/qXq+vUFxKL/Ay/AP79Re9DQ
4CMOCtIHD7GT751pS/txNhLS76vipCXi6Ewon5SFqiKWkLTYy7m3t6P3NzLHA/yezyjTABG76jp2
7fQJESEy5Ur8fBjKFSZHgwc1VKikl2Wd6YpWmLArOzdz4PsuF9cL8RIiEs/3F0LEOMcNJjXIxMRi
YmONJHXy9KfrtxzMQlPa2g6AmkDKLDJ8N4E8Jhvf9GcPobtyEuERe7up5QrmJ8jbAZr2DmEf+2EV
DUq3fLG74KGLeIM+B8+XyqktdfjFNTtcx1RbeKxIoDcSI4L7F4QU+MVfk4Xcr9drKPXuU7qYrBIy
7UFCnCvy0f2BL/W0YVikd/P/caClDczK+26UzaVYynv4qr/iAomM5FMNAruGxTadG7nFNeZ/ho68
hR4EqpsJnVAIeW2mED3aoWIs2uZMJnV9wIB9aJd1fuKDosyjgB7DrFmSgiBjf9NipccwMVyA6Ihn
AjyNbYnuMGUBVnFbnR2kglwWDdZUg/gSadGBm/aR9Y1gkcA2FZLjElkCDfw4H+zn0gkx7qyuPvVb
Ll3n645T2258Qwj1ckxIoyFw2PSbNnu0rgzEcSZxxEth4GsCBBZOTao2wbupUobbzaahFR1l+kqZ
hQpMQ1p7CSgmMbP9+7JkSDaMX/5QRiAwDN7SwSMOV4jnnLPbJjj9OJ4tPK1oMa+jInbgq6/kdPpB
Vx3klwJNyC1mAbL3qCt4oWoDxzAZ+3Ot6MF/OM2Hy/eUKPwUKMqUwaxhshkKa2vvJnu3oLKz97V0
6eHL7Dqi2VSODUt4+dSP4VPtXdVONHRNk8kFu8mVaAXul37g1r1PSo15rjNNlwg0231ujhLCOgQl
Y7NfbD+2XQLrcnpKRRXLYN/+BfQByAHI9oMVRtnAMuKVTow1wUfoUQkjKQ7jY3FrOqrh+zA+h5XB
p58MtixgxxU3x2jcJKpR8yQErXpgwfYhhCvj2Iaob6+OSEtAVyaC5yFE+ERjZUk6Txg3TtPXUoDz
u72BRb3BJ4Gv/air3Pom2YdxfscYzPWK2dA2Bq9IASViN2QNH1LUsm5vuAiLtYmegD4NIeHWL1l1
96CgS/g/AUqNxpmimCx61VswJ7dI6ZNvwApsZNoSe5epvWmCGOvnYgT30jC6678DVAAdez/oVzzW
FUqUUOlcdnk5kGNZZZSKu/2dcGjqhvZ4xMRImyuBVRrc8upLAUjf8EJ7V6uo56e+Eihmar21R48/
2oUDL1uVK9PWJlePEGPo5WUQuQWOn7VrtYnQskKbOgI6HVgZkiJv6o0V/jjf8/hVYNKCzZbdr8kF
kc+9cTQHBdcRASWBIYTAewZ41MWHNMpDR7FAehtnvJavokpdir1laZ1aOloIIMgsUz3vKxangT9K
5lF0RPnPS5VroMmr7r9Vm47zWvwO0dQGPsLw6nH8Q7KlCbmek1cw0HZ33Ww869gCh0TsaqLVFtpk
ksIH2dWgWnM17d5DakPMCfbOdGirJRa1i34cHfxz54eLkKVlJCVHfaxjXTgYdw7ncBqozdKaXAeu
5oanRZNcVi+s2wszVZZiLfW+CjK0zSdlLcTCsSthp4eP6LVpOTyFSPMFCrdUw/vZkB1c6rqPj8Rx
1GmEbXcUSGcmK7F762lXRYb15xix9S5OrI3jRO4orwexMFiiyJt/Uf3asDoI1vqrd/r84DOHwpKR
owYKy4BPiuIE54DZHU2qaQMuLUSrtx62O9o9Fl9TH+eTCfWv2q15qCTXsNd1APkNsQGqYA5H22ht
GxdGmCVSRk1dB1vwVe7+0Oofvp1zW9CHxoKmp+IlUl/xGZxCxwkGiKNgRJ8Z/kzPSvsPDAzrZuyo
RDjB8FLeTZpYFXvw5SvWZML0lad02bSjJihnju+LrkGeDksqV0FNe9nL+QMPEj+rKvLsnQNKL0TH
9FhK/wAgMCd5E6jKDjB9HtL7MDjyeEpHtjD+ZYXoSW5fgATJs3/KklhEtAI7rRKhJVGU2pOtgL3o
vqEkvZxm+cLT8Wf/bbx0Uz7o/juFF4elIHgnrC8RX1ri0bih/5U5ZIa9AooUeq7kbPvs6EYre95u
HFA63j6cUAqTYjs/PqCE3TOXL4E+qiCIir7ccYR+BNnOmPfHHpq1T1ikKeJoUrlZaAdijtHq8Mna
R05WhOb/N4e2H/DSAPgorfA5l9xBidR+vE/dveZIpSvNV/2E/8oYzTVpDt9d4UY5scfURgNNX/sL
KwAXqQQsZXsIDwWvefCghN67wOmScp25o3UenKpXTEj6v/3Gea2OevmF4VCe4WEPiXW0MQXH5X6s
IsMB7y7jR9haKjYWmhybP6suH0wwHU7LL00XOhpBjCWnhaZfoLFlaIJqXBL5Y+4d0Jh0mHU/jIFY
jFupkHDBviO/HqKZmSPBioK4TDY3z9L9Gf7qVWNAFxfYrk9GXry5vCpuMsWQEi4JvvWKXLa+qmYr
QHRD0+olHDLYmkpRvYGid8ZgKuYkNI2tlU2dZWiyPClh8IrdJhdUJ7snaDwuGwvFAUUhvqdwpZRg
EFQzmJfAJlA4Ue3gyXS0vva2/Pclo1H8Ye8V1yzquPF4nEirIePMQTghjROTI7EvBVaIM2GS1cY4
yUv4uSZ0WnYE1j9rPKnLBVs/7RxgFhqKz6BCWeEqszP4+tgO8DQ8ZNNh4mFdMLq0E+QvChzqYLzc
g1RtDGa8226RT5GYFMkivAx/2es5JXWV9xz+SbWxc8uOsidDEfBiaKxX0aBDnwno8OlUfoSMF2/W
8AOtBX+mtLwU0c6DIOGb9y3G6mpWk+GknRoRMv6AyTGx/RZ7OByXi/lijYRWiYOmH3qFZyG9aLTt
T//kQ9t6FJZzNbcJHbxAevhar8AP6Kqx1o/qm5dh8HxOK8NYU//RDxldfUHPHT0ll0LlALxZxDnr
hmTAAzKgoBt7b88rfy6kreODK5tCB6fabOx5Lx6irj3GWKxg+mkP2chXBe3yENB2kawLXBdCkCiZ
jclNj1HSo7qj0q+366Ql1eAAidQQiJh5fL/gXZqIMw2UZo5hJ9aMb6oHHrDP4gocJymE7qpQD4A+
P58KaldJYiNnNt6ria0JIOGc+u5TDjVtcQJUppPnfnou3BX+YQwvNJlocaMBPzbrasvRQ9Z/gKLQ
YjSLM07j/Ri5GctDMc/SYRDaU1m/mColZfLXSeNSfqv3fN+xjLmfce356gAwUWOUMEdB6C5J5kH4
ooWrSm69UQMIVcs+0XJJEMakglb+FEPlm3uu+V2o9Lk6kHFloaHw3Xx21pAWfdZbPgqXlHtviK33
6Cq6bpad7pUrDURw+a2xvhIdGQBVbFSgolhU7RxgTuVXAeLJMS5SG6PWdN4xfgHOr+B3XSJPOnlx
Ag+mk54CiBwxeemSyNzB15bYr+tX5nN54C1ffgJK59+RB4EKANPAcUGYRJTmWfRRai35cyALsNdM
vF6W3raCfutSsr8FNvk3UFQpD6dlqE7knGiyuJlSas99Tbwu+gDge1BI3/bgxbOxQhBUzi2HogG9
pUUnL0YX1Ojpx+EzDnt+sBwhwBbcMuOF9wK9Gu3w7AX8W8zLli3bEn0pk4hD04aFBrZ/xirKD3o+
Dd4RsDcfj88+Sw3fxei6WKYrGOwHEXjjj2jSnjujJy9+lpyS0KTWVFM1zxvgsTishUQ85NMweWJt
KKIBGpB4i7IdT9Yw9QQjfzsgdrVGtP4fdsgwgsCpr+n/5Ya4J35DocfjG1t9nhoWLvIs8evixKui
AOSlD8rs5mqQy9J8HWqvuC8K+Jlrv6vPOrKLk6+wK7RLQu8he8a214HzNJZNNSTKt8TakI3Au3G5
+M24QUb3Sx74G34FCr2kx6YpmLaqlaBSvW71yGRJc7LmF1SxHAdrcW9XUIvijsXJerJ+J38Zq5Q8
MULIRbflFBny+4gkVf61+waoRcg3QptWb3u8Q2Jn8rRJW2Ch24QFTHXSk7g1W81RQwTk985HgIkc
ozkmmuizytKUDoD6nGuQxLbsUUsgt5j+0KJ8fVF2uJ7YD5Utz56eT02Clda9JBz3xg3+42oCj26C
EDqVrTNIGnvob8kVB+4U21kSTTABsloTb6E8Sx9ft7jDJO0pk0B263WC1QyJMg4HFu0MZ/0j/F7f
f27mnxzF3jObPCd1T3z56uk/MoUw9ZIqLwjDEmUe1aNj0c6o8wv9wXlTr9nIsoiEwvjKy36lZK0z
g5R6DgHwxth0+6q3Tk+R0dRMUkC5niaXJY9QWVUciaU4Gfl7X1savO5r/zMB91oA5DxENjluSliN
JUgq49Bpem9kULVYsPYgbijZf0gO4n+JGzz1R2R+CyTULidrCNhMwY0V8VuwAI+/3GjWT+bo4/de
bygQihuHzT6C+ruJHIdnk+yMgNHxsMrvoUq9KnvS/KfwDYz9ViZgihXojc4g+QzslJJgLWT1B14a
cWZJ0zNkzW6PkJ0W/yt1ZjLj6xtWHRZPLrpUyQhjk/b24LP55+PhRvLnup/OaX7ueRopUJ1PA1h4
NTaGE1Z38JHuBUtrkUgyVCmc8aHRddgP6TNTWEfAJfwtEl1geKUO5Uml5G88NW0Fv4KasWWnmtS8
isr/tgZq/A0LUff2ETIEUJ7moddHOA6BjC9jS9j3gbHx8UEowuKcXGebT0mAVOektkFGhqppZssO
yzbGeV07OhbTzqVHCJCccxcCsEoslMM3MUMq5emDHkkV/vmTVRm46osaNz3AesD4NotwDafEjtO3
RFeuXvlVTahK0MToPVDEhm8KEi0ZS55DdkK7FWd5+bh4e/0h8tBhornky+88niM8foVq32QwkMsi
rMoImhI8tI5NYSNdVa0TpxbzzqDqmMx6cWxfmBwZBWYiDf7BB02Vhi4QKJGhbno64JX2Vf8Zknl9
os8VZQITX8i62/7ixDhDQHnhMQu5CMXs+mu831Sw4CFf2ehh9pQRuMIw8V25uxog2V0c4gftg6ji
B1O2VwEJfq4p8Yb3Bbbl3uSkwq0tUY7n9mjpwVJFw5tFjjN8k10osUqpjf4Xxdb37s6UZJPW3GRa
RVnmxKZ6/B/UpRU1m8UhuIFFtVb9T93JehPLOqTycxeLNCtFNPbLrqnB/vdaP4UwmThBm8KWJ8Yj
F0YchApvZkktV6W6e6eGXE6hcAHeZEgGCWb4TcfsQo4V2PpVtXiCeyTJ9Hc2PVKWrAH9sbV7gLPU
oxk526bqdPqcabPhNtGd1n6WfcPwH5I5a1HZ8Te3V7qhbwc5pEpvPDp7wtq5JaDvx9ngmenVNlcj
3nNj54nktcb89k4Xpm2OiVDQliN2HKWSYj20+RpjivIj2b0tOmAiRXhjWs3PGkTIK28TJfrbL3A7
YAn4vgDRIFbzDdI/3vQ1eQlwpNwkGkA+3KQ/TnwMdvHiq7+z+5gwCew5JO6yHJCSZJ3qCj65B3VJ
7lytmsQ3ZMHmNullw564M72IamkO39SaRahBAOYSS/s6twSKxtJP6MuEEufVPwTpRgg0Gx16a6bd
OlOLyfhDeW4Jki2rUAB9DixgnDsy5LGZcCfHuHtgSb1mglLwZTwmzA3I6i00s83WGeZE8ZmZNuvF
287Vf+yuWPDGpCe7VsyVIrb7kAAeEhRfCwe4L5VuRO/PG8c0vSZvoyxzh3AVLzFWT/ylR0105B4f
V60TqAFatk8SVeez5e0uiQw3w/LrMVVEoImLNDjM4aJw8EFe8qfqkvIwUdOM59KEAtITA+jkItFe
iUvzaspMZjZPF/6jEQhev5VEkTyamuNIUkX1DEvcZoExmE13TBHL9uekXBPLSLU3qxlQFzzwuhCF
jJNC3iAANot7x+sx1rUGMp4IIS28sAGLkb6ysitohGCaIryH59jrlAtHwgOT7fQyyCvgD8UxNtgN
6RvALXzr1cwwGyU+ReHnI5rZnQcvOx5e3IY98VbPOFyV7yDF4jCjLoYroaKgeZNS8jZr+gW4pdZh
nSQ6MEY3J/fGlaLBXKQbsFOjbppmyVQPRJtqnz1a3TsxslUNMhgv0SpaFjRYqrzO4EJsWY9GKuRV
0k70KsUp2wIcGjyRgKnsP91sjuprgj99M4AyDATMT17578rCwjdXj7sYxwPaCuWbRNjtKsO8AZqN
9g2kpE319vJWTf5//J41tYVST058raKBoMsnp5A/Ofq4uSkoGUxForbKjdUq/Njxjth9Fsc2UYWW
98e/niKbpWhVMc9zoDwZkix80WHHIiVJqvHSJOwERLgBtI6zhGNGM0xsD0N5cYX68KNv3mymzqWK
TwKI28/HRNwUkru5Ps+rS4fiv3QQ2yzHGpzlvKn9RpwDGRieVpRNHsy4woPlkGpfy/kGBtWABekI
0bhDPGASphNgyjG1JNjHXZ96S4QOsyioRL2MECY5jSmY8TND+ezqRdMlhBfaarR7iWszVXwq5div
AEqlw1cz7zCs05HVjnQVdp2ysm1KL1kzbF3DuP32N9t31ITHpHrUA1y0Oww5/Vh2jdSj37mKHXyd
A52hburJKmgT4ed51NDSG3pBJXVx3viza/9lPFwtYDEi2JkXH1MBaw+pQggzkcawXiPvZ2YWQnFI
MnnzRdm/igO+JrGRXVYGIF52X/Mfc8xNsRfJTDBnB2J1krNBzZAFBkJvWH35FJMzVfY48Db1MbGi
kxCPRME73lnzkCKI9ubqaOuXx8IX5nr1Y4Pu/IzvGnH+mL4xpLSajrKwfYukt3v6ifraxIKq+0G6
o1t0K6MhCO+VtaSmw4XEZvVJXQJKjMy3OMh5Zxg+WCN471g9rhsJU1R15p1mxz7kaN3wDib39q+R
f15Hz/BZxUqVVyCJmxh3QyZ7/VpM2h+lZDF4oqmOb3oRRItLM7pL8NVOvWONupgZ3vDOEZsCX8Nv
U0arYvImGclEIPKxzXYKF1Wj8iAEN1C8/2vlq0YgALktYoAdU6NsdSf3bVZBlFJYTC2OCwcya3Mz
B7H8Ofx8RZDypf4sfWGqR/0ndqvUMLH+LrA96h2+ke6mDD6OKZXuLFTWQnxuCXSojtxfyg3Wvh0G
n/ZxWJTp6TXgZZH6gkQlv+LiGw7HeiEkmG/0BvGP/Ms1zJplI79YJtu+0buu3WBosvoOLDjSu6vT
y6d4ehUdGp/bJjuGrJCJVDpy2xGWvzFQcD1O6ydpUYtt40lq4aCyuETV1/cPBcPvwbYN9SRQE61S
2KPdMSaec8IzTGpefh4UgQFBBvEGhpUinB6P+SerNl3yvC4SziijELQCJqTinF4YHmJRcy5bqvy1
phVN3HDYj1/OLt4aYxTr3E1yXXmvnAmagBWuQfbmtADAmpjUQ9i+v0K7JYOWHvTu0beod6CJvRbP
8EWSFBQdGPNMVHjeitmuLWizvTvlCoLgNurQb6kqweab+8r7bndNeeZs8RhXBmSV1iI7aONvu/ZK
iGI2kU/VXFNzg4IZY3XuBZ38rca1g7zI1xRbYtW4cnW3oS53T9n8fntaqNa3mllK7gT8F22GL+cx
uwMdzRmMCa+tJqROTi/nOTSEFzeXE4iiXpYQ4lD7O/aWVtyrkgeJ2zJAXOLudntl36jC6cF9msBS
KEedv/Lf9wr9T+OM6BnzHY4DaThQFHsVcgwgJKnKc/AzD6aG6Fznh1yqnh47ZpjmE4eWvhb5v/5X
GwqSpil8pQSoRTxplc6Aopk7w9eMbzzHl54PGueJHGtB+fxJAnsOlw5rip7e1BepVDBwU608GX6I
zMyHAxPG4kKMJpQTz61tK2wrG893CD4TNsly59e/iAZ1hvqPB3xpj7QsGnHubVcv6B7Ejhr2HLnD
MVAadoOrXsw7NhT0XCNDe1Xc3W8PNBHDHrpBTsv2ewI9NyUzhZujfOUK02o02vhL7ADHaTVW/wQz
1/Q9JBRSWMGjPj/ZuuNz5p+8zryImZAmb+ReUko8kKcZgOc0YfIRt8MCDqytDHQam8lZaWHgrc7p
kFSX0S56PUF0vFcy/U83bWb3to1RFlzP/GHkdspzlXk1aCSjfQmf91g8mhOeFhFg1a9tp/9sQzPC
6/TVXryb6Idc2e2qrRU/sW/HKMAqHmD8EMa9yxQ42JwhU65D9ig9gycDVG8fTmhyoWYo2sTh7JK0
jVdtSRiavXngvMBBTL96rmgszIwQC/J32T5nVDg7NMS6TqtovFJNdyANjwhy+viEuM/cZ+MZXXBW
mQzM3H30aFkRlxcNfnk/tvRYnB4QfxmxpbRCBzzz88qr+8luiS1FKo1Jl9gJVwZppFAy1zykRfoF
Kp6e2qj577Jdqf3e3gvjCwZPP6oPIIXav8LooemD0yc6P2P4zDQv4+h73x4NEMJ7JAg5PcRhTb1z
I/qZEmlr1BDjR+qqJOrGLGDw3KMjiRSmWrx4D2AG7ctW+cpTjndPMNGKSVmoPhNsd9l1rWsl7jjD
U9HZos8i6hzL8pmgYAlQlepmFTfv2hLLqSFycavyihEH4DeaGRZ/M/SWUpkwKz6zwg8ILxexe0yb
ri1mPjYszmpdBs+bLuClKAoK0bBhVjsZnDw+tanqealxvd9xGZ+zlLqIyvShyxS9fxjYprvspNFz
ghU8iVnx/IyHJC2VPIc3UAikZoXyW1avA1CtECfIGY6oJ6oJazqjNd95PVFOcUpmSDu3ZZqLLAie
8a+neGBBcVEpMvqjjS5aBnk1iNyZW7NOk5PsmLxCB0XhV8WNkmIv0oAGRAISXKSjuMMxRpEZfQoc
VOde12q8wj1fHlLxnkmPEUzuhX6xYs1m1jqv1uRgBOrIOZZm3J3NatT0GPSKmpz8n+o2cR5U0/ch
mWJ0/QCxqyZ6uW4PaqAcyDnodOrpNu5oTgtFSRH5CckC2DpOZ71mU2PLDPfdAkeYMiTo3IhJEyXh
3zVJWZ8H9K1J7LrQeDUOGCxcQj1cB6AEVljis6JbF6jYwWjXZt6UXLhZTrsj9pBDvvBRMrT8PCg6
hfD0wdonR0hiVyz/BqcogSC8GnTCmwsOHksjSeYf7dgOzlAwlKEBOV0es14m8gd68pOZWdxs5i6S
dUJfqYV5hHnVvLJY9bcV+zq8dSdwm2L0X5MHFWnfvfhg1VxnXDlik7oC3q65yVXJwX5h/3kpQsa7
f5DY+XdDA/DaYkODWZF5/Q9T76GlNGG1JQ1L8URL+g31OASLbV/nThTbxo32DOUc6zoafGM5MVa6
cTYACp5Xiu6b0CEbq1+lovvFknrH1Q7Tdnavpr2jkyc86eUmJ2r4XaqrEj8x/2ul4Xz/J5eGQmxA
AZDBZUqGr9T0ClRt2JiBndVh8mC1TEiM9woc9nayG2exqabw3yUVWAAAGBAD7FWGEYPjxaOLS8cz
0YYtDE6ewBAMZsK7/nbJNHheKwNCxW7WNwaKZmzu0wgUQovi/GKf03Z1bmvAY7RimORB3ElP2pfS
KYWd3vdfSW9kPHrZwxBqp494QwjuGwqOHjKH0m/xh6XTuvi238qjFydVhH4dN7Vg7Nio8Y/7RK4g
EGFZBdhqqVi3w+jTFyhwmXdR2piEoQHv8XYiQPvoUrEzBIEioOfxm+q/j8Lxb7Gz4uvf+6a39Y4i
CjxpAvCkJJ0G+q8op6zfM6Fx02LXLim40M8vveeR3OHlxnFh6NyUXj7rdpXCQqfLrM70jtS4qM6g
8g/UcIVT3N8zwsnkanYeLrM+pMvhqCpFMnauvnAsK7xWNacogqviopx51bm8gECAklC11Q0sNXMM
FKAlgBl/irCmphXqiv8yoVQxI3icyBAPPsmOZExshfMDDEYha8NT3n0rhBjOHwssFAwXb1UEQWhC
1HgYIpL9o1fMD8ZMDr6cPiaIhfyGTbDwvT+fpr2avuUIWn3DiOJhjooLk7t7rt7eB7mssmUyDmil
MBMc20Urlq+cOu+cVy7C5N7M6K7JimrfY8UO5L/LZk3/Zox3ZXmE86jq5Ec/AOZfAtBWGvGQnzOs
yREgq945Lgdx68a0SPPy0z1CtbOJU/mwRoTsbr2An4V82/1DEbRIeaRP3/hRSmnSJhghG5dP7Dxf
x0CMDahYv6rS9kc9oj+ASYmOP5RUQz7UOFDCiiS1pRzKzO9KAeR2w1lve/lnv3IPmzWfbNGQwFXV
7/x3oVE0OVkxfIhSOdAWeaGRTrIX9Dkq7DEJHYPyF9chZMPMRcBKrWd8C6ig+CiD2Cp7aeHrcVVQ
siEkvJfc6CWG3WNnJHYHdCbNWDlTG8vXB8f0XA2BbSkm6MoB85z+Dwsc2R5MOj4VMrIs1Jrp1sJI
gkaYeqQDUD7+Tt7xC9UaRqaKKdlxOnVNzeWwD0Xr4K9o2xfBbhmNtxY/A7HzJbVspVR8s/vVUFx+
2p4JmF4AEDADd0orW2fJQi/jtMo6cJFLSd5Wz6h9YA9dwUtvC9tUap/Vlasz2IkLEpLr4vct9aUC
TbLA5CCQUyKtYoU7mStGbvV2B+ldlj3Co5lcyLJQ+qGf9/e9urqUEG/RF21PDbeyZ99SH9xAAQoS
FXpL7rCoi2mrI9Fs0U+ehQvcOIXNFNX561lmUC56CB5v3inKggugvBSnbmCFUGUEeKousY0/WjK4
2ufmHuaEOIrwQxQ0npl+hJb30QFXNHDlbQQ42DGMA5esBk8H8n2JoLp0zVdV42xZ1yBhlfdL0TjK
3CmHSirg4GDW4Hj5i3z6ReRNaCSuq4xrpT9TVtDFUj/9bB1KlXRoZ1Zz+Yi6jBQg8n/12awtRylO
o+gdlXyR+aZsXNVHXLaVgvjnnwVK1yxYvsG0oj5gcG/d0AhQjA4JTErXk6ibl2PrzLqOot0+X65j
FA8Uy6+ZaCY7zU49oJQgsxTb/jf7aw5Bkr6PMV9SLs19QZPCe1mI9OVrSnkk1Szus6Oy8CrZ+5X9
m7mphoZUf5xw7KTZ4ibKqyWgvhiz/vs2Ka0oBSSP99fhF9iqvSdb0W+6buHZ7hX97phqXcC8RSQX
AokUJiMkmgm1UrTNz0AVcBUJECQMzfiMEXJGN9kLm4Me8aTJ9RRMKirWAdojzsH0gZXJGGMr2Fuf
JyKe9Cb7RVGvDIdJSi7MOYG8fnAGeZLKQ/aUt2WXthuxTAqqOld4cIr3A5QcR4Uwcq9OYUnYK8Hu
OIaYAYME0jidbbfuIA9Gz/dIn5e6NY4rH9EqpNYoJrGES1/r18vUFFeePlXg3c5vmFJ8FotuzwzE
OjuvWQJ0e3j9eqZxUMqy8i4AG52v4iPuBuYTVi2L9hOIiQU+hrw+Rx3J6kZDes+lDmg3YiRCp09c
SR1/NqokUk4NySH4Ia52o7X8zDuXDtKBELoYlXwSdNRFIFBVoqxT4ZYh+RnVkEqfoDgxw1Dj/LQK
emfPzyvtzIuVxrsoc7r6JGKzCZIWfu3SHy1YAmW3eRn/v6fLobj/Prhu5ItoQKDrKgoIZ4IYlJyh
PGO1d64jKr0sgW6547liow++HohaXbDSydm4eyZsqypkBDgycaMJMFdXu+q4cD67EvT3w93W7V7x
OShQzgqm4+TsAIzK8gYjphskBDIQy/XuV776YMl0F6fnxbBHY0zuuQdH1Oyja8lkd6LhvWAWEW3t
6uTEG38UWVJRaMP0Gq09yqLx7Iv81NQnvOEN/D7OQqpXg4cnpGN9PBAKvqPRDO8UdtdFUYKTbiiM
EWkFkcUdnzL5ddmIM5fWW3A373PawCRxExuyuwEI6OqLxOXpLTL9APsiIHNBBafMyj3flGomHyRJ
4isSnd9D+2wPmw3lwkBXDymRum9svGrHSs1JsgABogCy1Ycto3RxxTT6XZiqGiqXQbEWm9mXFL1b
JwLKO9CJFbtNaN+8djwkWaqNP3iqcvguBp3I2Fp7d3wDRZH25ULYKRX9l/4qM2hu9Ef8aFVbNEeB
PfJ0PhhqEeH/iuPwtuti6DxI3d93x91JMur+198tbMm6xzEfAS+Z6AqT478GTKoWl7MEbyr6chGf
cGoL0qZ7ixa3Ykd6lDLThyWc9YDwRPD0RTBCQ5ACRxNLP0GkaEszMK6pfU+z4Hjz4xO5gg9jG7fm
QcQeO3kHoQjQLVGjaXQMgRKV5wiKoROjWFc5sQFV/wdNZJJLyx1fJVuLorwWTWkXpGn7Zf3lsMdZ
RR6tTk0dgbE70afJvXqWW8xVAcq3oaN4giaAors0XNpGX8xCnK+zBqEEMNo0nv8T2wzDUMMcKlMy
EEntEgti4c7tgvIdkvCvyIRg1RkmNeqz9HUpuR0ddPwXjkwOAEeu9thIRRWZqNo7P1vsTrApRzRN
W+PgcaF7/CFBY683ROd/ZhPUJjaiPFnvRzBgJsJBTJEaXj2f4f92URXonzBplR7DnVlwKip74ZM+
RFFD1ktyLot8IyV4f4FZgQOG5Dfm1h5exdkAZA6LC/y9ZWiG7p0lxJkKuOEDddIrCOquaKIS2hLN
iSDPhL48wteAytAY3VUUFtc8GOji38eonaINrWRX1d0WDkt8xobNDgDBJ2hQEKjIxs/KvRNZ+3v5
u+D+gTEXn055fidbg0QlqMc0vjqL9/fHj1ri9T2qWb/Xv2l8mB96feipe2bNgEdrwbjd4KYxht7F
00Zhy1AViyONjuWT6vQ2nKmWRKtEz4MxGmqX+wKSi/M07eXU8xUPuvfpG8ImHv6q7pnhiGlSlMLq
fsOWvT1WdnnTLZdJuVje+RL31dUxFVUIfl2CVQY7kfZ+Qg3t66tgqdDxGRqyY+qIlGHYIgugFC9d
pqfOGjG0zIHb2FHTq+6KHSjRUGKSx6fkjCsg8IzAjiuXZ5n+6GC6DeIS4XuMBrCUCGqVPvGa/zPR
/r2Rn81gv8xvBqx/qEUg4zzw2jwU/ATqIv8lOqFKCAmYqBZQYYkqytZX7DdZy3FF+AknDh1anrZ7
AGx3tgzjPpJ42MzJu/hWDfVzZIRc0ZCXYqzyI/mUsYmz+XnThM1WQCeTUZIo/Ol08pIU9sym2MHS
gK8l7vMoXcrRJbg03zqy2WGtuAbSfYSWxNUaU6K+BtRQIA48//uwiHlMEFjGyaR6w5yOBlssVv2D
bXDblRiyH0cOGZniIdJAqpiLeEEt2WKIlZLEyOsqBxMSiT/2XmQtIM0EB56/QBCO1g1/prZ+xdrY
JZsWLJ85OaWbsFYzhqjTvmGeqv40JE2S4BjJAEpwiIKetiDpZ+PuvSFQMsGtHh/ooMzDXG8n8nOd
jMl2KCXxaWtPDwP2gqBTQdVm1Qo26/FGaAhpAVszUBnZRfblWppObQZpmsOtz3A2+i2L8rerxn5e
yGWkfR1ypNhyD1Ay85I45hJAGGw1iPc9taHXDC69iH5xKzdpV3PbjREPmkMvmLJ06aIHamvjf9Vx
C+nrB5tKNzcqVl7dVDC6uBGE5xKcYgUdYvghvQjPk5w0LSimP6beI+he8xZX+WhxrhzQN5Lr37XU
HmCm3ml0/jmhZDh8Jr/GyTKnECvoLCXTq6n13cp76S95g0geMKznLzfnD43jldQCFCg82LlOtCM+
tH+1PBD5FwcmWiwPrTOGOGSnUyy2mD90IVJ9BjjZqL13p+JsV0ajFOn9Fg8kp38xthDWXToPXhWw
wOZIaWyJOWqyc7dGkPIcaW5lw5shVhrecvO2VyCKjclbvu+4gq5QzoFa7mClHpfdpgbIQCizoeLm
Jv0Zl+GdNmv8pVgc0aoAiiEYfsTZzCu8FxRSuOvIAagfBMMkHn3cTdsCji52Ennq3qLLvZbSvlJ/
RqU9AsCN2hY9SpvAQ/KjNAiqQDRewxlr6KK/OxGtG2vXbQGeaDuEq/poMIT8BaF0DTePiSp6uztD
IKfGAN3AQ5aeRQST/nDhQ1v3/VJ3Bk+c94PUGVOuoThnjlfFzeKbezVuetyvkw2YkDNP1IPVrRPt
Enq7mm5S3VUmmWEDJrryP8WBTu3sgovZItArM2o9T58JOkx255HSxJeXfl+VFNHZ3x/g4cXCS7jN
CepqvcdnwyMoIgm/J0je7rmZJYpE2hqWz/f7z4sybTImcLI9Mv8EdfnA/Cx4at+7CibMKXx464h+
XZ8E7MTK9QJrXpVgp/3zTuTJjlFXlncdlqVhrz9RFXMquUtJr0jDQ9R9+Gm5IAr7Gkem4oTuTG+4
qrzP4SAR44sXxQSn33464LOOIIqQ+JkxGTtkTW7rWlwIjG91o1D0VOTBLu+i5Ift7QtHDnyyc5et
yz2WhEHUtw2THqQWNx+QRBH96MBb5VLqdgS4gAlYFxkQ07xDM5XV0nKUfER7t7KYQvpGsvqXnEpv
2Fc90r1vbSfZCUtdmz5mDjlXRcBF/xgV4nV3pK+rn922ByqFIc0kRsrWXxQPSo7QPvjDaWIclptb
pTlrLNMghPyMGaGMCY4Ey2t8IAQu8xTf0VSHHcsnQlfHPgZyEqJdQyGn2rKJVBeQGyAEavdfmrc1
O3OokRtlSP3uMTTntdcCMwg7U2aWIeXOSxRkhLujtlerq6uzkS/oUakuERLsinOUclLfsis5osax
OqiosbCFlMNymwowuClSxXmnDJeSGk3d9fEahxopX03msrxD61Y5wwCHS2zn3lt536QPwxju1HD4
8IgIUU64mx8d2KO//VX+nXsqRasyMGCqSc8RdMRs2zbdaX8vTseGmqzqunNxdAy1Ee75WGmU1O//
DxjXRNbajZECq6m91VdLuC7G8dOmtT18BrmGWpNBb0kD2Ux077v2FU0Ui2fdeswO2zaOVIaiNQt2
eULIDSi1XDFTXw1YUAl3GPXtLwEwj9/IC+bqvaLQNJbY6+PVB0t+rq5/Po78lRGJ3EMI3R4wW7Hr
4Qq8A0jN5pnna/xB+s49GrJzf4mYAe6qur96aW3IQMDY+vI31DRxjqLJm93tpToBGcUBjW2+CHQt
5VLJew+sbjFEpxBlSpuhJuI3P5F4WUlfqmcaEc+/KE7ZOVNuHmrGKVqSWdDVVEU4VF+jOtQr3DjS
1iwscAZJurYEXovOACEzt7kAOLjehjWdm1sxlQwD27vYSFR5Nu1k1biYhL6u5MaOgv6sGblQsFIk
7kwf1IIqQ1uuSbom8dUyolP4+5AgyU8loG3pcRR5JbGJwswu8OEtAGBokvQ+jma1ZwoDx30MsxvU
QdK2R1X92nIbBllA/Wj1LWJpzYjrl7RfHon1kSgxnTKyt/cLPBEFPfRfPvzgKg2woYjNMGKxsIXX
AP5TzQXfFE7rg04LzAZplaSUxhvEZ/Y4qxn2NbeREt7VebE7kTd1NqFq+W4iSOzXExIpUk/wdSSf
NlbyVSv0isozaqEJrb/pOaSwMnL99bXN6UCNNBWCjkLriafjHHd7g27oxpyVDuEP/PwUv7IQfNK9
4Z4I+ZORgcspFtP8A6T4bZJAEl02MiC8LIXuj+8dl49YIyRudxuXY7cqacnR7BxzS0jnwMMgkD02
ZrFymF+uX9B1ytW0Lnprf6QSzwbF8FA1IEmbTfM/aeyyLyLcSr9SFJkpy5mp2yiPuvnB2x4GthMI
VUfQ2U6L/tpYJLheaBlgoc8d283bN1lRodud24WyQSUKOO4gxRzQnrn46+ZYiTjq5H5UjUi5N/nG
HT4c4NUOIwK8imiAuKHABvCf6YOoAa7fU2ASw0yPVeMfZfnrFaunLy+LD63Jvw6mtM3VsrGCHEHK
fzNd0ZOpek7obn0yVTVmyGzgUSEk1cDXplEUwEX1qPcRu046j6HScyRPun3nrdFvEiVa/oFefjjx
E568iSOeJzRFdPG+f42WOuKBPRZh+RXg0epPhBC4H/OMenIInOs7bMi7lZcct8VI/dc8qRDNNKDC
93OKtv2/HtdIgK+Mcaht1xJUzr61t8h7SE8Rb/15L3IF7XnXJwZ51RmGt6x8bi45mc6FaKC6I9r1
q/KdbpC0GWlR4olvbO2UuP0ldkWcaxx2lgS8Jcr3tVlt0wH4JjokrwCqqTBT6hcgdUWFo1lcW8dl
pcRNTtoPjZeBoJwNt5PwZwzb2nmBxWdH8lsl9YKB0aSjhFatoc8d7dIvqG+bDDFP0VDbw0YXGiW4
uvvf4iVrRRBsjVhtWfDCy5HORVrrVpjrRpB448GcOFIuTMkl3+b8+NygWpu40tMdlFqVFvUdzSD/
0MHtn2X1Tl2+4N+rri3u/cIXIbORsBl7lLHER/BasR4N3fXgiRiW3dsuVISdSa1M0Nnsp84RVW6N
T9zqRzv138tHULm4PI7rowMQlwnKacCYHDJwPM/di1XP7l6gZE9yjQpst0JeQY2MYGlm63ZG/17v
fEyzTBeKxHs8yat1rUAvinogzBCrAgoroG+lyx6tmWOhm1ThtMFgHIs3xc+ksJfdpZDlP8tmUTzD
+zETv+fzQRUjN1BoyjVVUzRc22UwNaWsML3ySlFT6QjztHnkbRG09rGtQFyaM/+q0Qwxo4oHB4TK
JJj0dNfS1Nzsnoy0IwHPoDRPqDnqpn+7NtdAElNaAtmL40qIeNOxFeHUdSBSMnnjDQLxqGoFigg0
gGimcBBi333T90ZS/dsrh3W8WYO3obe/eDyqzMiaZwk4I/wDOYjJg1SgEbvq4ReUiwK+uqDS/NM5
FHWDZdwjyO6esemMc18aep7TL+3gpgCJB8gzt5mtcjLHmXJKKe4BzVsiETOzPnpJFqIWzL/5SzTL
OvXHHB8av3RU9XkvjggT+MuIiLZ6sLfLoAnksNF8V+6bA6aB/LhYgz1FHEzvbsKGBy5NweWvt8+O
Jf4yXbcffvNaPRxYmbTWwWZCkFO7qkOrQhFVpW+hrN/GeJ1BgqUv24tTOVRvfFlu1MdzsZp0rPxs
bBc1iHP7wNqyr2fRh/aMk81WAUz6mPfpQl27eZkePlCjLqNkVymsc3SC5z32u2rSfCGSNV9lPLDT
POdCXMBfKhiPnxkVsDM4FVgsM97DKkCfrteENQREnCoHfpMdNV56tS4bKW7pEXmPp8acNVLzv5E8
mdlItGPiiuSJOVWGnAVFhQ/3ayXNbXoUnQAPrea8Mhuo+W3BEf9UCg7wL6OEgTeLUw7BLyc6rcBO
UF8196JXO1BXgkd5r3bSJ7nYQ+rov3EG8BrVX94v+GLMcq9i1ND48R733WcsmGdotXYH66vhcRO3
/R3Qu6PNJ6lCb1MPp4ur+i9rkYBH/UT0BZ/NQAEbM4Ar2QxWiq2xev2K5JagxQLSZqS7+YAr+lUE
/77BgSSjrHyadCQNhYSZQ1XeAPa5GZCJof1PpK68EkuLGj0uVVRc0iKuwnB44eeHtlyweQTBQXPF
yjo6dLPP+2i4l+4chuEdtJ5ClEFB1lXJx2g7DZAMYEvJZD2aV4K23+99nbsL1DZkhmCS/766a6tR
tsdDgmEdBbz4MKG4phqmUMz+hqsBpoRkGpOP3FZNB3kghE1izP46pIYOcJLCCZg1Vu+TFl+FcLAq
DtuBzCU6mTHr8owPWgWp0JY4aRpPgPauSl21Ihhixo87HNBDzN9w3I+L8wMHj+8wLaMhSMYtw81P
0x0Pt3XhhrFs4+4EhgPcByj3LnvZ6Gn3forEoiytCDSdRcfzEUICgfus1zlBCfO9nJI4aXVftUJ7
lEZM8AuMoYb2oCXOa/pjQTpSKjqwL1L0icccpjls9SB8VULIYbeFnc3Fzu593du3wNGDr7sB6Hzt
Im0MxJwV/Aer/kUjf/uSdzOHAFDuvpK/9/fo4BjlJ3kUwoLKOyxcebm0coTMiloV88z5QGSla4Qt
JQrIU37ETDdRKcX1RyZce0DcleURF7lXBsRFjUhkdRIlJaGUj4oHQrM35N28MlxjbMZkALSLZqIv
OVv65nLcZEJ6Ae7jLPHtufNgydpdAuM/U0aD1zq9eurqJLsxO9eAsFiZpbhRc5kqUTKyWmKtBMwr
J2V7zZaOfT/EXqvvT/O2r3lIjAM/WRqujyTGDCDUdn1/oviNhYeVzjl1mthgmvw13AEfwzkNdxsH
/sgkh5wJz6wAbft35l9BJ9gtHNSASgJq3+x1O+/EHBW7fBwMdB8tlhjKL42zgpHRHVCVsDjF9z4u
Jp0Zm6WKI/B/jbb70D6xHsI6M4naRJxtlL5hUw08B3nP29Q/lkyocrakUyy/5ddZZLWhuGmSfrzK
Y7oyuYE/R/3vrM6ERmUxBWbycGN0BqncYLJmFlj+Q3SHn8KQr6c+DXqF/cCmZoML/+nNP3gXKYYs
lyi/ueFllut5OrymCsOsKyTqmQk7V9E/9uUgEQs5yLiHetyH9OVxgTB+VjXyq18uoL0rMPF61BW+
7s98Gpc6RQ2QkT2q8BNnCQ+rykWaVq1jCR653ITubTLXnfgfL/i3qYCkI5T/n89vCmCYUSMcKjwf
ZJV9+IbZ2caiYhawghjcvr4mlR76GpJsAe40qdeRzwnHEhdO1g0qKR+N58Ih2CsgKKUyaOtuRxo5
o/kos2GftUbg5cDcVDYFST+BoxD1pPd7oK4c48ZhLRHtu8Jl3UsLQY0pljv4dtQCu46/8+b0o+Rl
9lW9HxbW+B1lMajZ6cPqHSWEqJch0LHySOjsuIj1QVjiWE2poVJmm5vZO3g49uTxwCqxXrPIwdAE
smw+gVO+TM0JnzbIKZEdlOZILTz80lp42rhlgIaGz4kgrrcfaSSNiHLshgeHsnNA3RBEusAWUTJu
raV3Je4d71j5+ZXG3sWLdhxRCc15epoMvYZDFYWEOzS+OPDGKIq2gdGic+iaLeFjx7pFHlPls3f+
XnT3jcxGvE9lECjHb/DvL2sSoNi7TykPXVIOS3qpBPT8p/BlnMMhXCZAAbz2nD8LuwesR8GsOMgD
XDLsEg8nyJqynNbGxsoibKE4dLcbqbDBqsgKc0ac3+oTLGPCXwTItlYkGqkmXfu37qKJiJNmdoBo
iqDyWbW/TtDQ66dU65JrDlz29veHac277LMQUzF4FXWoFVjhelIEeaaKkx7BNPqvanaOWVZVTUBW
GzZ568TdFYxT4Sr5ZwCYCpBAZJk9VlFrMMLCUkWPgIwTdU6rpUMNVQZ+6F00/yHrhW6RUwTTuOAI
81mxJMQo2E8Zv7O6xhj0aO6cn9yGGBCosjY5UTR+DPGs94cq1z2kt44KGa5KB88E9vYapWALzijZ
LCysDIAKMJUpjv1hHxBFHkUvYla3EbAK+5pVe+qjSjmoCNgXcZ+bgMsQ9dHV97AY5onIMA6IzXIc
Nb24++mHjW4vLC4KdRqS4ppSqa163XzLXDdOc0ziaCtZJaPNc7U3vMfvnAxRZt2iz9Kix7pp7QOp
jS4Y620phgwRohXa9Z8zpWkootUAhp+CxPt/Gy5QSlzIpzfZJMNwsyCBTJ97qEkgBsYJf2iXdZKw
QMgYUWC6OxVtaKHvtQVBiDjrRG0aQnE6JdNa+Zho8k6oU1T2et2owSDN0EDxMBvEAN9eDo6rkEc2
tabZU7/fe1FDtGCMvLRI+weAkv+4D9teMSdT8Ql6TrBqcshF9DkGILD0Ln9Da0nlIURezk659Cfs
EUYYr6MxNQubWPmpwClJtp+DLONE0w9+YxEry0u+s/Evy6NHG9kU8M8S4+2BHIaRmTtbBW3t9xlc
0L2f/9e3mFpuZyUvgmUSoJdjs3EdOebGvOxaEzh3D2cXtUuP9lnEGqt5dI2kVWDyswLCbZ+q/Tt8
uempbTmONaLseTyQ6aKRXOu2JVcfG7qZMuoIuurTR6XWRe72WhJybxmATJ4S/r/vyNlj02KNYrB1
o5gqMdIlOOeVo9yI7zLPWpNlYHVp4K+PFYpTCtSll3HJrMs0hLV5+JasG636X6FWFds091Anek+l
loH9nJgEOpNmYU4M5V4Jg/DNcNsDsN6/zTXMgPn+E4w82W2MVgzHD6BKOLBfiosvjirgoPc87AnI
CLI48go04kl0bvZe1h/txGWoaQEfKLCY+C2NjRTeFz1XK6lZK7TNgaOpUhrRyxeRFLTfcUM3d1z2
HKj0gnaMhUYWOkk8X2LCn/JzaiGqtW7gHQinDMqaPfFBrp6K9DFToRlW+rGAPCPzoPohZKijEySs
7YJqh6YUos+F7pdIFoegffVlYAolgEMq6t7HjMepNcptXaD8HGBqW0gGFMhlbJNU6fmDnQDv6+Sj
ckIaQK5Zj9s+RxxFxPOSXUgoE64WHhj5XNMqouxGQ4L2rMQU0rFEAKocy+sjG1+2xCZjfsKrez6f
/DzxBcHPoGnk+09i227kdc0fgVW408lSPz1Lbt+hL+7k9NPZ4WQh7QGisTIBEyY0bXx/v7Tj0znN
xHubTJlg8ITk9Nx8U86LR4aVmT+dEDPWNg4O+qKpvqHNrpSANVe+Xk02mVwLsbCMHvH652MnUU1d
6yZMoJfVPOVxChlDyZSVSFKknKrVzHgFEU9HO/pvlufg7YB4bLkQeStgnwJFA8SfuH0YuSszVeh9
8pL2mpuCajZk8DjERthNzK+PcM8aSW3mHMt/HyOIJePFQDTVG9ryfQk/ksyq/BEIOxZZI0tHGM02
bEEA5GYpVj85SBB6hBhzAqkWiMM2NxwF2UcUTr+1Om4RK+URh52EL7l7pvmd0dYK6Ei4zLdJC9wa
mtxA4qbgOVHtRvcyyijR+9RCvrh5s+fIKjusvfkDCkMP93Tt5H9T9HstP3RHRJtxO0lins694syb
UYEXSD6IfIeYD5Nz1j4RgLinppXZO2iHulBVM1Q+1GuyyFgjzcsgYT0+Sa6xDKbJDhg0sQBUIlMs
4RbVVApxgQrAsy6WhzOHx5/FCzW3KDwS/HxzaZwOIWdMiTclImSa6Bxcu7fveyZlZSquJXjwptVS
6QBlz4zqTHGl9n0D4onWz5Tkd0N3ZteJTEAFbBU/HgAZ0RrOX1NrRwu/9OZRKDOM1g35myDI+faX
2LxMxta4l5aw27PMQX42ePQcspf5gcJUWtAoSk/Fm9WacjC1PXAjNU0ia9krdwkjaBU7VGi1lmwa
iFXppnRbACKXsQZ6oH9x68zahYWh+jpcCCSL3Oto2M+qFG90/KonLt/QF4SD4+qugPWG8VywM2B7
hWdUWaGivWgTx/dXH2VKzDEhxBHeH9o93OxDHMZCwNNQ7Or/ZaEy0LcrW9D/mZQ791SdXAm4OQDb
VOZVj5tZ9SATdgL8zykxDboW+zfsB6IjHd0Vv1fGXouvFgQv1BIKw5+v+n+rVVbbbaCc+hR34ZUh
k6+8KSJ4/QjdTx7D77b2gFpfcHTTcIbr+1qAqDFMuSxiQOVIDRNxGEHXsDgLF+VoWrOEBbyvP0dU
7sRcOCrCO2ht/l18RHCejsRqjYjG6/bU0hkGXV2bCnASkMEzioAqTV7/jgRoOLdyDjEj3o09VChe
o0Lh7iUtFdpvEUC6jPSCvOf6QDILTeGyMqLG2Qtqmls9kHpg57IX8r7GkyUK6s3AZmCf3ehrwijU
QMsZDM2QR4eOgc8g2q8BuieFisq9Roe90ms2qaAoaurn6M8Rw9Z6Xv/o1Cx4s47ovKXxD+Eu4d2Y
ei/n85VvCVXrHKyrrawctd2x7PydbpOlll3oCW+JkLWxHMB22tRG3EN4bsREpztO/6ZYE5PKlH40
jQl4E+uIAhwjjP5k5EAy3Z9OzKeXcOCEyhR/jP7Xm50FixbwT4s6h/irbx39AVEJDE0BsQ5wmVI9
VtntCoM91KHA6YXV9WTV3iec9cqDh7XehTwi+a8c4HJXduTK537bP3PW13zdpvWyOqjyF6ZeFJ2M
qsahsWyMHsU6DkxkNPUXxUdXVwp4dWh/gP84/fChJTzxfz8vj4dvYsz2ZbLPDelkiGxXk7wHr5s5
FLOyDDRM6MweX3Yqm2zgooD+Q5XWQlbrlhxwj12yGUsKPAEqKncfsGbPTF2iT2nKnNdS/EoIa83P
zEuxotxS0P1YeBLYKQc0K2Px0PCe2Rd7zILsT1zSlk0Lid3PAf3e5mOSSkFskL/2M6VYrY7Q1cgB
GJnNxuw59s8ugxncnp7GD1866xONHa1xz30MCbx/gpnsmDl/OuuMrJMCXdjbbGRuVVn02Gn9Zg1B
rVweiSQ+n7Jq4TACGdXXpfaRVqErocWdSLpqBhnAMKZpau00RG1WzXJZX+qWZ0ehQ8RggJkquwnG
01zFmTaRdcdpffvGI0KyqnRCuJTRqstYZdIWrDGWxQVthz+yBfpdriaJbp1w/SqsufTNT3MDWyNd
IZk6HSKkuj7w8+3dDSZOR+NGNvdjV/gfmU/nbEqFNZzgD+TbOAxyO4fnJ85GPdLVtFSJs9OGPwNA
OVCMaZnO5XslfFcG8SXwJv58+IeqyIP3kUb35yDdeiyprJ7fLReAEykbKH56m3aGsnkWL0Hmb/+X
zYOgu7SU5955X5n4kgLpHi5ovuwnbXgXb65gMkc5KAMUNAIu6jfZAs8chpIdX4OucSa5huaM15/s
/9B91VAXa4fJ8F3ddQRA3OiR4nK7X8gX7S8Zm94GzEma566YkJd4/uW0CbRcJC4FigOzgKtkuKmy
mad41+nk7xprAmwvvqibsjIVTNdTWFsKC/A9ErInh4kSFcr7Yz2BwZGFPz7UmJGX08gZANuVlzhW
HSqJHPgU+wtROhl9VonGog7gKhWuitsnQdiMMzTdzdXRxy3cM/ZjTo6fqdi1ZjkyiGX253AUEaJQ
dwbCjd+akcur5kn0RzTIJ+N8PV82gEX8hGnrTi5c0A8GvvM3AbL+6yLDSLS+7JtzWm6m9YnwxqAj
rN15zuSsk3+wpYlWyvQckmP33TVLXirYUqrBIgOEezqVdvwb1x1QOQrG1iSlHgG1ChiQEAz7ky1k
go20WH4iULzYmjKETbTJDYWZlnsYRw54lrdLpWh2uUFL1q9sKT2Z5Ta99hpa1C38PMHk3C3tpUjh
Qb/OoAdIMAvv//ubdZfafQbHBzrGJBbTWmwN+aWXbbVw9zhAGLzRJq1/zVw9DJ4JiBKNIircR2p+
raq/YaVZvTu7seenPy57acmcGZIPlvfL6Wqh89o/ZbI/bctG2cF6SoIdjpYZJORKNA3h5eaOChmi
MHNQ8q2S8rWeN44hRBcgMKHEPIKYhIOQi2FQ7IknKz+/Shzose3Gib0xtBFXOTU4sCzK7ddRWSt8
TBcWwR4p8ixw+CuIIXm19kbqC6euxHE4FyhB2V5stpgniJrJ62b+tBuDaw0QB9G0bdTxVP7weRYC
1m0qioIaPvKBcXqIY1nWJG+nZ0jI4GCZXBA33D2sq/0a/xpgNwNQxNUobmrGIy0dgbBQMiPHVvKp
dRZkm3q2QruuQPEMwDN8u7ZgxshaBV1Nw6UGtJGVq3njykz3xKzq7MbAftZyyWia1zutTDBKqaTc
JxpOXitMvjjzIv3NdPZmZFXUMl2C8UXY2relm4uU6oKjeVgJGTQ+3D56cnXc5SPN/9x1j2pJP1vV
0aUrenBzWavSJ3zCcmi0gh1uL0ABZa4tRwfti6zJHIna689d0Eibxk5tYtpzSCxrxNquJbWdltnB
xtnKgnyqAo9YtwbzEqxFoWHluav06SJ3GudrixQHoUUKz5trhFKXawYZeeggrUy5LQnU5opx1RF7
mc9H6mnKCG+HIOZdnDbXtJUJamauFKToxR0AKcVC4txBk4f4yisXcQBn+KTh2U+NIV87yN5Fn6kd
MJJ04h/8wYiKBpxRITM98dJ8ThPUUZcZlNRMSkRx7Z6haweSHnlLqWXy96daPaA3B0i3QJ7RD7b0
on1pe55g7/g8Jttdr8b/BLpINIWtZOVOP3+GSoIVRJv3e0w6dtzCB58Zvt4nFiv+TdHNHDzHrhrx
eaUiMdLzNad5upcvAruajtnq544xQLU8cYbAfkIsRNPqyGN50DTm1OKXf780Ecz8F66ZARJQYD6b
sm68ZQe3qI7FQlVoKKD73zPLJ0xLiDkTmGUFHJiAI3yS6TkVf2f9A37h7u4EVBJKVfWi7H9FO2FI
fKpmvOedJcsP8Qf2GKFQyg8G297UPeQDnboOyhT7p0Gjyq2uCGfCE0m0aGNZxg/yQvMuFYVM248g
QnCuQopn/ljVyVnF2mFVSQNuVNOqSviEoLHP1dJl6To6926xkWzbTa7tX0qgadJGQbdJWv3aCegu
rSPlj6JkbQcoiRqRnqJ0EIcjBTTn+5C3/IYfEw5z5xc0FbvO9V2FEnNWYok7f1TymuJpwlnPO9g3
0Kz6yQ9ApYJCfp7iw1qzl5OcK1/5CA6NB/ReIIwUt+pcCJ1hkRjKHbyghBm8t7z0WI6i3Orf9vZ9
CtnM6bH2auYZoSUhrKlHQ53kMEMbY9OnV4g2myrRGJO7oqOU1bWjxpcioUeilola32gvwlTb0zJx
/+Ja2iUKeKlWOtZ7BgtR9htFDC+ff8LBGTv88cbrr1lUqd9Kg5kDTHAmNUBtwQzTliuRUDfSYJmh
9YngxgfIvRRoD9SAFP1T0kp+Ja3HUGzj8jYDBUhwRsaXHnp/GPTEwQjNSOhA09o6tA7keOeHSS65
wAhd0NDxbgzbIzTXKgdcrEJhm1J98LFMwroDXixd6YDblhOa00XARYRcvM2t6K28yTDx5oGUDS/L
LUEub/LVsCebG72jIdevK0/NkkhPP3J1l7kfR+vbCJAxrqAQrIEvFlnoVYfyln7qV0YhhYCOwmWF
sinJBDzu9U1V9Bv8wtHNj2ytf0tJQWuBnwEXzap7IVCot2dKj3+I7SFEgbUhvooq6F0YllUpwjnV
knV1BK8zUJ3RYhIaHJMcevGI3+t/zpgQ7SJ9DQg1l/6wKO7BC2s5MlW41CZI3J5BC0sDetimqp2s
EEVX/nLsxiVApOMKndC0QdqXlLx4MKuMHp6zOLZiTcLFJmRSHIYbvfODSQmz1XBWSsLeeOfQOkri
aC3JHhfQCf4IBZpT/RW1DrbfuuC1b7Fl+DlEMXmKr4SWob/XAdTfnIBUc2LrmehniXReW3zqgp0U
MusPwwHFQuieu8Yjo8XhJLQ4AXo58aLO6Jo1bIIo6GqWUPdfYVVjX/p3Mmh00LlJ3KrBPCsg1obM
71gtF5gV6SwvLJJoLrTDOUH8DblbpvKA87D6tDTObzgwlCPHvcsUvjp7U+XVTgXtNWx+oZOces09
XkYY6qr9G8OuMfIFncVMwyhuV9jcak9Wh/WbQ5CIs531zbD8Rw7Sbbsk3V6q7fnonGtHr3KfvrCB
rIw4r0i/IXlYEIIfvhcbVwjqmUjXoT0V7h5fNiYRM252Eb/py5Jbl/a6OGwlC2E2eOIi+oN8Z60c
aqCZze550JAkUlqG1YW5QjLMitNj9pV1oCilyh5VAKveZ41tl6/4Sz6V0GX4zIrYX7TqW9i/i3L8
+Sj4rDX8aB7ziZwHisE8v95AmTa+84Js9cvnWzhKc6d+UX6SeqqMhZHbINe2RUAUMeFoc6Av+bmH
8DligEV8Gcsu6V9ucjITMFOqF86euNZ6DeV0ay3tTLGqATwsIUVDHy6nBi8ub/mPmBDLzSomj5kr
WsJK52Xtu1mUeO5L/SOxr01km5IoEGq1XS5FwzpV2xsGwbbXZLV7tuifYa+XnCWZ03nNzD4ecXte
aPkvsaqms0vUckN0YWeGuXt+21CMvKXZKBxG7yW+l7T1QAWBAa7ll0mBv/iSTlPSYCEkkAP1U2BK
f9/EP+JQk4JBnrmDcfcceAzKhhVC1qxSfzxWSSFOti6Epnqm/lJGpPaL8ksY7v7125ACl6kN6tp7
t/g7jFxtuTdPbns6Tyl6NhTuZ7QgW2WT0bHzw8CME6pVIrtYVk5eLFcFRAQ9o2oRScDBvdvZHlQp
g8j+dRzVN3OXlQ3I2PjOYBE1j4APd5SzMZvpgXOaK5lnkRmmAzO/D2yKFki2RiG81wdj/Cm0TCuW
oBrOchGW9Oo6L9XBqP51UrplMC/q8dYX6YLJOvvK+sQ3XYaNiNrDvHcDtr8+v77VT6NC0Pn6UMj7
quAOlnI+Wfd7NNF7X86b/d3BSgC5Q8iGDlP2QAe34rPsHKHBN14bxeY6GBQKF6jnJ0zxbW/25mAD
sDd9a4JGuK9MdRvPWCitn9KRW1dlWt+iC9Je28g7eGPDuILDrjC5grV8uSdTEXq/p8RbObb3tDtV
I6pHBURaDJaC4G3XQDJcqrH9Xr+et/M2pzLR0rzucswDnUKecHpO9b/MeqXSCYiCPgEbuy0/14d9
wh2WLexRMkmBpplL+M1CcY/7dPWpgcpqyZgXjV/7T9JryDge0ED7loVIQbb7+bDM2wtbktrFd6QQ
tvXCnkZO8toohG3ImwtDjV1y3iVjig0VRtULbyLe7An+2YBuFsqRFRhFGy97l4+qUQ2r2olZ03QO
oyNc+2fDckyJ42y0yGT8mif297nAHr8Sgne6tHvwpHi6pGjCz5U9k6Xmp8atUpO50wtQ5n9HnECY
ytjk2IgXKVOeX58kG5KD62zzHfGkJjumzDtI9m2jZBsjTmdqWvAWaDyCt+uJf43XhrsGpaNrlPON
+O/lw5hou1cryTzg5rtFm3TVv9iKDT2+3pHwaoYKJJRYWQ5FXmSwy4owJNYIXlprNlWof8uhuPYQ
3kfxGB+VwYP1yBSG2RvR8EkJXilB4hr9FUNqEIzyNN91zQnfGrJDMpeVwqAMVOILaNX+1AVTDHOo
pxcg9y28EdIAyS0uKnKdMjp547e3krJttJCoN53d3T07j1DAR292tj1s4uvLWpKA2d2rDG1qKzwu
1Q+3XLBuZ99HR1qHAaeiarUP/FuVf5MyfG67ogOOaj8iW5UONbBVHc6XuJoxnW2LQmrQjZcEFoO1
SprZYB7p6CHfLdYQQmSaeObd8Ab4vMR5u6u008DbHKHs9ASbIsv7UkaW6ZwcA51p1MYEZNvHVrTC
FXmoF67XNY0DFluTBZJYMzfFZOJdMv5txS1D7djcddFPzi6guWAyioD3ilV7EWiQGpd1fq3sN2a/
qvk0moCSaaBpjcFDxY/jTkWcCK+DRLZjUEVz1rCjQ3sacRydVB0cDFXRfHZPPiSD+d9X3HTWe6+p
2N1dhJ8X5OpfTySzs1ZKjNdQr5I+3yMBk3NGEcCGXbt27DZy/GauSGsY0S5SLyeBW9wIk+Mg2MGR
HSy8Pa4zj5y1jNBYcWNnlr2W2pcPiiRNN7qtgNGc5hBc/2YNGLMW1rEW6FN9AupGQlFteM8T2as3
Y/m1bqMd8RV1XyGN2nKU6YWimdclII+19dAzoc0+3WEVwnS7pEpc34CsGu/QmtBdZYyyKplNTSsU
PueBcbC93Y2QmCkW9QbXY20FvNDWuK+2xQuxJbSo2VRE5yDerm64rooXrRBJFCQMAKmOwWdv6RMZ
buLF3m/nIEEhmwaAyQgRd52b4+4p+G/95dmaYI1axB+MB6nIp8r/mNU98+1FGb9yqW35W93zFomU
wSsoxC6YDHguAcMaGBGtGrl6n1ztHdVTvPP/hi6D+fQE0bG7zdv9puTepLn7rKRHuT183lSSvlo7
UeoQ52+tjeSlcGPp4xh/FYCqdSHF2vVVdai1vAGZ90JS5eTtfLGgqThF0EHtJMXd/p80rKFdg2pE
0/Lp6zHJJVJzIviE6Lbw50x10FsOEdTYefudipBQ8gK5RUaxJ9xBXYol2We6GMSDyduG6fYZmldp
xXkwGioAM3PDrf4zRzHTV51SzUyvmSgCuolw9KYBvSls7oZxYQeU13ZXgzNNeuRceRC/SoCe7r7g
0VVBcr7Kwn8MWYeC/JXKZDpX7rOGaNuijlrE+EXSfEjiDvxsKMDlRWA0F5JY8B2cTZ4heZQNCmjn
aOmt2C+8yHK7Y8mlxzvxzxBl4iTbDDWUkpvi6E0xZFWkfNY84E5gx4hrjf7BkEccqvBlcndsxQ4L
e5YvXvCJjdCE3nmGCal0/8cZv894jEeZNk1LZHyz9aodb/0E4UxQvq+iUWGCoObUMS10i7DC6ukx
xjozBrvvVb9hM/HoQhyeGq0b0adgQXst3n4UU9V/To30/GhSvF//z5zPpfnbZa9MMYOhNDnQ6T7j
D4DGhKCKmhr1Bbr8zhY79AluHuU4FnLeqmILO1vWendt9sJLE8XQStpO8wdfXG42IbmAg4qEFsoL
C2BKTC9XDmUjcy/Sakp0QaTWBAsTzCOYILR0kP4hz4x3lOLAEJrJhlJK1yzBU/5HbMhs80+UrrR8
eKdUwAH5wL6UXRapc40CJavNUj3nVpXwqRo/4sa2mnXX/xdsXSMgURVxBM17NE8h0tO0jZor2WZa
CMPDKN3KzDrfTvTWSJSB7302n891wgkJXkyWcT36RW+8/bBHTUGCMwV5B1xlC0ZB+lXMeaPwlxFW
qlUCWN8M/u6j5lQ0lbrXSj5Xfv5b4gdxIx0o5Ir8d9XJ627MFfwVkMY7XNDOlg1LOm9FN4pe69br
Chgi6gobodOYdOYknjDciq36WTOj0vXO0U8mStqDTEwjtDdFPtOweykYuShp9UAQMHo8oRTu1Htm
30ZKmKg2etpzrvZf2Af6OHD2y+N7LHyfchiqSrDmoo5BzQStYsFdjMz392k6RSVDxySgsRMRskBm
COQG653j/d3BC/gZQn3j31a0r0J8zrd3o2Xa8XRsMxEqhAaXFKFuYGJpr4OojIhBiym0Lp0oM8pR
s65mLYjRLiDfXkuXrhjIpkS15BKHO0RpN52j1C6UBTPnYdYedgQtp79An1hTqiCxbho8qMkvQqCD
p+P4C5SK++QLKHloT+m5cSZybdEgp2ZE2OA8AcoCP4j1Oge4B5BJIWc5m+hb3DtV8geDTRzSXVfD
M4t3xIy3FgGbSBmC0rpIXTGuyKSkHb+HFhmHH8ZTS8uUPBjSb07bECDzh5Qna1VaXIdFQzD1qXMm
Mzzd2dfyX2ty+I5wyrp9Jv0Yc6tfIhf/9QvI9Kkph8mGvxivMrloS9J1AwSuwgz7ZdTz0ksth6lx
SuSOTSicrmvPsd9fT8R6jbplAqHIPzERfNh9TmJKHtro3W4zYqZ11j72jAM5J1ItnnoaEyzYrCSw
GKAMlxtl5Qj+Mu4RB5w0ea9jSjqk+LIK8xfBSyRDQLi5KI3FWnqgid6zUHk/NrF0IzZllf5s3E5V
8LdFUNlmiA6ZWZj9DpPD5PPF9uE3am3wqcDminxXB7vHrrmLKNPwuUxmmSeduwh1W/hRp9/KvJu/
vHJybaRPAXzTkIaHOdtU4PugzdN8R67etvdrWWhOWKlQFZb68mtmOeCMC/AUEezjIw4MctcoADrQ
N63JaW40ccs1BJx7pCpbNYtyTKUeyu7r3YVmbFJPs8FbWWCWJV0Z91lMKKdpP7WVOR0j0rf4sDjH
XAmeu/m7D7V3961Mna4ZUZfZcJPcqcS4/NXELELE+coi1EkCv/v7haYUY8f76/GdT8ix6cuaP0Bt
EJQnDB4oUZe9kn0gXrMjecKESZUIRA5I+xsFOLnzWVztdr5LtW5WCugFpQkYBwRK1vag3Q7YeC9O
ZPr03mCfoV4M8542uRvFAXXMLWny5xVBGiXDWqq9iCMJK9v1C6ISexqyIbm/wZDA34l4Nac3+ckG
CSkEV6VYelAjYp3QRkXShpapzt8fTPXGibsjf20I2zoQi6ph5ptiKl3Hc+LhVAABCiQyM/mwr5td
ZAmsth8HeN2Zt4k9qLrx4pj9rki7h5F0pXgAHBS+bkKaernZj25MDP1S5gkwzUZBXkqJ1ZCYZx01
v5NmAFPRCODIbnxfOjphgkQBtTj2alMywGIWXkksX/DLEBL8TOkiradc6ZO1d1CTBIG59md+f/BB
NAAAcrzGUM+T6Pc7lXBp8gZQlA1PwiCYXdQQmCckvXx+UOyqKDqyUYm6eZzDWpwcaBahtyzpVxr9
PWhltK45jWgtI9Vjh6yX7O+2iFDkfQf5yvAve1MFdKRagsAe+qES8kAuXCW7ADMk064cU9elq69s
T5fmX5n/uZv0otqzo+jgSyl3wGmLgyPnS5pzY+zcuyr7iW8dMu7WMukFIyeZn14ykQB06C23UOuC
o9ei3XXBblY2ppFaWJDLMV1kDp32Ms1atbubFtpeMh5HAYKxULyj3FQvBIerhssR3dm+J96ev6jv
La7qb3UnipZlc6CyOSYRRlNgmiVb3t2sclsDQyGMsv3irNDy4ZtH639tjMjakpYIuDjwFXw0pOFQ
w20ceMXAGaYtBJZnutEhrskCTgMQicoWE2AOHG+/8qbR/NrhDjl+f32XPAWBYmr192lDZ65y8iak
LQdlhUszUVM0rEqMNOregNA6xwp3rSDa4AKSa2vc5SiQ0S+LPtz41uXp3v6g+8t9j3/P+DYO/Zwg
pkmw4ds4HG+JtEyj2gfX+O1fCASUXmZxXM14K7Ej1mlF29WPeoxuDVSyqJ4iOszL+yC0BxzEjl2H
CItE3y4Y/yxZuHxpPgxwicH0nRvfLwYUl/GhYyA4BrfZctVJa+KNhSFho87TLTN+EQqR5sT284/Q
ohLCRstxp5Ir7Gl/bk/Z+E6ERPhmfpf/548JnaktWRHYb4q/BYNyjfB3RlVR+mMy1OyEv47OnK2x
5CPy45WaCboqz1oiwjErenDiiZiuY/l8zdZAnFi4Hckip0JnDE+HIsd6iPF2SVls+x3cwmtqfjly
Hqfl2DwKsvQCW6w+DglenjYLJ7X/EianeviZvMBC+qfKEdBpcyDz0NLRqWKwy0hRVBAj3JlsScKC
oIEyIN9q8pSq41pV5DKwZICMBSAu96fxwEhbo/oNAuI9a0OYIvKfn3PRU5Mwea8cGKJkA4QRJsFi
AWIic7jQKVkTKK9ed4U2BhrrQCMfYTikigGwkgfZOr6MNq3K2ItkMQjZzBpY2HHKVMjanEjCdwDO
3aiemAfLigrz2/vNSqB+tzRRSv2HhK49iW8ze8YM9fKaOMfDHYGA17y7/TOjrGmUlJFJ5xNvqSWb
NnHzBsXVubY9J0TTiq3SBZSJcutOmlSJbT/1riC2rwBbW2+hfZS9M/5OGC0Lc97IEmamL2d45Gya
9shqTXnq5V1xN/CHMav9k3H3vu8TLncgk3bruG8/99349HIYddzcTz62igQfCTWRSNhxvNqX7nLh
F6rS7BH0CZW+c6J5YW0KgFcgj8VnyTD2MzZtWqKAehY3uTjVllBoX6NEVhFabMWB0TWoDtI115Zy
zYu4CRwHWdnfo86F9WvIQ9ur8qnV+3lQtzxqiq6NshiW556QvDMUYt/G7OoJqEaDpPzeteWdV39w
Ilc4RxIdRpaq8paWzUiIrsoYlJDMFv4250CWCpd3Sc5wdFGrmzFBVucKJnqSKP8BULNxKLxAQrNq
vCImgItspbPkNQP+U1n1eK7yBej9+xDaknz0LB/PXsyTN3NZcRgsdgU377fLVWzai8lt/j5ry1Ju
mxdy5bGzpgT3DuC1edzmGI1thAXTW8413HQCn21AkjQK+M15cxwGWn5QmRM0wXgVXwJKFb9LO2If
sUbfVVhAARHCiBrRPQHc2nnR35p22rSKFdVEx2/2AgdrDk6xtctDBOA6pmqJLo2sKs8gghIEw5Ri
Pd0Xkfs3gnYMHxAyd2RXZQNNp8GIMnZTi35pLAqcGYhTIkVv/QyTEG9ukgQhH1uC7RlYeazCnqmI
N1zlsE3nSJ3zXEqDKZBA/eg4JCxmkDb9ZyAIYGbvDg9x5kyIsXN17kn9buDvHD4Nnbbog0cGW5vV
IjPxMTxvpljND0+FnYzR1AhuwCdKRNuvmhk3FDbga+BXJRbYMGP+Qz43tUlVOBNdW/a2TRrO8lI4
85tCiXfbITRvoET0BWEianhbKzU1uTlbD7EkumGJMHOHrmbrrP+SfdntUFkQZ+UictbNDNw8njdh
nOI4AY8ry/xNzzP9jh0faseNBxcSX/QEj6i9tSxY/zlCgfULPtahy421qt+t7vQ5liezkmNnrgT+
1qCIXrkUEqOliNdRuGJ09nWPIicdAyo0Fj0E/98azYJbZ5KNh07wM3g9OiblI31kNUdX/QH0ecxn
OiVl3l7x4s908Kqdur82n7sTKRssCma98FA44usw36Gv/gM0Q29wKOveTeUeo1PqMkjHa1/sj7DJ
YNXWqq2rkss5lbj1Q9Z5HU4NIjFmnOfc2lm37ynYrteP/XeeY++++h7D7//N5f8S3hEDF3VYaAUa
XIsICMs3FNril5XuPK6wycB+QO4zLXR3m0kUETlqTERmSyGUib/eJSGK6KPtQ1dJf9St5TYzp/4Y
iT5XNJAZiwEQwIXVBOsLLWd3YgP0BwmpTIO6m4rMaZoRlutNboExt68DynuThOEzlg912LGqd04a
Qohre8SaLe3lgkTOzUdsFw4prg7/P4wgqhAIEvaL0StwJgLe1Rp2gwTKGpQ0laIyxzjsxL7aibYz
cFjJqtOvbb1D3z5G6m5SXrKhQB+aT8+q82dI8NptpcDIMYAplf0VGQh/1XWWDAXm8lQPXDkn53rT
UveXgjpmVK9yh9SFy+QVArN458qds5kSc+8kKduuZr5XlC9JMmebANn3Cxw5jBfmdex7ril+DWMp
VGjew4KAjsKyior/NfaXpnwPI397b30T3uJYkOmaJ0mhoQWbQ+FUER+DWSnisPYuH6QqnxVDhfk/
r9yQ9zoUF+/vuUsspdAqxtJY3vf5ROLq6PIhy6l4GtSexM37GeaHw3I5mrM887pqnpQ+b5WxvD6b
0vKAVG4Ay5u8igxLs9ZOvB+pDg0LPRyqpjZIADSuR3qhE1n96tSeZIAgDcREk5Ukgfa2WcQTYEeA
lJ78b7a6Ex55pjiaqR5ISC7A1iJwJz2ixX94wKMTCKspfl5vceB1MkRLsyrR7zQTOp2CZ+5FfXkN
s6gBnibLghbPCVlFVjbbqaGjeF0A7ujNm3VrQ1Y90+3robuGCjX8aGlz54Q5u4r8i600Nk3YRMOK
vh9RvrljaADD8kT4YSS6p6vH4c21CSS6e3Zfkzqd1g6fBygIKCBpInAYM36E6JBNQqVsmw0fcR/b
qn7zM9kqxKVnUh6O8xhrTFLuxoCbDi4l7mr64lUqoN1qil2s+IEtv8uu3v56MbdSm6ilDp3fBdhG
HMNzBp9pg0oNihkIuBImVe5XNOdGi2CLXSQzdRXhTog6mYrWzTThSO+QHfVBiFSntRwZ9VM7XYyy
aOaGnCf0EOWyeAHlz+K2IAclO4BmSAAtf7pmrZUq0JQ7UDEfovg2N/yowjCZDGwgdmDDbXcaiGi3
Huzc5u8EdHIBMFRGRc54HskWhtcGqaqlz+OalAE41LiWPveu45twexrJ5M0kN7D20iClq8CtWSay
W/i4D4e+uiHNrLmfOZFg3ZXIdtsHTd9DCS7B3C8/fR6EqRsy7GEHqga9GfqYvBieDkTEfDG+PoWg
PidwBFOMWESIhGCU67ubZFnQRiUEh61yuOunJG+5XkuSPHbk3KWpshOPnbW1CIHWWDewBhaUVzD6
lBrdCBs3azBeQeLeESOvtEHqFZAoWsTz9zcZu5orIv2wLsoWDcWgmQrlEcRoiszV5HhQpAMOwSWZ
+oEaC1M3NzVBrw6EdFMyFdZfa+tjs5dEtfMa1skeFDhbu3+xVmbM++lRDpe2jRP/PjJzqyUNBL3t
zaX7i25HXxLP/ySOynrQLxNnB5PTmeT27NR9I+HtObWZMHGoAjjwCBw4/KRrgBFg+9UKsv9g1jAD
nI+dAaHz3/8cK5vai4PDmuwIFdR8fw3ToVcIL3hl1YeSaqaO+PL19PxRL6f2MvmCTQSiEBGKJopK
beQZwkR18Ua4DSFqRZ6b4JCbBat/3tNb2oBLywDhsWoMO9xggylGnIHvYbsHVzSLap74CvpB46hq
I/sBNhduqJIduVEdmy9vXddUnfmwXbYi/DWvfB1SsLYpQb3ruhHoPirocvoYByeO1Pxk1Olp53M+
NKpakWPp+5wpy2fTxcMj83gwcmiCpsAX7PFhmL47zEEOxyFth2KbUTZ+3QGEn41nYOVKu7wWJwV8
l+yRs18Wyf2kSxRuhADSVJ7T36+K0i1L4/2JhfrLgF3zQ5I2f1+4eM7pOS5Z2My/jXuGbGIYXF9u
mAHfGGKALGTU48kSFAevlPBAuXd/W8Qr2EvAAiANAZbtIJrFQMXD/HDVDDYrD3D/diOYA1AFXiwK
aLk0dwIcsLAQyUcvMOZn14A8CfX5SKIPIOJnnyNNa/J4p7cQ/C2x0+ZhIIMhAZlxwUnCpKudvdSI
uCQXDaMw2qWl7vjNux69OpZsLUUnkGzBWyouDUOI1AyBmrmiXICXozIaNWOLU9wVCjx1O5HVEpQV
rpFjiW8uBeMuZDpYTo6OCb5JbekLWrwo/0qkHWLVUFc9AXYnAz5xMSRFigP1wsZ9qwUIFKJx05V3
bNgxipZ28nwaDncfbr9W3KqXz1c+bUI21e0j464SU2WYF6sXrgRlTBKSkuj7v9krhtKcSjwAZO5P
JdFWZfeF1AR40SOURHoURoD0jed4cZ19BVT6utnMtIlFcFzbrbmWPNZDNb26MaEVm2IVq3YP0jzZ
o2TqXxF5VEHWGBDSmVLX7rEJ7oF5LO+rf+fQx3X/K/xNpqLNbmvjZTK5Houl6OevintnAS5JFYp4
JE4FbeSGXLWjyLkd25PCaA4ECmCNEqJP4Omdv99cYqvP5OIkeD3QcKm9VtSUp6Zmp1KfjmLnNaRw
PF6y2BD6sTpIq/aclYV5Y9vMCuDeE6MlgUFDuj/xnbJTjtwz+0V3FQRfNxtTGAOmiTv8KaSf23aD
WMsN2BhFtpab6+zbQRIe01L35zP7Sl2Qh68+YYSeUX5K0VNC/dPc68iIvtoiTrrgc9vDh28XcVy1
iJSj0htYL1mc7y2PUjFuqm19UHxKJQkAyp3wtUMhT1cmW02U3GHqD2eSsMpLMQNMOjUFKLk2YgC0
vzl5ILMPrw6UfXOqH4+r2GzQcXWro0yOmwL3AdQpVXzotkGjSFBoP2m7c/R9Azljrhlanjy893kV
rCFC3drF90yi1ILfgXfltcheSF35H+bBr7S0UwY7l5REOvQ0FPXqA0u4dD5lEsfdF5dAc1y32VyQ
oDbFEc4sgeGynwcM4x4T8zOrFcOl/TNrHxlSozkiE7MkXG1Z03EiCFAfu5779bbR2zzcLtFf06Lp
WFeF1T7DhKrMom+/is9ILpI6d9k9D6BDv5xOAHmpIK/qfeGpEt/yYpZYg2siJEV4P9gXpKO3p4cr
WluTyEsJBYGqr20k6v6BVcLGKRLNWavXDIqpqns0yXQSnS09IzTZU+FZIo11IVlRey583ES/ZEEN
Fpzhs5LAiqyd/R8ZD3Z1t+u+0u3EnUyUdNEQlB+UEBHRuY3X2cDQRwP5pCC+vtBUcWRQVNZdKoCa
t+XDECyUYU2Q56/FDrFD/CaG/2OtEG0F9gh5XMkX8dM6svYXjYKlemPXch8SZz1q9wFzsfxmzft4
IJlJCEaZ+s5WNBXMLt+iPRFz4tGgeWenrsfETehLcRl8diaAhHFV1r24FUnVp3GKI0veQb8d8j1g
KVQg37bAMvTm/c/voYuH3zn3yQQh+7zBMozE5iwcXqvw+BwAIR49URodV2TycMYQ+l0HE74c2eNi
69t/q28IVsmR8CbnlfySxhxqnr+oQ3eG+g8ekf25XG4Re0+/cBO+TxB/tGDRMCg0JXhIuRWWE+Fj
M6kVln6ls1uvhgaSxVs+Q8P428dyAg3vF4JNO0JEXWk/dACAAapBLusYQeuRy/qu492ypn+2UoHL
IMtKa3e3bDo/DByGHa380Zk3yGElpGhCRQZZctlCtiKcFLOy5s4E3UT7yCaqGH+obxfGwY7gC+8y
lHpvgNfkm8zd43XU6E7JbtrDeJTpl1aA4ARluOxuFe1yZnVRvIv07ZDWhRHCDThHPw5/5oEHmOER
u+Mx1+yn79LBVsvu+QG6ApN0ao9b7gxiJm//cdlL/ZgBhustiyn71jzEJo30tmJW6im5EflMi6ws
hWCLF+6sosiDCb2aEI3hb2+/oiJSYePEV/QJ2LyNENXfbbRleQaVhYr6U+b5SCs/87yCuUrsfEuL
mqwi6WFuyhuX/EugtSjx9cXDGK/NOs1QwDPRqv8Lh/EeIPZXN/qecMnr7qrIRoX9QNv0KxGpKOdC
W3ZgBPGNasniIXk1D6IrcS0oFkzCR7jW6N2lAzJ2W6YPIaLdEQxW4Faz1I2nGNvi5GX1zc4ijLQL
pHCt0We/lZjcWDxaAJvdyMH23ZrKRQNqaT9X5zusRuvh3Fl3fTnsQgl7BLMFrn+lGMVm16nrVSZF
1SjTxCrpmAxBpS4bgEge3ehUSx+ucbhPSjfoFMh57NXHIFNLPwyE/G0a+O9Vpkgs9wybCEuNdxrZ
YDEft3kmlV4sl8n3jIj0kw3jTq7GHmV1DbBppFvzyobmjDhcwfSrF0vOkjjV/xZlFdDQ//dgkGHm
VYe9dw4MWt8A3KtNkwYQ9RTjc4+3zadIrTC5ChYczZgdeb+4GnJ5r5DXqMCoVDzNWjlnY6MyqcQ1
UEs7kMbUDopvI9NPVpYKtVws1CWAN9yBi7ktpYvlaboT/cJCb+fkue96/piNHmfASGnHGzrVaCLs
B0bPoU1rGgTEfugDHtn18IbKpSwMTXOI/mCgXr3YkHY5vi5ZPeGAxEzD5Vie9vp7dR0oy2eqCReI
KkbSf1h+tEyZKrJs8BmSwWBrlTmPECGtFXAoNkm/bCetsjVKpE8GKI/wGO+u7C9+Ea/HIru37/5Y
O8GYMWLAYDhtPY7iKueEy2Y/4B/aHq5whLhY/Wwn9c9tfZHa+8kErFcTa6CZxSHl+YYzpIX+3NET
jyubpgFE41lrJv6DWNeSc6P+EzW29Ws7kgjOdYdwpB0GnMiZSovT7Om0uY8mpjNF2WrnXRi5h5j4
FiOeYXLna+dDDbf3OanWEc1jdxGg+bQVhPQ68oH85uOd7/ilgDmNrOVh1JNOAmTYNKky0bDcsxjH
ej7rVjU4LE9Ri00M0hVRdAYDdmFtwrr3GGf6P0UXs4blh8R2jkAg5xqIDG7DIQo3R/QhmqhZHLhu
hFncXFSu4JdlYWfi1DNi5Hk1aPWjdhIaAwVsxyPQovFUWpvhfv9nDcm0D/Vk3xdc7TmGRQyNnxkt
nD0jP87+D2y6lfJMse0X8E+bw7uaxoWCv8aKSAA8mXDWtwaJpWrMYp1GXQiHITCAbWmpEAjBX42e
feMNCg2HiTq1AcloSbIr60MW2eKrT2p47HlZmrVeP1j+qKyu6H/CK2k+m46Vg7CEQ4PRjsSF7C6/
sx2+rXiz/+SqKXpFsunnmbGyrFjgp8s8jlT4OG29OXJQ9RMretclonkGp1dNaJ/GDSXrmC9q9o+U
hAF/PMw+2TmOx71LSXyM6f7imnMEfL4RxIX2jgoTT6EoxrxwNBCaV47IKQk/La5Kplz/QVD0BmLc
DRNLjGLiDYFuhE+n6B1GkK6MwWDam23e7Jzd5uSfkSRRxByekUWFhOG35Hlx0IyGXXzpbI86BOmY
5FnMaHMi5szNZWDLP85YrYoEs4JPi9RerjrstnAcxH0zNkXcj+BSquWUJl7fIwdJ7dtW1hCrK8H3
4DXMLbs2uMrx4epoMHF+a/27asujfzWs2ayrNFFKO0T6c/z/BeaM7H73zE8M+PlIMLAPUAxspJsK
m5C2WVPgKq7k8L6WxXlQn2g2SyCyqIy+6zwjtzj+aYoV+Synr72r4KPjWl7EVGBX2zrJnfuyLIQg
V2+z4PROKteoRl3xGTVmOx7PvUMSF/kJRLEUEP4ADpGelmEIq+nnNShMW0LhBOWgtzcJXrbTF9Ly
YaRBxI5q3D+gxNTf47oD93sEL3uSNWD2ZcL5jFQncqvUfwXZuKywZ3BcHAxVU+mTURtEln2ZTB6y
LuzOLGFNVhoBUtE0ZcPwW2ozloG/jxDfoDbOL/XYvZ8XyZQStw6ZClGtQbWdVQ8bNnrTOUUnMaE5
4cZ/8cSEQulMg+r2Sgzh693xO6Chw9ZJu4QSW//9dNxQBDrixAsuqVQO0q9KExj7145LygApTIuw
cKGWmS1BsthFoBj1rmfsDDP4UoInICPJoy3w20H+XW1x2lKQPRenFzC44LbwXjqHJcK6+dPr6a5d
rEgZYTD5O42otj82TexeSuKT/DP2Yzytpdu5UY513KLi3IYvuCKFjibaaZX+kWOCW45L1hKsQxnN
e8vlpUat2VcUhutYMBNvJoQ+gUz8E/j1KX2KUN0UcgFJ6bG3HCFFvIGc4I9wAZvLvCU5GMg4lUAN
21HEQmHS6MQ74LaBw/08XZkhdBs0kl3pvHZJ5aNfwrJpd0CaAvbK7dNQ2KfU3kuJFekBT1h27Gdd
B5j6pxISy8og3xxEJ+xzcT+ggWHjL3QoC6Xwl1NYoFwwFRvD0hjY72IDrHzzhfsdd5OaHCzokhS2
kdJWsi9jy6JxHsRWscaJN6tY+Ge6OyJEiW0ioGrAoj7r5j4L92diBq50gv8EGNPoDq03c2iNue47
WSf9tu1QDghNnAdeRs4xdYuLZcNjS0J3zNO/UsP/4fQKQ5aeebLOFNHvGt1P9fek9WqHv3uTKUBq
36XeBHus9PWJve3rJ7d2NRXOSuzQBWFlheAyhWDYx5tCSiUNh62VEL6N8eaLsDMGMmbvn5wJstHP
5IlTt0fRRByo2Js5RhdoSbq59Gn/eL9rr2x2Lq9oECKxGtz3x6wHI36tCYDJimX9MzPWb0FYrtRr
ZKw/YOXIIzQDEO6geoaPvf5dY5KtgdVLvXhQp9ltRpXMFAusyG1+qYapXCsYSpX5Qt14O9cOYc7n
xXVkVHlsc5rccPb9b1VJiey8ZCG9JRSa8grz6z/1xT3fv9yd5fzkDMiM2jHiYgQ8axwsTTOYNKLk
vdZRD6X9c/lGe6AE1Zy0xUJ3Em/nbvdWRJSfQvf868IJlAe2zvnCSr+3P2t23GeNcpyEXo7DWDVI
oMN+gxkdQuDA/nT0GgYga78Iic/6qF9dkQgNGcJO1+ufg30VHYbwhrylZr0mG5KilnWdRKyd/8sU
aiggbDDEtUvOpFEkdbKGrioVp1t4khcuW70vz5bAwdpzXLhE/aq0GGjqwsQ2N6Pp7OYhxEC90Mt+
Teihn9rxp9OqkmtM6eBLOi9TXUoZYNlsMS4RBinanNRo1UIMTtc2iRQDkYbxzjMWfKVNbzv0JsJp
0F3l1XHIauktPh4wUcuPk2XdGfbm6XwIMBFvgBujO56WOQ1ZCiohxTdHa40QNOFjuvfwy8vwrzH7
M9XepybsMkhIi/TMV7gTdnC4ykQhCTkGzg6EraNGuPEISuKcRy5VIhrXz3WSyQGHKeIvUWl9hOYJ
AzeW1RG9LufVzs/R2+GT0Vfz0eMj3/hnL22VIPleUtKX3QckRZJ9wmpjbz+wlPRlpZDZ2aNQzXfQ
ehanHH6jZyt9M3F/ez2eWfVeu7TPmLqwuV6NvWrD+90b441uQmSiDYDLOBTRx2nqL0avxmPWZHJ4
/WzlJH8ro6ZKriSr/aFMwazM5yN7YEt4XveJFwCzbaKGBaKDmGPdFTiafm1LDtuMG5TMKYZcaeDV
19ZGP8R83XhgE7KhkuZA61ScwmkTA6+V1vZYXlLlZiYFqeyRqt6dSmVmy59NcotinS36hqWQmASy
RLhF/sn1EzmZ9R5bBswSiALUThSsDVkZtPgMwMe9kw4pcmXCwL5aA+YJBirKz6TWxsmaqjoUn+H1
+LUSb18+xogXxLy7tcaVdxUrU2UdquuJyIOsRkV0zIkAsniewhvTrah4jDtoUPjiTQVy2URUa2qT
GZNXRup7G3Rf57lwkIvhcEBaIS5TjEhPCgsZnmsjKKrWJ9a2IwOIBdskZTop8/T+2HRhKjfkxAGa
e3Hvh7d3ETvCFzRRzsxHko2t8yGMjzMztyJlW58jwrZDM6qjWJLSNi9krU0g1NZ7ZKmS+Mlw5gz6
ML53HGahYOkGHF/WchKcbks81ye76RtAr9/csDIroMIEfGG2KCDEauL21lCHrPt++RbAa8afLV/f
VYh7ulud+9vdutea1X2nmOaB9mSD4rkYpPr8OlbaTCDMPypFgvAgbcWbxKHzMGr+NYgHHW8ZYP3R
czyeUUIS5ZAwMP9mOOG7XvC9bEH6jncLfLlGy1qimdC/SUsoUBq+bXlvzHm41WuSUAR8I/90MpAV
WHter8FE36qm5kiRb56uSPlID9Fmd6A1dq+J+Pe8/xWEEsjzJmuYLv7d+uJxyKdIkJWApQSiinTq
dFi5VdehmaKRcg4skq6e2bCjJLvcUqKYWXVexuTS7DjBs+SZ/OImfQ5rkZ2y4oH4WhRUsJbsroly
FCf5wBV8goJ60weSEAU/MFqm2w2B8oZMU+xN25vTlJvtNXq1sVJprm3ymtKKZyGqcDwjag2WPTsZ
3MiZXvK09EpDbjow+11k5xXr7RUEu36wXdyhqoEaaOAbFAwbtdZ7uYve2LPgmrYjguzFn5iCjdBs
BEvk/04bc4YrktfVYLiFguRScgZ+vDwR0gXnJhwyC780PfeFLR3a2/Hu9QSt6YZGfkFKLO7vxApC
BYrppILDPJI5/d2d5nCN5mYjqn1G5WENH8DNgFJXwyzg57TUGqxBgJkVbuEQy2TAs5rlOSaE4WQ+
TivAuiOnkLLeyq5GwgW7fKRHDEnzkzFrcrxFJfKQUtCzwEh1WXii9WWETL+tyZbGezj5PATCSpyD
QmxcwPwszVRXjtipYrpiw4RTOCPgf0IHbVY/5wMR3w2Bd/u5qCS7noj3RwW+eCwqBReaJt5KTZLQ
ygaSo1kzcGBMV1YcpI2W1qI+Bx6ACGgNypFRHQeWkUjBwnYt26ISUr4DxpBNvtypLz6To+VCn81j
lKtd10FzosswUxLX6FRq97nS9PyjOp2fCYylxBEAmu+8Cd1QnBVIW4pdfSTx8ZjrplHPRaENStDg
jT+fetqR16A2jvfOnUxWmHiSYqAUDpvRu+bSyO4GchaAATx1wczWVYooX4jS+CSyublMxuYETWrq
oFfjuUHl0M3ry2IBlMdeVSXhDbg5xiciXdWXP2kTLsJtlWkMrTDBp3B3VfLpdPI2ddY49euVRZgN
HTcVPogx1W7oBkBDMl8rse+ShJm7G4bEoGEdn8B8VlKnE0qC8xfdpkVxnxh6usf7K2GTdiPrFPEm
equXOLLJHHKcZG6KYW2wipaoQ5tIJSXJ4OFCuekEmPxIB0WR9W2zvkN4/u51OCVC5f8GouNye+lp
M1yJBIe3OywuslYKj/16hTvX6dTA+23GP1tQmaFjDrWwiDBNoH4Aany5CtupHME7lqsCCAwTdgeF
+OlGQhiQVD4rrEiUwLeORNhgEAHMaolDJGxG/tAW3Mp+IQAviUbHXesBXR9U6W3MtF5v4pkrW3Ek
Mehhle2mze67lIYXB87nMJcxkjPmyoKZZaRpi/JepiVqdtWW6ahV9BR2qgVZbOe8NWOxux22cqfj
2vDaXQcgzeW41J7D1tniTGsobP/aRZlewRUhbScmUDJvrdMA7SpxrMwxt8yu8MSsZU8Xm+z435ZF
WsvJmTSK26Ga2/wa6CYucfMJs1t+ZoQRlu7cBEC9RO3J5omSpIh1y6ko9fPAZM7QhDjm4M1spFO1
ioVaZ0+FrQoZhu7mwX7vwzDY+e6GcdM5RPGfocxB+KYMlqbxqPYalzScx5LlOOP9mpV1qs6+Ysl5
4wEjPEefGNKtefGeHDUBgL3chrhrziDFldq2U8wNk0L8YE0beg0cYDCiUlQLF70YRkJ7RBwscMYl
5SVf8tlUEOEWmB1USP3SMR0NqIjHnzezcCISVCbGmUNsJHhtpDmufnfRhxs4ef4CjgGHzEdfoSYf
H2D076eOoOgpoke10l7oS0sD8Yv659y+euzFC0UAnhafeBo82FUrPx0SCLlzxG2mSf4+IJDkc6K7
5WHtRY1Dsep+xB+8Q/HiW+s2T84vnh8waO7ZD01GqbTYBuV2p+N2wRLKJ8hz5+veRW8DpM2w7F88
cQGEt8f5ZJol5/4fNbkiKbyJC+TRXisLNwiLY+1CFg9UqHouMWfHPv+sPXgcQjnaTMIOUAuQ1eTh
aAXnpXeolW/x5diDRlFj/IBWy0eeGlquuBfPXJQgO7bPEXcgR6aAIaeObDnQxvw2N5mxMymN/Dx8
QWN7IaOovoGSOvWLANdrP9z6otrd7smC0mHRdGwc3wFVT1C6Ggy0Cgdvy3p/zoqFTcVj/jDr9Yjc
YDmUI8O0jfjkTbMDAiPS9w9z0tT/Yq1Jlw8U92VGYZRBcgq3cMqw4NV/25tDHogcupTXOX1Aw0e/
C+a6BBJ9qD6NvrQ140nBNWsODZaYICmkg7Ay89JY8PPhIIEvBb+wmcKFtsC1V0ODUm+3ZWtOKzzn
Q9D5U4Hczj9Pji78y5DQkI+KjRvXvYP6e8nkD7cWyyNhmuqq14EV19+o9uqw06w7rd9BoyB9cvCx
XRlzdKaFTGVRJfxQnCGqVxJEMuME0agyZKzsBtSB2mTYCdJFhlKora8xzgepdMNz9vVdBUQey+Mq
UXzfsCv7Hbu2VQ6Jz7GBoHEaBpHfPMKF//YLr4HY0TtINoTh3DTE5qBrj8IoqIKEhFtC+2K7gxce
9L+yBBXlcVZKqqS8ria/dVVqE5rt7Rme94N3o8yyxt5xXUSv6E4bQTiiJdUiSCeNfXZNNOOKvEIO
4DuvuOPNyBhAmkbKzzncslS4S7VIrjyE91j+uTu9fUnuIZ/ufVs8tetb0eSnn/WBALfLgxL/a1s8
/f8SE1iqotpwYGxiX4IZoMTI3qRkqVGZz8M3XP8Mc7X9+WJomZMsGF2KdPbGExTc23i45MV+1EUv
h/0+aiXtqXLsALZX4bJ+chLmR6o//ZMpk6KBpDVnko3XUU1e/4DM14H4MyMHOkYQDzGVyw23MAT2
vohSc6MGfkUrt4oGwN5teo3v20bXPJxm6O0sY12uxSBW5y5VZeN8ctcyusdFcxVXKGRbarFW5Ig3
Y9+7efi+Dk5m0y0CHOWIClX9yQe+g3PPEiZh0P0vpQ5Ef3yfJpL+zCoAIaaggrHpoYbV4RtjEewP
aPnBVIE2/hblZ9CGmGMVrlH/7xAVadbTGMuK5valWDAL57LSSgbqULgyS412XdakFp+6Z25hJoyu
EZHy7g7TGcReh5btArtWDt7PJcEYXw5fwboqrTheqxtAy61OWnhzHp5uRBlrG9PHuVrr7cQ4NYcP
fuEHc+VDoiyV0BTy4SQDxRUhtUKV+W+0aTisK+MfRyZ2K6jrFWlZsRFldk5T/Sab8SOaVlbsnSq1
u7v1DFtwoJuJO4zvvE52JJrK5JlSVqr0uOGG6HatT7MFWyllnbU9tj9RfYhrv4p7Tgk7jSY170bE
EHCpaYCKIT1ZO0Owy++iodyMZwTef5yGIRKDvRUibWujPIoFyCE7TMlGyNwit4O8JC+N/RZxacy/
m9x7LzWNHFTMGkqaT6tdnWrfASLgJYokl+t0oQx0H7UJzieLsRY2roGbj421B82Sbz4HD6ue18f6
Jp5LXYtF/MDtw+E0gVJYkrGcAwpZBBku1WV9ZtImXZMTF/4GL8QuMMuBnlaSAsNhnylsIR6gpE32
jA54EF8pBUHcSKh425wwZgF3Y5Gb8q6kmNV7BQbeWqTUB+HMb/ouX5IXLwxYCNANLEUB1pDe6RgW
zJCLFdkhgkevaIwzY2zDjYcoIhTJdTKF+IhmtCpGvN0/KtIo3ZUTsufXYIyXHelXTcCDtJaCtQUb
hcX4S6ppqCpX+1iD1REjYgHeRrs/QZsd2Z+NPiOzTCIgvXYmYtslvPUbkKKhv51Je9IpUjpVtdpR
QsOt30QXdUUK+iHbUqkrDi4Ko0uWeFDkFMFaaZN3cxo4XyI4TYqiNJjWzUOtIB9a8JrIKAC6OExz
dF23byVMOu1GNLXtihU1hSwfx9MItdOJjk4ME21lYJPSpgKwWbJrqwAEJ1RwhfJlfWRT/YFAoogZ
5uajHdbdWlhVNpGOCiMUuGwo7SvKSbNfbweWWMdAa+tzPBiY8GTrvabnZn4zqy1l/i6Y7Q7ml9je
bt1JsHRRxQEYXROumfHRjw0kbH6E/32R7FYBbNt2y+XhxIlD1gQ98AxeOENUhjeSnaeC69hnBa3Y
8eUKztej5plepqnWIiUMTFRLf9+wxGeDo9Aqf2vsP7vhgMfzArQZ4CYys759wMg+QVmMop/+y4WE
VJK+Yg/PckfSJPur0Vlzft3Zedlqu+ex5R+VnT59jSuUDRhajhomjZIXyixjwyKc3i6eLr/VU12y
TxE8tQtDPBo/KRREoFGER0bC1KIzpQH1QAYIwu7rN1fuIsoidz//anmjcsc8HPuRy+Cw/S0qM0K+
lw5n7czwCgkpX0660YuJafIMI1RcGoHIJe+YVe8DDumRTK3zRJqjZBx+qK1n/aedguZ0IZDWNPeZ
1SAmX/sqLMqrgDBtC0OJUFwzJ0NSSFprNigRJnpQiFZsmNvtpQG36Ts/RYnX4TN+POmB2LwfZgS5
pribZi5tQAYn1CXNEj/B1qa6oFI7ofGnJIsNdZE1j8iOBIAWbYH/4qKL1t0g8++E4V6f4KgGeEAn
bEde+W5hp7QNw8Vf++Oc3mpvuNYdZtPZXzHP+GCJj1EMilzlOq0CNJPfZ54DTD63TyJdPFi4UGzY
An3IqxDXTWOzE+abbpk6c9BOd7zRkc8j+ixn1QjizYxBnqqYwBsPUIKctZ3MMZXzfY8ngf1IrEw1
//6I/rbR278w/0mtgz4ytyHCuOR6wOIi76qFsdXSI9t33vUxAoYQgE3qYChnd6l19Sbi6wIfhbRn
qyYOiw6cclZmbsHZ6ZfdyJhIM8sfgLT1pHUiY0jfMVP97dnt3E8Wf6ov63WJu4TYxAd40gSMNMFa
vMakW4+GfpzNhXQkYu4IC7DKi+BxAUBmYM9HI+bx48b/QbQa12diigdypEVuFT9DqZKmI9uuQqHF
MSjgCpnsg87K8KTODQagFs30vrbKA852cOPFnTtsP+Z2xPqufUPd6arBacF65VYql5q9gpiYVcgJ
XGoxrzrnFJ3opADx5IJm2HLryxiXub2hQ1rXcw9iYRSuHMQl2/wIgn/mpoQLEF1QySKHZPJUgl2z
hGGl/G9Fqdd4/gr4fQph0EcYdIAf92u1MeNXZza7l1aBcK50U+CBkiwIk91eLIfd8CRUjWlfIb77
cR49G82TdkS2rXI5PmB+R0xH69U9xOCcfRgg7URmhJ8AQjIaGLfljgY9IXGbHhPIXdv2VbTlHHxN
Y7VteadTnvTRfNPh5ArnJeVPk+lowv4pbd6eYpLlg9OQk6XW3wdH0TZSZN5RKAUNijqjW179fNXI
b5fPn/RR2zBNrTW02ACEeiETewQYVCj6Wplf9VsbWOo5/EjXXDvi8m4jLRa8MxYdDvT5s+89nbuV
R+F650aUpWhtbSF4NEnsnVEZnppsAKZ1KsHCnHOLXWo67Xe4Fq4JuG9ImPK/Zs/3SzHGaoo8eWIO
1GhvEZ2uzGgCnmwR3eSrI6/fgwc0Gdw/+OqU1EQrh00x3Zauj3nAcP6tipfjYMqWW7cgIhYYRdSe
8Ky20DBcvLzwAHg7pzUOdIr2JShmRx9rqL1EmgofNGR4v3HjhaSii3AZaYJQwZXRo8VGdIg8wNxR
0zqtbsRTwwL0C8sfvI6WQ31hWJfflE/ODJrBFmTE0aEZ7Sl4amT4zQ8uzgWdHzdOfy8WEuLZo8xA
MzmvyObT1a4YRlTu7tzBLoS0cMV3aInauI+4eNaWO6C6iDWTL14sNnkAz0+L2fITaYUNSEXdtN5j
SWv9cuvLRROn4eqEE84SxaIzbObDLWMcrbxFzydoJn+usvs7HxP9ylZBgX5upUW8ShzF4lHOZGJC
oavlRXfPwzuylSjjnaGv6yoBHV8JCd1NpvWp9o85RrJShb/CW8fzzszDVUWKf8B+2l9AND0g/k0A
Sd5BMrlf6ZJi4IXXiClr2LyQmsMW1mMY9rjl4uJ43d6pAhXcgQUNR3x3VH+dd8fGQ6bfUzuHIwct
LbS2/PFa/3mIgU5CpI8HHT9Czj8tibCV9Oat3yh2SR5XOLk1hjiW6k0eGGEmFs+6wU2LL/12KY3J
fDU45fpaMQepje0kTdIQe3QTFflygpbqS+Ae5fUTSj00emVuyNI39bhc1NsZJXZqSP2hViIZSMxz
PL3PGxabkQVLdKmKjaZnup5kkDK7nf6ZaLWsx4MX8L9zAvG2GXdI2uk6mnoILDgypzhlkP97vLtA
E/LaneGqNfYpUOuyMygpzftbmI6Qkk3ptYkSG7oz9JkSvkdoYLRPWju44/r/rHVrbGmQQdiJ4JDG
RNfpkQEavpG3cGI54K1P8gQvFDR0oSp4a9yt4vRBg+jUJUeEvVJJ0wrNuNqrWrhAZyKAICdhQcMg
8s/DyS1BukgMLcgnq1sI8B/z/LT9nscilIzxkRpUaWBWFpDe/AcS9Q//3i4LCHRs/iWJ+WW1322B
z8RCwrhvS30pOQY+M/v5PTP4eJ7i+3srPvr81Nso9yzbLVY5ishx3xoAcHWv0aacWTlR7MN9XCEo
ZNiDxqDEaa2cxjh3MmhGAHdOj91SJO58vUBPaVOs+I0QoQXNW48wKd2WDnGtAkgvCfkznuHzpg4b
ryIyjs3pjJXfkOpbR08YV/7cvcBqcx1V9k2XXTmoZUMYLYSBdifNRSb8yJMYy6vjbMpVlbTRh1L4
UF6qEUYKoYsXHsZGMcYERqkQzFQxPrcSrLfsnlPeSmd6GsMTOBsXF/JOod3q6yhilk8MuU31/BG5
B219fA1l+klVb00j2s/hAAGbmn7kThdbwIJpiTDdvebkwlgRaWsn592N0Gs2sXLJKLAcu8naAtsC
nB2bAx9zyTniHvMpCdviiNy8Vpw+g2ENjBStFlURwxfMfpnH/FLGyeSo7gYMMmkshCncJBmWiSZx
jXoJExtkbwxE5GLT4UMeD4W3O87Yerqecc9XgB3kct1LLf1LRU8Km6+AwT0JL2xPe0YcpvCljq1V
b4ySS3/kgb4jydiOH65ldibb55zxfKRFOU107+haacKNaBVElOcUsCQsWH34rYxycJp/5DSkORoW
82RUBSvfV+MY28owwypuxr1mPN2lxsPmVk9TGHZ3g75pFnfSfN//C+GKiqnpY+nS8Kg5suMahRgm
jzJdrg1tgeqWAm7LWkTfmwBe6uwCwF5R9l+F6wZXfSqHfwVhpfyg4OcYG7OqC8r7LPUElqZLxU8u
R9AM3HUqFu/T93SPgoSYAPP1ob1yNMjAVHJN9uvdreeY1BIxKDHjwyAqn9L0UZtzES0Y5a6qIcAY
C2r6kDU3l2O5tB08gZ0fz+jROG/bQt7QfM0JRrqmMLSLy3thsszT3dc+j+YSNT76A4Tt00PL5wjk
wI2GRv84UH1Bbg+OsynTfYviDB2Bd2nmVrdqleCK78Ng2+Qgx7qzEzMUs8bGqg4yCEbhIXGEuiph
8+S8jiEcEQ8B1Qnf8a+8YULbpg/Vu111Jnw+k5iIRsEGNUXXVM9r9Dzk+hmQi4KKutoJlrQRfBX7
UieTZ+nMhmhNPv4cAirScBg9lCklza/oXOnKNZaGQ0f8cIi2O6Bll9PTKWM7gdkZyL+nVYAIcW6Q
nlBzGOs0QA/oed+AtWjYhoYpkNUMYWP2Ay3jzhnRFZD9nv1lPdaJDdQuvDkta9f6mO/taAcgHn9W
EfDpSmm7Lx7YbeS+CGt4Eh03INoKpB4xBxMZBybXym4CgsNuSw9mOgEgV5PQEVAcxsIMDzrWixhj
qYFKk1X3F/0HNsOaawdzhqeo41ICSgRGwhneUbymtfdnW2pe9JUxSapVGPIlr6OUqJxtPpUgs33z
Apu9iRkGTnln/LzD6tgUi/z24saBgmdTdAzGuxHxWfCwfnSNe4HY5QdU3iWPWC7MhUaS/cO3lNmw
vV5uJptu17dHHLmeMN+OPobQrH6odJokpunfNcLAeru5U39fG0ADEGK+mqWUZM+ucGBZubcE2uvr
LjZArF0U2aRQQnfjRys/g/7QxENZ2r0Fw8wlEOfIQOhFTUc8s7E5crUO70afIL3W6uJ4TFkdyXpQ
1Sq9XnwzoHBKJljgPYnGrgzbSqhoC5X9SIzmlhx7RWxnB0j7tB3UGRngGdvsNMUzmt54wiHIyLK3
uN0K3aZM38Whqq+xvkOnzam9RH4rHiVFG42hfstor3GtRMHM+HDaboHuxq6G8UjSVgqGtAUS4mwN
cUjf8q75p16bO8H6RKApLCRvE82rYRcT/qqPKya5m5Cben3GyDwReh64uRHdnprf7oEJanPwvzb9
qgV2+qE5SoR0SPep8ExZxWC0nauP9krCWlSEet96FEbzDE3T0uYRstLnyNAWjvpTIE9P6f5TMIJt
N5a5MGLtBD6eQ8DPP2GeJGtPsoHXdHZjGSxRwpou75lpf+qhUEAdkNOc+QVqveG9rOdrThs0Z2uy
RiNmQkBFG5Xum0P0kluCaavNIeDQ1AWNTpMH5K/xtmgpuyb3vD6RBfU7GmnRI45EdRQinFO28/WG
4RP17Y7ZhUa7qA4yUOSia9m9Dn7GgoynHlNIJlMeXrvjGG3iw5vIw2Qy+v7fX6Fr+CpQMv2Wo00B
aHA43D3MHAnIpYGvEgKJBUvw+mjKeZ/ZWnGGvq0WZ50ax+GbMJvjYLfE/NHgo4J4uyx6vxoXUBt2
hpycx2HhFWqcj96J4ozbguegSAtHNUZ94Q6WJJIYBq2dW+nl5LOtgaYj3Sz/yV67FDB2/KRNxxHs
7f5PMPj982jlTZ7oDyUjI+1xyo7Ref8u+gAO7K4BELSlGTV5wICDAywI1F3Vp+JFqMn1NMCnNCV/
dVAYdS4SF6p4st3FPlwZRE6UtLR35e5UNFSyWM1i6thGmiJ85fw1KdgR+x/5Wr0PFn/y7SudqnSj
wIHyo50de+lqvUYHG7TXguPTS/rIZop8RlGdAMsA8GPhUJzAkyXTChnKcJdHipB0GqceOrx2t+a5
oJukTc6+b8sAhHDVZUwDp7NYUDZ/7F6AlBf+ZNnoAoZGozQzLc3EOJ80JxlujbKt8SM2epCWDepB
tqNjIBVjQLhSaEB/us9JgAju2LVdoViqPIeWpJcfh9e3saJjOERK7wVC2wbvOZL5SFvLirBin1WZ
ohDpJi39gL/BCa3Rb+wCIXwc92fqEE0w93w2HALcpLCCK6zaRJHh2Ckc2EIUgR5og+AXQM2WtfWq
YOjuygC/HVLdoBVATyxJWbFo4h5qpoGvJc2cwwDxhwFGc3xozFKfy+ul5s77h5InkkUEX9cimLCo
3odqhWXwuexQvow1zvQF2nlTWGvgjpUwO2Z4C0XMN+wyzMs49DcIaTh03Br9kbF7VFbDpp+dV2bu
dl9A1ylcvLrTFYyW3KXMwRmxjZS7gkj1xKq3VQDD73qqEPKyV+SGp8mbY5okbvSi4Ny0s+TvXtpr
D2dW/OUfdO5h0IOECljiLdAGEDDzg6dQOTv0XWN5mDJDzRcHn3SySLdCHw6q8hS17PFA1bBHmJbC
rvkyq6OeTs8Goa8vElPgHg8taPRgaaP6HDzBy8Vyc2kcJ9wmxvxZlkwHb30u5vA0bGGpvWg4MrTa
XSQTelgcF0eYX1PcMZysoFJy/IL3smfFVvIiBunKFUNTbijakNZiTvVZemONI9XsRN5XNtl8E2bM
om5BYRyoYN0oEqlytHt8AhCBE5mjO5dVeJVzoEw++8mhLOEVlM/NCyz+ijTvRQ7km21sTHGhRjRL
I4n2XuO8oxe8qOK+ue5xsioFFshR7UURGRgdEk1H/xnGGuz3YYu9dHI0+R3uKq+zpnUNXpgUKNF2
LuMMJB1vfqyYxdG00t1AaUgGnxDTxrAY8dYOT1l1PkAIYvm7D2RKwa/+RL8Rr4Q17j3WmQrgTqer
hFp02LlX9bEoybpkBN1+qnV1ut9PmPn4YyYLfkUtmoCgqIMyomBJWUrvXQE//yD4BXz6hc8Vwo4O
hsIfrNX7H4k3H1d7vKimPiY4bwdvjz3WdasKGYKGROHdayS8aNy0AViWjmeyDvX8IfLOFtJNqCLY
f9kYgSUnZ2Y51yw3doOu7lvgvkFk2cZUpP1IYXIThLP28mLbnv5dtfhx6iDau7HwmAkedWGseC2W
54Wfl0R37gon1jSW3MgNsG8G+HozDL7SWvYn415oijyCa0ppapyhmoAEve+IAhgvO3pzuZ6lMob8
uP8TznnjRNvYgZLUHZOm+Q0egMrtirTUCHjPdOgfdWH9y/Qfv+3wJO13Bl2oUozH4EGD4n12RJt5
9Uhf8GF2pHEyo37lwra5CHWwyrniGFkZgRMSQVgnxUvkuJW76YaNBbbQQ/AvEhoLYiCPmbLTDtbG
EGPev4JYTCjf7yeYaarg6aH28br5mJaXpvvh/Nfudh8oLcLjk8qsUQCpdLu6IxKK62ziUUeUirLS
hGeX4SZOt6t9jhLr+c2FMRyIf5jAX8bQAv26Azk0pOzTWefSXZ5eubhrjcBrLOCqeE8RqN6SBRno
otVn7QWH8IJWLsAWQPBYwl4OSdAdDcBCLNyePKR0W3FLMS5HJjvVbzNs6saQFVU6zRvT1iCBjhUA
x48Wy48LRhxi/TvIYrSnQZGSsGuMmT3x4RCNVUBh3oiqYtuW4sMnahsx1RfQdsHR3TAhjRrNPdeK
ZDgm6ucmfCA6xrzEMfvT7aL8eeuZoDqFoYLTwczXpSTO7TVdObk5sakMtEMaH48gMUgliNoHNFST
HRak1Yp6quWEPw3eGBslzennY96c8eUDWmXsvoHJI4zKMXBaCsPvYW+qnD9zAO2WTag9nOZ3vAOC
PMfXzxlMS6sIBStG/x+ZYreDNrnRrY6DyoPttNjNj8pu8Got8U3gMOSjNyUL2qZacHdbZ7Fbbtfh
0T922aXrfe7/z4i1BjXfinQkup8kw2xO+EJJRCNDLKP2+eOWkZId4VFBACy2wIuuX9Ww/ik8hbLM
vBvfC8k2uuiB24Zm9PKF/jBiju+2Hcf/tVSXvMP18UKlELRqdcboNEGcdEA0CGXcvJHH6zeRFRWv
stDsMyfCjTSfAUbZm8/YnrLQoWtzxYhgnvjlMBgXbIG7zC8RNxg06g0dt9cCmlDLRdbpUhUjX71b
8+bHvKd8OMyCgRNjx760XK/ZZK1ItS1pMnOgg3UxERBys+VXn4oM7CQP42nR7GzcRDGWpWEUsOfg
r1u68AJlyNm/oB+mHL70SqT578BH2SuDHFwUUnsJ5F661x9WY+vbN38X8E/O/OD+A30kPe/jhwck
tAsURJakONb3XZvDQ3yGPhGUbcYhTjtJNwbrQIEw5etG0g3Uaugc/nl3MHb9CMeGrMM/xkKFJ75C
CBpkw8xiDIa7Td8Nd3efvcIW5FYxeacrbNqO3KN1nr7uZp0RbdRMh984ncByM1msAO9K9WZuF9wH
lFvimV/4SU+iB62uEiwAURxT/3Qezk7dLE8R/h0niH738Bj0hos/Xpdk+DYDkCkTCRZ1F/XwxbWR
DQFIQDDHX4kaPvhg8bAxifW2tPgSTwQpRq1zzkeV9chsOaGgelKTJuy9cNBN2rPC3hFdQvAwDVQ9
dBAwdYaU9HganAjLy+SdalQ9CyJlg3v+F7sy/Zm5oFOb0SZPFSaAi1B7ABlu8tWdFz83EbFfoQzW
SS6UEf9iqFc5DTqhwRxngn2pnXa3AXT2n3ZnPlaBxmEsetT3t5XhIXQSZEJZDxv9r+/Hw3g2nspm
MxPD+3sA5KFOG59y+0iaGZ5b+9d1/OM9BK6WzrwtBjiv/kqU4dHusibG1Db3XZPif06IwT6Gi18E
LXRnBYLzP/+Q4RThN2DJyYEI5xiFAA94+yt0DTAPCOXtLpXoGBUSfgvzWi7XKF8WgChF+U9Ek6ba
1d/xPtt4l60JduTTEmwjdapiskjVIwi1rOesyVM3KGkoeL6kVLWCPZZ4fbZ/hOXF0vk6QCoM49O4
PoLNoxgLMaBLWq+jgOth21qLe50PYCoKba58SKgfoBvE4YPDdubwxIpRUpDMUG92KiMumFVOgUFU
WlZTaqTHLsJatZaJpa4ERF1RZKZLo2Sx0S4r340Vdh4r5IJ5oV3D0CJsZLgXRYwQZyw/RRTDnr+m
MRbWUNT7CJJLD5KZYTSj9m2LOhQVMbd1jXhnJxzyX2DeRyyiUEVIfBKDfDQLFoLTw1uu/t/E5rCB
z4N2d/hjJU+FeasYNe/8/Ab11w1eH+DL+qpKHP5zlGfj3+z/6pRqiD+SGNwjuMOXtBWUswQYCBUR
n5ptfCMCoCc4vmkL/mt04U0+c1PADJWyOHYU2xunDL7RcRZtl39ypyJqrXsSOrp4tKJfozyCwGdV
TMVlva/K5/+xi4/cBZJeIJRKEwHicQ0bqAKXKw53lzFGOmBNGhUAuzEm7vrt9ZHG+58JZYP/vC3V
e/AP7YCH17WznCYo9ORcplJhI8BNj+p4FW/0rQdjMCoabT3Wm5vWqeRhBR3uzs0HbOvq6x+HMdtL
Rx2TtRRN35CbdX3sItpb8DH2QHrwkA6w7ptwcaP/j4eSC+cTrWobsJzRQY6IeUejXvOMqq5ShOZ4
Az4feUijIxCcmXGBZy1f3j91xBvAPPXWoEBUPZr2TS3KeKw3/L9smUuneSZAb47TCRqf8dIkN0Eg
NQvrep8DmaCULk8kHJjiKHdHxV0QFKUJOEQdBgNFlvWGizVj13Uoh+93/ggGz205Xg7aN+xCKTBL
GVyphkjW2FiNZ9gf1Walp+K2QMfdnZcBfU+Rpegjik61iUQFvYjsxBudRgwW4KKNFEyZuU7G9SY7
AkoLJPZxYFe7gC9bZaWD3jvlRs6NyLYFlmHf8EpEQ5jjITxcl2KWhOnOTnSuI3tYSrJ4aq80qPCn
UV0y/F5dnn6x9Q+Nu52PBEVmXknjPKhdTsfPAs10pY5umySEErH9rPRpP6I1wIzD3KXlzkKRsMma
OeN6qh8DY8z6uy+nYHCJ99EKXgl+nqq5NxG5o+z2LUTQR8DmC/1qfSfpVUzF7eh/1lc2Ag/b+K3u
shSm2qdFTsUcVmNDuTuktkEJ5niKp5QnF/Pu22HZ4OBE5Pebva1KDjPZ2aiLtGsyOFSw6kuvrerN
3Gzeq47Nb1I0LWffajmI1cdhO2D9nUVvqihDMw4ZbTAqbK7Cz9xbc3HXjNlk4sYZiWjuzCtFo24s
rP9t/Ua3Eh5tysgMl9M9VzeKvHDCbaMa/imOU21OlW9HmK6cKE+8s0FAXEMRngcnkeo0nZVj77BM
ZUoX/DwGYXxar6JUQrTwx9nQfmjo2gZmK+9tP8LF0BQBtlOfZqJ3EKgoRaykg6jJrkgvXwsSapGp
c0UfhG0CfrL4/zH+hVtpP+D6kLoFFnd0KvGy2/jM+/KurIIScKW+tC4E/ZkqrseE50Gu/CGidHlL
kw3PlZH8+Qzm7UHgIRBfpPgUTcIlGunUzKEyBWDcWuqilRejPuc32x7bAD//mOrIrKBFVUq1oIXJ
3xSGak7tOYWoIl2ffd4Rn6sjlMHexLyAtoEuv5EUuWFKjG469S+CRLBgn0wTOuQ1xX/smEi6CYRE
phervk6U9HihOmELwxLPOA/nAMIpxYOte77BobDLCqlvEZW+wn2rblkya4k0s239PqMvD4K6uLYB
epff6UvTaQNDtflBwG0sXeFVDga6drrF7lb3UG2IJsKvf1NEgiVROBFRONUn/Uce9BE3LQnxI+Hw
HupFWOhahWQQng3BEfM8L/PEqBoaoMPJ1SCxsj4u6e6N/q7a6GTr/WVc1rHtHQQaXp5+0skm26LW
jMRN1GpopcNo4k7g+EU7Y4ub80OIC0wvtAN2KmLLV8nWZ/9ZK+SqLx//5yIBEcMgHt/9ypCbkU+h
J+tee15A/lwuMd3Y8Ky4IcQJfwGCqbP0QVg8o2j93GSfmhL5sv4yburqhCXevLQmWhudE0DNw3/9
1Vgz9TgpKydelgPv5Owl3G4tNmY6e8+f+QXLolPlsWabvYP3ItCbEEGhVwfjIEvxtoWmSTkXTD6Z
mcTvM88vb240XAVjj9TQdr2umkgdvPoAxTMV9CPUslPeGpZ9xa/4HcmS+rUmGQWhAaEiaF5wEbAq
fMcQ+1Qi2lXOS10FyofaIUM5Ju4cDugUZXwTJXe5D8KjQUwlXYrmSSpQYbutSCEpK76R2rCM52XX
CRrPNXTTZPUorQE7GoNOkHYKKvfMoXVmIsTJUL6BkfqTWyBrck628NHfQpgwZlfkfQwmi3dy/HyG
xIdUeNgdxWvVAYpz4l992g2CxvR9NsSKMNb9dgSsRw9gv+bcdBR1jVI/n+XT+LPvAnBxjgHLLT4X
sD5oleHvvB1YAdlVA3ol6G9XeudmzcF5/TW2CvDhpvOylgsIsPzXoMs7VB66xIM7aK3dIgMnyYZ3
klznxxxgdwZq6kqM3mPj4MOkDVTnsmoplknKAFJh4C+wzu/rLdmH1e8dyJZ3IcQGNDmt0LLx3NWO
XwvcAkaQdupZQlzZ3lufzDmmPjw0SzHnnruHCrUc+x9QRDZOlM7q+nMIiKWpRqSnK9AuNVOjeGi3
bkHxL0EsXOlhuq0x/7QRzf55M1jovoUZvJXGO6s+430rCIJo7pqSL1GhkBycaVhai5mwzbC4Ng30
TbSxDpqdMqrl7jWd03z8LHEPcbTstxMWXwyMSTED6WOgJKTnAyWp7TS/abVSXHYop8guv7Z217iX
7cnsdTj1MC8e+O6CAGOyed7IVhJ3d5d0meOPU0nuaU+KCkcacUqDI07LG9jjtIQq5xQahoKT+pQW
tpvXFrob8u1K1bv3eSPydf9YagITJ2NZ/7LgxL5Yf8DxpfZj+NEMWJ19E+Lxb8Z0OjgJ4JpQMnED
H7FVRq02UJXd+rTaNtRhZ6K6VxZdz22i9MGL29v61RaGVTjN4wvs1vl0IaxoIP9qIcXHpHRfc+Ax
20hhfvPzTQ6WpQjQpXiuVH2xrYnJkbEmiL+TJHVKo8DEsWa4M6wCBpPyhx/alQHtCCNBHdfPxshn
13eserPOVNOhYT7KfRknucZ2ZruXB7F0zTH34/M4Hz+dWP5dZKiTF0sn/ZUWUHwgQKuHnrDtoc19
64kwJ9DvxQTqZomrZu5IQbimCuyv8wqON6J5fRW0jFTfpTO2Jjk5MCyIewmVwJZT4Q2GwzSsIwh5
XlPcY2Mo6LXdezotAUpnKZ13aiJyHxvMdeiJhnttFjHlvUyXKPW/HWqUM2qUjHYSRdfSYBzK5Zm+
p7I6vqM/r5EaJG0L1IcpSU3ugQPmdLK7LqSWrkJa3Y73CojzfoBVDpA4lltcnXeTGo+7zhNG6tIG
AbhK94ThCTEYwZkLQyLgxvS9uOYcCfu5g7sdp8c3GlcH3lKr93ViFBgOz5+TA10nmJAajzcEjbkm
caI8PpYqX/sdVuyPK07iaN94BidFyMAL8/dy03/PU7bitHXC/Re9S3jmOjXej34JPCoX/SM8StAR
RA+6j5LzhjsiTDcX+A2df3YmXRJFZHUiFT6rnJQaE84ETqOgZqna1ibPFMFcFyKgNwgZbZRanrPR
bey76jQLEZ4TTd8WoEaI7/+DGdFZ7WxyUZOE4VjU0z0TJtgoU0d1cEctZ+nwbEDon6IUYQW0xn2/
GFkgu0WumZ38M4JbDk4CZYoAbR/Ghm52gsHJ1oeWokxtv4c9hzYM2R4Y6JrFUNR4Fw+4uyPGQpUj
VKhYHxj2SXmLmAayI1uiDL4ntOyJk4xsG469Yqwo6dCcdc1zXNNGhk79kJ4BlnZMMMnnohOenNRT
xKflJNW1anyqWhrN9FJbiGesxMbPvjFUDuytsCa36iDk3dBOGTPhoLtjT98TKpXev3NeTcmDnHLi
rCa4Cg/5adWXB4xmwDJcjR6AGcQjZksLAF2yBn2yZVlxB4k7BYM3GYFwiDOB23UgqzqmfEJrL30e
zv/Oq+b5SZRbFZY5BwKcI4rS/bsVKwEXYSRV5WZfzm49c2jTBUSM/NzBkT0Ksqez+hLOYPppu5Fj
5+9wFl8kMk+XCcd1myUzgw9KzoXzDwNqL74GVW7MMQ3+tr0fpQY103g6Bu1JVOaFKuz6Cs2NMd5Y
0NvfpWW3ssRrJlzrHbdlagEGS0MI2Uag2ZyYTljr4aYWIsqsu3ZuUNSuIbLRZcbwGhHF6dsAEWoP
wdaqBIpVkK8PnTZ8AawebtVppjN1ivbHsUsi1eEbI3nqIJM9GrYTl255t59bkpeyCdN24xuPbzaf
0weag4TJh6vF+70+8M0KIMLHo3x++5dOjyFb8BFzNoUXqPsxHQshh/LMf/+XGcDWgput5+os1YHS
x5yL65CwEx4EKk2fWXNGwo24jKO7XEVXnrmZs10zdZr/1XuxpxxDsbf4NbTqzOxRvUUn9fn4NBE/
ax8LvyJfTUjwn1AjxtM1nus5p0ntDEaNgSslrNsCUf9UwNhSgSXuKPm2S2/j1LNFe1ZLYm/x+rtG
6hYkBn/vN/Y3oWwizKrF7qgVnAIHDJL1IgKqOoYGL1O3usvQMlCqWVBg4CBkRz3bHqfn5aVMkiI4
hjIMhQXSIEqhQ6rinlFo+PPbrAfuyuI/RovwkpBefUtOsDnInC+/uU2xTIJerkWDSo9MlG3/uYc/
mt250BMU6zr9kqS94k03J6iQ7FeXGzbsomrxF4+A2C4bTCeY5zIfzkrlDAK2+EEERpsp4phjSivG
oH7Ddo+vOmP3xz7SuiNcVpMhmOucayK6vC/lM0T0m451jhJKE/NleU993vgHzy39dPNDo0+PNrXK
daYDZVaShFZei+Ezva73s0/Xw4gbPpCwE0LHl/0eT+mE+DVuLfmp5H2S6/WC/8FnNnxK+IBBCHjR
HilL7Vf5kgkiJiloLIWjkXAKIrplM0hsorP9TjbP2Jm6sg//XPnGhZPCFkF9h2vfwYkP2Lh1xxg8
AN1hqNIfiIZEm1pzmE0qnd3e7uNfBWjEsi/cIIB/Lnj4FU9QwTYu21y4Zmy/K9AhdehwOlQrzR3y
qorwL2uXnkEJoxKK960Wtodhj6RsUZrI5JEmc5Vyu0J9zzUkh9+usd5DJMPMueFiywxB9PM/yyRK
OIYzhfGEzMDzzK3RJ2FyHcZgYiha2ioYNNNKPxvNgoT9heX+SVm872gzmL453T4CxhP7f1k8qGRF
KUJ61ZgNPtIRd3W97Gc+LCRHBpk95ETce+mONjHj3MojNZPpm1M520PHyfUeYdxbrubu9AxzGJlM
ZNAvg0dXwVSgYNs8ATYKKbG5BNQrvjtUALzOfl+DKUXlBNAGhw4ZOHs/LjPP+qGVcgn0/9ggh1K6
3wi0PfXpydpcbHoUEm6L+hlLQzHa1XIO+Z37UOJzaL7+XsUDcPZi761s62rtwRS15sz1mJM6CcBI
d3knzB80YZoWXyunu9UEathw3R9hLEuMioh9jPwF2L6YoTpOUFPWQiPj4FARmTvXYszwWlFAcTp7
AqBxQyEWvaf+EXrNogC8bMhN5pRRcMlELVwhljYBQawKVF/n5DECuiQo1+mN5BspgNkYQY7Xy3zf
qVoLVo4nZuOAKy57jnFifW9cTYuJ51RfyogM260MXKvduNfrvGFmMziYUVEX5CdgMR6j5xUOLa7V
2z75hABXX+jtpMle9ogUFlHSi9xrbiS+FOCj/FmQ/rHIX24NtKK8otd5QzuGIWtyKLRgHRjgAeye
na3vNH51EmRojiByjSWqx/YF6/DVrjFhQK8quN4OpR5NTgmoo7h1Uj1Mo5i0WxnYKjxjBql70Ymb
ln8DWURC7LqDA/3md+vsa9HmzPAeYVTZ85qta13M53ikR1aMzzdO27fiUcuJbyT9wBO4TAH+yKgM
eBUO/8mb9muYxW4EbV2x4nAonTQNh3vXMUXs8spBj9Z2IiEU+AVESaumvDkisU+CPjyL0cwEkcng
BOEH4/ejDuN+FgG1mQHN0n6W/C4M2dCQ6usxJ/hUbk9trUmR6f8/7DEhR050h287EhEVGNkHd7CX
uEVjUMuOodrlAZMDt2EIwAkB9ItwE7Yawx3ea9v5aBMQEruZOvfpjXPDrbeOm+pcKSCPUb06/tvi
gbFwjZ1z8lVYKjY8tlMWY5BcbtTrnG/nOnWtYHpRULTwtB76ApR9jIBP0T5xhAltMVN38mfni+9z
ZvvzMk2XGtScMixXwL4nPRLMMzs2eoWpWpbCxzqjy+5e13isXON29Z9bY3FSEPN7ZxWaK4B2TmAu
GDh9iuOPrUyqeGA8/fFZ2HyOkUrokwYNXbM23EY+hko3/jzvuFL8HLVRpf776zkNoPyH8141Puyi
/Nsmvq2f/eLYX2sg5g0CDrWlrP8t9N0hhA7fEk92D/l+wb9we/ltsIFihyNKcC20levQyp16PInR
xP8QJ42xXjcT8Y5AHpenStD3EVg+lMo7LzWzKR4K7KAJLXHhMHokUqNDiSlWRpB2oDPmhB5icXlY
0xrB2DDV0vSb+36V9JYspulTaoJo2UbMSQ5uwTIobsFeNlmmMdKlImq8xXGlY81PreduFDIRdM+7
X9trbfQzOCsWBdkS9vSXU05o+DN7UZf+hLA6Pyb7TEehelnEJsLhhqi6ytSuYVIA2RaF2IZ/JE+3
lAEtY7r3cjnIT36k3YbN4Ffe+SVJenLp8dUBRJzkxE0os5qZMzCWeTQPKbXQCopBUSJMFzEF+dmr
E0jeU3wC+WYAn74bUy9mduTjZcaj/fP8ZB/QTC0ZeEUVAR/3I5G3gbyQJM7NGOPE6vMNhVGeMstt
AMaHckF8EWfVVJCQKzC2rdyszxEHkCG9/6PrJ5K55I6ZXh1m58HCHcTb6d1OJCG3CLoy78AgQqyG
LCimdq3gQ4w1/EwRrtA7oYAxUxipxPjbDDoBPh8Jb9rG/f20kR5PTTHEm1Z0J9pr5i4KzQZ1Hs8M
iRurJUnvnlq2cb9W9FZxUv+RbZzerD1UoYtwoIDs4HI9GV0HU3R4ZpbH+od/7OlbNdF3kiuAY2Tz
a4AVXZkB54uUqFuA6qWONHo2uxtYb5SpaZ7wQAY9TrQTgVjFGuUYU8w7icHuj2NDdpvJoI43PX4L
awtDpRFN5zgBCqQsnXIv1ln9FdEnYianAiFVG45bmtDarbdJy6e97FhCH2ynVY5dnRigM/I8vG9l
LF0kEhFlkYfodskip/OQubfiBmuzVqnoU7Mb7DNLBay8juymDVm44Ph/60M65RFbI95L5GizpoN9
E3hXSgxT12fgmkMqKUtrlj9y+3bU7FSuCQoKh28Nkw9GOIDi9ufl1KHG5qP1Qx18sfTC837LdEyX
Hc54pKvItmnymyAtmOdeEhLwoYcTY/LNKF9q9G5qf2bp+m44xTMJoh8z8K+MUGZOl9vW8LNP5D1e
VY8freS20IwChYSrvzHnFZqzz/JgV3x1fBQDGXi0OChdyMhmjLcRd7jV2aQIPQGas03Qci3yZd6e
RHAluqzU4MwjhyiQvn43kjEJBM6MAT7YPIL51yPxu1ex5c1t1JFTlubsF8+6eAsnhi77miBX5GUY
LCqXB95vvwochXiVPiDTUmGHKhokblSkNV/r54YjmgWSdjh6fp4zsJUPU91PUX2p+i8IftZY9BF7
Yd34PHy23ZX8wCM08xn8nqTZ1qBDCEpbKOsN9AlCbrQTJYLF3Pkvl4gbWsS3i/0hEGRsas2Z2Hyn
6zUQKbq6os96+NmUbYKwh2Bt8bqKNlalFiYz1mw7TXNqxppx6yhC6lnRBAYW/4ehmUvkrtoyhLiN
kzYIoOnWylnurl+U461qoOm6lcj/pnrAJdhlRnmJHqN62npxJiYgtSo20tms3VfDNHN/mQ0QTW9h
6MqtvQLAgA06eRgAs2nWVCSlEMUrtw2XlrmE6EHSRGyXBBX9dieKaw5W1RMAOVUt4EtxNUQAVVhx
QA9b6FAFD47dTD/rYLMAeeObeABCvBM/ADLOmcO91+EQOvEWmhRay7U8N4d3SKfJNZx8mCqbrLSn
5ZcfUcX5U+/jqeS9TzrbFR0WVNHg0gAh77UnozZUvtkOUL+J/gqG3dGsuDjK9jn3fsxkqj4WhayN
1ESUtGpgAQVwfKjUAlfBQptgPb0BZe3GOPxwPojjwnjiQJBqwWPJ8OLHA5GjFawB3gt7zFlQjiLS
KxKtmo2jteKE6LoaWzBVDSDK3TwNsIip5JH4Nqr/RKJR8u7En0S+5r0gvd5Uw6o0fXuS6ZFhsx4R
VLRrqr6ZkYDZYhUkgfi3yPaguewNvTs97XQ0dj4skBG+uQzqNpLp8N5q6tYCYvhLPDFjA+WY/PYa
7Oxr+s83m0DDjyFuWQufLYkTddgYv/itbdFKdm20b4c70e81kbYL1NbbGsxAGHQFeLvF/9Zfujif
um5ftNZ3ShR2wWfDsHPcEr6/I1o6dF7jbl95MD+NctMWnkvnphEnpq2pjzgwww8Y7aRFYd8fkqMa
4pC10DTeomOMEXfPUOK9x/zS0M8tr6cnVSKSH+Rzc7fGA5JXRQt+ckdASpJ4C8069I7FlFen//Qg
cMgqx3cOV+OBwSF3LL6CDAjj+/cJH95VwVNou6sEBiDu6kTYhbXebIb6PWun2zec7CA314i+Zw0G
Dmx24Sc0kKr7Cm+pL3FIDD34h+8umR5RPVKClWhdLysyLFxfQ7We5aoywNiq55ZcwW+LKL6akZp3
h17ItVrh+zwnJq1JKYasZDw6kHJB/t5ogxhtlz31+78fYbKEw4d3hhLZIeVRfNfQUbc2FCEIwL0X
qLjYrlvXOXmzb3nAQF+usU3Zs1xq8YIvZgQS/Xh9B1p5qMXnWIroyrYfZAi6JZHPpU8H6Imqc9Mb
CU2pqr/civwCArPUISNxFzmE9OXI9dyvWikeueOUt/EALS5UEpK10Qi5Dik5esMGEwogQnqqJId1
f2rUf8RNCqGaNqHUGBIqcLiz9fALA81kKYMllRigVzGbMPocJPJ6b4HWz0YCZREv4xY2fwG/z4H9
ig/aD0P9BH0nbKlt/Tg2tdlSurVN2iRCAqAxd/+DCqlbEEmN0bkTLXSdtGz6qRx97sJNE42b2Dnx
ANEGZnX0ibcorOXP/9Z4A+YjOnRM3QKSBzalojfFS0ux9j9M23wiXw4kqHtGlg/VG6edHptoSwUp
k6pQqxaswD0NTdzNlc3I8EeTqHf2p4zsrU4N3KUWqyOUBOhl1swB+NXZYXq/AYA/y5DE6CTFKy3o
KsmQ/EwQeJPahifShuFnpS5qYXx3LjcLPYKUflVuWvyqAnKwM9auaLPi2wL1UZhC/fAygkK4c+d6
72/flNBa6raRSIIbqgEzMEPp6Ut564jiUCBYq8QEGQEEzJCLsV4r63+vGHlsDwH1Y4heYfq9NB+/
Ppjgf8M/E1Qlrj5J+q9V4HBKAAysYWrOKyeMTPYHDqEdNvrNM7HBjqWA48Dp5hOq+iZL2XedZ6cK
aMhS3BPWLhcG2Fgu8Q9jQlfnPAkAHG4bp+/8LJLruLgJtD43s3ErrNYFPEFVMKJ7UuLRXZZzb38C
vYB2np8DEWldePG/8SzlsL5qqSDTsuh77Z9EQd2W/5VMidI5fpoELJgiubEY5FvnO9kT7XIc2Dmk
dUMYscyRS+1Odt8LO0XK8RlkSvQ3eQYInNKeySyuTsNQNRBlmaaQtyZoCSAMPZCbAlikiODFo8m6
dRSMJ1UrharyD5yDhLxlHAWO3yu29RySMCQaQZirWDRx44ctLG9O7HAC0cFBhDKawuIxGukDCCp5
nPF1KFadcNMyaqMzy7PLmS5yfyDdDxSlxPv49LbUfv21u6iEo2uh/763KlNJFZOQux5fbs1o03kM
WHlTwQ401fv+eurUyAJ3HhnKiE1HXPVOznJayRDxNFt3xLZJit3FKu8bRkIpD70El7mOhaDWkTDi
XZaBYGorxVF5XyYhxwBmy4L8ybaf1fqnLhdff1DbfI6+gw+y7DlgAZ1kIZ5aZw3vso/oJUc4kog+
CyJxOQLL1t85qN2JlvTADNXt/+fB6yZOcw6fsywXI1w0zfPz8Azh/weRZm6u/8tsU+5AG/EZFYuj
b6DQJ8meavk5XYY4G6Ku/A3Y5I9vsAoViccCwIDM0J8GmIcTHq/h6fNjGVTd/g3J/0W/eIFPs9qe
gpTbTxuQURkqwAsB+hguru1Ut5O2wlmvERHab9ftp9aZtnczaE9INPIc3bx6uaNuuXq2DG7UOgFN
hJOShi19jnr7M6vzbIt71kzSbdUHmFNa/9NsVV47XCzWMaPDUvIEBs6YFW9tWF0y8nLEEpBiah+v
QDb+KY1cW41tw+siEkzCxxfIUmiTq7ubIoPE/mVtvzGLNRph43jxVdYF1NdIXXlZ3VX/zJ0ZKaVk
+RuKg3UWbG5U1Bl5yqcVpkHqz6Y5HBfljBL0lQUEn5jA90Ad8bKbTLNfkW5gdSddebvh5Q9eh4T5
hsoCMdjO6Eyc1eojLK30gT8xR0HPCIz9ATzQJm7HTcoIVguP0KkKt7nfEvEgyAwTnJb2QMzDQm4S
o8qTaIN40bNo4ryn1fgyXIjGiONRl78qq+EVbuw3OgnQQpFfmvEfk5/4yYVjJ1RonNq4/wVR/wh/
rGBZ73cGlMLoRouYdmdt5B0iVRatFNIkFOKnQBKCpQqBMyAtQ/nY6rTcP+PcTElDFbtctiuv4t1S
1HnN8nhzkfyZQ1deAQ1PkOe+76HjgrUCpT1ZSKP2uEF+6OXEjuzAQzL8yNNJ4tB3scvKk6FlFgQA
KeXgx0QFLNPHHhq4UI/vOatOw4rQbvfxKCAARq59ioJxURl0uawdw/AbYJS2W8Sb7GiY5lUPW83K
L7Ff9NaUnkCX171ehr5AX/qjRwjDL7wa/YGiEtXfBlBjrb0x6q5hQigeWuppUlKl6heS6PgaCUnW
i+MN6Zzu6kM59iP0HFf/KOp9HLLYeyX8P93dkwnQ2QnZbO5E+hcMpWaaCHa9bcgd01S5bLPYJAwX
Q6dH4calQ+M/CvXjWZzQhNEz4HP3zvy7S7sHj/FTEQSIk6kbB8iixLRF+mTnOZBxbb1Ai5ZUiMqB
oNwmQf020SiTyoKdGvF8R/lg+D0sCVDaFmXzdGzzhS88W77pEKuOwyiwrgu1rWCgNvyzuiliAz/w
Kp/s07K1yAKQCm0Z6ukRz69ib8D6ebTcTqwkLVPLT8FakTokVQRpub5nawHAtHucWppzKJ4wTRuu
jPgb6/aD6BSyHnu1FJSGeHOFEDZvhuxSUf+j6BxqSnfpZcH6HsD2TQUMmrb+9irnHuYslPSCn4eC
En3lBC80jcAF+OjVo7+4KmKipwCZ+PUEtJNDpKOeR2FxnCMzZtBinqQ1F2unk+6oMFET5mVwKqNf
Lwk3aNzLndsSYHdhRCUC3zb/MbPr2HwwxU73rNqc/FOf4mdIz3Z84DhUJnMy2CggdrCG0pH3C6Ot
IHSEnfOR9wYjjkub9hQhIEriIT/FpFEP1gGqj6N7akvxDZqUeARtdUsu5NSYiCLAK6+Co3wYPjy6
cWx0oNOweGMmGVpDs8afzvRoodm0GHbml7p+Y83U5O96e96xApnQv1Wwn+zE+Q047c32Jj63X8zD
o10OsXpuaNXmcMpKPwFYkaCAZ2yeelQJ8n89yBQHyAqD2r/3z41Z4aD7MwRDwJeNSwNdVl3sQ5TH
OMZPgAtPU8MFX6UICHnI2QXPq35w8yblYYVECZRreOJEh3xc/PbCohRpTNUjYT6GPXydwVRMrCjb
0eiQeCfB8NNL7r2pKTf9r90NEGjpo9rNQEdA63mPN8ePFZ9xaMGft41YCN3e8IpTZ+bgHQ8M4rM3
HL4wXSyAzOWX4xnUztBJfkmST6pOAED8kWMbquCdb1Bi267YcrzxD1BtBmJR/ak4rrrR2Y33f92E
Ij41/yiUY4wC43mGuKgYl3dkC1j5P1t4a54T8heADfp8X2Lh22wZ36rHYn2wdo+7ae5RecYjFQ/i
mfxMg1apvQLCZnONukyJV+6WHTaoX5v1mluOxYdUKkDkrxoWH6iKCuNXzf6dbQY56Y/bMGcw9dVn
at3YXc5/GbXpRTjN4FbbZSZKsRrpH1p90uluk2lSXbNU7b7BBdNGLwDkzG7A9b2Qe8HbkLtwpBj1
RGDA7aJOwGJAXOvzRAk8RnwEf72fJjnulCYHwO8AMk7R9ISpe3P1t9xDZzsXJdG8wVsOHhClAd80
n/DkbjnLKusPomFg+PbUYzhNkhZ49/BFNhjvGArV8v6c7x5G3DW1ABVNiB+Ea/3ei7ns1oyo9qav
B6LzLSqdHHOC24Hqj2D2RhryQC/LoUrbeQWAmiex+Od6UvdF6PxtQFuZ6cmnH8t+7v9AKttl2vuB
yKkBBHI4snWFajDlLv1jSpluaNybWYWa9KgggeULfVl822y216VKWkc6zmZmdxZ7V1/AVn0kTqnN
C4qcKTe3qxh+elIX/oaU8YvoN/pBSLFFXQswJHygI/DBthZHfusWRcz5YhmSou9/gH8yRjxZY1m1
Y0rpPI4Erdr0+smBiKJCeI8hfy90D7uyHi56I4lfXeS0WvEYZfqD2lXC7VjU0jq90Lyn6sPRJnRE
oli1hWDR7h7cBGQEeTrcbwnIhH4SLe1WAXVbnPt2hWjg8AWUdo++1BPqqYx2prwZVgPjzOYua6PI
0QKVZh855j/59oZmuZTnXNBGyToMakjTbj1l35WFneBoIF2CWjFh+OKQVZPv/pZMSBYfffKzrmUx
GdG2wr5mEz6JnfDWkAZ8glK9UhTX+7uNFz5qTInNezedb3uMDPCNUWR0eth58ygvhWvaqPb+GTWK
MIPOSLXixm0VYf5dZJqkvypitq7vthWDt6ZP1KrXWFVJXDZJelrqZSeSFDigHAgC2BfS9zJvUUt+
sMAIn9OEan5+4U3iPrZnQo7h8nDhaFafP8OKV4P3EeMG3xRkqGSmQMHWEhBf1B/86oOmnt5cxLiu
LUXZQavs2nY1NhJ1OFnD4lhh4pBhRXSbqVyO41l5b2AsOlGuNtRneXfo1pMgQq04G+kE3YsSpgDp
3gtW0PG278LVX/xILH2LSd7wWKIUHN86PoP8mImjD5hG+E4kbSjjNmGt+RNLTgcQEAv1Ob0gdaSc
GIyHr1qq+ZiQnFHfY2e6XdQWKK5wWeFXJ77MkVgF34tqKm+pLDGYcmicf7cMzW2bflprAfsNwCk+
u53RCmIrDBx3m/KIvMYhJrdryxfclYHb0eGibpRTGxldSAay/DB/1qb44WTSNDM689/yH4dImu/p
/jQvtEZhREIqP7RnOV+s3pYmfEYsKo6YWYzhAr04m5pR0PgYLW7lNYq2QS1QNZ2vnohj2uTE/2PT
n/Hbonerw1Do6SFVnmsbA66w2uc6n0Dk5200WOq0mxiYAf+W2pZU26vzl9hyWEjkEiu7CztvKPSY
5BvPF15kYkCwF+VMd9S4JLAJ13ik3dkWGuEOzWuXzU0wk6Ipdtqw23Cycod5Ob6j6P6nn47dEV83
+/B3xQDbwl3a3A87qF7KBevtheksanWeWYeS45/dXWprEohKiHtD7BhNKokryesJKkG0tmNvkJKQ
M6g5zpWBnoJMkXz8AkO+DT5dT34mnyB2+sOnWVw0zd/4yU1Xqsbjw/zpCXjl4g43z9MunZo48oEG
xj54U264LM06WnfWDVSAmQoE8f2vEAHt6TOv8WDIq8RrIKAJO1fgIs4oXrLLqJtYzbvTega7b7tY
5v7gWbqzmzI2hkCy+FyokE94p13dsSSAKEry/wIC4Hu4LBCvGmeWT/zsVCGItLQMsm17SIxjR78V
/99fKXgo60NTyh7plr3ks77p9v4B2NpdWjgqNS42H1+uS11P+RkwH5w1XWDyFhza408ByNwvLDTv
msxKPxOYBOKu4J4Y1wEXZ/eO031iZ9fkkvvV+4Ix3MZ04IEpX0N23Rgd+JM61LN7rKA9BLYqhPa8
uoDefYeknQwF15XLWIHIyCOr1HM5aoEooaNMneq3vPxxbvdr45hQNOY7g9YX/e3B3HcZo3cIyB4U
MSUw9wB5A6QSM5+i8J9/imFXjUFp0cZq9ZQas6thMbRKqwWAvMsOlrhQfwTVBTixuDx22pvgt2yv
5kHfWBt7IReJixjAWsSna64z24ehSq5kcN4S6H2pWyr4Kpmjsk7rydyQ2WJXgYh1eeWf/ulqG2Ko
KXBkFtIfliG9/UhXv1oMlgGbHENYjM6nLD2gtybVEurnMPQ+KsHrNTr9aXbkX/8vTWdZGA7GEilX
hBLZpDhjP/TRQmf70NOGZY/9miX4tj0eC6ITETwjeBhBPcDjzdUP9rOK+obnKZhKOjta73uPf4qD
zPzEXZeYtt1DbluCnqVXxN/iQniinIUXBKtqZOKarvTvxIMUfWJIiO2BeHTxBV92yGlcRpoOS2Hd
YmI1R0EbBE4q350wqvzTTXbkuWHg226ZCGheLZvHouSN6ppvbmBi6AREg4xDdePd0isEqZuaOClq
M1PTrwWkiwxFQotdZTgz2l0ZcrVZzlb/JJzl1cCfYdlqqtMHg0WYxRz4b/r0xpOWAm1Uu/dgpvbg
E5N26jB0qnI5TUhEHq1Kia3do2c1jj8NHMeBUyzWTano6/OLX2bNqeBv2y8UZj4jbdDwfeh69JzG
JvZg2Gsv3UVG4BRwFS/raRWJqYBjabIvePlxGNuxYsHJxnRScZS49WBALBXOofE4rhweLG3/Cq2+
Fm5P8QZS0RmrxxH6HHu6Zgv7xQiLeaHlyxfVqPsG6egiaGatAB6LG76mKpPkOwAJB6R9ec6LGmMO
yOiU8bMvvqbZAWvCowHgT+AUWpY/VdU164/h8KJkqR/LRSZeyR5YZF10rFgoW50OgW3UeWUOgj6s
IsfRDbrAYT6vU1rUjfMF4CnpRnZtCvG9BMAEYaC/n71z+5eZS7/7xetFFfkZb91PwlY+tofGs0qf
tFwcSHlApG6sr32XGw+nhJ+MwyAvKz0zTMTLJzHpZFB9XDr4VtgGRfjC1iQYlyxOAgW+yJjrXPPG
/A/KVZR9VrsXQH3fVZwvQ8+W5Udl3pIYwDMQ8eRmUze7RJTPyb8NAU4jWWMLOXC+A2Zf29skf+fY
aRvNmGJnbFkDw7CgTG923yiuwvZ3YrqGlrHJuAvDO954m5wWmtnc/dIBKSq3QzKDtj0BMtzfJwR7
4+N3UyhrpgH5N7l2+xeiruJFMcuo4du6tR0YmH8MrNHrfE/5mVxeGASQ6myqxck+4UymDax3T3g+
V2obg3AFHW0lVa0viI2WCf3cJq7Z7exaOP2P6Aefcx+blvgnOvahUsES99UowNWienBrjksrKmXa
PIjAyoXftklsj1N1/vl79xFKo9dOYLPEYqjsqzF7d1ONkBdBSjChgrGUtrqrzkPLrDck9Mtjbr4x
/dcJ1GLnbzptL3NPG5LKFzLIVE+RM/9J8O8i9OgimKN0POvTRh427Vyf2Kxzc/PTUnLP0xFsqZZX
17nUBRShmJ9yAbY5/T+X7T5nvYFEKs4RzbE/h+AXZlCOuJch7cS3MnNnf+GOkj4914PF+YutgPii
6ZZJZzgD2VrD3a0oy9gX2CNUa0J3+UjUE8qGxv5RiATpocW9faSl4+iNRQ5zUzKgzpNr00ojSpIX
D0Jk45tWa9yD2ccA0c2KNsOol6fcwi37rl0U8S4UXTUeULOYtnnuj0ECAojvBTdvlJ9kYXX2dYt/
kegZWraCYTGuldTwitML1PkFJdS93iflXYBMAfq9aFsbtdi8pLLmiqBqECj/e5UJtUIvUz1hY+Vz
EqoF/1EmzzmPjF1sLlCgQoIu/BuOrPNsVxgTU5KxrRTkEx8EOVuaxET2kCBwX/XeXrObiJc+b4jw
n1k6D3VOb7vU5OKPGxH2YtdOWvK0wEzDSeg9her6XooNcebOWoTuuCuYU8e3zNyQqwoFbXS1r4Rw
EP79yMgLoYBH1pA1c4oe6xLuCs1g3qnUAkRBpkkY1b6cPzfZxjixzb94rRD8N0Mp3j9n4qas4lpU
0qGFRdVfaO+Ym8//LpXbPXqygKwbACMiJwYlP8jttWJj6dPyPKShVwWPNDmxYQjIBlDkBSj4eOUy
7NddQ5ujrpK5QSftWSVOtWQIWyEJqSbdzjju6EsLl1baaKUveutBFqzChpUXiPxAxAUXJbx6+uNT
GfS3c/1fInp1EkL1n2E446kZrq2V5vL5tYRpb99+rcdHfLdDHsc0YJu8sD7QShxrOel7JN31c4iI
QCTEIVPHKqGova9tunT5nlCfOi+gI98rwds11oYRsJ7SKjieNI7S3qoaBhkGMcJOCqaGJsvB4Sf8
jqifPy1mFsT+jHDXGFTuMyyN4AXLE5hoT4a3qB5sXf+8LGzeHxaqP38pHnA/QfbxME/rnG32Qm1+
dJOIKalue2juANQa5w1book/OuFRFIoN4aBiOj0rdOwZumFxJAZYw3PpQGtbGtgA/0bwjm6wbo1C
C+Hug4JO2KoDAkwJk+4zDw/OMOpWXRWFTetcK+ZUThi0IJinE4BKubY3uCzwXCFaDcWR8sqkrOjU
IzIRTRfqZ5z/ltLnNHEF3aliJARZZpwUFm59bSvrhfBCu7MmGNC1CfzBCaSWahI5uV3K7OWYIsxb
xUJ8WHVQQwaRsbK0tLDNVxftRSIPDvhBemXdUyfYPIglQoKDNVtATPqo5Lquz3DOzUYRd+X7xytE
6YfKlATRCmgTo24DuZ1fC/gyKrRpnw9R1P2TkD/XUnZpmjLV1l6D8YMOBZLro2/LHU2ZpFsiSMrN
hWwODgdKvJrM2JjneKL6hU8ZB+HPwr2b3tEebPppfChMTCvrfOLZkZrPkUWAQtnSWSvt9icTEpVn
SSLNIrFj6TBNtcv8/YP1jRtavUsq0x3lXRfjsvjMvaw3zDkEieuu/UcqMKA5D+iQ7bPQmPnDbakQ
r4bNw0EWGy9dVY/FXKcidwPQ/gMzxx0Q6ELR81NO5MFySJR0mJ5UwtEoiNF7QxS7jghcil/M8Ok1
8IwFLyLNIyLodCw5ARgieDPX32UzP1AVaQl65jOA5IjoqaTadZGb+GBOyNoQJFfTCyssQANjtgFv
8wQeR2WjN5GIkL1TH9tsEkKg3tU5oAgHn+OqMrhejGw5m3ivh6rLsh8PA5hWWki2Wi4XWiizhoOR
Hb/LwIhf3jDx1o3SIfbu5YpkqH7yDPDXYqLAd5d/SmuZbzSf+6cH1z4OQ9LuIbbM1bgyKuLJScNH
d5wIhhxG2WVte0sR5U8VdtAbnTb8fPoyUQsSAzhyYpGr5zYBumXPhEHvZOS1R2kF6qP12ouTB/yJ
lSgyQWbwKw3zuvNdRmoiiYwXVN+c3Faniktj2rrgTUprHomurEr7kMU0JIBcodLqrs3Wvih2ZcVL
Sc9uJ1EsOMfEzaIEwSRzyQ+oen9gLZcQclcKR20sPB+Zv4RqftVrDbRQ+DfS1lpe0gmDIAXelfwK
raCHP4q81UZXQ6cb10ZTExC6jJdFpOP0xJ7jfru61d1a7WShAmgWnTdZU0ncvTrK2xzz+ywZbgis
1nUlxzBkF/eU6sA4id1pIfn4QJ7AslnjfxyRULm9oFS8Gw+Dh7ETEW0Agy/sIWg+WBQhza8lfTaQ
nu2o0/r0pPOneXPr61dcqgzglh8IZFtK50vQnOvc+mLmIhdP0qGb6nN5G8k0co/M8g0KXS48zB8Z
NT/m3VsrxBpVsryy5VrTuIsU9aK0BtZE+kaR4lX0lFiWu6bhSKO6xGMG9KQ79SH32Zzh+yteiIKg
krP9sAwsTE2CXZdfSt3Mir+/v4TvPMNxSlsfkWVxJaJ2qfMggZJYAbCXJGs8zCF1e+B+SwJNTHAY
3i7e5wxezYo9WHmluHmiUgZa8rZ5ym2XpqEq+sIFwM8AHeBiiQ2mL28VcoC4kob26EVI4ocLw7ew
T/1vs/UHl059A81yplbUxT+UrUbebQUjsb0yskNZB0dWFGJMGKvVxA3up5NJmx/nCQkVhT94DEeE
rQ5DdqexfIujt+EXfDA0PgXi2CNE299rMt/N9VRK7JY7YP22qdvI8iPL1TP5o5mY9yz905u/5NQh
zcEZf+EWI0VfWgMdYFgeiSdsp7IH57Ju3hHiGRpTobnQXuYXxLJhWJjHhM+a2tgfO7Ftue69d5Kw
LHHeI39THtCkRX+8KlhK+XZnexD34MD/tFaNx4llOmSexKQr45ZLwsXpJefF8aOLPu43mYsvvJtD
8JZM52/W8Bf+EKlwRiDjXbK8T2s/DtATq5CDx2MuQtmw3T3xGZ17ufZJRQbgQhr4qIE3SUwZ8col
oKx53XTR7SuyXMA5ShRhGJfFCR3R8VUkGI7WgYJrNLfEu9l8E43QS7NdezaiwUbq8qcUZUq/HXT2
Ecj8pHWeDV2IEY+bvpgKNnUtDZTluwyK9fP9QzoSO+BHk3/bQuTCFc5WAbNEjtfjW7gMCuWxxBcv
0MosbrcNHv8MGXbP/y2cplPgkvVT50fpPdpsP0L9XtZKd5s1YaeQ8tgLBA9nOqBH4rvZihJ0gz9H
k/lOSM08GmG+bpjoCLhyWt6xIyQ+mtKUypsP9y+fNJzfSnn53JaQx0X/aLou87FGkGYznhOMHpZ8
tZUHk137qapuPmZXScxb25LJjlYObEp7an3j3ATgGkVFZkM8CMhFXdBkSjrDLmcvlFJubwchd4Am
ITVJuhpnt9Ydttl6QpIRH/4JyPTNULjtAnyj7ZGg9vomxJh8klGycn+RhoezHMm+VoAuwby7tVGj
SiPNIRkCSo77/uIeWR9ZQLaVUSM6yd8sgSzNdR/AyB0LSNk2mawdRzmA1pdHC/bxICWk549GSEE+
kDj06dopiQq5ez8MdP8aDGimIf8exzd2HQv1rgzaxs92kPzDPhF1Cs+VS94yWNA84mlxBeZR5RIz
3Ynf11wPwzptdCRlKqU2gK707vLgrzaTcLrza3emBgqTfAumc0ggR+KIHvzI35Y51dFhVrZOrxGZ
dE94KNiCL+Rbc6dIqnXysQeEsL9tT/QFR4fuvEX227Fo1lLU1hvpomUEsmCsafWbJQm95AyP/g3Q
+fYaMI0bgceVhpYBenOAP5KvP6OQ6hSVdt7CRSXAgeJNCg24+b0Y7yC7uprHLq44Si9/RNKhAG4D
9hTg3U5SFBcchHPHZ2d2iAbQ5vVreH+pPjznpLCmrEqxAMgbV9R6vBQjHvyW3bsK8K8I09uBBYRB
3DH4uCKFhKXhzQvoYwBqYgiqK/I4fD/R1dAOErdO33tdHnS/dHQS0PeNf2PeigEmquuaYvnMFQRV
ST2QtC+01KhZgwBu9zmaH3BQE3mQCkvjOM6Ua/7t+ekxitynKpCIn+OLVW97DVlvyXBKvq+xC5s3
iMdbyseunGBEm2H4poJltF/tlWJGJEjquEwNYYVjgCftdQC7YVrZ1bnNqDC0oSAbr7g9nKcpdw6r
nUYl9V90yu3WZKKIVE5K5u4537bJmQoLLziaCooJycy5VEoN9WsezJC2Pbuq+fV2CSfEmBVe7bl5
U8efsbcx58BRl3SY9LLL1G4r0VmW6m46xpjHoNPWL4uEBebQsaKboNZ0vrbx6flRvpJEckFmKcFM
B7zNbZ8qCJPy4tIsOU9mtbUgHJwZaNQquuoG/Wi/VRxoq296cB9RUUovUekxTgmV622wvXydm2Mj
cXacICJdYcHr7uL2oRRU9aHKUSdwCY/uiR6hBhN+VPglmJoxm8kUXCJYE+TknZXqDIBlNt7Fs4Ca
w0eIr7NqeTVb0Qk3Scj8qPcBa+UNYDoyIRp7+6jc1NthTp1KPtf+OqFPZZdhssWF1Sxng3/dbXZO
76d8EvRfSIrM3WKcIy5CghJ0sMWHEwel+RycchtpGJJ5ObFc8chHS975skfEVq7JUvH5pYVH2kO/
wL2DfSiRNbeOu/fAB6sMYoOxLTlnAyF7dIG2mYHQKpXhMzpKByo7VFISSlWpxVtws+xFkS/yjAOC
TRZd0xpUKXpGO+1ewZWFadd395p03eVjctSEv5GmaCUXWsTIPGSxGfm1t/nQ1EWUhtv8UP0X3nfb
VSu2cEeZ7nXYMlAsVSTV8jrfGebs+4F1lBuNwnZfcWkJMIMasv/TwTisITiQuEsWq54Gtxu8OCQ/
EiZNgsibcg5b3rAH50b3mIkeExM1GdLIjImz/zgx47uANYMS1J9jXlmvdjnpFKJaWPWBdxHkoPK+
nBvj9gXfPK8bSeRTB5pKaFC0e3PDRokl7O0QJwOg60cjOWWam99npkVWfRhkOOQO5d/u0jfCqihs
craDS4NlxL3IrNpswFvfTZICBMJ6M/dZKo+Ed+ig19kPUE4+pE5Ml986BgKCixTJVKQ9RlKSiXfB
oQo9+9/BmznwNS+jmu7BLsod0kQFQn3khwodGKSx4qRigNijEM9A/m+OBtWqfvhcDKkpL77QC/OS
ACjVqLPg9QxIj4eDxjbcI8ecPzFwBtf4cE/bp3cmf49+359kNCWH2JUps8IQIvFRe+ausoyt48rS
XpsZVuHn+JEyTNr4Yg15o41LpYXytMLMIXZydCCIgQsC20a0gUfmhT+M72Q5CGkSo5U0LcdiFrS+
hoRpLu5WJURpsd8hrXHsG6rHyczaxLelG3BGSX8GVq2fUlmxry5liflxEMvd6IzPSH4LsS37Lor3
+Qav5RFXM2yRBW3ZfL5r2uDiA+W1p4FBBNFogF/En9qxsedo2TDc05ZZI3mRlbUiurUw4+fz1FT2
iL/6csNQrDnykZEOS1IVU/KNIg0ZdnTWXvH3fMNPqN39u8LZ40sKQwmq4EZSa8c8oKSF75AgAVo9
HY5yR3MEmYL1qAbaYH+++T4ua+EndQ7+tk+3xhYDfOgy8Dsuq46Iw1C7Tbxld4/0DnJzSW7654xK
akhtwxmHY4qrBGyFHEI5r5lwgsCmLBoHg18Ej+Qr5UnBs+gIGKeIMbOGAHKsC/4fGGbaCsdDoa2A
BiOHeXC3nPO91VGz87iASOBEtmAb/24FEUsLMCC01+4knnJIloxeHtEMH/sDuDpx3tnA1sLbSGw2
Qa7ePN4c1mGkjiAzmYrL9GN2Tcvsho865aKnXVMu1I8wzQxm0MuRSt23qsJ5eB0xNTh/4u/5ar2x
fpqmeTAwCHyvQH/Yt1JtJogr/tXPqB7io7EfhmB6itSOoyty59sB/NOvHRKSsTZTs9e021JOxo75
hZFZbiUUDTYq4/+yu2GPdpDtbJDhDA10GhkGvDdl8mke/6l4e0ggVVHZ/uH/6CgOsRD68ZfJy4ZL
hlm4/QMIvDxqqk9r+yu3l4cfROb9B1f2RrTMRg4bDToH+LPuM5mDcOIVFoAtUQO+GUHvwaSJhrp6
ThN8/QjnCUnGIFDMWQU9UCvI+lcCyGo/Eyxamz1vlS53/NzxkkK5B5GFoyEtxi74/Jtz3rtSM2Ru
2Pt54cMco3fDp4JJ1+XGUDMP7Mb+AF6VOZVq05S8vM85Uh8ptH6Ykw5CI6mdAKIOw4/M9zOFdtig
4zfgNZ7L5ejXs1MKqMs1xXuZG47loPXApaV/gvEh2r+Xil/YTfVJl4J1YEDyOHZdCtomXFKLe9K6
78Qgw0OoMVztgLWV26RBzVNVdI7bq7yKrSQ5pbAEpYthw+wwxTRYj64BeFFw+6jq/ex8CAZ/lE+n
utJEwyuvVXXPLf9YBjjHxmvgf0VJDXV+tTdBh9/3zdftRTKW/mz2zg0DjrgzbI9+tNUSC7gv7K7y
WiER+pindAVuEC/I4mg/BznvIMtFH3y+iUyR792eT0jr2v3VWX1dHe+DokvBgPmoQzD/oBY1PaHN
JjOFInK9bJYBdsOuCWNY8do16bSXmNZJplwSY0rlzKgSXkopCapc1wn7COfYlhA+9h3J1h458Tz4
qTJ8TrID9tL2doRZ6aEaB4wPTpBd8RqzxNOYB9HB+u9s+j1vdweuQ7/cM21h0zwW+lR5LJq8BEfO
BVD/RK6cyKFH9rmitnUkCXbIHvqgROs2u9kcMfORXEgZl+eY8Y1I8fouVrnGLNn8L+ISwSNJze/M
ENMLBBVRGmxj5mbbsatRoQ5sO4/K9V1E49VS1s77zrsgYhW8kE8cpCOIcJXoOK08tGA5t/9+91F7
fMrk5DkmPmSl9F36+Fi7rXcuGtECrP2S6k8iorVoDczTDGVxnm15YGucc6dVZabo+4Sej401w3Hi
ARPaV/T9FTXWem9+BbBpTM6arMdinQ8uAymwaIGEtP68Z3CrBE4co0npu5YGGMyTNvk/IEIaC/th
zguXO5HfDQ5TRrqA8K1nLf1kkXdWCqv2N15mgyLW9ejnB9lfyCHLrYG/8HCSdFSXKJSWKYs3aTIp
Yi26cbBCcbPhML6hb0dnv/eJ351i4viseQb9es205q6QZutPHRZwU9mwWxmKTsRr47in3DG8q29p
P+O+FXpM4VREkFtukRGm+ha7waGYWbPJoF/Cfc+Tnp3nh+wOVAa+mZA4jomCUXpvzftCKIg25nI4
QZ/xEcNyMBpVDzq+zmqQB3c3RwC0W6qec9V6gFgFaqPgoKMKutEEjGf1YxA5k1zKUc8tV7J255lS
D9rN69krU2zDE0kTRD+JX+BG3R18XcoGii64pX4MFjQHg5r+5EJ6U+6Mj0bUGNWiw+lMRnPR8Cu2
UorfeCQCaPQ2guxbZt9liEofOXKqdS2GiDVjyO3y+jVD8PK9VAvGAKCciHXJGYGkP67QzXvyxo/d
rZdwQFMLZmFR3HQHfcvbGZE2Oo3sFmXvfy688kYtz86DJNVKExhh2tdrgPHmfV5KlaI4DjaSuVDs
xHnhhqf8ud37IEmrou1rxXBQ9uHXCd/POgmhQhvAPwskFYhEZMPuAD6KSAIIghRLhAYIionD5Ch0
AfzNRbskn979UZCghSD5SL4FoF/meBJOgWyZ+VmxGG4o7vuaGICi1T6+qS/1v0xOuLe6y4U1dBP3
7mXzdVQDDzgOpmynS/afzwoedbp+Deo8ZvfQi/GE0T6CXhk6MeXu27MzrNVtfFvFGUSZm+Z+cOZw
OW8Leg8aVDha4M63Ysx3EoZ/sdTyr0KCdfZIh/HDJ7CGKcFXNbT3DplAYOEiNYyF1NIyYNBV6AS/
KVWxsx6pb/sSkHqGn4WDBqU5bODz0jjozqiU2Vb6bRpLlOadNpOyfuRy89PGmRGMEMbBiIa9hzPY
I9Khi7lleZ+AKmzleQBtRTP998yse6LLBavkvcmZvGSZjlJh+Z8oGBsaAhJsOKtC1JA69HfzUezg
QeGPrmTCz2dIlCy3s83FzqFbBPvLv6vaOaghqO1/L/9Kfr1VoDrZEXhthnShnUCsXtKG3Y14FGzZ
WhwN1M53vRI+U/0G/fMhzXzr0FXn98f7Rgd1/USWIaWYr2asDPp9ejKxRpB21EL7tSIfDyDL5fLW
m5zUqCQRDsKY+tFhWk3hOQkIo/cJ4LgcjjJIZ9Yo/3g8HzwnRXgw8LyceeJEzZ7fuJMmKNZ9o5xo
PGg14lbpGNwm18q9/Ix+UVHGk2Pww+aMgIyWJNc8qDC2ZQe7wx0J23VXjN39CXk1xXMaQPhgDZ3S
Fk0C/wb74ljbJ7P9mltG3gXhOInCfJx9UHPEOvJjEumUo1TamtC9eJBeJw42l+2YEf5b+9ESnwDE
SQ28tzsZ5iG2f7OSbas/x8haLo4WbiWgcBhouVPOaYuGbYPTgheOrml6zIXHSuXT0tL7Ddj5Gv/f
rQnC9xoYvBcUb32bI5rkOMVnKQ4qmSnSW6fAuWhADP543HKPDbLnGeAfsukXriMXv/YyE2UgbUNi
WxJBWHGN25A/kIzRfQEUr0dVbW4SheFLw8aH92pljJVo+gzgVU/Etgz4YP627URYhDn3o4eGa/xD
f9EZpibVu1A1Xv5cOCgsbjE3AFhkbBkI2YPw40mwrBhtmofJBT0RPudi7XthBMOgWKztADkiBHDr
3aHKlP73M1At6OYXub5ZXfKHvKSkL1MqaxLxVFlqpStmp46zmZ9iZs7/XLTZ86imYA8p5kTHfk/N
kxbk5OvR5Hl9P/nP8pj3NWABtT6UedJyaxzxtECrcWDDdYqrxQv7BqeaxMjv9UQSL5xUKzVlqJF5
IB9ddw3Wd3JoplYLMqBKkCPQeA2y6fTBeJJuXYdV6NPFWwAzAPm4JN2K5MQOHyxwusvt8z0IfXQp
2wDZ7zfQrqprQ+ieFYvVNZ3ElAou9qBhPmCI1FXLZ6kuoOvsCmrq7YcE9bybRiqJQFspu8EyYHwd
dEeIsiV89RPNrElIzuolDG5rec5Cou7FmLaZBV4pIbk+9eU9/M/4Jzl3rj0udfLS7DrFJikqAwI4
b4yypqu+rUFFZq5mAFVQSZsXlfZkHNPE+YH/IrXy0mcJufgC5KsmM+EfPzSLw5JKJeNB0H/dmAgJ
4ZP5W28/U2lJmq6vRDClI7zwL77ypoJVkbULIb652OThEdR2ut13Ups86OwXjnzoBvbJvOrw5+B4
XaKw7p+RtHXVaBUMaRPDHJBkmakCwSAJNhLGS3zymGl86DRWGWIzBdpOn1dk3jDtQMDHvE7Ozz8i
K0kint1yvIv/Cc+nHmG1Bk1y0S6zJXQyq8+72UtSIhbdjsTHebWj+oZb1BNLLRS8M+dEyghtnMeT
VxvgaohWnLjBCNP8GFsdbCIxYKRu96wI2pGCOudgeV4cIAZ/AHAd7wkt/dXb8MNIhw/k2Ax0qB5l
tBWJqQOdm2Ie8XZ8qLTCMyHsBuly+AXzx1+aQ9DJoQc0Kl4zawJdoZPvkj+ntkxvbgym5CbulASM
vR2DSstMXfUL07YQInriL5kqtQ4GnD/yLAxHZeEVtgqK7Kii7fpn05iOqRpJoq8ILQFPgA72jNUw
Mi0uipZkkTd3XeD8nUVMDK0kQYgHBYMjwm/msekQgpgbRYfRv2JeY4ITtkZKn4dzndatf9DTxFmy
E15OMup3qcmkTxX5VMQDikehBauMZIs75MZToUqcayI4FsaxagQKtEJ4ceVBWZtObCqKvqOsp8q+
KPBPIHVcWgVNYzsy+uPwwb89NNSlapJ+YIdZrgJZoifoKGuNMZAywttaO59f19DOLvdKyFc8RFMe
xkxY1FrowrMddoCCoeSXhIuj0s29DSuEm/Hl6x3bs/VZe/fFpfJ8QzfykRUOWTaLWek4QV08hTMw
oV3v8XqPb6E/0Uo6IWY3CsBwn00WLKGxG+GjKPkdrc+jfJ+NfwlYSnmrxhLZ8LvKRjOUMguKjutl
MpFjYkvCkfqNT8/bmsjBNMwyuQWlJZqyhlTlnHGkgmqyO56/Ym+3nM47yQIyEdqmrqMqPEgYustE
hjyAoWht8fVMQYKxEGzfBh/YXUrCG8pmZVvQBRD525vHlCmjWjMNk6dwJs0o8hnXV3CfsKiLPhzj
0oiE9drBkzFwWfYjLcoZw4pDn3O4Ntkfmjl5VXDy0aAt3rPrukqwJX77GT6ksfIg0ZHCCfxhmTBq
ee9mU9vWVQOmpSvyzqJT/NBGvqOb5O1jKcYQUvT6bvJJAFGtwEHUAiJ+We88hvC9aD3VQoZlwe4U
Y2SwJPsoqWE+208fu8qbTpt3qWUMuXWTbBq6kaMPu70dm5O218TY+cXFnd4rbOiA6BwlQwL73qgw
p+HnhCWbvHdoW3HvqBov93Ig9JXz4Izp/hvdmRQJjB6KRLSWRM3oRAG7jiEEfbJiw2LeyhJcMtw2
zdlV6i6RTxTAsl8tNUQckhNogycWbvZPw7ENy2bknIuY6e9ewqYl/DmkBwpv7sPtH5Ms2BskihWa
R1OV/U01vNx0E5S9ku24vvCeJ2IBYi6MUR+wndiKpsr0NwyhUpjrBBDePdJ/EiioSNSgxZFpXfJo
oTwKEwYuSNReSQaFE7IL+GXJz2sVPYASUHlwqUmrbXYANnMNb9CfmdRdylR1begiN2TbBMHeE9g3
T5YpMsKC3qYisY97TkC/uznc4POcj7wSELVLJg1E73BGD4euqTiTKzXIV3LAgFyXcluef2MbXkpO
qsePRa84a6yannJG0nXJ3l+FRp/X1dC6e9mziC1YT/ZUo5jpgNTKejjr0cRS8RIxd1zhI3195MRX
uKvfJKpIwiDVWRbiOkw6Aj9sMxHZPIN0BdL/RLIewRL789501a19BXf1kLzbiJFRwRAnvLFP1Et1
QV6ekZ3Y1aCe6Gg5QvqZrRbUXgbuhUnITlNtjPDa71uQU/Iwf0BW9GIVQaKjKm1QBgxhLdC+GQfN
BLmMVFSOumpCosf7phbGE8n+xMVA53P79Y0v8CcgCRElq7fdnOeJr29ECFwz9lv6HCEATh64Pb0d
wZu2NGUa0i5ec/ynPqhU1J3he/YjQ+qyccoq6l8iOAZrWsLqrF9hqgPp4TDVqS7yamaa03B/NLmb
+/Ts4b0M0H74Vowtz4ZMi+iaH9e9oMmt9HxqRspGmty8hrA7ZeWEv4Lh5FLGPAfFoerfMwWVsHdX
dyiCZDF98rMPSBHQ5qIzq7tFIZ4VJ+OBNT5GraKsZxh40VFyyS9W+Pb+Q0ieA65xUOLMLfJGdPI6
4FlGHWuoOo17zJH/v5Pm4WZUr8gSBhM995SjWbwbX2uwt0APdr+WLVwMjwdj8j+hVPfL5hhjq97t
72XG/tKWpwqsm1CfAh8ZWatjAP5AnRl/OpuFE2p09fBZ7rS62SppZqeTm9+joGAnRohVrzIRnuvu
Gm+ESi8BJwlLndVmfpoM2voXjrMbLWgnw0xpu8G5aBLg20RRVl1te/kRzSGJ6+WFj6RNDQ5HSKTn
O+xo1wwiWLBcjNwruTrClqbnT/7hZ/9wBzjjqieJSN7NbjAeb1EsaFQFTmfEcQb7I5NPpGj6aNcV
r5OmBzXh1f9bfkU+swKFXAk0COMbqvllWMhvTVdHdHOBhr0KN+LFr7eqQ50NIiYFpPgM4/7Jiie0
UCT/JpMBNxsGlx8Qb9WO5eDz4tMz1MTtCWOcYpI960hpJg/8QAyBSpPROiBfbuSvNBL4LsQuvdVT
GC/GpNt1TavOionKtJrRa8C15nirWFph/7TWSnJy98KWCjkT6269ec4VMkO8qTtwEteGXGSHrQp2
qEU8v305nGAVBvttATWK67sqzvRemJwcLRatEtMNEoajsZyhj5dW2GLpSYWHYSy+McrhOaAlIFMU
lXINkMx7N6Rzvsot7hxyuJ05adFoa+exMUX4IJwBPzoJ881bnI5ZrMHonunNYM/FMFxSHbO64Cai
9WKodYfovb+EFv8p4OsDsajNAI2rA0x/AoKEYdbGDsN9/uctq/E39wonmmbCgKHWj/Gp/eZkcxD1
zQJUyJkSkKkYEZdLwvQ7hfKcd+ldfZsSECj737kmtRdwjmNIIaio19WOrlFDeivZ+G6+bLKTYGb1
3vsT/+FzxexX1xvp3aluSN9TzXZJZFrdrSoLvGywRcuw5UfyRduBGltT8d854FlTv/fhIc9MfRij
pAOFw43oF+proEvPDyeZxaXDWFt8VTRZVB5+o7n0TfhQYuvaGBGo+zEsZF7bx0zEad5sLJVg7n6N
0SiGrLM4g1Ry4nqI5/LpnmZxBUlbZGkz6ca0swBVdgSG5EZxTV1XzbmXyx/QuTwCO1+kXVJx7iUk
GVc2X3aPnXFyVj1CemUxYEJaiwZviFqq53c9m6ugQN153nMLTWiKuRGwpWWS6YoeUYrEq4n+VF9n
jXfXnc/U/9h05d8CgdB6fnGiNc8wAMzz88xKI+Y22TxWQAZ90owPhL8r7g41KuTTLPQGbw5qmOb+
W8sVwYM0p6whNjZAWxSMC4YTYWqzVKHzog4Qf9E6lLvO1pmDPfjZjQ76ieBO8UnUyTPNElv9Ltfu
E2n8rTiIrRWQxaPbMAhnc1ayQQ6bDn86Igz0oCZrdl53JIyRO5yjyMMAeDgvWGdPmOb+vTOUsC0z
hCE8jkK6b9m770uCKAjeL5ZVURjWviFSphAL9eHCvkjpqjt01a+SQZkuu5lJJXMzpQ4bZEipNe1n
xbyTEeb8VF0ingjFrPK6ncPuquD9cg4X4xLiNWiX86d8Gz6aC2q14xUFjIPk+48pNm6R4G+creC6
VghXgpJus3T1FhzGM9jULXM5gkTU4wfRvWwjN0vY58XDk/O3JsvN9SBXgmD9b9/tcSCwkxpvXIez
W0/JAIQdGYq/WtEqkulnOa9HvQ+dnbf8h1cOpEk8i6t6PEIMOA+v9KuH0bVqoHmwysYr/o6iEYsZ
qCcpyolQGOysKUEM+n9+9H+NK44juhctyQCYQTc9tk/VeD0/yO7A3txoszDCeaUyvZnevK7T0Tml
tS9KuMp5OPrqCz3o8fC5+0pLvkbXNNbqoPrLs5ICfJL8jeXdnsjL8tE5Dyvwi72pHKRR9W00DI2u
Foz4pZl2P6crk38RFGHyyIz1zLwvCbTL4WyXmOP6PbZ1dS4xZxFZUI4xFxJf3bNmV603yozADxYY
QEEWoGX0fMMUD0LDvhqY3nO74T6yubMs9A22IsAIlxRtRgNipRgnkgO7B5fkxCWM4NmRZbH2Qq7Y
+zVgZJCBd7zWjpi3xBB0uxPTlQdPi0zN9uuSOpFFF4Sp3Td9TjCwqmaq7oppoFc6ZVTif1bkF/Z0
t20YHC1Fo5PYN7SprZqw/tGzqpbV2t2ZSY8CM64+c694Av7tmgywt+RFcTljG43SaoG6h9T4DkEH
KIky/LBOedyTdk7faFSpUgFosjKnUIxk+ObOCIre6yshDRsdMf1nSBPBK3EhiPG4cvpqJFsvWgQD
u+lq/Ym4nQzO5uylZmhoMVAzlUgGFC6/fuwGiKkZmWiE69SMtE/XzUjS7jh+SCriHJlyeJUImAHQ
KIzHJaiYJZ/8g0WqAgpRwHRA818MyKT/VvbACneJcpeLXf+3MOHwLC1+8oZDPq+1J4PPM2dQcPGj
JSCvEBPdrmBHS6WgYbvebqjMauYdK8fE9zuBPlKVjpdP0JCGo94kbi1aH6hBgZHwFUGx2wn6Xozo
qm25nnGd3Qb0CCZhbB2tQfPKN+WZ6YV7ZYVyi2Eb9+bPD2nvj5NcBxu1+ZtNkBP+0z28E0DfOrW0
5jQoilIbwsXOkJISu+remualjv8I3g5EsnQo/Vvvka9zSA7j6i+7DwmtmPNbHsg9wYE3/FjtVHAN
bL3n//6Zc0UAm3jKSahES8M6nzqFVVPMW2ioFgGOJC8xBQNH5dp5zfWJGf7xGYHKxyiQ3HJORn+Q
sb7AexEll4YGSS1w83cZ22Q1t27yjpL4GQvEvIe8yS5pnWVgIsnzT/+DGrZz2FGPt03j0NqnaEF9
320HdqKV9kDdASAu91GlTVv7u92JIbm9vV8j9g7RmbGrwrS8Yz9B/gKfgisPY/CpS3n182/LNkhx
lmijjOZzQLPiF67ER0oLBU4G+f4d3J7aQTSLOk4HK5JfBKXgRXkLG+LsN536H2cNz42lKm6ULzPN
iP2u2a8NyzXcfSi0Jecv03ky+O+Uf6GjEGSJfgU9U3/5DiepiFkL+TNVS0AB8yeuSPL6DgG6mRox
28OGiX67CcBywvq9izuqzWQ0E5R9Q0KNB/S+J+Eufdqu+ZoivgzdxYCtJl3xrIEbZJfRMseErhgB
xQGT/J/QxUI74ACf8si7d8dwi0NOciir0FUG0eBEQvZiFzLxrTUPpF/m9hKNZQMLDUOgHk39H5/I
Z53RXNf6i9NP33xtjE85RBhK4XECOztEvZxpgMgYuPny2pr3f7HWh3bjtyhXCs3v4DS0iQBY6Kv4
VI6y/aukKxfuR70lxRtkpl0rdQI/4fjrRFDXYSUHTykBzM2vrKTEvh0MkCx/w72NT2mLl3m6LJ6/
0SlJswLULaCYvTh4RYEkMwmZJD7p9x2fcKGwuBsxY9KhaQLL7qpc5kncKZfUtAWH6lRpKjo59W8y
gzWeV8FoBOdTYE6H80D7CpiSanPcqehW/piTEnKh7soxF7Bx6h/LbRQRQNuv9Mbpz8JoCPlL2UFm
Yf6M41ZD/XnhWFJxQJnKSnrAnstJ4R8gTVKqI6a1BNrXDKzxrqrYBY8eJsPXaHcqpZcX5eWouicm
e0LTEvMqgoI2vQrdGVZqS+jvswAeRBLa3alPxuGy3OWvwTjLmzX6dIlN8L1RgP4R/j9ITcQkHZ+F
956B90ksZnmB06Vqz4zqYNCvj0iOUtAt0dft9mpOUrg8lAx6RzUXICUIGJHmKsSuhazFrIY4l4Li
+GkCXtcCTBzaKgAi7DsVry6+BzQTTiti5bRKIt/98RMmVEbt0Ag1PcBXYK6AJLZYc+f5uQW1clyH
NFYNStimGUj+eXoH/Z7NlOyBiCu4C3a/Vk4YzFbxCuUuBuLrXKR8QvaSzV7GDFTPp9HdMt9khQQJ
7L3ooq5WGvvJGt/XeW49TSfdk9Cpb0EH/bg5RI0TQuURP6dmerjgj3XtPXvLcyt3bqhrVabgbV//
18N5nf0Ici0geuXBqMHd7GQzMwWDzXJ0Si/cl4Ymq10hPb8Ejii+dJHUPHqPmZsZC6paZHa7TVzb
Qtpmik/OVg8vUn6C8u3zS2So8gF0ytE+THe3OANDHoXr2K3o4H9VFphMK76QWhTwMEFgK4RI/lKp
KNfb6mahTAyIH7wzCbGViFa2L66RA8rOax0nXC/0KocIYHCoI9mfBYnhoWnWayxTmNV2DsgNHn3C
SVJYkLF0eGDPw1oA8Ifl0eD545K27vKnJdL/bc5wypwW+6vVJEdj44qQ7TUm3mmTNWcww6kNwqLc
bMNUcXXwnwWklJeY0QRXwWqGH6RNM1WLxONjk1QRGOc0KFE9EgtmJ8UEUGUU3u6fN/2EHfK3aCVc
FcefLBhQ1kwVzhzJfpkdjD22YWOh+8E0ra0+tkLfKFbAOy2gDSDpT6DbsYdiWDTpRFwusPXNM7kB
l5Q5hvAoloyJ6rpaENs/4YAyN4Y38XhJC1Zu1f4MJZ7ZCwWCd/7V4Gj5Z//AcuSHryUFdJxsywz1
j8N+tufJ4sHgWBYptFyTTC+G8goPPqTAjr481ZpPJBH9aXgmQpgolM6tvrKutgppLnik07QOFe5O
hrswhFE7chPIejFVFVtFlQ0Mb8qAZH73reToxmoZEy6Uzaky01MpDWb3bPK0SUY55i9X798E03D6
10q/Lxzd50pMV8g1RQWbQtp0zltasujvSXJMGgq7JgeFF4b0jzqHEuf5RTOby0iZJp9bi+luNIXi
q5RfCrGP/RYz0/E5MYqeoE46vvwe7Ccphum74+x9lVLj6uXkC8gc8ATKaM2GWi/ssbgDlkcnCz2U
MF0yRedloWL+Qx3GHjq+JzXJxFRbzjYeMp4BLVZICV4t1d9MK56hC3njmOz6cwcEWIcrxghwF5HV
7VUWtkVQdZs4rQsUkMGh2kgzPerpm2d5x2Gul2eOJjh/L+MW4pKyny3liDMDUAkUGOPXqh+0ppyh
h07D5wZte1+0EEV1UAPob6/Jd5vgziM/oJPtPw3JxkqQ/apvi4Ivxo89VZBgrlvJx5D9xFpYDjmH
uvla4sJM8Q5OkLnBzggCXWU4TJFmAqcqVRJOqj4JGPc2eJIn8+vZcuNVluk8KvQAJq6JqPU1lghC
cdNk3Xo9nQFNrNHuvmmobWrK/q3odPIvik8VqBaDa+gN9W/q+nVNNBzorJHqKCn1R6Gxh1Egc+b/
htU3/A2WB81L/hLXESFm49JhjmQYR3AQ/bs5XWO04mZMuvSCo7J2Kipi78jo0g8CJo2w4vEazyGP
E2cFwIHDhsC4LJA8GbNnsbfIAy80E9ny//iRVJ3Cz4DuuGPyHD/YFfUV2/6bkuYuks3/szNXpw1F
byYI6B2Ja+H7wCNjhAlraNUPaP1o40HVhqbpUpP9qWe5UEM57Ua9O03hEnZV9/hBZEK49AcpvPSb
gzqWWfc+rfRCVxLx3r4fRynNo69MitvsmNsdbbM/r+3cNJyzzX6Z85PMes4aMV3WRPTFrEf2d9LO
yVqF3rSHoFWp9ih630qgqksl+N/drfyJP6hKxmJWnBGa7hOrw+mzzxs1DLqA7xSrQUiBieDctoRW
5dsEGWKZUOdpGP63a4il2qi15PRv+aIysNzcnP3ULfihKxnjCV+qWyMVNVfeH/Tu6Kr4K0TIXDrT
u5wrXziEnpKJ/G1cGR7/5JdI49GyLwmuhfAUGetk7esyByQAzI91KQwRaUIqNE5FJRx8LOM2hTmQ
/QLBsewwDfXv/GT+YdAqZyNOPmBszCtl6VtQ9+SKj910QKzIUjT6KteG74cPa50H5OWD8OyLv3ef
fFtaM4EneTT8NXL/V7nZBpNsitR7b5QzkG3nmqMBU57pRQfh61grF5FZosu9NhcI/y2zX7BQj6rn
39Ki54ZKli8NmsKpdy6KmOrQefK7YiinJb0KkrzdyKTFKFNpe26XHPBTZVBLaAdOeOcLFqtBx0JZ
qySwMIUrHVCU2NSbosBojB6pl2BWRZJ1l+vT2HeiDPVsXtt6NzmZRnKtFz/+03zYBoMjreiCapy8
Abg9sPzAB4MO9Pz1E4NYQwE+CPWCsbCvYXVpbglikq0mlrDDr6YEKlbGZhROK26J+ZJqN7tIMVqN
aUkJjySvvW7f3eRuXjc0YRMdNEWhkHmIDYAZ4cqzUja4RYGq+hsDrffsjyVf6AcXaVVYaKnbf/4K
9MhWviky53AdC3EEQyN9+njaQP1AW6DhjAuzed1CFSVKns9ToTB34eReykVHc2Ga6aCVnckQ45av
DOAx8/MsHjZ+eelejIJtndXmDz2rgzGjzTMP4DnpwqOmXS8U5v4HycbX7hpQI89AcJUXCBxzm+Mn
hIwXSJCOi4izbIXYG2vS1zE5xpSUPVsCZo87YAbgS+MaVYhX3DjkG53i9AXeals1XBdbylka6Qns
zMYb/j/FiScSpDgirgls7VvdS4lPOVWUww1EzbMR9+6zfIIN7mgJHYAMjrqW8l60S0dTlnakvTHb
NE1dCyp1Zi8vR5Oyx4StZB3zf3maWBYDZ0wLF31twyBGfLGipgZl93ZPKMKnT/Q9DgQlLvMahNPt
w9rNa1h14tmMbOz3gUJUAeSYMQpE1gGCYCArKWi3AjmJVjTjLiY4uWORPYlWC7swRsxaFUsKnDgm
GpNhu7lj+XCkF3bV5j/zzBro4BlIYDiernejrFmKcaC7EPldTYYDT/G1jAtj7ykKbqB2eeII1Vtz
BlugG8R3dVkuKPuPc3z4bRG4EvCpuxDTwyxke/4umlYAHs4TFAvZYM+DB+YgZ6P7bpPU6hYrASJx
Xqb4S/pC4zMu7GQjbdHpAJ4wxorRxjSEmVw/oB2HlDJBIanRmfZsY4mHQQDpmbX4bomLOIAykRUX
4lo8Cxk/BSq/IB/rfptZvdUmYrF/CHPwxyDPMpjBKYVxOkDUpjykP7UZIofqZ9vudO6k0LXylh3Y
anF/sHpgMzrG9I/ku6/XfIeTYsN/h2zE30W2ZhSkS8ccuIAIgiIfselmhH69HlF7puqtG7JLibJH
ImctkhJI0/xWOiKTXYRCrBUXNCdKli7zFsd9kCxNI6hjIpdjUtWuH517yI1AVxKNmDC+FexnXhiS
kKf2z8qYG6KiC+HUE9j5oHIzhNulX/Jroz9PqlyyKWHUDVv03RugvFrsC5UIDNGYONBPa+p8WEfJ
IvitB+3ZnPywMk48urUeCAeJbF6rN5n3MqZmyb4sCqcKHbYnc3YFT00nDUuaDOMnwYzhiwe3OZtb
pZ2K17NFPr3ZXv+2U22+Pj7AC8odH0V6wSugakN77j80lFNABX/ChChC4cpC27vjonMJSuHmSRn4
CXm92mYM+LcsYzllbUSvsEdxTlk9jDYP3tjyQgYDR+XO/xqJuSAvyR4A5xBr7udw6rl/vxWeguIl
fJQlqzLPYU9aUpnD5EejCaQd7Y7wdXvUMZY+1lICRqEJJVBtsgk4aAYZ+wmxhJW6hmwWqqwnL0zJ
vn9we5svqiwT989rMEtQxC7QQ53lqXssTuC/cbLWCn8zbLR0wQS6FbG3PzrNJyE66MLQaxUL4AO8
PfIgtmrWRVwGAEIr3GQ+Kar0EgdbLXH5OVSVgwQVyboP0ggqdh3HINcMqiW3DvnhMtX2/fP195Qo
9ieMiLZnirdM78VUNCfnRvjzPtIHQKJUZV5T7jYtcmms47bWTaODVX684L+s6gyuTSi20iOwuwYZ
/VKmhjaR24cTVdXLpJzh59Wy2Rgl8d+BwUsUwbDvz75vhzjPAQpnMFE19M5oob+/CNiP+43qykUv
t//KRgrYMs0Hji4ANKUytgrLwM6NpEaWgOgSbsZjEtpRV1Y1gXIzJvjvmNZlXkCzK7lGxHbUBTIp
obWQF5MQJvz3lJvckXd6SlktqlwBx5Ua2UcWe7ModQmojocDKm1/T/s2xB0OBvwmIOGo8VbPszFA
jUDLBaXIwvIJnPNDqbUm6KXMILUei2ExPD0G9O3355LqLeo3+dyqb18P4BTspsuALLGU2uf0SY7z
1zCrNKJMr7mbHX39T6FUswRHaNXt/up+5qUuAsE7nedR+t+LiURDW3sMSYagXmhncB4KL+jvHCO4
uRqT3MEArDkARfUkhT9Tkro/raxMxCZ6Toac16nnZdEplDUOMxKco9MU/Kd9Cz9RzukVbmitu3hX
8nR75yQ+pJAZbh4rDEXY/QLFEFj9Fcqsg/UtowABzSc8+LIYQNMXqEAQiY6DBe89p1b6NAGHwEKJ
+J1wuhATvM7Fmpz9n4axLRVHUmxXZIX7W6qw/NwmqpnHPxM8Dh9L/6WJ1jK0PW1SQwPt/2niOmma
sRRwP+yL+HqOeDV434+ncegvDivkxLi0/GwOGxqbHpKvFdqUkN79AzsM/1wAAAcey4ny0bI8j8KZ
owmPriVi04kStpQBNi9vJl/NslONWuQDUWx9ulYd2yGEwbwondx37Vu17DIrQXOwmTJI8Lu0Y2qh
U/6bjCuUyr/3H10nuqcPXIvwkJ8j5dWWSPyXWGw9DcoUVc9fFH9KmXwWkJznbP5hcvpRd1+qyp2m
LIWiKxvreiIiOVtZUWD88FVHp6ptkTyT/0rGCBHHVZ7RHWUdyLNWaoNII+9YNG3fU235ZVhsrSSY
DnO7G40Ero9jHeqixJKmCiAVHrdCB6oDE5JXm4Q2NS9tijPN9KD7XbyGSnN2aSmStw5sgsQ/iWBv
RMloi/L1H7bLnR72BnzDRY3W0phTONcxdI3O9SFOIBjfSXDUFY/fAkqLU2kyeQw/agwuhBCCUfmP
CN0J42GOsKU2bwX7eL0lFpcb3Ukq/0KPr8d+tq+IRWU5c8Xfvzf14EgTzn5iTk6+x3OlwpcjvvVJ
4KLDeyLuq3aDtEcDRWizB8xwqNjWnZGh1NcjdbpUuBel+E+K6FrfgsvVDGa/pxtuETiTfqFVXFtZ
aCtE/2zLh2GIJwR81y9LKiPh1RmdgMOFzq/kjtM6UOWosMHjhH2orpOMf7QJW7faYRDfZnzoHbzP
a6G494n0rM/mbG5AwzWHjqy+HmamYXu+kZEM4mKBmssxQY7uXvqKyZ2dFCtyt480SuqabXG/BYLE
gGaNLcgP78cc3wxc1p4PD+7wPuqCZFHbgyIgRbfHEeUDlMzpx3ubkYfLPzQxv5SiQC+6pRLuNJBB
E9zNnz4KeHCG7POuFz5F0l9Kt42RWNgMsh7qJ2vCP6RD8KjNHapHpW0N9VshfV7rsEB59GiNWaQY
GDfcSqeBpAqIWSy9FNuNODZI9m81PqOQoLloKpoyZ7D8o5pTGYyI7cx10U4SekdcRJHgLOT/uGq7
wQSm+DVRVCi88xdQ6HwKHycPu5VbnQZ00F8d7UpRv/eddqmGu1nbLfCrytRT2Ah9Xjv1NknRol1n
4yQ2pfQijiVlsmT5hVVM2zUDQg691YMyd9ZxoI52ya+D3BGcr+QAGFoUk1l08aLisKPYPC8Ir8OT
WC2ymmefEUoyjs1/h4c2UecSvC+fBiYTPxpWHeF3k0ECOoMtNbQ28lFliXlIioqRVgYisHK9jCWX
qBbJYJDwEQXZ07Yz/4qDb9g9TuJbvVFdhUGvurjadRxKt28jN4jqs5ZMCC8pDj6cQRQsTHe194aV
T5BzpCaVnvHmFmNB0HBpnogmlCCk25X1BQv4Dr3ESYw1IXjDJ8IsGbVJYV1zqEy/g9BnQLs5GEv1
CQULMJWr+Fk3wGfPvac3uIffehyiqv/5K7WtZVXWVfEleJqer63c7CinWbvMIHWq5lPXWi+5vj3I
kFgK4N3y1Owjdnt4GuzMMmKxIf9vBddzQD8KirjEH2xl+bKtlwVjecwhWvsOGC2tGaMxc5QiHqXF
tKjohNxYSLSQXT84hbRiI+p+dCUCul2xoXQAxmWV2z74lO1373ru78X5o9Lkd93i59TdMq7yPLYM
FYO612cbI2kXo8vYV/JlGw0XMwdB6kqk/LolqZ1mvKK+3HNYcIhNgYFWrOaDPV9BNLCH+6yjfjMY
1uxB1ua0UlK/GzvC2gCbYOoyW50SxArpWIQIIeMgxohil+3Rc5J/n+9bYIwfpzSStA8teksM8U/s
buylueJcDUm5DC4vZZaUGZr3a8z2KDtWJkzROxLiNnysYJ9Ll91g4Bo2dY6InuRfmgY9TgThmFp4
jcifJdu6VxMnhGbu9lmSkTC7sgZq4f2KostpZzqeRys0W29ZNA/OzxCxFc8hnKVpknfjRKK/V2za
qQXggOhhoIu4Zl/wnI+e4Y6zaWpakegZT0sHqt1oFySRCM1jo9IUcbwGxChMYuqkO2WjSBjPRYKd
e366m5w414nZnfpr9XhNEbDriZPqO6ZaBlt5rN1no0giIs0c9prPmm12z0+CFL2X2Um9kY0VhfPm
zSOL2HX8Bj+0ayrwhIZFmGacvuBF/vTXBEnck9fY3SrxnA7cHpPmQVlIbAs7YNqocnGnep1zoN/Z
Yh/yZph2bevi9pgONyGFJ+QOj5wGx5knKjblJy+dUexfxtBjKAcyAI+ZWPkvOclgMKTaWu8Dq748
j8tm2Qq/zbvkMIdbZmlW1iX3b7FeW7Fs+e5APsyKzPc3xXvCDsxFBGUg9P3DUxk+SlXQJEfKWYaj
Rv4VjhaHJh+e0lArYIZFH8kloIxVhlHDLfF26C8Ox3qvUzxfz53zprIdkAH2y7r4ngPr0fhPIIoR
xqpeqdJSW1tfG6g10RBebvDzDJkTiguy2xrWrzThGLzfT+DTIs77fB0mSN4IdiyXEBjFARxQRsLe
j3HiVkla8wdxlM1yOWs+PSDPYXBaF0rUxr6qT54LsmF3d9N3Xco7LK2/KNp2KUaNoPm57QrqLXjP
E7MB9226ZnWsXlSPj/j576KQjPqEh8MvDPFtU7+G1fFw8D0eqaQ1wPAYO3GukUhLAofF2lLrbsir
0Ilxj593Cp3x67o46bMYQLO19IzvtfCDyeNzaZcvuFpkgSUCk7qJt6KP37ixNDLDbDxfQRY8AegB
kGwqVve9N/qr+ouACNzdmMkxK1Yj0Ly9wgshp5HIZbyOyTUTYej1MuxfQWU58kZlICxWTGwzPLP9
xhs0k2xJPgiS9x6wmvnyXoqDTFUM8DQEofv/O7qFrCsFpJ34qwW6UcqJJKo86qzk8c46OiF9lnAK
jwgAwV+dtSdd4Ir9FJmrcSrPmvDRx9fwBuUnuJUnlcRnLlN3+pUpJu3gRGM69ILiMuAiCS+P99Or
4U5zqdbyicTyPgzpV10wtSkr2idwmyimdJMIHviyQUWvXLwxY40EpGKgZtTMntU11bNuyLrMnMSB
/PGOdgJ+qAn0kCJOlOLoyI/3R5oiZ5S3OSlO0WgimuN/Nex/AtdY5dkOpzISE7TvdGpA0v6QLo0C
jrPJz5qqV1ikn9NGNcvPZuEEgAvkn6OkDbaa9eW4kgxfpaC4lFaq0n+tQTkzA8CojeP5wIaHgPbz
XnK02swuIr/Xifa+rt7+b82Ypn/D9CmO9DK6eaaidLqn3T62aP+jn0UKofU7zYbbjEjSRpRe78CV
4OVZ5PpF5FwpU6lu/iuDdY61cG2g8gHBy80ppWXYSdPG0uaC8Mlw8UczZg+kB1/QS5NXuyiO7ZJa
1oeKzVLMobz7UK1veODP8rKmNT0c8FB6pW2ai0puEp2mlTSGMLNw2vqrTEOTO6yLZge/uOg9qS7b
oxjsbGJIKwR/qjCOBCzSzGsE0OYnn6ht4Rhs5zsPVkJIKZHSX5w0Fzg9d1UlbNOPCmBAQqxU9Ru+
IOW0d/wK834axtyvdXu5E0c3jnKr0MLmosX4sHnz5lxfW4rA4QflKkJ5ln0+hIPKcK9LOmroJd+6
YgPvm1Ukkd/bWUyxa9r0sCivnCBo6MJ6FhWl25urvrgFtvzM2RF6yR7Xt1OkINr51V0+BbCBLJbX
XqhKA7cCtq/acNI+M7zQIde5hEKOIzdnNNWDCV7Nc+Jpi3Er92o8KZRVpbYNxWk1HYzVRvdsG4MM
Ajf8G7F3I03mxYxZlS2GGo75FkysOwtGDRnDGpaXLL437sj3i7DK7C4o4Bh6NRCR2Bn4jEIHE5NT
D1/YbiCoV8Mf1Z6Oyk49U8MgIauRx88hfpIOIESuEfU/dAFaDWihWy24RrQ+S+yWp9a8KG4oPF8Y
p3oTdB1Ajvq6h8zr3Woj9jHqAGM+MzI2B9FJ0loPjYeuyGxjKBEQb/p1DBG6Eiz259yQLyPZQMq9
waIY+9T0DvsMrwwupPBnsX8n66gp1m9G+H1jV1nnGu+fnEplQnvTXCttbYTP5Q5fCx0KqLG5IN/Z
NDcClso81niaj8OfKoFTQtIfoi08OMyS+OkkAM1foE7+x4PANDAckHKJyFB0GG9buy3Ulb6XltR3
GYm3dZeMcPJ90oq1VZ/evy42q5CiF0kj46kGIZd9Mnv46z5i89sRSnf3Hx5My9+cRuRjv0z1fCWu
eU76I655fmdUSab6/MuHf9TEgjJ5IcWqUovzx74Jj3+a4R0R1iYYZf0hQzk9T8i9xDD5hUG/OuI4
sQEKzxuwqEt1S0pzzPu9AjUZLqiDbz81R+afLwThAuWbqPsfAgvE8DYXHN1id9vI6dDgbxLeK7Yf
MvIzNgL/iK/ljMKNjxqxaZO9gyQt4VmsHvt3R6p4D7CBJeZMCR5NGX/bs2F3hnjf1jpJNun8UJJk
u28zS+GWwGWDoFUcnQTOCJmztJ4cq9y6MPMZyn4GQpbM9CAGvJEtZcEprqkABVy3FoXrrNbNepCp
byrtePZB69tzZoq+zK+r/iKeMWaR/a5miyDhgWNJsE29qvCxVHn9i2zTrvhbwtT8EUIAlFdOEizf
aKWiQl2G4kP2kAZecheFZ1/w7eCNm5n/Y4ejkYxvEWZWkzg72p1N2Tj7d4gTFteZJh30I6b/N4YM
h0IL6m5IXmaNX/WOKn5z5M0dIfJmtc/ejBTTNkXnveLojJD06EW43+vsYN3FTS1MJVeW9M9LHlrw
48WDWVPZ7F8CW7ltgLf2xRJURAF2ZrpZlrYQlq7MV84WsdHi24BSv/t4G9z6v468bUiukR7fUWQ6
17efVsJQbAj2CGCNeBl/nwWAqL+b4z+vgWJ5FHQ+lt3OHM1BTlSXuJSrYKvHRR6kVxhM/70ehtjF
pAlIHkMkmdQTpaJAQUo38q6iupIZ1QrMboz/QeU7x/YnCnJH3U3uPH4aX9FiE46z8OHp+5CBKGSQ
gjR2WbIT5s2u2FoDjGZ/KrA6I9XZQ92LtJaeGMKa692y99D1SSDuBQOi2woOst1FYpMkIvWTbrFc
SVzPTWkMkBGQKv5t8Kf/eBzFgno7TbzEyMMhSEoBV5cegw+THf1iTSfwP2tZtq3zhL2GYugdRWD6
ON+jPsNaRnjHQyyyTw8jLl2KfQmJxV+T9ZcOnotVGMSwncLPTY39dzpmFhQ9bdP7v5ejV0XYcgtb
Dlv2vTrBRhI3W0hMoFKc1w4DURaYQmNQARPvJkY6xw4u7f35WF/xajIHLfusuBzIlv2sdpVxdGM1
3IEmYDl2mTOCI/ak38L0p+b8ox3ayzfx3+eCCxzhaIdF/g5lB00TLLIeARKpI3MLdSg0K1l8PWL3
Tqsgwb0TObOx92pcyLRTDtaCf0NpNmudubcHNyMa47mraLxdWEfyF6vUcC4UTJZSS9ICw58sVRsa
JxJFxnNDwhIDAIj8+S+z446OxY8l4d0msmqH4bGjp02sdOiJ9LDe9Fi0eaKvhQeUhp3gz++LxZif
8r2U+u3cyYbgaJMieRObDxrQt7pQKyasVSyX2ZdV4AvB13FiMHJ4nJbtJ5DqQfDku9GuliCPjLo7
4mdbqsvwsTo0Nlpgfz5P789+aWW/YGO4mm9Q9tZ7KuBsWut6KPUhq7+4Jytnyj9GmQJEvHFbZzi7
+nNrVMXt7rkcEp05twuuKBNRRWhXuey274Fqtxl3I3x4oXi++AISWVJIYv6R8lRRqofpNO9WYJ5g
jM+WEg0HESZ8QYFlWsdMzbwLL3X3Kx9BXwcJkg0q0zWTo5E67JcCkCY8tdXsQd/PjW4rZYVxcLqo
KW+dJWOkEZ3/7Wd0Zl7eaz+u8fCHbxmeaFaYvfyJpji9rWxn9sWSpdwKEDzUfuqPPzQqjMU34boJ
1O682amCKeVb+RUFQkVScK9Do7EbicHMujU0sYY3umoBV/AvGYAW6hZ8yD1FgY6pFR0QRS4/+q6v
6Azt4SN3M06z7hxL9q6CpvMGMS7Jj5ofhPiW/u1S/rwlzLVVYMW0+qzp3odF9ejdWAj7y8V4o0K1
D+N/FeRIVtPzsFtFAjClgsqw3vpXzBsX/f1wdpg2c+PH4m4DWGTFM1H84EGHd6QASUd7fxZZuT2X
lrxQxLe9q/hT3HFbVS+ItToIA46rWQxuOaMSkBFhPNA70b02FaXI/uBT3EJou9gEahCsogZZa0pV
C6EVZG02xWPVpN3omL8qlC0vK8WhhpSCuOdW/tGUHYCzt3zylA2qOB8o03X+JyAOv8N+UpwNgs4Z
u6n/Qhx8QYMsIkP5rNRXOPYNoECvnhTArCrjO9y1VhpDDyU7NWzPl02vzGFarDaiY9wm2IvBOHO4
C2dmdmwBhAKI/sFW7RxM/s6AKhEBqeQIZon9vv2ftT5wYtgCHZqG4oZnXym9F07bH5VLiQexJrxQ
LjBA8UvOwCDHvORM2rObabIzR6Nq0qRqa1dJAac6WJROh2KS9uq0lD6SnZutV2IoG9avKAgGNzxI
ZiDNKtAUZ77MQec2YSCzKWtYBaw1dQ2Pe+H8XfD0XD6ltOocCzf1oIGGnTQAGWl48pzq38URNEyv
LPX4FLPMmlafXNNh8ZFHneJNt75CEo/snL00jE8Kl3RhL+JGR36pXszUjCTzK/qf+74ZmvfkNi/x
nE+cJj3ECRSEqScQYNZ7nqkiqjJN9pG+/E1i850BWxTLch0Du5CQtts0db5RB3G18a1NOVzAhwMA
WhiQrOslE99SniiOrOvt4O9H2ytCfXifDbO7d4YMPUXAjZZouTrwDo2Q7t/gqm+sOmgCaK87H/Tb
Ej5Wkc8zz1SpLDcZlCt61kleXZOI/6b14QPB/eWhlimQ9VaFZP93svBxb2APlOgvLc+De+j+WKal
piwZILVSXf5Kj+TMhzUy4HJicTNNgSRTOEDmJH3foFlARla5E0ZreQGZ4z/Esq9E++hh7wTQ8BML
4sd9M6S/jl/WhGMFMD2jr6Ph32NjVSAciSWC/FeGLfEbVqoTvw9xNJOjCF1BrCIwy9BKLIy8HFQC
WU2pEbI7IavK47RkbGJkq1fcdXZIwwcsq8eZrQYlXioo9REPupS1wHFRwgzdAjwzrw3U4s1d8LG6
h078OmYR6M50+y1nFpMPp84HxhUqF/EnOXmcamfWaePtJ1lYoN7EmG266Cq/UTCGQsIfe1a3+vRA
YJ3O2SQE3XtL2P6hRZL8HzIZRhjxuvkz7krwsNrwsU5F6GAGC24sSRedQ0KPJMjQscgUjH5+mrsC
pJOXGmV6qRwg3kAujkeglODCzRq+yxSz9FmSFkZcgzEKxpPRmmnHnG4uC8e+z25eBorp2ntmCJsF
Sl9L3yfQAnpfOyuIqKC4Enx9WFl7s1v0mk/JjW1oGxygsQ/OOK8lKF3axqb+cX/O6EjJg5gPtgUO
d7ad8Yilzbx1j/Da2SrCYovgeFGA4zQdjAGObptomMzDGv1wZngbFscGMGMX/khhK2Kxywm3U2OR
zOaW/OEbyOKC/mhKHuKbZP3lVIdjvJJ2u264KkQT6Y2Spt5/zyAu6O8rmE+Y/UrNKAg24TIAOOIs
2XnMtlivCB76MOpyps0FO4H7JMHKAemohq1lMG7+l1TRN8bmsYqwfqIGIA8Q7dxpnTt/lDozT4n6
n+risf310DyuSg9DEJPvQuJp8o0rGqmt8BlRUPEi1Qpi0Xj9URBE/WHhff9OYd6o0/UhwAmE8uDY
sEW/kb/GtH/8M0EOPA0NZ6Egv8x58oGOfkG90So0nmGUclhwoKdOG9ARZjZsZDy3U/XulBxP6UeC
beFlxxvSZihwV7ycJ4vgMzkD3ocTzIAH+uwDogFVv1mobEiAIR7deVg8va2JGJcdMFbfP4cWH3AZ
Azol4euimz1bcXgWP9vOGWhbjilYOOxec5bHR0lmHMVa4hUtENkeL6pUZPEDpffHRHiRCAqLsP4Q
zTsxYhNG8gbfhIsaHt/PL5ZitU9Y6BzFPgyoO0dwrnvwpTScqZ+4LBJUXnf/Bo0325j8+GqNv2JW
U5KBYuk9TEwOD0+ICN5J61CQh1i+irYFqcB2zfOYgIiGdaYMMrewejh/TdOEoowUQHTHwQw8U17H
8lxAqyQj7/JnwpIZU3M7SB1tv4xSCytCuWRNh8E5i/bmuIg5YhCRAn4YymZ9Y0Z/FX4VSPgSeuq0
xujiRKgAfit5E8hRwUYJOkJMWD97PHfm2JAwWgSXN5P2hRW8zGEqlXdMLyU5kx1dTDH6CL6x5min
ci6l8BQ4Kugn/VEj6x/4G6o6483tiBxa5v8rtDFdad6AKW5Llqr0L+to3U7er46ZgUNXuwYssPIJ
xBmMbXuXwJYljB4/QuB1IOVK6bXf0AwmbgrTC/FBUv3XzJStQ/iaEi4yiFh3TWKF0MK7VcYQGi7K
R68yoU0XjUvUODex1fUyuY2+sYi63L0I+QSo9tRdELWv52hM6WHFOBBGakd/LQfpka6mx6ZqgOYy
oeTuXaDuZijcMfTTzb7J6TFJTmqcuuXlBP9AjVz0+rORhkT8ehDP2IysSq3C4eDlx4m+6Ml1zf9s
TLyiELkpemCtL30/wG41HJXJ3uoLBbGxR0sctLqJI7C6ukInkSsocKuRR3TNc8Bwsnif/yD1HG9T
abSGsn+VOT+xOyBBwMiCS9EIcBQJpyV/KkuFVTPIvd9DM/OUgN9hRWPrYj8UbgDf8yT0iPFpgJbo
3CT1DgBzNM1FfiQQELmAQXFvwugsI2nrEDgWyGcYvLfWF9nKMJ4q7dxskSoL8mQuBuwDCPuI/67m
NrMd9Hoe44rsMC1MXmjyivYk0j1Gh/woQ2Fbxf1h5B++UsfuoYb4DYcdaXzB1UoBdrw4M1DO0tNH
cV4lNV+CNMy0s3VAzmM40Co6Re6ED/X6TsY8zoGLFzOrEjPDaCh17XmjG35FRdTdwQm8YfhIKqJA
6LgZxoi4CiBUXk7ATchPAAJoAmwIKlDNWxV9R4nrxaWthy8be3M4bhloIiOTt2T78o2U/5JyvKwh
sKpxSku4fhGd3ZAxizUmZFNuqofIBn2VI3B4fketmkzRUiztL/TgoWP9Qbljtaz3jCBb6yhzP0Z4
Uy63CUST350fxJaEr//fyS7oNQmISaFbWmeP1VijdBbBhjRbbxqQGL+PgnSuClWmMZmmRomDWr6r
lrl7SB6XRN1QmHUWD81jtomjy4LIUxDahzR8/o9NmKdxrq0PhwmDOLM8xEb4OZevwFCeUIXtNm8d
uPLZJSSabVfwm1lOqLMrk2NL/KU8jKzGy+XCx7XKy1gQfGTnLMXJh43KjXXqp1vABAUuK/Yfa7EG
C0JmvIJ6bcusV1n2Y8s+M346AvW04fLyQkSqQz9yVtkZbJYjhWgoHJPV+8yuTjB/LFoz8nNktrn+
ZUALEslIoluvwdpAjlwJ7SN86EinIeF/RtCZyiqZPsQ86Hpz1hxuEM2AiG5zbMo/Qmy6yuKXpYbU
zLr27YheMm5+UVBfr8geC/R1qHchvY+OBC2Q2/nxUQFysBnCZhE6bcmG12/IhoaUEn9hZsKLXEPy
bv+/vYuRdMgvRzZSe5IdZg6tifqsMziveW8zK0kmgjB1nYrwTx3SOGgdvAJs8ZPN8Jgw7OabdF46
fsAaJEZsnTwhLofyQUm0Demo/DTqW9ajxjg653qpsp/OpbwMp6MDSgOkGY/K9ps7tFFqCdgLWCXd
q4NbXEENdFCQTKSygBfcEafya2tK3H1crJSjj+KWv5qphQyC27jdQiVebVvX6Cvms39rSRgFQR9t
Ksd7ejMwgYBaMl3IcsF6HQ+fUmj0PnnmM106u6/O72Nd6fILJrw4e+sDd14MekPrQTrNejltsr/G
ngAKCtcHUNL9GmhRYgL1Ui/21PgFYWvlN3yghUY98Vf8bym2j5TRRoTdGHjLhZxPv+hoD/0qsw6S
1B3/H6TGWKSR+C5ekeKrbnJVGjjZkU1ulMC/onzxLNC3Gc8REsc3Hwpbx63MaXsE0TiPaRvoDpby
qaNeU0p3UEtp5vjvYb/LNig5eNF9yzGw/e5atZsVibtfUWjjDqiSBwro2NMe6fZRnfL/RVXQ+FKS
RDgWCP3hj+VEzXf3dVGLDTQXpC7ZtSlTh5+ekplYpvuQtyzzSmadPvRfMJ/kjMbd4Wsy/8d6Sp9v
VXkAZaBqUlUAQWt9+p8XgsuWuj/dFZW7TMin6UQRXBQf1jVAFbgmDtwXT5FUf7tBzwVuf56t5KpR
a7ruEU9dlnrr+n053dr3Vu3wKAdkPQD+B0eT+DdOzna7u5YVVMzqaDaEmbiYdeMUio4vkRCkk6JQ
j9+uGle58i6lPZxEuLcbM7aTuM/fFEApyfyzrrRIvGWuHCTvWkPHjPi9SMyqWAhLOL4zuAEkF3Y8
zGAIvzkg0Gn+3mGOFEl1odsYx0r7R2adr2wBZ2LCN8I1Wm3XR43EqB5KiB08dm8+p/3F/q6kIzFD
iOkkBfhG86dbfi6ahsOfVpXBP+1FD9P3+PSn3xszN9hJ9VbsIIhM7jjqhk7rMb8ec9DkFqkuYPVo
59v7szI+EAq8n+DVHLLJOk0Y2KEJAMBSVEOHl0IQ9nXkvtLgrDWp0l8Jlrrv4ggXAQ87F8Le7qXR
Nnj6IqsTlRUWiHcy845I987Gi/bopS4+9rQ0IgnDM9ZqCU0iH5EOrGdRjW6IVHThYkUDMDqnRDom
YuBM7AUsdGRDsdCUbQXLIy07Tc8uUplB9RlqfAtaQe88Kk6NGwPnrJDCL2tQlo/eTl1U9iM6P+8X
eSFrPuyREXu1eyWDKzcPohMwWwueOz5w2zd8xBPTZNgfFAQL3eBz67AtxKxOxvH6mh/DVSf3m2L+
G108a1uRxBP1tYYslQnNoeFdCY6yevF7ISPEUsJpmuZt9oiTifVfb+PmeSKkDVg4ob1WW6Z/InyH
AS8I0zYI6VsFVXtmrwp5mI3saZA2BVjiSkINgCPD+Cxtsw4ohcc++AthiTGxPmggXuko+S48MURR
2W0tSB7/qS+Bovh0wdhFLbDoacOqKODKaD9fqX3hcRgvSYx3wxHAEDp5jECjc1dTxz/7qHWW5HGX
EA/Kjl5ZK/3dVJsXETf8QVw3U7IPhlfQIu235VCIL3z+G2p0yY/VdnFfYpoJHCoqXQrGx46p6ize
CYRfZIecGFU9YKIsEfWGCjjesSexLI7ms+F0okcfe0WC26H2nICm+WUE1LxA4omLEC2+si/9auBZ
ChKAOJladJ/eJYRVY4nkRurYL5Rg3PqQeIj0LdEoxSDzPvG7nV7ZK35XoSpU5mIYIO7vxjQ+KoE1
/OXvWZcipXd1IxNnLvZGnOxHzkbCUNr3sGldM6eAqk4OGPQGmtH3IrmfGGyciL9cwdGz4x2CqKFX
DyrvdME26qWrV79xApeMT07C5xtDcXX130LvYNCnOFm1+0d3wzuWEN/vEPgHEFOdkqF82pG1unCp
6+PPpW75U81TLjzNTLI0bHtwTAeLLufJtoEpXQYupVBwX3r8shw8ZDCuTYWlOn8mjCsWHFEjBqTB
OM+Is5JxbefFpfCqdjh7zR1Eid9R4W0km9FFr9AcfCbVPP9sDpWGrELnGQurOyelvpq1CZJjLs3c
jUObBuDzL07wPNS6LkwX98dMdufn6A8C6uI1SQsevuH0S7s1DCuBx995JCxJPCAFwdDXMSXrgp3h
piJZSHdoXkO1ON4UgLh096xBW1CIV/4wV2DA58brhLJ7WPxSSTZK/nvNK/jjor7cJP5qHf3kCPa3
/PF5FSZbLWe51MuIQS0753abE59fO2d5+1K1VDR5arTQWIeScgxh0ZL5zJE0kGXrxFhcJrLu6VXL
cUar9k/9PpAMJXbdLuzVCYql/fA0g2joKQ3ygetnXgsGC3hrLTrdgrl2d7UXP+ykARvqH0b1ZFL9
PxqeZw48hGuyMT/KJGY7BIgqQJVVZP/fWMZvayGdIPPX3VjC1Skw2LTBWa40zb/dlg+USE8ayIQq
Y/nJ6IzpkJ1NnkA/Lt93Z+DzAH+SnH8xBuLyywLMG4dMPBE2DtxzacJ9xKzIs+rl/fwAm8RXz8B2
1PO+AbwPd5NC82D7ElpISdq35Lae2os1YF95K2VMAjl7jc1wDx5Cy2/uxlvlMvvHODkPecR4Lx/n
zLmd6S5qfsO+RrkoEbckEoakM/prOV2jjbibsmdIt4FqGagn33080TnpCArm5HP5GqK5KASQGXSK
kJsu9/os6qp3+TItLHXDVbuSJMo48/SbTNxxRkhtQW4RT37csq+4yAA9h7YuHL6wFjplJ2SEjo17
AVTgi2sHjKZxrqEICz9CmYVUm1zVNibs9P7Zi4MV+AkJ2SthpnWU1QFBQDZxYcefzt/ekJzVSWPd
gnq9WjFLHEjnB51iDLxiL1h9WsGEsIeMWQExaDUHqcjeronzbd2gnOGThQtjKQXSPCC5bgTl40jJ
mX18xj2OJBIPOSdbe+KusBwyEyd8dHghiGRzE9pN8M2VohbNjmWWkFAlSr2Y8p60WwiFzNv8Tow3
y0WbrwJAzspGZ1wLJIPBhDFtvWBxKpVFspqg/+lEcjSm9j1D0MiP+4lGfx9c1794qIfYkNtcqFwh
YCTQuC1qCP+eK8eUUdgOi3aQUhHqB9Kz4qkCVxBB9nGZf3jz7/Gk6xTuLev9qIV2dybzChkSQB0c
zEv+99/2UnymSY+oa7c1e6y4/F3kzG1OgfLyC/Firj91jYwfLaivKFBAknUYyIBJS3eaL+rxMrvJ
77feb0aRwtULWyvq9eM+wlHkw2/lhUoiYEEdohwP5MWNgxsrcvDAL/02bgg1N055OEEcc590l6eX
YqLGuXbw4Onhqgkf/D+HArXaOj+N9EBbqF9NfOvzLnNoDHF4Ac/k7PbZSHhBldEw35quu2Rn4rE4
RIPAOTDw+6V6EchbLdZilgb2l/QROC72S3VoTu7AihVHxbtDioHfLI4MZZTMwy4XN8ZgInzlxPUX
6vaWnSJ6xnW645mvr7Nov5gx7zhfz/qd2Fc+ErwWIdbMHqnJDE9OwEx07WE1HU5hZQBDBJowzDtL
KcPuxxZNy7GM/4stcRsFQ6AsM4XEYHLQmcwpoqoKdE5rAa8a3/kulH8bp62vxv1B1gof4wXqIccH
350SoxG3zy0/6pbEo+EJYzSFxZ0ziLXFvFNPpQOIKssgJBscomFhLD0SmPX2BPQK2QbTI7H1wfvA
8jDyAhp/YJmQKgLBPjAv4zbjgyuqmjBQX3b5o44w7NUiOnAPH/Oi7yrh2KvITXK5M8FusOIsudSp
5i6cX98IwLE+r+u2NR3CtVuuOlX7zUwJmF1YTWY0s331aIFpjoGwQOR4c5G+gnnuqk8Bu6HY3wZj
b+g+yuTCx/goT0O6JOawsbuD7VkO14v93YM6qBfG8p0MnV1PxLmnetF6xy2YfaTHDOfxehKM9HBu
OJgMXCVUqjWpIXy4r1+C/QXwD6qxKovx37OjE3he0OQu6mK4gNrHZzcSl0Lxv0N9KkOoBVxCwSOt
WbJ6yqnyjxLBI4leWSbpMbwewSQUzHvEBAJY+SCzLL9JhXys6x+k12JA3Ljbac+C+q7hapEa/gPk
Jr7TeZz7u+kcm0u202zTD1S1Knla9UJGzks3JBOA+coPp2gXrLfSL8Q8Krl4LKcYzb17O9oM3PbF
Mx3DyFMMaPVBy6YdcmGtRGgZwdRRlEl/TbI52oCJvxIZtvbi6n9Vb+6ozesOXznbYsox6uKFe3NE
ah8wWE+QbNtRJSxbBXvmhwvPXKWv1B88GHQAADMV2C0NSx4I7dgdAi64zZF3p6yhUnIoPI3nnSYH
U30X/Ehmn9h9dvbwEGpNZAxorgIk813CfBjNDfzyroYtFqNSwOA+RLqpWj7UwNzVgFDN6PKX1lfT
i2dUo9difFF8qzAycxRXneh5+YNlFfWQ+mb/BA+Kv4RFpTd1LVI94w4xKHpjCHs3AFLQw4VXYnT3
Icx+wAcFEAWZPUxd61vSyAfHA+yhBKbzAwjLiK+puwIjHYrb9XpMwyBsK6kWNmkGU0g1G9cwZJXF
IU7Y8a6d+dKJf+rqspZJYlhRQAsPix7D1mJLuvPRheaiKU80KaufBrkrcJB3MSfdselpj6K/2irJ
XgfmG012E+gJFyP0wAcS5bbgeidOYJlmZTyzh4zxAzGBD5+JloeGJpgzrluUVM5rG3KZ4/WPpJn4
79uiZGkMDh+dGLiDoCj6Msi+wOtnW8giyO6tuj6NFUoF3EDTuyzY+xHRpaUo8tVMx037KtrOVgU4
0WUkysV4sprnVzd7+bGP6ZPsHQ4qNCpXyQTHWrQRGcSghNC4zxoweUecDicCPk/37b10Wy7iP9kM
6DN1Vjl5W3MzBXnP6ucKpkbNdl71oZNTM3oCxlaSE8yT7Kx/JOvBJa3iegqNIMny0GCSopwhR8EQ
e18bzxsG6CY/edgK8OI5fJHTT/9X9xErbKmeCmYBbNGqse4k1yfz4z4s7TRbd4W9QsjcERIo13B0
CWjuGlK3QhdcqS4pyooMDbZZxTGc/TNJR4TVZtzr2fil9+KRyv7zCWHRlSa8/YbJMl64W4GDVhzk
pL0dy8rQi9Uqozcu/mfnV917hHUQfK6naP5vj23YR1Hp2hiO/cT5wzO8kih6F/X03n29dSweVL38
Ngy9UpLN2s7h1d7vqdQzYWaYiXjKF1+7X3KdEJcEqI8c+qfMrs8o1TYcrjsloc1LwTQ8GMpmm+nV
EflrW6SeeILLNeRugoicSNf6S7jHLaQymC/cjfUAiBHEz7Z60KGty4w/i8gA7HnOrWq77+iP5xg4
0sfret3UD8cev0h6ekih0hx/C3EHMoWHQTJfcxssLKQs3apip1rSmOfCIUalsGX5U4oiJ2JkmxFt
jT1kTYRh6F+wAGjhbxZ9vpoINrRB4WWipBTtRq63LQV4E7hqWdxvUoga7E8LD3LMoMnjRb8MvXeH
JpSP/B7PNFjtOAwoNVrdz4mxs2v/XNXgZw+sg5ku7nmV1WuPsVJZcIAu6YNiScEQMnhm4yrBHppw
+4ThwxTTg3xADK3LVnpQYYEZqy2wznjgDmu/qzNwtvInfcwsxLukKX1NHSigc5jhe0Lz00RTWeVq
05Zb3DkXwGUMC9WNtFMxWZ28ZKeCYfEYofBnvqGsg99vv5PAhX6uhAM1ut295lVIUXpdTUQnO2Uh
TKgNXO3aPt5cIN2U40ewDQk3RgSUn7uYVY1dJhetv6WYkHjyrlR5AUomGCqsSVfLxZKIefAzvCq5
QVBg8mIjqKj4IZvJ/9Pwy3ePkr8K5TjupGTzY9/dWbfR+8TQt6hcHjYs7VreKmEhVCLhdysUFg01
hMiU1eIU5u6HLJ/yjCFvYouFHmevn07HdYepbv7wMbtz5u/u3HCC/1s913PsNtPHaH0SGL5BaPDw
tuxGFjS6O1sW5HTVgIeKy1M1UTe2E/fb+NL/jsmboofS3xKNZFR46YoRVZQvf8yvbkxVlIXW/bfO
67cAgqGzOyuvpM07LsnPhxFcQgjmHjxk1qhK54Y3x0y4O+T3AYiPYEqwlkZbxigOLHN4uu1ROD4C
tpyo9l2fDPl1VZSUWF0Wy6zzqcL2tet7KwV7NlXirovCxXixzGbhcMsUrEPJ5byZoY1ITwII/fJj
B7WCwXH3Ygwo+5geIIlEARWr4fHadoqzHS2TNhWAsH/nIx9zEQwu1Db3CsM/dhlEXy1E301TEY/0
3/oKgL6IOJnkPmQpl+ODGGOuYSFWqQH/tAalCUyO5nWjV694xPi0ElHvSi2KNz6LzIXHOO1pSnIU
1h8MSsiPY0S+/PVPFLdS/qIJAgxINMkYVORoclhw3rAh9S3bEPdPkMEhBMINAvc3N81bO0bKKCJ4
5jLKx4EP39i1M1/+7+z5d/9nO47s0HJxhhLPr2K2kBosDcmoDtVaCHEK2/ErJ1Z5dIKjsM5uDPxK
1u2M6qsFzbJ/s6aUPltN0P6Y0enCYmOSMe1/tflqjdQYeRo5K9v7chH1ntH86tebNH3iQcv28HEL
Dt+AfeAnZh54qDly01DbuNeCvsumo0xfAlSQEKEYNhkxQPPaKlWYDfmoHYs48I6xUFJlShoIsHhW
xjxqg2Ug423lFv4mJ/DmD5PZ8O+ah5cfJJu+E1olqgJbtvloIEk9+69buS4BVJ+zFBEbK9tYulBr
xO0sAqG4eyPT5WmisQJBZU1CzJizoecTuum0zIeR+z2g/E22LsphxXcNgIcajft7b3h4nNwA+KZL
9pLN0O/8nW17MMtyObDS8lzqAus3HP6ZK62XKNGLB8dnk1Qfz6ZMVzkZ4XgBOTJV6G3qWkKLbxWx
5uiweeFboSkAXoKkgSw6WyFUzogFwwr1dita/0iqDtbXrjF4bFhqqe3kNESdhTvTDNk9qEyhvIqb
cEM6t2I1ugSa/mDIJ6KtNYrkT7OYuKCMHSHIBmwzxtlZDVayhpokbrHvhLwU4DLhVVAnvb1lEmq3
XX3hRXPm/YGaFFH+5twaX1AMV7f5uQO8IGL/lE+KFe0Di5L2WW1vNxQ0RxaT4Bv6qM6AtPf3qD1w
hexGX/pi+Tth0cImA11GH2OxZtpTyPx4RVEc0/jx6tI454/i69bpo35lBILBK1lYQiKJLpMVk27g
t6Gz/Tkl9TELwTyYIB/G0RwKXqYyQOg3hOhLz+qjcv9kG5Irwrn0eo+PnUhl13H441rUh0+MO3Ve
qzOm/i+srRUDwMrLsJakKR15caCiZmbfuzI+BzhURv4tbf8IoGfoJHMeSDM63F0M+nHyGMMcLUi3
b6ZkAN5HfFYzJWB85fsceWzIMXkVHw0pp5H6PaOHwSqtv0NBPKRS2eLb95AOEpiXuvC7Ds6CruZ1
vrevDyfNQCzMuP7rXlqTWqBrOFi9W0mmeGM15Z/SRldIQ76xkeixDdHlbL1j2jM22bc7cUEZ1rya
+/bxBesmXw/Rmy5jCjRZc7kf1FOJkdov/4AYYFaMF9WvmMXeF0/GNe3yYB5AUNfX7JEGyKJ8aG9u
z+rlCA5Gan64I7PL23T5XG5c8tCy8JiqYhHrHTeoyyTJArPPTdgS6iAPsNkS8DPUIkK2cq/PDc8t
WNCcl7haO/Ev7M0NSRh5fErDZQCIQ/C+cYXSSyr+TbBj36XZ5aBUUeGpD1LIzs4tiVC2F6ube/1U
a/2rPV5/v+hGfh/Zq8eR+IuSpB0KIbyAjOIykZtqToOj7uFbXdDunZ3XSn8XGcqsdK0GsYw4zwyf
O3YHXMcLN5bZh9f9urTHCqaRNHsyZarja2MTJ2Z1e+0ArZZNpXSWw9jVDwA85ybhcFBLBkyuShWL
USSJBNbasHy+I2Shy7tjinrXcAT7v8uPtAOCYfqsJ5nZ5N5LVAFAF3L4aBWSvrxreP957PpyR5/e
AvudQeXXOU3et1EsHyzLSc65y1gObV5uNIesZ5C2/LrJ/WcQwfChc6VSDWvHne4JhRB2PlZAmIAk
3l0If1027e3NBJPGhr9SAN3r62gXGlIr2PHXYsOLcUxfEXwAS+Hf02Zw6O6lB7kSo1D49vOqBIhl
qucAxC7hwUbKjXUMOmq88bWtSbs4EdkevB249fpta0lX4e7sG3cTsv6A35TUYFIF7No8DazHoyZK
oqrMkIm4bpyxWWVk/8EzSSKAzLtb7vfHzxwTk2tWB+5WDf4TNlEUCOh8ppe8vow4Fdd6cBVbjZn5
dPuDVHJ4Ez8KkyIPtWqpO6jcoc9sJrShZ3hFzuyXVc2OgzXgdqEm0v+qKJ3zkAQGw+dwyN7NK0Xo
07Z92sTjapnbMCjKz6ceVri99H4H3jjspVeAzcMvvC4uqdDNWtsqkhvjH8V4N8miUlUvgIXdpzc+
wNPhj0KkIWAYZY90UssWmkrzOC2TVS/maWsI/ZKaxbYzdsN4QkBzTUvOZUoZbmnoww6+Uuddr+2a
7MwO0XgbkssceTScRIzdEubBqFNQRl7uY0p664mhyYeIj7pP2qrc2vFWPPYR+CA/p13XqI/KFtP1
Op9Ahl4beJiM/5uNN3FGe00btCjYJyhQcZAOujyYueX7gu5hb1ZPj3OBJGaKSG5mLN2nay2pBPIH
kgWaOWiCp4mSuIRB0GtOU8oU3diAvcPlJnStkrCA/S8TlGEEP1I1IBtaf+CGZ9lZHu0J3zO3xAXS
gQAxGyeZ8vHfcM0HnW1dPCZQycQyr+luZ+57wlySVR5/CR6KRONT+cUkKvk6ti172bXRIfYw2x+C
lj9RPmseRgAyfu2EufxNDlb4pYZayOkqS0lUm2Scije6CUaIVrmH7S8a9LORjbaB+VlqVsJrVKoU
HO12X0hp/0L7bJH+5Bu16sU6/bSPqeSzoRBV9SsLief5l7TGM7DYd3j5Hzw9LIlYmf/TVoRd089R
hgPjGRR1hJ5vpPsa/vUq3QNJByk6ZnSkIAFlEGz7A0mTh1sMr6SKg6LYHLkpjJZiFerrHsGxL23w
e4xpfN/NBHwiJ36q3mK3PN0r1jVMYNqgQb0YdA4PrLSS9Z2I4DzDz67eVbWD3jJyilLpdvsNYdM1
lBA7Yd4oaWHEdvBsi+HhLbh4s4hDXyV8u88ClB38F9uBmzlPVjJSdEiukho3oZIqG/lyYhcL5ORT
ZVk1cw4uE0r0elIBK23Z2xT2K+DA6MX1KhuOw7lUXSDkXdpTvM801C/eLFriYR3OOYBm9dDMMWDo
GrW8XWzB3OD7Iflkfye+xQ6SZHODdwtkyvAiwclPoyBJ9pbmEvJQSYlEZ2kesDZ9KERUux2Xf26i
npYlP8ZRJRrhNGu+sPOFou/u5bykf0c94OE6YX1PcMa/+kRYdzT89dmxoDwAUyWCbjXz9FcEtgpJ
mYrXJz9BFmMT9nhO2j7QquiKAz0Wj6k7j/PyhiRcj88NiLK15PH4vH4nsNIl+JFo9pKkw5MHbBPt
ulymaeuOL2gXNDAwZd0o19jD3eMkuyMSXQB1wkXNnk/pdLkSTpFiL+s+XLB88LgpdP7Ft/UhXYwC
i4kEhWO6l9yWYGT9+FtP5CLydFNumuQKMl0Y6IMoUPv+CCAW9Z8h+BOdwrzP45QfTZ/lGctPfNCq
hJEvsv9BIMhCa5xm+oCu3NyHpRRr1yzhvsVmjHb6ekbmVH49WkLJh8mivYojWNMKuvC/0GhhIuR8
3vC3G6GHlVtF+fXPjDxre5zKpQTugfjWsW63q97f5GklXrKxeY3r6PSt/Bz1rFbK1XQV33m+HBoa
Ys4AIQdmMHa+KxCJpc1VN4QIK7S3brSkFZszYlZD+rHwzoAGQDOz5hwt/J2ZeRy2aCF+0wr3O3X/
+CaJ2SJ+H1bGZ+fUqwOszfOH6/veE9LWJ4G3641ZLpu3Uv4u8ZL2qOORJGh2hZk5+IeiBzR+UvV7
y6qqhAfOAvJYV0PQSbNg6s1Cna5Z5m67JVNrOXTs5vHFHXclhbn7MmGfVFfGkkFp+F+wh9qUovg3
PPd/djRxiv5yUtft/xOn2VimTN0AHkqAsufnSjr2pzKQo5+s0MiwgXwKJ5OiOQ8VeswOV5G/8L2B
4tQSwEy/CJvxs5vRTZQWChe5m8xHekECGfniNKK0nsjyM0eJ4nLSGvMSh/dgr//LFJrdk+Gm2lCu
eouFd/1NTwebLCrIeEAnBkKijlwi6WX4o9pahWG0Sy8t8gwv9ykAkmfT9QOvNYXpmPZdVWRH9pRO
YjeS5IOqsXgaU5RJZqVrZyhPi0+7XDETHGdn4CzNbcmtpPiDm++VWDI8BqFjdWl/CWglNs7nW7Yu
5WL/BnUwxu+os2+8TLulwvMblwrhMFYUlpQEBF+3qahBfM2lnUJfPIwgXeMLDKf8jSEhNIwm44q0
2/DLw4hwK7D6xBtATmaxzhHUQYsrekdmuyGW7x/FDlRsWoMENEqPVtKl/XoGDRRQrHr/NGDVHjFg
9xPNtl7Mvf7UYeQRlCEIGzj4Uqz8wZ/Du+PLwTN/v+rB0uYA5A7IIMWe5LdiKkvHJkcE6UZwekw+
OpeAta4MBH+9hKN8A/Hih+uO+HBh8tbMkQNlZ/DNbfAUFyWLO7CCYx4sulKYybgYPCth58g28j//
ppmhXf+XL/QxzuLmQBHhQVZsdN1wkpl0P4aWRwTZFebKmxkTeE24DuqUF59FY6+VW/i+mRV6gL8C
DIGQpNUlNVJSke8FjpCv9JJldNaqCPJoI8Z+s8KQZMvHy67aokiBFRN1kMeLTBVBmdJ74w5StgmY
Y7o7ug8+js3DUj6cd0nhq63TlHV/v6gLZ+1mAPJeEpX1XoxD7+iYx5R+FdIm3p+nruM0DJSp3RXV
aJmc1NZC3GsP4u6HhW1TVtsd04eLSLbBycc6RUnE0I2W3UJy/hpx04be/KFXfgefDbMsnzHrKAi7
llh6m4S7Ef5YdTfkAYMeCv9AZ+w6jlkfAmPyZ/1inqwmeeRA7cGJAB5eolX8pGuBKBeN8kLm7N4P
mEVjFiIki3R/+I3XRtH9cuq4EZihXHJUvcUAQ5A5GbfyuL6/1sH9BgOT8Lm8P8tqunBau/j077bt
TSbCnYKRCbUAgsTxzNLwpWh5+1thpiyPV+DU7F90Tmbdm0tsM6OPaXdqcPMb6WnlajjFmUCyvqWQ
0gmx77tKnkkXp4oG5eSqQWc4PoWijy5u3j5I/W3luhYq3Iyf6/APkm6bgNpUxjm3zfmoAIbN6qZ6
JFLwn+2X+CKdfvGvYehHBE4v3nvEeb+16EyKoM4i7AsiOQdnp8fazqrsUx1dS/zndjA0GIKrnaB6
bxcvWMvh3181PzKzUjGwtcXp6hyy2oIzAB6F1lQhJW+ezyW3Ow4c+I9c2thKtWclGldvf4QSOplf
UNBcoTO6/fWr9QhROaRzCA1kzRKChOu5xO7+dQkpu2iL36NOBPcfP9AoM5e75pZ40x3kM4CGE6Cn
9LK+t/raPBuH4FFsRy4jrrY+Ly/4bRmCv8y4lanAU1mOXCgtDhLgXy7KZ2+iTP2QYAZVwTo04IsS
DBGGJpVFEDT8WK+aVamjNrp1FYeLhrhmFSw+WqVNPtX69X6a+qLewtnptS5+R2C+euUgnkorAc1K
DGk5YwibM3wVG+BxlNUneD/tN+w6S+DowxEcawnvn/P1xPOV+bFRS9fAE0C5Wj4l3AytWG0otZGp
/RogWhzjernRapGpE0a9di7lQ9BKcE0/nWaVo/jxOVGLZVr158bIVIfxH+ildYRu8hsN14jiIlTK
Bb+TcUer2v/T15BAvNZcHUKtBwfWe4Ad+DGVCJP84GtdHO/u+pF5Tn6881Ji15J4lNlj9xIT06uR
4GyK4CeYtDwhi+uycCdd5s93qFmuLNOoK3uMMy8A2Dr/ivgwdaQIyyN4761trSmjXVUOqvRr5uWG
oaCoZV5c2FdwpS+QxhDBbTFbIpRnTkA3+UvRiq2yajq4zl3ASjq3TMaBT1PpazV4qaAN8FpuBo9N
/fJgEFMXSnGJuzhgPhGEtfr4pLht0HgHSOVzwdzcI79cxdFeSS2aysEjxLpbSQ+pBRkOOivAVodg
KqTMDps8OK+QCxGdQPWZbnFnC+olphZy5aPGZbSgbBPY+UHiA0Zr+w2Lg6sWPd7WLesycvAXyFA+
duxGBKLcq/d/3+8zY+FqwHZ+IC9+6I2yUQFaAvL2MTaHUlSStHHhtPR7lae4DPuOcp9rD4KgMcA2
JgAqjYyxo6lKLQttwDJmsNrFvddGiDKdmQSioc6wxahx5NtAsBU8LoUYlvkoDCHDDR6bZl4f5b3O
ELvol5fV5TVNf3jEa5RykkFoNwTjBm0UXfcBJt84ypdWojcmyiYdX/SzC0m/STQ3mNzTkOOXZ/4o
jlyFFz6dn4knDoRj39oyrEpZWQZcCiskB0KnhRorUengm+TNNsOsllx0HO0MaK9OPSqnClQ3GaiS
pVyVBm97LMvfNkpQYBPn3Fad6TpSYlieVzVuszXPzIuNIisMO2CqtcJXneXE7D21O9z2cBk6M/mH
yw0SRBirAQGjo4tRGS9e3+DCpurFCNzZ4B3LsL+WjWKsy4xTl3s19fDLWCe9oWreYnjgGG/T/WDz
0vXmdKM8iqESpOwFfZIB8EAIhqMhLrac/1iOOtPXVNUQLnU46qd7Jh5CoxaXDQxMJJ7jg2FKGpAY
1RE7VgZ30S7cbv3sUYGsUuPW+FcUVX0rKTcBCp8ZOLo7APu1uYl7pG4gSudC97VCbzouS55jQzAI
OjXskxZrj4IrjOeH/sL7yYgPN2XoGhakTcyjaYXpyn58DyJW3drDe2ANWssc3qkWGZoPn1UJcGpo
X4ppjJlzodE+bCn42IUCpGiliCjtYqW94DRAxFSIrg5GgOFLAFU0hAKElyobPkX6w7Ec0vLHLgD0
7C+wb2b4oQFutni+CpYHRQC8XrK+RlMYKLHpmbDSyd1jTMkVqTtru8x6FhUAuWVeH4VPz1ylWU1L
Z0H18AhUIqQ28H4JS1G26acpWVj2WgpzHxpgsUrLkwdOayUJLvWU1894UhIT/OxSUzw2bTHHruuY
FV9IUh7WAAOZELfrioDkUZGgMDemJjTt1aEXHFJL5S+reDY9lWBfVxDH5mQYwUP4kfKPiS7v3Zvj
6wlbC8A6PAcKjl5mq/h2eoRZM37svyCKwUYbYHkwwZTnJxhsMk/hLHAwozBV1aZie/2qsix7HVlr
zYyq2VaOauQ7YiVm+fGrhtcUN7U9380ntgYB4eX0kpL6rGwaSLJClHD+MKhZP7QoK73RoCQ+PEwY
FpqbWi0jU6f5qM6EZwhcIl61Tr8A/8zdDoaCOl2t1Hr8MLgqtK7Ryj+UyAYq8LIWGyZIwatM0Ow2
88hD7fVgKKsMGdAhmsE90VtAHGb0pdGRqJLQy2MAh1ts+T5oOt+DmRdoR91CRVTZutBtz9FHTuI4
YSILG5mBN+0mvA39USC0gOC6VSoZBxJz0I8CyyE8xRhy6ahGpVDRg1SkbzCCYVtAcQqk9iudnYha
6zb4EGZexi0VjMD/Y5Ipj53PUk7XLQwnWCPU2yxd/kmuRyrSBOtb9s6eYBLDBazCGXfz4LL5LlSF
yfWt0bqvRABuNqbWVtTESdYKe4zPPxQHtKBGapKi8N62sBx/Sq79REEqkaWbOIZ+xMZzlInz1W4Z
SESxmH5EPP7dgWpcDIMT612rYf4OQm/DaBORyQvpECVgEcBf5/d9wVrLGURIwgIOIve52wFnvFtv
1mFnSQG85y/cUFOJ5rDAH1nFrVMqN0JzK/Ef88SdrIHok7un2f/tkSEV6FTxBDLZB0W5XnOr+rT1
TWcQOSuv2Ul73ybyhLKLDxyNMkvmtgBISiSIKQ3aA52D5eClkOvdopmBvdmv4b5O8eWoPosPd6FS
B5xN6qrlaFw15h6oi/EjWbJXF/9mWZN9ApoDq08HAKZoWM9dLKywQDeBZK7T2LzJ/APAx1HxkeqH
LfHoB/uFUF1IFImXd8huhkY+taRJhEqU/B348tfdwkYHG3vwt06JN5pdqLsFTMDOowfJgmTlmnSY
+iZCKrgJGvP1DoVdlEEZgGm2zgbEVm7hgLh9LwfqQOXeyeXkkPOAFKUFtV1fVpiLqbXfxb1ORc+8
XxwMGsXEDGBWKvpyoqUFJfOTwzyFQV4fWlV+mC6waOo2bCexw0wY68H3WhFu/9xRES0JYuYBA8kt
m0UAHqqax7N7VU6CzACJvRGFvz1WuFIVCDDHmjntCOytjY3h6vcG1GQJmnL4BV0KO5mnJBjaaM4h
kwQ6Q0f8ISq7gwxH9ByMNudkiNBIEfOwMqoPpU7dFWnOg5M1MPSAPNGwmvrINf5WxToPRUkNmHFF
GFudZdXMadZ3MHiDZSK8y2GMvkxQvmyOju6wf56T6Fx2Pp/IOJP32mJWTQ0gCxCK2L9E84+jZcgR
2P1f1WMy8sktw3k3xi8fExb4VQiWV9qj0xtCqZnhpht1HDsNlb6iHFiAilHqfY/DkeHTXKuaxwfH
PAJUYP5QqHI0fORf94mRIE33c/krPlu+ykW4MvJ0oLbMBczSuZDw7qhw1jLMSMTVwD4dKeWg0yMP
1E3APACJv9kalOJ47D49c7hT4pq2+LIsDrULLKfnJGpRqpx+VuXrkVT9u38UBjAyhliFWKULJ/+2
/uus++4c7d1RVZxso5yx+WV386Gu1DdkDXkpvY5Ul+LWhJCg1t7mc9jUpWWP7+SUeDFO+riqI4wq
a6/HoVkc1/0g5FZTM+Y/NTxR5UZefKqZDPszbGS+ZPhAMzAmQ6Xyc/L47WO648rzH5KWoA+NDGRD
Ze8EdXWmya2ui7kpTsYnVl16fMrbHhzBHVylCKwW+bzEnn69zqnyoRw4WCnSZk+J6no+NV1dfdMB
xb99Xx6RUvAFpjfHsoxoRzwNvniSwNSg+88n4yumrXzRPRlxgNEKxZqoN3CN3xlKUWebXslmBc6u
9WhdnBlq0FzVBqiwGmnKibrdgXE3EIK1cijHaAWOu9Y3haqqRE+0aiEBUdMdhQnvgIIlzYk8r6Yw
5HHXbUZI/hrBua7gq+wg+l54EviQYP9KoydVXNM63S52f1runPGr9qeohWB+Bx9hxt8/Z2sjhHKn
MZrfNxKX3aZc+7GtcUKIRQu1QDTgC/vXngEFM/FFUaqZLHyk8/Tguw6VuIjV9Dvz3Y6CigO5uf7F
eV1lSW2NvVNuoBmUnNk0WZTyxaMnUT8yTX6mHs6aNBZHoDHW/oU79Sg0FLaRmo14oMzBe6wrL8o7
2+ioxei+EaNmmj2MB1Ce7jt1HEJXReLQgP6Ssn0Tm4gOeqnSvR2CpGPGnlFFxPXuhOGVvEIbCQ9i
NPpnlXssUhHMmyCMeCNvtBkVu+/Sd1uYdZw56+WkT4zyi7035j8UORrUuSjofuzUKeCNze4xHVG5
50AdzrBzIVhXW8fP1nLD80+DPO7uu3Xr2zwUtaMTtoZCKhEKydiimnzv7tOMdT+m9htfjZQCRZut
nkH/nW7xB7D9JRx0HGHX6XTDwzp9TaKokw5J9V+zRKx42Jt78wbLCv8At1PuQKmQL4ufbhT2PYzp
w1j3W8bMGtkPCBMjp2z2tn/PBG4ej95eZoEWk7HKHZp9c/WuSG1G5EVaPNsOPvcg96Jkpmk9dzJV
WW+11kHV49UgGskkH8mDe3ytPu5UqfGEm4IAS/2RmpPWPio05TWPGESViRpXnCQsuKJtp9jdPcHF
BuxZh/Iugk8HA5UWxR6sudlLr/LzlxDp19Q/PnPov+wqD5vwfBW2HXypzceRqqZsNipoBHSfuP2L
M9lcFb8DIliJxE03IjlI57HZ/EpB0u77wnWYZPhWiCb3HGqlY6BP3EDlEHwv/PRQ82rlB3xYLM1b
Tb85sqHZ+LUWb0bR/T+0tOd7CG7l7QtHr8vnvticfTdaGYjLKfD7bUiZkkTmdE3GOEhRZ5m80szj
Ny4N5CXs9gknhB3BUdEWvez5BgKwyGw19ke77aYqHWK1fy/x4dJUJEREiLwSgACs5o/1gjCpGfJk
tQoxBNyxtgHwB6KtdPtQDaJA/xsUNfxFanXvbJGn4suGnPsWrAq9ocgJPifH7IAwp+g+MhAMiAZa
ZJnwp9fv8Lf04gni/IIcXoohaZAb8+roCsi9zup1jkBWnSubVjWarHwSmPZwJpJ1w1OWU31+FqE6
toUWu+CseWOE/ztjPYI4aY3sNiY5AarcMDXZKdJTvzSW5NRlP9WHjPLhbWWBD6KBUiXcdFEDl+Tb
0qm9oMFRfWYa223biTp7C7xn5DYBN8p1qHfK6VyHihrt9Pl025EUYKVvdnL94RJ2NCdqYztGqE+k
jckM3B2X1/cMVfm0iJN5zJKu+gtks9PufiMEzAMo62P4Ab6h/zxbzqv8460ZzG1aIU8sPmmRRCmW
p2ru0I/6GxzhxPR/48cRaJMZp7tbqrZIfjQ86GQwpB5o+WkfU0tqcpICpZfqw7hquPAUzcWRkswU
a4MQYXojVx8y/V6ZJkVSCTubZir4Ty9gBU9qTX4ianqgj/v8zNqIbDQ+N5vp2hUns/asR0jIwzdl
Dg/tGhtgmHWHcSroSISdQ69qGGSjsihlA9Lxl0qcf2ZPY+vW8d+q2PlTEkhUINPjH1pPNADNOLwp
DbZ2TEC5Wm4Jm6Ti7fICaNxkhGwEj+lD3Vq4gztxKTEi57GU7EAp59hJXiufy1UAF6ALRiEl0A/s
CV84nUQlpQc9ZHfphviu5Mipt+bvd3YKZyfu2yms8YTkvY/lY8h4XoijhMjOUyqIo3IFOZ9aKdkt
lpul9kwb9vVPXyTfqEyomYP64PUXxZIH8lTeQuIlpeWUjV/Oi8z26wkwiSNr1GpFE2j2/n3OdjOP
ssxrFbZYcA0tVC2HI/lIhVbxwJoA287EJYUJmHf6VQpKhKfU+tgZKqgcyraFGLl2y3fDYp1/jcwl
aFNi/IaWv2/ROW00QDCvmENyrWyp5E4S0cudUe6HdGxg71Z1E/FP/zE2ZmNeytGhQMEYAVoUtAyO
jUCFVgVuLuyZo3G3hVsleMEw+dMGPLHxAb75SOFlUqxNj5QB1dD8i0cSYdr7BW6ElAIT7rOVFeVR
nLgM5FJt97UnLnCbvU/aMcbDtgSv0dxSFLOknW1cAD2q8TUw6p95M9xiSo/+bWGWc5vTGpnsEAMS
YEyD924X5ZgG85KbeMh2SE2A5BQ7/+jw3a/cVRkagbipvA8O4h3rpQnq5XvKmLuTW7/8TPE1/0Ck
7P1BukIRlDBTC7Xfv8m2Q9koFAKXEkdQbRCRBzSqknVbWsC4orOCttzPq3dwKflVse39bUOk6ts6
28YQkk8ZvS3aOsyGxZemdpIAljtUjtbyv5MqUIul8ZUsJS1gI9mZA8sHW61iWpoVD9WBC2YxBIGE
XihRyA/Z9BlAy6zZyK1YdqOnk7sXx6kqCaHXU0SAQ00rEmG9NFT4WvXDaZMQxV9i/nb+c0rpl6D/
XPalyQFwf2nyQBXXteASZSfdEs2s+3QiCujBRyy+G34gmz2LyVJ3V1zC4k5grpPZ55Xh/LFkUEp+
yU2GUX31yWkCfcKtovcP2OR77cDQd8F+pd9NDACeuj3fvGqWG1M0aXOjCuRtkFNFeT+oNAygm+kt
XdGrLNFUE+mO1ZC3jlh7v4VxcbG7fzqOtHUqqOcsWdLjKpBJV9kUkNxw61f3rSvNhCkCm7i/n3jk
CcfP90pLimoBD4PsuyRPYTteEKeDuCGazuHg7cDeUII/pUz41nFeCCWZSWjlH1rh+VwMCX1gi0j+
NTHsNNidFlyGGPE5bZsd0nFvG9Fg+jXs7ootTE2gFaU9KG3o2xIA1ymwnhE3GxhTf45OFVlOsBxs
c1rmpHI4/MWWCYdwqaiQ7Gw15EU6OKVpZvOEXYAhHkfB6aZxKNADGLrRIuWUG3nEByMSDpgE07gH
f0euKuRnYlLy62xZlRLuQKehytg1FCbGcUxQBRVm6xhktOqmacibzuR6VHN+FWQlys7uObKS/Dwo
2ZrRtpey6+LyJgLzWgMR4xQEBd44V7MG80hlqDcUu+4OF2/ovegR8HeqsjlM3gOxL+Tbmk64Hs6d
DENoObfbDR0XPr443pOqbDRUFgb9g6K+EYYKZHOBbkoZbmJ3De0bLzLheAjhPYI2YOxVIeKe6e4Z
DfvcXz2jLDWK3IXs5amGJecqTFVgbwh2HQRAvoNKJTzPb/7MtKXcbHCj9xKt/WcW+MbKnweC8E9c
WpZo6uJZ6iMkoHj0vpZlZFq3pDxmNfL++rbotBzomD4pe6rUvgNCkVHURU8UCiE5KSPRp08d7xi1
kV73Vvjynz84ZoTzpTHR8TtXhDRK/XXjRGCfh308vBVh5aTHsfOJNVYwqPpZUUAuaggnxve0liZC
FDG3hmR5shjeOVYM+Qn4Se6w0HJnvKm7oDpcgjiw3lq7MtVdGq7JqbMMiG58C5A80KAvz4lC8Koz
iJYgL/dZn6A+qZ4R22P8MDNpfwGWjSRoW+JJMjUXZ36komIkEubBbttuyRCoJR8Ei5ECrUKz6lER
zwNd+RSXflO8aNVS/PrP8l/1HCqYkaUhkcPFMsopzj+C8lN+Jo2aF0XmblnBWJZjvFQ9CX82zyGZ
FINW056P2aSxtzEIR2tY+puv6dr8A9tsmUGWtqKpCqD/WfXUcBnbvfszyQ4sJTbUkIcLIz4IzQ8P
HEnuEQREzVNbwyxNOmE3oohht1pSjOOKLsRDiyyi4lpAY+SRPiXATinZco5ay2ZKhqXqCGlnQUzw
R1A1AjwjXHwEfxvvdhPJeA8AkxHsXkJH5K4Gw6HLJX49LIn4BpS1dhGcf5H8yDJ9J4dSjc47QVvR
EdMnLHimx+EaJIeGuRSUCeR7CdwEfQvMi9Ekjxk1CwFoLF26Npyv+EzMktLBXKhE1qvX+76LVENe
of77ByxZS53P66Twlh6FUigicc7v8CXgnukuo2ER1sg1d3WbON/y7U5DBCzk7/JN2/dycKIrvo7V
LisGTJ9TQGDZS1JGQ5OFQiZhhT/lcN29+P4yu9QIP9Yj7W6Bi/LnJQsU9Ffu0NqDMDDgdgFoPNYX
v6v6OcsgO9oP+mI4Zj4ZIslExCWm5wxEGGvPg1T/Hj/BJRBGSeaLV6pvo+4LRk6DYN7CkU9VHqm7
3ZIR1/sxxXGYNhmHh3M4hl9qb4WadLa0ATaPjFpk3dmypxBhotx2IKqNwidLYhYgoybc0Naz5o9o
sCUi3M+CguSU5x32mjTwQCQww5qhy7HKPWkV+b8EbMxfsY3H13Bqwf2M6bD7UJDE7TZkc3nsVKlm
hAKZIq3N3lDIMzN7ATsliD4z5p+nF2+Q/yalSJnHLFhkce5EmGaPfx1SslJgYPxWxeDFnbQLPPgD
W3Teay2OX5/xRLB/KYEMQNMkgIusvUXeF06GvhRzQi47LesaS3KaoyPCqRDv9Dn+H6rNO6LtCrgb
VNuZiBsAgMvwAgPVgIRHf7bZqxrTMeUJfRxMeSha5dycoorgUZw1kgnJJeTuf9ReQtJkU5z6WcCV
q7xLj8+z/CBf2uS7KAzCpexnabYUP+fWvAsifQwwn5FSVzkM/wuBWh115bMNCWaZX9yan2MZ2IXG
xSuzpLNf6+DvL8+6VkYqQZG/M7Wko3njZUfpy2WoZJZaHPEx4akEfi+3LbGiDnqm3XcnxdIpFfo3
mC+1dV4pxUDgWthbiy/VCEDATWVfmeA5Lh/hVI4QDO+nbt01bJh4VIkR2UNaiRvPh/iPcsOoQiRz
dCf9FlwAivjs+89cpR2HV2EG6DJKvheDzWkHsy3YODochM1sEri72sZ+D1baLd1twiXMbdCNU3XA
DBf4+rJVNlzd5Y9ytmOem+JtvJQa+NVOutHvOLBpgRy/N1k5sxQ8rf5d/inilFMp0ob1gsPo/Ubd
NL46x9Xm13Bv9HV4zFlLr6c2xVtQl57dbOkgyqYfy3r2MI5ss6ehB5Liz7JVHM4oH3hg6c+PYE6G
FWBbwJ3R3lozpt1CebH6lliQmjKZ07H5bIO0rrb6KROHI8N1N2JAW/APy329vFjzEs0BXTPNBeru
+oHa7mynH4QLwGQCh6J75gHD2gsqnL56+AlQziIOfmtib8agVcHLAN9KPGv1gmpIbanJKpk+Wt/y
boQOoCqan1CwgVfHc1SBJ4+46ZVkFF5hsVaBtmFzL8f6kYeyCHmRHvQ+Ml2BblaI2KE66aD8qAkC
WU0dxz8hFEOj5JBWlorS5ZIgcwIcreBbFfm/h8lf/qPSKp7kt+V1ADSltp5KHmaOEPRF7SGtSa43
cmIJjcTt8a6vkcygWsoAVmjdxi9nG/tRKycCUpqsWvUSqOIcJpaVX3b+P3z/gJWe8jJK3t6PYIW5
Qb7++doF8umA5Z8ntHlf7lfNrwoqHkOHCuyH8GHnzH8V3kMXwvOexqQAPpTw/EzhYt7ZkqH1175B
6iYJki48PD5aTC0r3FK71Dak0faCj8I8wYRIFUWoFfXP6rihSGiZf0a7j6bYim5iia5tUTomwLOk
ntcrIMCIclVBYQEMTQlpQD3Nu2C4KE/BItHZP8MydPQWSyEfCS6UJ8VzSB3iR3dxZ9IOO/OvDCgD
rhZSRJVJ7CvWXPIiZJVMJI4IugK8kp23UBrTv2py66lplAzQ1zDpBe4y0nKD31G59aI/O6gCmJzR
GwLV8/X0kpNbTvCWfMj2Bzze4iQfYqch02ndnb40wLntH7AdHvKQuIaIe351DYpz0b1F+dAZYMYI
yH/PckOPAZk6g09tKFwTPGQX+TRIBwm7bDtre54/7aoLwheBz4F4BA/6cwXppWQkKU5zZX2FinuR
AkztiDEeMzLpMzK+S6CASas6TTRtNLEqzaO7ql6lOSdzRWPZNCYP2BFYj86cUxBd664ttgupG2Qv
0LMEZtA6OHMyEUjwumVMH3RAkBAWh2J72o+EsmlkQXNDDrLpfW068GkEqDdlqjhW7xFCZtXwRLcF
vO3CjwMfEi5NYR/4y+/6tJKmZahwHclX+qk1Nk297CEndtJ/HGEG13A6sY13xXPiRkv1DFFj7R3N
GtLndsmVt5dlYO2Q5FisARcBxnhriFY/MSO/hY7/AiSNqHxYP+aeJ3oSeVxvq7ygVgzgd87bQ0JF
bxxZPsfqZoHJQsaqAFi5uLY7aA6ooPCxRAmoSdMV0t3f/Af1hk5l9G4Mud/S6kl9loW/UBa5Lc8H
Tw8Fe+VKjVU7OOQ2f6TQb2IE1tzz+qUn/fFZtk7Xv1Cir4zkfQ/mR3BlHgUd+zGLmYfkf4AnHSZJ
nnj7xi0xkVirvrj9gV9PCmqrs5OlWLpm4eQSjmz7VgKn5ApgyYi50F60hxV5eO2wleRn8XiTQC0H
EA3d3hFuJzlDRShi72zHxvpfx+eYyobeMGkzw2Z3JzwVs+quNCIxhUph1vZ1TQi9VuM32lbnVlnh
4ScXxeqNdV467mkFxKYD+tp4avLh4t0T43uzghC0Pl5Hh3yC4uJBAWEoG5HmFYytRDOlakPVsVeH
svPjVPsoVnIOL4mIJJ/+pT151h3LPQY+uCWNxWTdplli7qiN788bYUS731XvazcqQvys7C/ggBtp
oeIJmxDxTwHC7flyYcM5aatIXd2DYV6SFE/nnLPCY3ygR9ryv3zsnlwTm5effOkZfzbT2fblMs3/
7wcJmnAGm7B6qtY8+q3I8pSceqepecwQRyWYRQnaq2UK5k5dWxUeL5RRiJbssCM1W+aMN0I6Gmw0
AP7TCc6wiXNOIHJHpwa2WgssrDRfsFTjenV1fwKb/ziiAFGRfylvuu5cpKe6KsbOUXbgKfHpcoRW
mnMBcIe1Epj97adR3QAXuAZnYw54gKfVDALR3zfuI5FmRo6/eA+a1MO/kt/mAjej79rjpSC947hA
szdybDker8f8fRy5E02YTAoGZMcfudn5aHWaLSGi+DlZ4gkoXMp7PkF0yEiFVdT2+D2obMIJ8ZB5
Echnv5LRnmj56sIAlTneTOlXDgCYrJyeWIOd4+/+/oSK6jrE71dHkTvfSeTUTLnDhKXwPIHreEg3
oas7T2xVd8It9vgfSussVDo18+SWpyDreyYhfzO1H8eMgbf/BpOysuXfpaXEGFyM3Z3VMg1UCPYM
qv09nVMsrwqgCS18jipeQbAn8VDL8i9Yrc29XKi/op3ay7Lu1C6bCj2nG47yAafKLbU/S5r3iTS3
uSpk5gVHykGqsyhlwljOsY9g0UkpjSofNopZPk2am/NzTXwQk27AffNq3CV+TX8MjRftyfjew2zd
463w40O6bXpwKd6uKCitHyM7SWkR63NJfQkc9oUPXZkBojd65P9OPbv3/pOkWrkf+ZhWgkCUs7Fu
QqZEj6Q4gEB5Amb0GodXqW0gtdf6donu/QFGsfOd8Imnblfl3Xe0u+d3E6kkfn6vFCDF5GTu0u3T
BCVrHI1OtJzB15JsIVSl7VZnsy0h8AodOdfbfOrW9EvQqtrz9V35nbbS5N4eLNeRBmdohLpi2m8Z
M5o5CWbBgmGqxLFDpVbs8lEjmrA1D39OCIOMu6omwBZulnlTwIgC/XNFNrnz1WIhSCC/G1GLR4XA
s0Ci4n2bSdI9rKUN8D/ffszuZOqdmDdrPnR7ogqPKIspfUhT5YoHFQmwmiiJzBL1bq7LXwGer9Gw
f8Yt79xoaQMcOd1BxeqyGmeCqX/QDhHXBFvTi0yhZvQppSXGUnbjM8l7vyFBXefYteZqBsNHTmLm
fmVXR/DOuG+vJfRO9PMzjKgsJfIEp29lGF8au1mmQgigA0rMCFkjj4pMujlqhk3k+Go/AJ0ECcKf
NUHk6fUGStAzhFevUR7kDDzGAsvPXA4Hwpo/NdK/unqrPP87TvrgcorjXOgRpfAPOowMlJ2MFJej
SFBUAA4As0mw41jySH+dTQBn7QM8pfTNQ177n1y1RsRVyMrL8f13bSd+cfrcJ6OK0DLvTrvYaa+u
GiRsMeCc3yXySpBmdhSOqpK/IJZ7gjH1FopnDi5AKmaq2KkId60sq2hrdXqgXuJjmtw8QSL38ca+
qIOd1h1IKRHyZjNOnZ47pRuSFP1DrUvyA15Y60cPc0s/1kONsp+1aEkK85NufqID0ZQ/RXIv39Hv
euRl/LIN9e80mLYTlmBjOtzePQ6d4JcM2sBI7oTWZruakynRr1s8vYLybrn4V02UOdYGXOUrNHqZ
qYJ9PidYBd21r4jV6XwJRMUiUr6/9XVur5jhGj6fDzPdp6X0XSaM5ftmesvXhqyZCA8u/bFxUqAt
WHYgSh3TK8ThY7n4cq49iBboCAqNlDpvx3uKI0sdfK1HUXEpnsgCgFdmZpBOMpBEePulP7ylAyQd
jDxDaWg9ZoguPEzEkSg83aCxYeLAGJYEtf2415jEk9U5Qde8VbYGgJC5J0vEUGTXhMSkFU6Vx/qJ
6DiW7QQtQANZa+XbGqg7778yv5S3hXGb2zm/6VodEfHHj3Cc68AxTUrtGEFw4nlo0KNLSXDd4URI
4k7sFqE4Ba5KRQLYqTXhIvC4LshLa5N6sCSRSKLO4IElM7EOp9JnRufAgADBSm1EMDLGMtWi/F2G
C+TUQzDDe7awzFdM6STgGLxgUHPUHfNRsVF7xKQGoAe5GBlUpjoINS3zG/kXxrVA30UCgBi+/cRH
SKkGDDXc6EAa98g1hx9+GU14jLwK60zZM/uQ2D2OMQEvezqyLgTj/MnWyiBV+l3kl+MysV83dV69
D8ZQy3es2V+v0tOMnJd7i36ha9KZTuhuo8Ptn3vGdcEZTfYz1vRiN7Tprmyft3PuKjFEkyBZfikz
UcrsDIbMgK4gAjYJ8wQ9TVzNBpVNl/6hWWvnMqjRPNrVZeAbxBvJncUPscF8FDTYBWF65e3YC8BY
yfVmGoYMONUtHG2RR2I9dGqNTtJSjEbSgc3Cgy+nRgFlscAmQzd4BPpTrmw0YVWjFR0j7hSv5zFy
NvWLO6T55w/YFd5D0tjcwqIDK/o+aysA/gURZ8dPKFG97nymtVDDEHAXQHctl8tvuM4FvwEtcF+h
DgFUPFiNs2KwQPXcC6Mdkc4OXmTjWdp0r5EZKFrOmJwIiymgYWX6Kr3bEO0ldj9+4sQUx0Vhm9gQ
s8aUXkujAOBozSP5Mnx4cKFSQqaERy2M8dlaPIgGo74NP8qcvc9Qo/6XyAak09FLD/xdlgCUgJ3o
0v2ggfsC4CHo0QHvJMgQKvMeR02y3G/sgJO0YeZIOOpvXWWKeP9JfwOge+L5UJbSIvet9OSEMU0F
AJ+0vJ2GOIfc/VvPimEI5vrX4BHrgtdKz8Ww4A++4usuZ4fyKHRR64+Dw6IiReRmGlB2Cn4C8orR
lGfkuQ3QcvBSOo06NeOzkU0PUAC9swf6EwfdRP/dyy1etp/miCXSdK17SgrWm1mGPDZx/3lT2Djy
v77H2wlXsYf0ddo8UuN2bduZ18xCSRfLldpJ3+himi1vL4V7A5V2ZqlCNPewj3YJjC+X/Uo59t0V
KOVFwfbFZT3CTu1SreFziBc/SEu13p/rlCgjz5bhmiZ7M/YcYMu3O1lyFBtRyya0FtZZ/yfZR3bo
MI51ZQgoKkyzH/E2u1or4hEzC0y3BZNQhBB/EEUv7UI/+LY8WdCC73KLOHlxmuVwF5+xd909ogMn
MZexlIBaSl4AwW8975UNMkrMHZuu5G0W4Wf3JwMgHXRHTzVN3LkoI2Qigl2u0VO7anSoDnHDnSSU
OVgtN9T0grWvr/uDRevsgEVLvLVE3VypCcmchPv0hzlWgG0MKieUP90o1VrZCsIECW8KhdQUzs1E
e5GqLHoW5gU+dGaH95FV2XrKRiAdeABVJImcqZ2qrk3oFm92jNQlKkflHMT788PbNnke8bxjwc5K
HSrwVlXbfCX6EuDKQ+Ckly9v5tO5g5+YcitGcft64zaRwh2OylIjdYy35llDW7pjN6cq79BI91M3
qRapQuL6agX4BmER8dD4JSY95eCYhD0jr6zjRwG8RLjx4eMq7YHObm/N+pCDcWql4/j2/NbfCCOO
cKENE1yLviC17Oj3y7ttrcpCx1UWlff0SuyLotYAsd8dBvONsyyppPXex7mzxKFHlo8fsv9uibnX
YQiBiPFXYSPKNV05yVYCBbx0gF12o1m6U4N71R9fAtPtlxLoaNdXxj/nd/aPl80CNhO1elAXq6Yk
TXyRhdh54cKQqYwTHKynfP77/Yd4RnlwTdp7pfxZInLbcyRYxAbMxuNCFtjSXD9Xy7sGoSpFXBrQ
OADBlEAtuWwCbzkFzWP8M5tp2Ijo031zsMoVpE8otFsIGjrTO0xvlN7BOxUm9XRCBVBZlN2V1UQF
7BwV0nFC1Y41eLI/3sToL9NcCZ/g8T36O8fc2sNPQDkx0GlVBRAIMlYZ2bJ8KAVa9B4o+s6pPKB8
OIhx6GE41mo4H6RIKRf0+VwIIvCJOdQ67tXbuAAt+MITcQcxQtUqAwsYsSNvsZ17AjR167gfbjnC
+CnCyXufnCEMJWuPNR4IgRyKPyqF+nsDfSXxRRbfnuW+X0eX7sCehh82bPqYHIhi8GQ5Cda0c4fT
XCm/4i1Trn43DjvcCGObVyAXQSbkG8LmMEeVxo+K9+H/1VHsTu0DXViYwRHsN24geMi+OS6z+fa3
RqQ2lP1LPdeSjTEKzpe8h8zTk9B0lmYcw0kBzWuvD85VbLCSxF0eSJ+FgNra/R6geH+YjDawdCbC
29WiIE2BznGapEd3oA1RaawrMPC1++S424PZCiuQcmjKvyJRiPxQX8Zd2uOVcXmsQCt908ikb9Kx
aUeSzqsM2z7I0dNVFauuGYIl/qAF0jzxIDVIuf2/oMd3laXUgQLEiH3MLADtjK59t/ZisAZwN5zL
Z609jOuEBpcHI2eM0GUHL6+bMA7yg1d+RbkVxDM9rsuhKkTXD7kWSIp4cQFtSNy9Tq57fx+EdnFE
LEimzUjJu66K5qjUvS6MsIOI2nauEZcBf/3X9plTU9dsW4C2LTv/Xbk12TM6wWM7tqtwc9dHlxxO
8BJPkQOXyhuCE84YJmi6mdQA+nFUDMRSN7GweDi8dbMaIg7iD05DwbygLc7lgdBvSmJBbmAcECbb
oOONZyzU2De3GNAXX94g4s69v8lGcZX+7SXT1ShhrKwc+2FVNg5Ve2gaCyAPeSt8iERscqGyXFEU
7K1OfB0UMhbGbWPFVNE3NP84Yv7ogNFK6oCN5C/4nm+QZ7nXE7IlT5LxJw9pJy/78YIyHtJTGNBt
kG2/Fw3aSTkX2SQ5ul81iCaeZGR6wo6WXXUgU7T9mIZlV+UGusjfJEqRE5Ih/dJSwe+cXXPR0p0o
umulPcgEFcCXHgQWv9GO1wcFnI5niivxNiRJOk5fNVdFyeFI1x2f/3kcq3IyY87FhDnfFfGA3jgl
lyP2C9VFeMLFQBsEIkRLt3Rh5U+QIq0xlJ2Z5+ZOBluDD8PbVkevP4Ii8xwJvaBDyptsNPWLLuAx
ELFILya1DR0k3LYuexWvtclFzLhdhDGeCSJj7a2trHoxyaO1P9AuF1b+7dN66gcDQDJIOtVF8uGP
THxyWOjFa2tTBJJbnt92WvRXZejdXgHWfYaeuZ2uyemIyrXQ3mwWA3dMDCZEPN1a0OLeiCkOUVeG
Zg38oDMfxtWf63797vTwLJlQiIBaqEWi62hMwHGTc6kw3WH3wEGyd2lsekTzGuBGpVRKaOfF1ie9
Vu95G9x9dK3NWwG8y4cXyCnYMZIe4l8za4+dZhJC72P4IBei0F20EtpPbSMqM46SYu8vtHAVHWMt
/lgvvOnn/ZC+I0m2RRri7ES7iGKhSNBqusO+oCafGFkXgT4WxfTiqZRt9ynhY+9Y5wqJUnivsB4/
qfMKuCCKgyRj62MRwqrFPaPDCF1MOyApPuUnpgruaV3Lf54j97Vk9Y2gVheEfZ/iFQyVoDmjZotT
RH56PEdMB/HAPQmJCiBNS1vkHL05nXBmnMo6w9sou+zFxyTtkoVZcUyvEzkrcOg1SKFg3BifeQkV
2Ngb/bTfBNDviE+q+B+8h9RytnCkj5S+5+/kWVG3EoGXQxj14PnFotras1NIQxpkLX9AZHPEIuJD
NiQ0cJlr+UYnYyM0BxRk6FeDvvG1T6SKcFsAv8oA1/4L5vKpH/V6KnXGaH1rQf1AJiL+RbSQQ+AL
H3fl5T6eQ7VDr8sCwsTsYf9Usmgr7FxBJvZtE0VCDmP2CeJ6irN6/dwZ8OHEGUhcSodQUpsAILeN
gLLPyHBhxq88bJ+TqxyPe6HY1JFSKbbV/FWCxks+AIFnEdpQ84pqvmM8clCzfys/iqtKldgsJIhf
L2kE+9CGqCxzQ6CpFJ8sVEagm7AIqezBBIb3RJRRVOWihN/7ri1fBBV0SFnqi5WX+WF/hB4OQoCy
034qtfP7yWVHOU/+aqXk0WF+NhJWVbEctaV7IVosDJ3feL9jK365kepysxt7LbHRCciIRhY3ZQOg
pEAfDvTMN1Sva9veDETXu4OM00oihiuMMsd+ceqJ/Y3R4K9IPbZmajZ4rJ2AzMRSWAmjQEYPfGGK
wZ27dq8mqxDZ6guVsHvZB1oAJKVeUb4LfC7RUMw/cPtDdTmkDr7PWbNjPmluqMJ0vLCpoRU9HurX
0MAyARyEfxWSAuZrjpMlkbZuZJjh2m6sQqzxh3t5rjr2pcoXQtDLUn+13+CUGUD/6F1CnJeV1B1z
soIhl8gqCZoGEQ2vdlBdVygA9CvJ9DEMLw/XnTFrVYMbTpHR1gSSXytyvnB+tKX0snR1aT1rLo7t
f73PmF4d3rn/6/mujj8otslTTSlMe0S76q+JSvT5Y+dKjREysMmmMI5qIgiijgpVj+gZLINtVDry
ACxKXjrXP23nJj7oBrYK3P1iHfwuyQCYLRsBk7Y+P31/cPjJpMU7DutycHKKrNrgb8zPLH26QZaM
MqfolQqEyNl7SNylELF38V/ucJQnlLPCTxkskI2tLrW3WyOm8VMpH60vOxZ3ugqZaAR3oV+UdDoY
j/oIQl0H/RHfYPZpy0yguqCPgiuwAd7G5QmroNkur9x+HNvDX3GmUXg5vaXLjbiM9eoNVhK85ZUy
tKw4TbFgGaYACnAzA5rCnn67w36XSdDBSq6uIQyUyUekqqnhqyWNNYDmCZIqPkAQ7F4AAikwYUVa
R6ynrnrV/giRHrvAwooQciCvMRblkaPt9TMQwns+xA5KU5hiupxNiELqUi4ihN8gJYKRLnu9Shhj
ohmntXkz+Qc13E5uXWPuWQeYFFd1RvoJdmK1JFsNgiANJNtGYwK9n1T9ninNFvFWD5TbvYuCwIo5
k5m/Tk2IxhLctz1/LPrbNTLqLDWYTf6kJhcWV8u7BWhRZHWRtUBzm/E6HrUami4xBkNfxe4SwJ2S
rQChK2wZd9NNnNXo4P7p+G+QuZtiV+wCDjiPmjomsza40SPSyQxCN52iC300/PaRZ/0s87Lv7mQw
lPPEVLO6qS6t+Q+dwqYai0nsi9v5iWjSUxz4nCSZ3Fa1TQHit/DIWyFcgeJSjDjQ7WUXr5To5Lrc
rLygajc0oA9rkmcpbedjoJX8J9E3KPISfyvwdqfurW3ouOn6UTrI/nyqrJUNT93RjmgOjTIk4wTF
f/Zd2zSoPcWMvYbL+Jcwq8mX8uwvyUU+2Yj70M5jSXa8eKP0jx375dFjKLVwsJSBSNaCtA4VFQbQ
I34q5CohSAFTIexIPYPMFy07FGaJ4tZMeXTg0kbwgvifRi8Ik6YPC6VN5k8AySKBxX8dkZKqHbHh
P6Xor+ddQ838RoSvrvJ4X9buDaQ2+YwXF5kqv5w7RzNGWi3o2Z/+0MudNvjSjYJNwcdRZpZ3fTe8
OpxA+sBbCToKmQG4aW/fvlxdG/bQ2zLJKow4mCOc2mpsvFPNR+kpBeKgYKIqJ6RsGtlOSGRsaV2C
VcMiXeb+KfM1JvphnoZHE9tYIF8ATPpPjiSN9pgHuAjEE4VTVj0bDmK/kqRfvk0pQNIEEs8O5QI6
b2U2ue5vpigJJ5ETw6oTbJBL+0CZ0IaXcHeldAIKQQg6Yjxu+XkdRk27QsCJqzUOzBvfy/5dwaOH
pcQyiIAfxo7HM9HkfT0RgKQMCuqLGl8h8L5Cb0oBu+KXqCVowtzidi/q6H6l8Z5JUwqEATSIGbFM
ZpGWRzD8uUVWmicKz5CVPzALYSnfuTfPCq0p1VsjQ9RM8wsVXD4chF5pkxhLQ+ZAY8ZWjNlaNwfO
JreJVwHxqPzvi0yvAK/aWhc4s1gUfhDGsIkCGvnB0SnMctfmhGrLvBYF56XNibcg8NpbzaZEjplY
5NueBsM9x2BQfDqGoYJkGcyuVslyLZznR3HpxVSbEJo5fc6mOqL/7ssjq0aJ/WEIlKbmBn8EOJ42
WMD7n7kjdd5qa1Y+DjTauACBDmJmwX/S7FC2UrzD39i41/9Cz0TA30ARSLO1ZJJ/vjjFR69DgvlS
pr27AskiporjNjED5+p4l4qgQy79q8hKkv+Rosu24bOcImNRUmc0TbFqfoEMTansJAMcOST7+Iya
xFA/w14N4iqHoCHVCRPDNQzEyegdGfnCnC3wNUWzh+SxmeVXa+RMRKJq4jGemnria5K9gYSDLFeo
brJSjvASlHVg1gr4be9lPeAixfWrbs7l4idq86VIn1oRM2mz4eiPMCZyeOl5k49sWHHI1rhIeWOr
wqKXWlkk81X8zpMAQEWpIEIt6dMEFg8sfXJnBpt76tqfMW/q3iJB5k3SxNeFW/iP/SRPV+smBYaP
RTP5QYwnjc1LFb7wzsmyV+7/tisPAWVL6co2UXLYb5QiA2dmFoVtfV7vvPzaFZ7BDNVBcEtdrKGz
1zBHHZSTfn8lTwBmZf8mrOOTHlWLfZ+nLGM+7OBm+ufaskLVSgzkSv+lWu+/QSyjhuyAOCFciajQ
b3VEaO6AeZHT8lnhGnHvrKY7GBY+PevG0xiRPL1Aho4uFjxDu/vwG+rb8b4qy4ZR3dmTdFMAoY/2
+7/PKDPq+t7k3JUsdSJ7TGP1dz/JmOFNLDOtoVB4imU0C6waCzUBCnp6HfCezdJoRQCcaPVKtN8J
9EOPxzTosgYiNGcTTBqu4Og6sxM9LbQ/OurJ3B/6Q1nSmiMH/g9H4wPvGgnjBsbbz4vyz/67fWRh
haFf0VtVfRhSqa4NZlnmvwrNWWMHl26IUnkHTiGF+XLmNscuW88Vb7tR1Oz8I/cm3lffEXdvNABZ
b+Y1pmf72CCFvOUhxDh5FN0OVLJk1Z7rvZf7drJLG+3YlXCkXSJxv4m8rJklf1zbwacMXK95BdE0
rFruFfv/+bfM/FJqEmqdgXfotOPseHQvMm4QnhwWUi0t8QnyHpflKyNJHLIgp3Pi9onkP2Mgd70F
GvMXuFFe9cY6SrWx9G2UcySfuWSyfar8WZs1vqC18RITzmhbTKce+i0/ezmFbmzc9LQsfo5EQ0EG
oKDtQlMzePk9DPA0OIKXY+12kbQ18lHOZb/iOhpE+GgDRJcXXZUSvMf5oalztREtI+53GyvmU0nF
fKp79BXQRucW9dso2z5PobEPHI+MiOhzEPefcDuQw4dhHVLCFIQiXpqPro1sWw7IiH4ojpIwiurY
ZvYMHm0VQQrJXvCNPItVTtQXph7v5+kmIMWmnlO8GXBlCmJy8U81qG8d8vKA7FNpN5gfM8sE0vns
W0ES6nfHYvvITUNDVBTdIPhQfU4PymId6DW005sCwdWO11ksF+udW2AhklrFCo48MNgl+CdEjd4e
SySu9ElnCfHMaGDqF7db5PGg9mUAEE2gXX9pX9+fDlx4sOBuZz9N23kdLgaRk9NnWkRhiVZwGWGz
DdFIIUhsePEBwlXp+nCnJgpR9sSd3QUqeQ/52vfNUzvGjMAC5TH0BFBrpFDNu7Jh27u5kPVIQFRX
PT5PED+M+WmK2mDY54f6bnNjX0UabVoInwJJt+Fp/h8hIG2d3goYdRkof7ZekY7uDP/ZW8n0nddE
zV+kw8gTKPdJ5O0KofaOvHwSVUpc0DNgqiG2fRmZ2BrzDbLYHpHh50C9OEnMK9+j11KbfMoBAiuI
xBRcVSuki12gUbl2xdwnsC2AcLwi5oVV/wdl8MAiVt8NzfJM9UYCfa0w4y5enWFZKhNjIch0PEme
cbZw+OBnfm6nut0+2WtzluFPZU6Um+WmT8oDgkeW4jrq7JPrhwb8+Mf9AzZIpUo3RdSvc2Hly3Ow
075lPNcol2x5l7bNflk/uvjvn8DeS3xNAZEnlhLpHvoIqwNbhFX3uUn0tys1zp8p2wamXnRPowXU
5LJmB4S4clW5SZdQsLDMjeBhwB1o1U7lA2vgA+9BfI/zD0BJLDhwupq/l/Bw5LQ4pads5x8e54aW
HlyYBf6ToYGkyNypved0oQD2tReVbDf3hC/zPozMnfWndhdVIMzxGNkvqxOGbz3iQAv3oyUUsIiX
04NhepaJKbizgu/qOod/XdaF7ZRQWNFTZ3nXvsMWPQV0d8rHak2iv3olNfW2+5UbGdtKAAypjydd
d5th6iobq/6oWvxtOkTQk5OVv2jQLTq5BFKC/T5HIIfyxn6e/7/7CYehCG33uts4vEVmq1Oep1SH
dfsiHUULQT3P+/CHb5ePMxOMumdYKUeu0Rsz2eQHd/TKGQ1GHiawnvSQSzLxdNOwYRGkZRjViHK9
7A8+9tuC0A+YO0eNt4hlD7+MWDx5YtpxmAdXC0koDemvCL1sYoSnEBgUozHGnvl3qMJeYOEcj3Y6
pddS2ChW6KcmtioxegkCrORWQAfVJt3HklbGO/M/HRIeTlQ28CEQyGHbZF2S7x+yfWAEPgQSkThR
AWAuMhr68wldSxtEeJJiHibrciCHCrhehlJhm0YpDoMPSPp40VNrv92EQ8fS6xdBUiXA11O9vWg2
iRrrXotY7sN2Nxb0Yo1UDko2V2aHhi5tmixsZSB/K2GBoDZLmxrLHT6m7lV0RPqVAE+/OS3TJ5jP
actJd92c21LtV/m1qoKdsC8YPTFdelPIjLqrn7zGY87ErRE9RvO1Elrl+W21oYVTd+PfcBvw9WEj
AfppNGsUIiRVR2CzRGa3QCLx26M9pMMJlrqttWN67Y2Ro0vImeuBpqCbvI/jjfJSQnukLzAuacjM
uWAKN4cZWkygD4AA7ZFbB+RMCxuT1hG254rdiBsS0+T25XSmC6KLVr9ox1J84q/V9tkHQsxPkaLn
hkbtQaJcMbodvj3p7JBN4NGIWnbGipf8L4QR211LxMqyBULIvEtrmSXSTuxiQm34Y4oMHP7sCDdH
v7FM+qLri3iupY5RlpyJ8UcOJfx9R/onv2H0TsZXvG/JRt6cVkV8dUHNZwKgCT3VnLNP+fqaOSrP
fWKz5ayu+FDHBTVDvXpVS1DivqRret8mEb8FtGm1s1/NYAmcdI5EAUpo2EsZTKnXTnhXq9T8YkCp
ShtJ7K0CuwQL4Q9HaGKEJm+0dNhZJna/6ib+JO6W2ExBgrtXLZWVbZ/dXbotZNsrk6wX/azVfos+
em1Wk9xLU9m9DB11W27kDB+jLu8CbojzsPDxAnb4qFPv2Bmr58aJeXu2y9ydA1pFoIY9AAmorx/8
jIS1qpf6h/BXTu+y6fOAtgGRpm+/FOkr4up5fhgVCE2M1LS4GXj03Fd5/2m+Qmn38TAcQ1WLKv5+
CK1Rps2MGfAwtm8qAc6bDuJOWePB54GWdRSMeKVh5TejARWYFvKoQUpx50/JPJMIJ9X8GsdNNknx
NNfqsFXGeSVmFhrWkb9SHM9sU5esOALdo9gu95z65dskQp5T2K4aKrdQcDYHATUE+9wvH6CUM3Sd
KDu9yKNxosPxFbeGHpK/Q38ON8LSfW3hpiN0yp1m2w4iUQNCfpb5Dl9Wbolh363nMDv4CQ0jD5KI
b8fftpdoWkKQKPVodLhgmD7w0dqv5msgoTMGotpyLu1PTEd6U+U5dr4L//XHIkvOeu1ZyrXMXMSb
HS6Owo2T1cZ2mdedJcO2RLeYw0Lgvry84d7FyUFfKLVPg5zpP8oj/Ss26qZeWf2wg3kpMMnIpBbj
4QfrOG4w71ZEKb5oXj9Z9AzJnnpxQqWhfJGciyN7HK++NSNKcpjKI2RmoQ2VKDhevTMB/mNMEf0p
/3WnjTZY+1biFWXfzA/fATUx/UKeetya766xoBb/vOFT59jkjBfcG9zeJJsS1AJbMqWMxxh0o4Qf
kUpI3gX6LZbwaMRvprtJ2uD0jJBid0mb0bi8ss7Cj3NxpOWUchWEAZZAk2ZYfA49qxUCqDOdF+du
xpV/op0NG+VIMIz9pYSDbfpGTdpbbtnutH4f4tjsMPuaz1GtomHM0vcjSPA6NxA55t/IYDOrtLHV
/OcUNzSLprTiTa4Y9wth0cOAHN5aBjRBgLFsp8HvQP6VuL8iNvXmi/+Wk9+SNsfN5MYE1/Ac7/nC
MRMGEbRCmvnu7tArG8kaAAoOX1ILaD21zmxr73qS6bb52ud8CCn3+TQOClYEbmNooJN0xRbwRU7e
oU4PjUtrekk3WI0QS9aq+Mv2cprFgZT7zU3eMDI2bNWCncwDLupd7F/iMsMaGtz5y99EZMz2BvHQ
cUUquLCgEFfvz2SYmfaXTkSXFsAWjLOGsdVSuRgEwm+GP5ImV/cmQqK6Jn1UL1dxXB9IHvQAUmLc
QX5+/k3HYoUZwNNTANSTa5qaKoL0M/rLuoHzU4WxodXbsNBoyDQU3MaGxjsg5Y544fO7Bdd8ZxS7
MOjtDh1LF2fervSLBDxRNSxG4k/z54aezpLYa4ugr1EWCLCRvBAXRmu0vg07sGpA4pWyxnILRB+B
axtXzkD0SKNktMSs8uEDkOCrH7JF9C9v4/ZWq4lJb8vrw/oTOveOHwwhoKg0fjlhkt6AkjOOv4rX
0JgsBIovu4bjlBeV3E4cY49CMz5VSerjE9TYU41rr0AF6q2wgZg3ek4nKMK125NVkVuBmqXpnAUH
jigJxEBiTK+i+1Mc7OrjPEyFBP2A1RyCgI610whaso9b3wbP/nXlWVqmlNGTVe7bmdLtdg19BG7T
iAZmkpKmQzNVlUA2/9ftHEFR3yh1wztzJ0dIQL9XoqmwD8YY/hFJqZw0lvxnFT15QRVBt77yJ8zz
2L+vaZlC3fLTmjaHTlsVENjqB5PYJELWjEzzYtyzNmZWqeoWtuvWKr5hNKJZE10hLQFRiuKGrrV8
PrWjClvRdunvDsuSavVaCcZBGbpyqmFy29jDHBcTvVE/PL1PCwQ6i2/8Pc45FvJYP4lyYV/9Y5nj
LGf9y9LCt4D4qLBj3b+N1eH9KcJaCXtzs2G8u7FJBs9TPvHaIGaoakjHpn1TELDxIJVbzI0L6NUA
zepvpLpwuaAftkqgUZZJ1goEF0zbOw5l04RrDxD3dQJu2tUJUkOO9f1WuY9b305g4MsOJ1NY2Xmi
DHGEX46PQ/nzLSz7CjZ55hcFLikaJJct7QKSMM46GHO7fztINOHnlQ56egX/FDr5TXkOj4JVJ2Gf
E2p+FbbFoaUP8xDwgeKwx7r72JxQ+PYAhUD1K3F6qKdrxqS2+CHlppIKBfNCTcb8avNHS/hj5w8Z
Ax86n/gMaNNH5OGItZDGh4+QSveo5V2RtZ5mLn9O+PBkhWIND4GqAqc5fX4OWu87PqCRROIN7S85
68s7Lz679gI7z40boWWoSiOLQ/SCKVfyUpGibpk9kx1UMNeUluokRYiV0xCfrCB7URa7X7DXOAD/
8rJBjNaWQMFBNCnZGWIBzx5K20WIjtCLFvgSHPYet2UaDeZLs/MqZ8M9N6boBoOmOviOJ8J7GGyZ
3knTvap2w/vBJsrwt8NRRzSRk2zjYUVQ9UtCRN6lXH0tnHwcdrqgjRShQJMs2860tkOZ3bRFZPaq
9GqH1olKUdslfvu6tMxjgpI5c8p8W+/uPe0gIG6+1vRd9V8Di2nlwohRsoJ5p2ALLdhPboe6FddF
UEIY7vHSTzWjI3SAkWGe946QKvd+nUSISgcpbzREMXsinlbruhZ8yJ3C5U8oXkzFpV7sHIw0yF7i
IoBce7TBwSUaTUBE6ywalWASPhwvARaeo3x4tX4SGH5BERCMWRWMLCu6RYaGXzj+DDaJZJAlNFO6
gvhadC7SZVDUYejF99os7FTGXI01SMCa3OAqnV0VfaCR8uiKwzXVF1eS7ufgdMbV1DU5pMjq6YsD
ZjmBgrspeYEc48VX9HHmAWvni/a2mMRtOc6qBlf8k6cff+JG0HPpAmdzZwro85XLEt0lWgD7xA/4
MYXZagzwLdDu/nsG1opZWZyYrLssaLbVf2qHF1EgTCZM87gGZrqw8YveVjWFmCqG+E3PN2ucSY7P
/PfNWjLSv0Jimmk49Wz+6OtJh6VgRETWBzcEKeikT8K1f+EPUrXVMYoU3R4aKfDEMriZeZwtchGI
kDFHb4/tSKdyeTpNWRUfonPksbaRxhgSmwhz8ODyHwBNqnEtLkJ9eyUJ32JgxSjac3vCgQ/A0yzB
4A58NpuZuEvJGuiQ7eN1ONZrAulrS3gMsIoEYSvojRFR0VPxEi6XBuICUOIBLKWXvGqf49yFCTY7
GERuJ37o7luPIO3/JQTbwcbg0I1kJjRggfGDqm5jAs1rDgNNigMZvBHQftRmgPf+9xZGXU2uilPk
/o2Qui1YFYr6m2WfHQhfXt5U9rHwv2hgXyJC5PPvUq19zmOuket6f5IyVSDN8qTW/irVcHPUV0RI
wZ2uF4QQkgnAqzsmcGVoC2n5YqowQYrtr/HNyx5vwgHd4duNdAOeUWFt3BX7wgTVFpz8x3pWRdJc
eIxCiSbwMClpzx740XO4xH4x/H9lnSJ5p8DJE5TNKeFMCgizd3lG1FqYX4xSXELV84P1vXuwlcXP
tKXRQvntx+gf/gQmTGAL2rQ/piip/+oW5brC5pkaje7hJtemIGyXGn+aTq1+we5mlHzCw+edc6vi
XejcC7ItocawChAOFFk+SGYl5z9cjbA7pYJqQboNMj7LVFvGbf9cN7FKG/M4XoYm2n4rvnUWxSBK
0z7QLIL1NPjJiWj5n6fGZA09BSKOBEjgKs99jiHgUNyKMiPph/25bZhjYhj/wBYJYeRUUJM32iJ6
dCr0D6IRa81mkimVUJJSNf5Gbux96xqym6X3DtXI3hLyRyCA0fgRkLCsDfzPXqc2aIHw96qRGX5i
Ak6nQsI5zcKKn+Pl5M4rCwuA1qEcoeBp98nFpL1yGsAo48Sro+SxXaBStADuk2YHyL7rWuUPYW9Y
cOhvhfIEGiKYPQOJ7YhDnuBRPghjjpMYXkPEzCvyV6NG8JoDuW1+2jXuRIB4Y4+k3aASIw5YgwRu
mOmwE2jrASb8BZrSiXZuYtnzuzrMxnyzwDraY9LWGpfMOOck5lx7NNQM20LekiLmf5uyY/+1yINY
4Rsa6etWIyQVNMs+be/YpkNoguzBKir6xuSAczHpf/NqfDzSc7ccwozIIMieUCqGXurZjEh+3uPe
CZQkxFwwGYi8i4KDvllrmP0mk8bOgxyUbXF0pZUJiV/844sdx9fiQfFCQYkgGZa4j2iLfwBcwzlo
zT35i6UbSiQ9Q9MFeZ8rRl8vl5SwB3oLSU5xQOty6nWoqaKwDG0DCdADUP0ivp6FA4PtIl6IdKdF
W6bAXuuHUzSX0XVRRLqLcOkSOkdMYVT+ncC9KgDzHlwjgl6zGRQh6shFk3rccUOPRoSdVx3jXue2
ERWUBRc3zx3VojYXndF8LqZcgyhSiEgFi5XBZDl5Tre11KooOlqknnntjH1mj010yx2/p09hTsTa
TxX+5DcgomBYjlz+ZirzR+tiXKq0WL9BPkQBPHSwvzqAc4TZpPkeuMiFu8Hkfc10JQTU0ti7mGAx
8GsxGxlv40QaGhqSeMVy7EwB8bsbPmBxSVLUDZgS4gl3jx35W/H6fPBNb5WvBxDw0auQkUL2e2Ka
Qamvu3yLj0eupMB2zYQxeINgxOfc2Y6PZD4p6rYAItC0s3K+Qb2Gu3YESHsbXPw+JHkn0F86/fE3
XZAbxzzOrRt/1VC8phUcRqVhIaGun1IiZotMPXViJcdpmLCWPqTjQeIFS+aD5NNUXaFSlCqFmorr
mvZs38jwMbtUg5QlmtWwjyNHcM27WDe8c8k03MYJWMIo9fG7TC8XP74n3tIVsnoeHTN+WO3VEn7d
IZDQIlvLYW6qgLrEkrk6VUQE58mpQTxtOIEXQ+0q/vfICYI2vpWxxeJ3W5QlgF8FPui949cKV/yr
6DbiXAi+jDnK5tGWH0TLLeBF4pd0WLh2C0RpGqOu2aJcI83K2E7ujaLP4DSo7F0UphOwg0wzo1+V
fbIF62PMG1/RA5xgrPGgnlbo5l0JT0cVb+HjmtJ6RSWyEDxFOpX8IK4c3U64k1ibnGyMr3h6XM2L
EyDQvgtp/aYTARm8SiN6TvnUyWFHEVtLAR+/LrUjDETHNoj93ML8LR80i4c0IaedEser4KpeQOCj
GaW3Fho7uIT3K4DF8EE1j/EX28R60KXf4S4ZvjiaYHOQSr+r0iO8r9etmGEUhXByUG/HCrn4v9Dy
QeT5gMuue1dg/MfG+k+BINDE5i6ZoLUOMmXU+MjPx9EpRKiZmiQ0pBcYt5Hy0Py0V0SqXKRYC2fB
fAVaDIOq7fj67iYLa//5GoRvhpXhsQHTL+DtIHIFTtF0I8ZZswZQ/mm/ZD4Gppz1nXhYVaQJqhTU
L4221g/XNlsXsSf8yYvRwooAzYgwkYfuOKI5fyBoDH5h88++ciUOoIEKI/0tXIRe6frjrxTLg+tm
ZJtjijBZZviuh1/W3wDiCXemVjOPsaSF6WeVfNPwfwZ1WGvgWTAe5ghtg9AGQGmhY3VMnFlhfb/w
/CeSRBwAtnmh00BiIp91ssPrX/gfkHvK5JvbPIZJE5OyKWpxRCPbBslS4HyK2WbH8zwWiOcNccAt
SxA+eAtsi6Kac14hAFNo7UBrhlS+go4qZmAlugJ8ifCGUGa8EZqVQNPjoIfydkemE5G2xWHqU2+C
f7VmZJT1VarKJMBv5jYsEQTDViQOvvYaKbD8SFZ41IATtIh4HdORnZiQdykTa3jIe2487WIcjuKO
ETjtqruERmhYnRjZOWQpHB+cQfJbBZwaFNDgYjOVSZpuVZs8sWW4c9J4rAIw2HdBbLCYIXykPome
jZG3TTQBcKLgGOUiaVM/jT/cxqgDSD7IyHhTdWuujrZLRibeCGNsCcXbiVajubRYryCXl7u08KdP
f/5Ox1wkuwJ8JipxeWwkV7tw/0S5s5yV9ZkF0piaF6X7sfjqGdzgYjmIkxkoFKlI9FDjTEJurJRA
rdod/N1Mz7HzkzBepF+B4s+lkbSw3jsZUGht65EuiKG1evvsRj/tWZR/zGwoucvRrEdJfzbc/X1r
cZFNcZ/EtJmSub51IXGqBMqFybRLANpCjsShC86WxrvIoQ7tE5POPF4ukB57EDLegtcmDiayS28h
eBHLQQQz320WlQ7chsn6wy93Nxqv/3wy58hwOWIISptXdrpFmVZ6XNQVf16mHwpYPWfmdnCyow+l
tpTHDn/h3OvRcFaWnX8+DIOx4A1qb0rbR5FLJwTC2haqEUU2Ik4CixiWS5NlI7rNfdfzy31BaEWf
w3J2jzy3LTenbxwLs0LwWXG4MFSh+wOg5NZm/uKv3SpTgevB+ENr6C8n8HDw3e4iA45G8+llEYS4
+ttiUPP2OrWlFbbtRgM+PllDk/PLhdhYYDzpsThE5qcP2pUJdfhoGqW/y+ul1XeahCajQhf4ITjC
zWIB9VhLtLLUUSjLR6zDvK6b7RNk/8KqYRWlsjgnrB1Qqo6T0vJsdWio/KHqBBxIjjdrfkeAvJ+u
78zEqos7vGQcwSNUN61VxCwFTOKj8giH66OQZlqatcLalISPNnj+ltqqW6fMqaVqeLkHou/zyQ7Y
TavHursTHY8Qn8tYJ2yBKF8qUKSI/cX8/Ee/r9c6mNJlB9LdM34RF5XxJB09mPpq21PfSChrABDR
DtFKKaXUHa7f0gPMemaz49I2Jhq/6TI2gK4FAwqhJ/MhnfOmb/GmA6nEl2WA9BPl6XGwpDPY0kNf
dmxot70LOZMEdsWz4YR2r4MXsp7w2a0dUdkVkL70wzLV9dH4VSrKb38VP3n3b/HonBsbBeuFjUng
+DnDubis9XGCGIg0ercpKhpAKC3L3whsH+aCnxSlVN6/Qg9/osnWIYaXk/sKuITlGbn+YUrq2uyO
9vLa+1F/zK7yGAeWnVZkDTXiU7OUE3XCYcRRuinwzjvzvbmPm8Yvatcuqx6FDE0UGpL+OSbz4/vS
48L9uq978CtLcp0sZwlrGeKg4hYejf6VQubOdA6QQME6/fu8R7Z4JOrcJSmcSXGaZv3ubLk2iHyy
kjZd4/+UC5dzHhMXb9WFFe2I3+U6t5kCZPqd4H0k7xlV4YPyBh2VuV2qDm0yc1PjBJt0VpTD7ZZJ
/mEuDgwq02z+X0CJ4RdLxzY3qSWVWjSO3GHWtbZ7NrsW26hUcnWM+F/Vo8neHt3vY9AYeLMUYk2f
UiYYrgYPcQXU3We4VkXxtXrR8HuuTTrgAAGhzsP64rV9AQF09hASNS8CjuKVhxlGJEcAKvlNoARy
Og+eSFDrFfjBn7B9ISKaqNBG19JPJuGW2p70H5Bg7D95SmifKNzU/IJGrHQumFByeMbb6QVuCaBl
ujPZ14mFpaYKarulOXtzz+7g9J5UE7EvdH43ZkFp+wXAZpu5RYzfLM0soKGomiULXOkcw0YhtF12
Zh8Ej0ci2WlFmidc4DHgtUtjwqzWCDXu/t+iE9e3dAYJ1RFwmz24uLrATiSA05E0vJoI8LxOIYek
Ea+aEa4VHoc7dgttao5622JxySjaheEY2Ag2LbV/hPgDj/1e20wSP3eWO16UIPVF57OG57WSziQh
uvsaSG743itR0MLdEnE/1d+mLKoh04PJFvUaW+CmcZ+fweDH4ifrWLMYwyKTeMChMfa+4GSaXT6q
rRQ3xwq/xfYXdyicnSkD4oR2lBVkc4XrXFshWB5iXKgSOZWKzhoPJi7yvo6x4N8PnXM4qPWsJ8dP
KBEvX/mvOOhEMNC+ZaZstrKV+IgUUI84vvBkfeXRdfrZ4HnCUvgfS4QqGIQ6vpy4VwrCgYyfu1hi
w1T7F3AJ4x8b9N07DHA2UY3noZs5VoRiELpHmDu6u30MlEQHhPplZmwo9QikjCD7GkPlS91cULXn
NSVKdOWPU/0cR9XQ54FAL7EJX/4SpwHPq9Xuko2w0s39KWmObuJatpHDdr/Q0SXez0aOup7A297N
C+4vpmdYtJRaVTZJuEbWR5KqBFOL+z6jFOmi7+mYL4KyjqT1adlA0a4BinGeiXMEu6N9X09INXhw
+2+JjOiCwGbfPDkdLtIOX3chEY9irL75CbZs1d5MiKCimKq+UDYI+iK6wxEr/tST1hgsir9d/9cS
mTnJTAMdAQQA5XvOTgCqDqh8bu0CzCtQgVtKPVIOJDAbfAgw1t1V68rzA1n1aSCi2HxUuPyY9HEv
81w+HPPVaszdNqluhMXPSGS8drtScE7n2H1QDWsEyLxQoa1FZi7bD1muX0pFKymG1ueQfA/7hX/v
61jPHqEUbeaELSrUhhFEN3tXct1MXZIhPdVjHMk7zSr05JcFfGUHamEYsHvMDYBSSFPiYmQden14
EMMONSPuSF2hgVPTTooEs/LdMH2XGUO3Zx92qngOkTcLIdeYt2duUiOr0N3tkYK1mVe3ZfEJ6Qtz
FEhJQ/glDCCRmv6MFPW8JNPmAwBUM++fRTudqdxddbttbzDWhxJ8w3dQePaNKzM1cLLO+1LXnQYU
n+kpU1wiyF6FdSY6psFkIgYkcAA0HtPfW2qx0cFxHRJkTdm0vbgAOLnFtwBaOf0hcDIdnRnoxknE
03IeXISTklh7cNrsc8f8eOxU+0RDCECHcv6/BK4+MKUcWJSwPXA32j/0GvUrvBDPRbbmO/xAmxtw
S2gJ+pW+SeaNycrA3QZnIX72xZE1SptBf5UDdUjT7DuoB1Hd7tYgCgkRYKkd5r3smRZy0YGNvNAl
g5aZNNYGpLovVwEYkUk6crClhgreAMj9ye3pcg4WkUF6bXzEfhpCU8xMvdfXZjPs84A9QllAMeaZ
i4syVGE3QW1u+wLt5yBNR4cynMpSXiAAW6DqJppwLJKrOM2foCP/j7IQneqFM7MDS6b5ODQZo3dz
nXV+41aK0twns0f7iEFWHg0drtbxxuYnb1lsmqhRTKHkLpWcxcGCHscDb1idNGXhN9EKB19y9ktb
Mir3JXqghXNzFNMjWphC9UqEIXuX4Ly8rwXAOudN15q3iW1cnyQkWX+ouMuZwC5flBC+3EEck503
RQU8+dEhdInrJiUE4gWy9peU7JXJTz0QLF215boJl6q6UDAmq0M8m42OACCTHWPvoPEjOQlsBXMB
ZHH+i2ojlMrEQ1xWJhOFijQOkF9zjv2Sk6Ppnn3PEofWXaAkY/T7wzQFFLdY4MB/sIO5CRBOm3fu
Oa8S7QUmoiQ/YD7VCtLq8c7dKUcuma80Xrf5HA8o0IWJb9LtbCKDODU6cx5y1sHORL+WW06QMXFO
7+FJo5FiC854f9ugiRdEW0YpU9wzDzsyQPxuLgnXM3HLMTGyy3x/6P5mr2iaoGeWSNoTwDa0RDew
6Gp7OEEcriTkW1K4UgYmkDx3zd5lSFLOSdSdBj1KyPOWaHusG8nUqz3FsD/i/2nneVmaJbLzJuLF
BG3R3sOS7/jotBAg/jo/n7Y/Ux9+0lUlrCOp2xryMLaPpTk21pVSk+9yaK3ZyNcPngdtgPP29bMe
7evGmSso3wS6k5XCslMAb0SphconUCUaKIvDeAZzUEbywD9rVL4hnBubvcmylP9yRQAwvaIP0MDj
rYlkz8HllttwOHLqql/HM7g/ufOAy32PIYHVvohcA407LGh7gKdlAJau8HWoutHsy8MuMToFIJBs
RDiR4CwvpvS0AHkE0C4a35sE5X8oCMvyag7rsWSXn4zY6QOgXJVsVzIeqirvjxInJ/b6pSXnlItx
2OyXzS784dGrQHb4oETWlcw3iITp5XzIqgYINRrNz8YFS3Zme9pTEqYxf3Vme4iiODETW/A+N/Bd
IdwH7JGvUePkhs5XwthjhTUfKnjAqwl5/VNIU5kRU8kyScz5xUjxI23gpVQnQTCkSOc4yJc/dYzr
Dy5eRRRNXUhzJkTZm+eHBfOpdW1nGI2dkJEGCw4Rp4AtC9UXi8Qb0QF6SOCVmgtb6WnuM7eOjVmg
udS01b+vvtJtRhS5rNpBeTXBZNBIe3UX34HG9vtxZ6afRIXy2zRbilmP2p8oRfwZPiwbYBZf9kcm
Fw3mQ4XKvSY8dhRVBdCoYa+/ocomUAOMdoNmXmHd+Tz2klyNoH0dc78rpXTY/e1tEyKqq18/n0za
PeS/Hgz+lzdaxIVgfOpDU4K/nL3gSgZA1a7mKT2b1lrxbOC1ialhp+Q+u0zKGxRoa6tUvqMYLmjn
92IFGpJX6v0VlFu8GgxkJjsfhB+7pSb+Eawf+Qw+ghGFPtJ0KxWM8VWpwipX1dB3aRSCBs5mmzTy
pAVj9kDDlexi49X+ry2d5yhfeQlLbmVrTstipHcDiQeNyuuD04O9eU6KI1V7Y3Wq/G7FOMD92501
vmV/vKqXtC68fUuFkQmJZVK5sTeTTj2aQha4hamvmekdSDNTHfiI/BAZr/39+Tql+18FYVYikHrv
R/SlBYUJyw9PeL9FE/w+I8bTOtic51rQCGWhkuVQKRdi+GKBCu2YdYGqcNvG8AhB3jzgFIMvFJ7q
p00a5f9iRXdKDyjQwous25UwA4urAWOvxz0ptLAkSOVgUh0/QN7t7BZihZWC8Y0yoNcjuJSCVJxv
kWtrqA4KWuZlbR6Narrh6KmrOXM4o01DIYr7S28/dynG5lks0Q8tRz9c+AvLU+33mcvtcOkAIZFL
aFrQoEbTau1ZRc8NMAQfAFywXSEwv9Vf91+E6N0Vt2du+ncO02VIvFbA7sFBOmbh4LqwAyrnHf+y
LDNvaqMVqO94ozgKWYojmzmndqCfyZj2lmPgvzkzc8KfnnzJ34dFXxwCdqQJuFzMyPvN0wwjm5r6
kJF52fl37Cn3ZMV4KclzH0b2tvjCldNmwPtV6Lwt5knJSsbGuoGBBjV4nUgzPT29BnGRy5/U34nc
3TOTIDNHoQIfGd0d/J2vJNNkP5S6bFwK0WZJosWp2/E0r2WOgUMuU1QAFjhD6LnlFWgwcfZP9oqe
VpHuVJOpNNlymQtsud7LdiR4wmDPKz/N1+JfuTRxruaYzll9STwuEoNNwC0l0FoxAsPlmhsY0nd4
+tZxYcCXoygmaQQo0dYBBl5SkfnfUjfsbBYebfhNCSSMsbrqpyXLBFOl/EzLeZpweUcHHhHeyIPA
jN8IYmhbpc/avGX6kBFErGgxGBDX1tppzx+g6Qd2VmPKNp/Nuylp/ShFdCqSu6Y72fk/MHcA5eFM
HsLQzZY3qYkv9bRsP8CS2fQxseAC8XfiNlvaS7IVHrPSTX2u0Wl7vA7O6Ukrwvm8K30AmWbL1/t4
X4ag+tZdh3NOUjWCHGVwl3OjSx3ZbHZzOXYfTT5rzmmLPUe3MPPOPMHoECSnOrDZfUgETB/aStK4
NkoERwZDyYgFdSE5rKEwzjDJ+/t0bfIyZJS4M9uQUXYghgOBT1vM+aoqAcvGf7KXZN55B2d5gNVN
h//+1Y0A30+wzU8u4yNEYTw0W8Yw3nY4ycIVnwkSwlL15KcoqpyMBaJS8e+mXSJ1Q4ecKFhG73WO
SMrqDuOeRbWVD8nmkpRgmjmPiCWw928mfLBmx89aWuSia+hM4mk3gvJCyfX4iZVwdKk2ZhHtNF6k
Q/nJ/cV3ainaSkzsM3jcCq9BiFEXLUN0a1G1rdY7Xa0H9TO/IZHAyBiKysO7InHh1XnpwBDT76WK
zjsXYZoClbjRhCzV2Qkcx6A2poEt8D51nGZ8M62mTwzin9ZJCVk2TPLa0CEpQxnAwandRuvj7sxt
ISKvqWktH6d8jc5jmoRGzwGERwuo3XBSX1g8KLJ+2IlZ/MrxaRTRTfjPHp9AvuODX3HMaNi9Pd2D
Ql2gghM0kfR/91GX9y9bJbq1/kQk2Ae1H/J5nWamt36LrSu/vkYLEEjUoQ7oGRKdpiSD9GqafBfr
UiiyE3PmXsON7d2pOnW50wtMwbIjsllC1BE5/Af2WkA3wCJoCkAfPK7nbzLX5H7D3EqRm/8itssc
0VIWIfAbV2g1ViPG/foAJ1vQAGGooOTdib6IOcRYL99d/lXSp3qxqtVkHTY8QUXSx2cdJwBpXUgX
lD5OiMi2xMVa8ucrXDpAw6VhZPl+Tv6CERJ8oPjiON7jUwbA6qyLC0jwGX/X/d6Nwao7XXAPhLVw
+a2J6VQ7gWKZUiyEbjoaPbqoYY99DT8FlgyloLOu0D9fB4Pr5WiBPLQ7fGGEwy6XvI3Ydt8tHQ2q
sLDj7f7kX4mjdah9nyABVpcYywqvsZCm9gxYd/M/5hnWtcT0xHPjOQlnUy2mxv5v+25i4+o3tBqM
OvEdoyADdz2FBsdl1uLLE0xVaYY8KKmzNw0VSRT4zqfIq80t/x/Tqop5MlY2ynKaRuCQo663wdSe
qTWyhRcK0A+RhR+1PhH7opcl4lQUrAJQs25dbeDQAOw4bg8ygVFqBLbCxJgLM3Fqa0tAvXMT9QKt
8jkUvQ7SOxCUDF9ywm3YFMIVa/gDO9ASk/N0o1GZINFoHcLolgq/X7MfZgDPCLm9J6DtZKwr3DwZ
OixQUvYUY0Qa8LrPwiQuVoxuQFDN5ITNqkwpUXIkexGsb5ngm45Da81OYk6sulA0tZ0oFiPSwBAE
G4TDhNO3SzG+qpeSqg5Ljot0T64i83kaA1WW+NTxvhqxUymRdo0jxfkYZkkGHbpJbisbEuNJFGbH
/RG0glWCiIquTAqI5Xf7pT5CsyWSU+ffaKRzPjKVd4vckYBbbNYmwKk4WkJUhrvof1gYhj3VebEj
i1q4EL/6gbFqzAlu49ovXqffktQlE23lDqooyw69wvJm84U6WDgceHt/CvXku/NvCw4AZfw2C/wH
X3Z5FxkZVoS6OOh7CN3edFV4LJqBksIB5mHRh4JN/3fUkOeYIi9vEawALYrttIiJJsEweM8nco6x
SkeToX4et43181mHG+gC/TkdU6d1lUxZvhnjNcyHwS0B/O7g4IrT0AUXiJOBECktHUTvhFfqBmMy
nYIMO1Ot14Mx6M+WGzwLHi3Qfx8BdpZ5xokjyRWyxp4tZ1Jt7MLsBsWhps/D/TQeWoSET8TC7/S/
M8clXd3dmC+4nRxMzkfxb1lMnWFlvycGwQSRO4BONOghI2IVzWJ/IV+N9CDyGPJolmMN9P6V1L3n
dcaE0Ebtqp/WS9Wtsi+Eq9Qz8rWbcnjxDHh6xQYWCsXHDUIR0F7PIglLtBs11lteu4XccqMpYrsQ
Fr/5A8Saacwl7jm6kOyisEdqm8Z9KDGC6CKTkRZqTJmAm586BtxCq3sbdjTfiOgVSuT7TcxIauE0
hItmB/vSdERC69QL+sSmLCpfW8WiIHrZT6YxvVZLTYdxKYDtMXUp5ocFUmhfMs9ydgUsX7w1qzDM
QIPIRCeE0V5B7WMeY6lrIoZhIsc1xJgzXTWVFsZyf5JKpmInZoFZj3/Rg0bGy110r7PspIGvNUnl
r70SIAZOv6AUj6pfsbiOkE59k4RMJ02TCuo9RQkJNImskkzob98tj1IknkoVaW8uA8lzr+aSIrhY
iXG/RhQ6LwVMMvZQWBwL8xJpv89YaxgS47dOUPFdxrOUAD5lhrXo2HH/OZ5dQhVOfeSXupBChuSq
Hqb7eLcvps5UjUwM+u0VYgk7viz4/yMeTJivDN7YGJVsD60q90PojbSTdYtSclyUxSzBtQgtAxb8
gd31mrGmfkwJ70vptUflIt476Ke8cy0v9hnYM8mdAicOalIzPU5tT2ib+MZ0Pw20qXeYcr9ryPvq
d7afo3ptW5tHFahlk+MaAlUuZrWdvZYR50OOh4rZfT3VttocE1CGHJoU8PqUT18Es+2NAK8l6XS5
iRrnGTHO3k5IN2m1exKG2lXFX6CiSmTfxFsOndw7mHHLSIOBtbpgwZLgsUFbpTg/JUbmZXg/0hvj
DUn6j0ob98erG7rS8KGpw985FDSzLT5QZY3q2JmDKPVs1ZGlCtBxM1YzIA1y66BU1CPvYVGXcXJr
hJOfgxSV0t+io6v64Rl+aML47cadSNGxaGOVqJAP73UoSW5R0kBzmk9QHeYN2JoyTFtEexG7OvoX
x7EAMBv4rSgZ48u6y1Ca/KATGxbudi8ppaYhAaA1uBesSB0c3dRQXTqGKUrYD+Dyip1FI7Lg/FhU
UlxIq1Csa9v4YFZ/SWskYeLUr8/l6uWNpCDyFA2jDxNenJ6YRV2Qu0GKWEjcabfb58N719GYlplv
cBkhwih8nbKFc/BW8N1ZELlcavL7RaYSf4h3wa/aTQSN3aK/xWXian3EKZTntpPFRDj6C/vFy3Dt
uM9sVB487TZVlwFJvM6suXxh+bGfVBcESLoVPmhNLIVGriHegW1/nFA2dRbuD2G3Hc+mMS3RP8m+
A9AU64aeW3ZJ8NNWdYTyNotdqoJbZH/6MLTw4U7S8Y4QgF7vdceQEzmkt0cyf+0fLRNPBt6RUrZo
E6KeHnIwvXWYs3cp7MqOFLbDt4yBk8hx9ygx0Hs5O/KKmNXDXiCvhr/j8TjVwqTcjFzbqA3TbNAX
zh9hxCsUeQfhmujBKwl7wOuCaWzKgI8jr4JIdhRu2tDlqQzF3KNLfonXllof1pAqBp59t5ykph9Z
Ovh2ZAHlzDTe2vS1JIt5vAWunJLOuSnHFozHv1EiuJEUHnR9tBvstIKnwcn9dSLxnGvKhkubNiqw
7PiMgNq1tmtaqb82jIT+INzsG7mb93LLYAsT6aXH6NyxrPsxEt7lZm4Kidh5u6mWROU8tbEiwlOv
xOElKf6RbufWKFPGgnjn7FTOK2qf8OVI0xeT+03LHneglk5+sAnohqjdCSIdRIH7Ke7Y9i0vB4EH
lDs8phiDmO5tMlSNhqV7FLjWUSji9p7VeTJ/RDt4bse4py762yB6O8TB3QY4zjts9Swx3jBc3qbs
CQyZKKHDDiAMkv4Zr1TB0Ye887Vhbwr+NJMUWZFqYp9PFQaWQvdsQs/1JdV86BDQCMLeO9GZ2hB3
ka3AiptrDvjZW4XEaZhK2D+6fMdyG/ZE8pslcfmhId1EyFLTnbk6xW4E6ofw61y09GiPuEw11Ss3
Y5rMzOmcvBxeQb95k+MA2Cz5ZnqaxSVzPSLAmBEcNSU6zkV4tnVSJMadu/qqk05S4WSvuNqGq9tT
RTKg+SvRoUdRR4LATWOBEVDP93u9KsU3KJB4r83Fh/b7wICacF0otxPUH7SxoUoxlbbhxhioI1S7
rIlxAbXxRBx5iQlkhWZHL+8sgqd02C88Gj2ZdoO566avaWOdvbxyNk/AYMr4i6VGfSEAZXEm0U+s
3VeS5JOYr2xU3VWuL7JqogXZkFcoxXhlyhglZzgfO+v1CWCagjnh4yYU0q64NvYBvwCrOeN/gizO
we6EhnlciSvqdnmISgstxC2xsqZqRurU+kttDpc/7dqbo62RXwgtNc+CibU6wB3iLLPcTzs7nQXL
dbSnE6aDC3TDajtcEMt21gXP6K1U/ka+8p4jODBMaFlcU8bYR5QEOH7f0SS1nvvWgS15FLSMQhZY
r5Ygvpi2Xz9um+HvGuKluOXECYKplghJnZ+x+JkbkWY8ZfqXI218h3RvAcdB9EKvkBSCEYptK8ir
J55PAAVqOuN9Bk5ulMMMQnSUeOAsVymALbxzFpRIycTcyKheW7H1PcFilnpXDdi6H7XNEXYyu3qk
Ac5OZsESHElu/NPdqp2+UlJFy/raqHr4veX7dtPTyLkW62t1/cA+Yu5kKSU0umTkQkCF/TqM2En7
7BFUv5NoeDjchG+dn6jTqQtoSqBEdLvId1FOgdX6hBsrbLbOhG5zQ9m94dqbQ+jOexa18qr0gPhF
IKLaWLm7J1L/YFCKXUCkc190itRvHvMgsDYA2ZTWF34FG/8/QdkL3t4VIfdUKGkeSD+K2unyCqTf
QMC3Hr2shqPqyjNQkUJKdKkyI0eFiF6cKOj/TBIATusIAOc8jLYNySLSQsjU2cQEgmpIdLEA+79T
qy11QbX4lq+NmfDiuEGjnz87426r6+pxhHL/9A9czhZKBX0AQIkJIfJN0PIQI9zq4gzKfGknsJhF
XmZs8mWpuwvuQeUpT7WzVAqdV7E5z/xUGSkqCJrPaA8F5mgCSc3zY1Etas34J8jIL4YdF9Zvo5eI
kJrxaHZWdiW1zZlkxpBrBCQlQtlS+BIleZ0gpmBx0E6xExSlWPvBYCYXP0vgI+2FQYVA8E5Q/POy
XNMMkuisXEHnGcKh+QY8nYtrXyX1KBS3EuLv7vVtPHU0hgKZz4eqezwaf8HftutnT2JACvOeM1XS
dZ22UR2ebaNjjfU7UleuOeTIQdHZml+eieTIgOdBB1wPQYNSa1HZ1/qhykUkdOWj9vLFYTueUyna
bpPdJjtDPlD5iJtX1886NObih18D7mhc1rgBPEitmywXsi+JUFFQfFJULrWo4ZfEAxddVgc7GucT
ZHsfPWJXLjNNNvmSRH14hxWxhFpMipsL35ledkFEwJV6wsVaGhYp0H0MzK5zjoP7YkLG6EqoGvit
VmVB+uMFIhPT9n0ir08sroypzyK+lprRxCiZUujD0BINlX9+xc9/ZeGzNB27yIEEhefs7lbZVfsL
4MDpZy9BemDOkhOm9ojIpeaJ1eEG18kimrN32MPbu1etLJBbZLa4B2+Te3x41Ut7X26lo+mH4QhV
5d8zuNNYz6ml80HrXL4ohzfIv6wmKrBLsWu3+1CPVWPPCvWasxzkEZRwq3qs40VZLyoQ21X0ZEX6
F/doZxx1j6krZn6+sbZGHfKPblpAuiN51Dik+2tag8AbA9tBrhY3ayFw8fBY/1jcTxKAAvgQfg5j
0+JTngpfoNH7CP0rq/86cnFVj1DLQoYDAO+nKhiq+gue9Daxcj30yk5Hq7Yzt8FIrKMH7ua/GEVK
tyTI6WQ7mAhaShZxarTblgLcWMHKNcmA74Eyg6DOXHejQUn++Pkr8Mcs7gDxOc883p989KWd5USb
V45YTYtUw5ICU5i3XfPKQD9UqAVBz5Q8VmUQe8scPwZarYTLcAthn0N0r46Z3yXyq7QNIzf1qSLS
syPcZ22hWJyf2lpGDDhw5ayAlhwq/S8AVYsS9B4xDHdig4GlKlaEaZ70Ibxapkk3yGVgDeWpLiVF
z95EMPhiS+RgCf+868irhoJbmrZgcsUNkfyeJLI8pWizZR+O/i1V9fJ8c4WFrr3ta88Q+/kwoLrx
rNPYu/YJaMksIcZsYZXah0oNeXo8nYY5KErupk8rJDnSrZAp3F3DclvpEbp4o2Bkk0KJ5IQ9A9YL
OpgWjM+OkY17hEc65RdSR6Irs/PIaMsYkULKVJjrqvm5lyFJ9BUgUPQQpgUsaJE/ypN67D2sStuS
Y5/SiCe502BCO0zQdEBNGaQaB6xIPNYfrSc9AS6QlcVybnDIyODVtKr7uiLfgTT4ECpJsIeGWxwv
xfCk6bcXtQ4s9xbvpdz6W0rVZus/aelgHfauchTiOf1O6TmsjwW2yk3dpSM9DlvAEaBcGcLNKA+W
KY+JiApCzQfHylJxm6Azv/xUt+qb1s1S7ub8Td1Nzh3kbQWHYawI5MDoV5b4CFTpCYTkjXVQqfik
arilvGBDJxA48xmNaVZhIQGumr9FvfZx8tbRucjp1rWXsIp5LvnSWKrc/7xdH2dPHPuZkMXzUe64
FoBWR7Js34Bc4YeiCMCTbSTWtVf7+dT4TAPZ0qKbjVA5bDzxeYf3sc2kkeUnsP4S421C0p81UYNS
hVoRYngjHdAVKtJzAaQ/ONh4iqrzrm3QTFoPQImZaFvI2Ft+cJlYGMJk525UfXHeurY0rcc1qMFU
1ePtCjnKBFB1WwzNiKz6jhN6HMlOSeJvXx0klvvFHiblAJcvBcg5ZkgLBpuLrlRdRqtThoD0pGLA
2wXjtOsk65OK3mlJ8PVA2kiTJI1lWicXmPz6D1hd8O7lZRoErYS4pIXbPH10kIwNZtFns/D9GJ78
BJm+fMQSUhQnqTzCQgljiPCU6MAKa1G39NFsiiThAnb0AD8HW7buOYl6araVWrzMejAmQEv0yNMb
3HTCcj3FRPqb9GUTtIyFTXBMcYnN+4JQEfPSRwClNlrPyID0YMIM+SWWVOlGt/+fPPA6N+QaNQJq
Ly+VpPyHYeO+2npUlojiJRVNJWRL60vYNX1pjZnp3ki+WnihxIf8beJYn0i7/Xm2JGErvDZs8DR0
Cs6GynNx7nT7UgNFNkO6dJpvToY1XV27KzovRyLZSSoiTdSu09N0x4PwZW2dOHh9lbYe+34Bppz7
xRNs5jOtR2kcgCh6kEJ/Ypr9AS0j0fO9AYh7W8pM9933ipVwlQFJQ1i91+mnxu2UhtZFvwj4XTAt
kUKHGwIQNm9lLBvkvFzWfWyI1zGF3QPHKauXKThM8gPwMw2gS35lt22ljZ5WTWMiOgQc07c0gxn9
aBXdo8HszBYCFfOqVFDcQBvggPmFFhDe0BvctVNScPRaPRjAIjEiMc5NqXrN6d4sTPZxsOTh2AZC
HLw3oltEHwmW6lzRmZ1T48Ta7Dnc0HI1gOKVn38+u6DlzOuG34n05VYqCwQiVYtI2DMOwBvLYedw
jer7j0zLYNCwyvuyphoVJ9K4ObsUkWzAtfCTqkefP35foDSOVQ95Vk/tMwrw3SEHhriXUX6J895Q
wq06qrMoTZ3nQrbiSnB5OmbM28BhOlNiHOVc4GKuMcR3lvLNBYbdZqnzfCK8MNM0Nj2jrNDt726n
L8MKhqvY45lVXC2PozgCA3zljJbXCqaAXfjj0rm+kvUGiSqvvb51NBXhfRTW5euIFzYyf3GHkXiP
Gka9KdCKpnnxfWzjQPFSd0qRrECd0Ep+RISH5QsLJ8o6+WvFo7MELs5jPNqKMT8b7JQOTP6v9o5x
EygKH7QO5O6qdINXR5th5Ikb+oOxU9SZR7KRkjrtNvbngLfYCKEg2E6FSzhtSQALvnX5dyJKQZPG
E4juahT5kkKv4tjrv+fa+4/QDQzz9JlpIgeCz7VxJ2RtF/oQJNxVOcuz2Z4iVOSiXyCK1su8Rd/C
M0Kjk0G9ZYKlYe1s7mgE6gDRknI1e7a2JV9tcAzpqZlDb6/AnswwvdUrx3w1gaQcT1ZbyWZJCL2K
n82J//rdRY89kMzib3BfXvud+fxFAhlaGv3787oneFANLOPRU/ixJqoZyz3RNY2Fchi2wbFrcS5m
c+7DuGCsEYrCoEbeOqw9IRrantq5SThWYTDTelwUxneERmfP6PwCdl3Uy7BkYOwrlbclTvehodjl
Xm49CsA2pdt9fczPs3qlvvHW0h4STk80APRV1Xp6pE38eu3nfRjkfqnCXNcWkJWg4y/9KoNpekno
Eq90xWdYNVI61BpWRXs+/YYDwVHrvikv9SzEzx3BT8Tc3ZplL9ZIuVDDEZ0kRyOSqn/mgXy9+YcY
gnVhnwZmGP4TJkHZzZIUqSkq+y553TxM66o+vrvgWzeY4dvY6sSrMj8Bp6/kd1iLozlvBBEjbZJD
DG3ADf0Y0I39CB/z7XUhGEyHfutY0Gspu1TBJzmaQc345MTEa7qKMMIjfmKxFMFrHhEF//pNL/7H
oqYzrSA9fabhOMPQroJBQgm+Oh6lU18eRYhd3SGPUe3dQFx0niLJeLV2S0f4UdNjM2ZSAEMqHNTF
s3cXFg37TLlWrevIiDill1alKqJmE9nFbCLIef8nw+TdTqG91NOHDbSaiK3dLs0QbsMFWXa6l+Ir
UropIjfkbEmG1ywdRT9TVoiWeBgOKU71dNqNY6pYwIUgDwSNYgPJOa8BXIThcXXlYvmw/dKj0rIv
u5FZe7+jJwwjA7fGWayh5xBYgglASGnK6oXGwvH59lC2WVF2KdUKVBpIepaGhM4Fbf7TQSACgApw
pOM4FQl2Kybqbx/GLUd8OsGbNR/Q2T6e3ix1yTG4RwZchZkx7+zr3PVjGo0qSrRF08LUAHxfUgtY
QDcEQ9jU/PFRTOw3/7k3JGHVhYxBV7iHgK0Aeezgf18roZvsqQGC78UbKP11EWc83OGcbwEZxKNm
/dFe81sKtJbdDLsATS2/urjiE0Uk5HCfStsijWjWhXJRZ8TABgJveiCEXr5ZtsRG7WHSbRwtr/he
fcRTumCIoCNZDzTny3+afutmUKK36BhcNT/qq+oQhH+6ciQEkr/L0euH7FyU9PQ46lrA4kocoYs2
DFwUng5IGAJlJJVxdCKYTP/lQ/9eELQb0W/YEcDWYr051pXIV6e0zquzrKYZ8eJEZjoRl4w6tlMx
TbMmLBbiz3vFLzPgG/rUIEXFE7i9w5DatcCDaZ2IP/NC8ulB/XOLdKzSVHM7UsAGdX7O6Mf/xj3w
LGE6E1xz2b6i/VmkhLGYcJogtyTxzfGtqc1oUTaAYjw79jj81eMncT7fP04ZsHOdAqmtfYuANcwJ
PjuQ4PREFrd65ypBWcXKlfqWRnGYjAISOX3ZznKf0m87Zcu1J+ZFib6u6WMJE84vgE/2KZatJG0B
w1H+gS+7Y4K3sbLtb/bIgG1V2JLl7PhRJMlL5ggZPiXPKoN3OyZbYlGtbyBR3dbzKwHwAOruqLnh
+HhT0XFUgNM8CM30MR5PNIwz3H79+2TUWsBpKoLk8Sn/kZonCeS//9KYeJJzBQA7xbSaX7Up/ai9
KJrxMA5C5PZbSJSoUu9tkPvoN/Fx5XItQkf2JkjeXbEQvfU36wilBePvdJaSn9nhf1b0LeBa5P41
fXxOE+i3JywYNaDoR3kgnzl5N1H2Uj8ymzWqslqyGxcptiYneAwGyW7bkFLZq7Ko0C4JPKPauJhQ
p2z50oqVFvZddSqfRNqHuAIkogu/2ti/YqpuqOTCj5JeRY6Gq2wdgluSx5af7qD5gOHjfqvsVMoL
CEuxqsaLwc8bssLRicxLj1dbzihXOjdnSLcpA7ENfoxYjHAcv7B5k09By0UB/V3FumZiEVewUfEW
uO7EGZbdJwpLup8Km7Hj+MYMk2CC0dW53oNIbUNpQQ1lvpm20d+GkmfDMADq8zoc3ZlQi8c7dbrK
lNhcxCiqf3wKm8A08BRNxoZWnanOCLlRyk+jvjpZhCRZg6eFStmUfOK0fnJm8TT/SpTFYN68yNus
FsuEt6SXoFuWwLaVDhmEwm/L6XgU/HvyW0tQN9sBdu3mDAAwwgMYMNUndMM8lqIfKuwwvYP9BLgC
WFkTt85GbVSCXHEY9VuTwUW3q6jinRcHleIvkh4e2hd3eF0wugFS0NCUTc6W5kfgtggomKXhCwU9
ysurPmGtiNWDL0staqXCzbjXSDtWptHFSYtwzJxZdnX2LPeb5HDelydcs8Am+c85xMd/w3Cmsxzj
LI+X+vAXRyOcHoXGO8tuHBqLDmZsnNMz1yw4ltQKmlwnZmXaRdNINAUc5Efdxg3fTLNUp5Z7aZhk
uMnyg1ztj7uGupc8OJN/ch36qH84DK0t68D6ILB7VjvjF2KBxcUo0uszI1RSIySJBv0Spi4Xsrnz
mr2VB2KxQLY86BER/HIVn7BFi7CfpQhfdTD3sLqqnCW+cOeuGPf0qGiePH18t2JevtaeAe2c/2me
BuCKqnMqAbkiFJJ04ROPZFERygWhH6vRpmea/kIc/mD8NMqKxZZQ4nVh2tAA1BeQGBGyRRvxdvcY
h8tIIBK2RxppQn72wzg9x1Pl4Ef/njj8fdNkvCDgWvv15cMLaLdp5/S7IQDSD1D7foVPfQFpWoRo
qKZj1yFOCK59slQzQzh36rSuzs6M6TuZwBLP5dPoYCABV+bjLfsvwc2KYjwL+D7/ZTvED/QD5cTM
Z1gDhSd+VtsCMYfHVENdmm9rNZf22gMXK/QFVJlP5LAV4GFPxqJyNtkLCy7PopjAzisaSyMTrkIF
BpZGOKQEwC3r/Z0b87TpiEr9FuhMlJSBHkeghSifdNAAcUn3iGgdbOl1PwzFAp8VUYVWWdp/oHC3
KIQZDG7S8+U4ty9UoDQgQeE0WZuF4Z7QDZYnRPLg70okOgy0jX0N8dHJ+JTsfzyt3v1zLq1i4SMA
1YTQiess4D5UzUebtm8RM5bc4FBnGqB+oq+Nb3yLuCEa6hzfnoYg4dGmBPuKWiSeaVoPJ9lkl//X
zRBEIwqpHPeHA1aqjZv50QSlbQr+LAR4YYMqcEiDB4yl0/lwHMbntHjSgzfq9MBbafN8w+IIaWEd
7pNR4a8JGVNc5jWVPBaSn9eYjvL26akH27dzusHddJAZq6Tcj6Uu/TxqiN7wFfNduumD95ENVNo4
h3d+ItWhY3vrpk8gWOQ3cvnRQVED3RbyKIfonJXWZwTAE0wAuRX1OhY+oayBi2tVgzFmvfPa9BCA
aKkA9wfMjRZF/Qu0Hemwu8luWUttVIgkx+XRidpdh5LG3es4RRRuDmHK4KQpr1dzbUVdSkFobowi
KLc4Cdo021Yka1F6IhvCCRjVo/9ek4tLhuQJsW9iAuTff1FYRUX7/Yjr+GqOCdmWn9i6TL+gQCNg
FuG0a8j98ZtD/hZd6wOYxt4DAWpInvdodb6G9KRSQgvEldO2lWwZJd/aV2OHclWoc3yAKdvxPSy8
+2hNfinfBCwcvAMJJ4XIDrfO1cxy5g+fVlFkEKL2zRxKBvntjqVG0QS3SPEb0eS8QpthuucWE4kf
uPVNX3Y1T5HINQzSSNqdyRmJpFemYqUoefb5aU5+uTIPf+BvrEIZzgvJlF77nbwviS3y/zo70q8a
ySSYsR3qCOdKL23FM8wmS3MoEc9kmWP0uhoNlul89AZqlwHq7lxnDEDierIsOwkEL7T4ULcHJdDr
jLNtFFOR6MO3ACNgMtcVyCvA3hcWYMLHYk0cOs6bOSPPO3J3xm8Xzel2JYCb/y4qDKnXnPE7d0QA
6J/MRtjoCH4ZSk+TfGRMIahn7hZ86meYbVI4fpSYBxS1YTbq34t+tLheLpVgK6k9AJArtKeStn+E
+AwEMp6kSG0MHh9xWCnlK8X6QmoyGYUmME37s/ddLMrrLPI7cCT+yVsg1C6s2GGINEuLW92QQdjv
fBvgkhDAEUbcHLHUC9XvbgAp+jbKI8ygrFlslqnoMqGzMQ5uuXfYijfMeSxI+nKC+P5s+XOXcQAM
R8OejnyIu/It4yot5WApl45iQ1bvAv24Jgw0vwsPBTxOh4deOI2K60Lm3U/f/P8eP7EF7/DQjYaX
hFQ/muGkYjIfvIRQSf4sAaD3j9y/lmW9DZQRTtTIXQwx8W15qKgROgf/0tDfsOiyBKFkA0iWVctD
3aH5CIHsOB0knb26aD2ZoiU08On9TwxfnMU/WH3AZl38WbJpnm6Mkl5chp/6QfaiK7jc65Ysz41Y
uq+WrxndeD2P1/g8Vdh0d7NY1Uc/MFuhBxXOOvowE199rWNnSxGgcDpR1lH0xyJ/HLND7Xz3pwZz
qbVh4Uj6mX1oZ9biYE4PBjrLHON3ruCgZYf0hK4VLBlLXOMsmcAHKhMEOmOH8WgkDnAqUbBOQGaS
VcqFlFTeGxMlp29KXMZRzW89n9fz54b1HYtYY9X0sDzphGF4vPjRrX7ynaNefYvauEpCVPrGfyJo
OUTWfUlgY20fqEVWUt7P9rAW3vl0exeYhTyP9G29L2Afe6uI8W0noK4A8RjV+pwS2C4iE1e+oky+
yWPA3gfjDLZOBj8+dlk0Ogxz+tWO9+WyRrLkcOrekvkzR7GHXVPqpBa/Wnzv+fS49iUX1LF6gRR3
HdZ+Ufgwwe5qJolV179ZcCVzjpuYn5Nve7Q/jPMb5cc0AgsOpWYfrq/5XRnt0e7X6YUZ/15G4DTq
m7F0YrFMsk8tixbZTWXNCnm8XxuNN7eI3OCFPv2LoP8k4+xm8dxQfmkV0nnA7xYJrSShw7lzuMM3
pi0DXnLRU3dbSFkL0LTd93kBavMsaj9O/GI6gsAgeK0iSjVg3Zs9rVZ52dTs3LZLxhq2s2Gnn324
sjFIykBZBv3jMrt8e+JX/2FRjev+4Z+5sje2uP+QVGuIB/IksQcQp+oRh7S4FbMBUt/gz8C/kgjb
XrsBJK8A2JIXtmkUdDjQuyCKwKoKteDxrc3wgvjzPgG0fMu/PCP3WBMwAHM5qqz+bO0xbuOf/Xzr
QtnhXvo7p9c0vtIHzDlIRsbmedsZ9T+1gUcNDcQevh1mHmodRM5yqMNJh4dkzXMjCJfgHJqsCBcR
zFVbO+9la01hCobv5Vro7iIY2syQotCT8ovZlImWIpq1lI1bnchlCG8vYaevP7Hfh2LTaEzb//05
c6EHrFd3WYF5APQb02vSdKnJ/cyg/TPiWhP87iP03/WduluPfTKZqIvKIQVShnF0U5tguyUvA5A4
WM+QjAGZH8xyZvsLRnaLZTSh2QgbLZ+pyH482Tf4f+/F3uOxsllOEvZXhRvZDmYUGkyJcI3IBHQO
wVJjgmihBkiDdIn1WRaLB4hoGylXyrcz1uCyKkoU+4uBaHemtzTxwHff38a6WD3lgpaZ8u1/kT2z
NpSrNz5F5GX+8tDxqtOdblva/5OfgFwafvIehFtIIc+yhxTDnieWowTBDdmZ8ytE+SeFWhLQfxFM
Rvp+Ym4w45qtsDT5BYZUOpS8W5UH34iwfKzvlrzQog2XawY+Q7a4FwMhGzX046YfLgDQ3tRkXLKU
x8bF510Mx9E4hk9XAZ//79q0DMAFIrzMLf761BoHXzMQSFQ/LWKryfHDSxNrwv0VSr+rfJSbdjPK
qaSw0MtQuBkgJHDvKTl9vMg0xJrtWkELbHYXpTedg5TfOFiq9sJEQXMGhZHn5PI6Xy5XHaFqIp89
cuwAbf/ZlKdfirGP0b2TCFVzx8ZIaOMp2M4IDgjiyQ4eYgfS0XmrVCRcKJiz/DcWZGNulW6lYHhQ
62qI4WQsqwb1DiaBUpR3iSzuo8CPhHsCcxixRmkDBiD1sMJ4kg40jgEO/F9F+eqikQ+iDYjjLHCk
Ova6ssFbpYqPdM+NwSk3fJ7UiwCdtICzdSrH5CYwc2h9+aE89kFwV7iI18B3JjYHBXOzdFUxf8xO
AMdRrPqVycBbXp9P9GSEbVmsWMlLgsW/M+lgFGwKiPK3kEYeW615h+bJP22AGx4gUVd6M3JpWfu/
Gnh3fbD/b+PuyMIYsG44ScIQGoO+MCq4ae151JRkjOP4z5C0C9628vDGSgY/IxV0y/bT7XM1GagY
AkqK66mfMfSoJKbnS/p/JXR3iTkHPoHABHde/QjuWwX5tapBp4jLhqAjVR6tY81recOUqe5kjvzu
u3neaZHXwckrwUpz9pW8CefLHMEGWHHgzvU1ztUzyAqO8y27xJS6ZYvcw6iYY6oBl9o8RHxOFJXR
P4TtgAJd7GWOAyOCDe3ZEf92zH4ZybQyQzI0M4nuRbZ3EaKoefkjdmEk4w4CjipiUqkq3MXGjPxw
UHEyf7sTbGBSPAcc5PHb9hE1atF6r3R9kjZOc7BJuVyyAAn0qX4UNEP2/U/Xhs/72n86exsa4DkT
jE1oyzJqC72c3TX42c4EeNvmotavaMq6o8rww3NbAoYAxCgFE4GolXrxF2LLIei9qyHfMF+qJ3Jo
4H7QGrdmu0m5/Wb+S2fpZe4B7pfAPYYiHBRowDYyIP4LEua20CoIRvWYrqenPV0e0BWUV7DfaFRJ
IcWrdvXUn/AzPWrozsB7HCZdadChYnMiOY3qa3dvafTfUH4SsxMD2hpHTw/vxFjL20XlJNeyELot
2HHkafL9zcjX5jOUn1LNoJ38IUinhF2cDU7XsRb3yb5W2m71FND5GBSsFx8PBu1BGzvuz7tkNFeN
QN7C/C5q7kpCmOWXTfXblGSWOFGh1dDrFH2auME2qjMj3dY+bTI6poPP0OwHjPgGWAbLiTiYovzC
tGWVVILgENXLLmcKdloBqPnxJCqSgUPH2/YLmpcmXYZjNuonxtd3TX11XHZA5CuvfQHzlfGk3sDl
4c4shU8MP0wapDTRvMXqucu5BnOAxA4+SDjelZSu5BjhSuq4NzZEn/MU5OEqpNvj9Agn6zuiY7pt
xW1F2CqXqXlEg6ptFjBwJl16ky93tBfKyKasXEmNdup4i/VCboXnQa9li3Q7XbOTpJG5s93W0bhv
Ke6TVqpoZM2PGp4XL+ORPSPsHb4WJ1AxnZF9fcsfMb9BTochLYdHfN/ZvlT6eML0jzIaz41RTH16
914zZX2OC/+qhwG025oHvI6WDOn+H3K2q1A4GADWlAUqQVFIzjmZP2hw/g3FXslpPD85VpsWZBiq
yfMGKz+81+kZKCOPsRMXjDJoG1FFkqmKXpcqQ9l24st80Jy+dcPp34B35MwJtMFLOwXsL3naJGmE
M2lpQm3U+snScGNeEE3hLl2I6G6Y5jMBnJo0hxdOFiZdAcl4pMIAa+u0T6Vh3G/GjPD3eTJPXrQG
UezZI8QHRfq6c++8ONOz/tyqMX7/GfpNk69RIz4cMcJpPhAbTuedcC5QtbeU3L2rYGpq7vUETtcU
Tpmvm64UGem8YW3D9NF0DLIetsDb31JPfIKZh79ielYIJGWv/KupR6pZ/O8tuQhBWAG6nhgXss4k
pgiO9Lnq0sBVs5NqrC3fX/DeWStA6MBf1LgVVdG7eQLHTcvTiyk3F8DF/youqO40cpDSnm2fNt6f
fbYpIQks+qjMuVVsee3/Na9OOd6IvNKjF9jqIkQo+Q5wdVb/YHIH4lfmRuo9d9p4u0Jv13N4f3g/
mhuQDW+67PBpb4uVXDIFRMoCoD+FPhyOOc3HgJTfTCiEqziDLPRJRYHmTQu/ZDneK8k1BB9Nqlzn
CTQerz1znf/eZMRoIJ39QdmjRzQBY5CI1BVGbmOmPMj/hyngaq1T5rYrE38VJuU5DWGuv6SK9d8u
NpvNUfcDqnWcCsvj0DLqUXaxCiZ/mGFL2dJFdgr6EMpQaBi9jTYak7TWUVq6Yx0pklc8aSJEmdqZ
TcRjB/DlJPidiF6tdt8z6O0rnDES8fPLDBQCNsxFmS789mgNZW6yFSjhpiZE/zyc6hIru17SaWly
k0preQXhGPBXeN6lYzwc3e41Cs5RCwn14c4pupPRzf0Dsvf7UpaWeK8GYzMtk6yO7YEglYYe38T5
PgWLq7rITsptTXktO41/vwmrt6arO8nF3XtWQwGRIp7AIxwMjxu7wZlEvYGReoZK3W6aDLalHDTz
WIrHR0mdM1aJo6EQ2aeLzsO2nKpwpS6bQHPu9OELKiCojSFIDAfOh1fFmL/vWaKUGqP/AliV20AC
6vMRyefK3Z9/G9jaBeci0drPjo/bGum9QqQD4ediIvLmYWz0eG+9THmNMqekHIa0oEWEjcI8PJrb
ioEef8ac9hs20cXc6P9+0wGGpJHXXQNR/YozOTe4bx63hyR8dNcJtxsRn5I97FL9yy+hskQxjuPZ
R9bgIC/SQHerC21ys5KkdnnWLR1CzeaZNLguFzUPoZ5oelkvSnRP8Ha5nLnnYNSAXh28Wy4sIqcG
NHq1LakngYGQ/veVard/933TLs0EaK9GORfwopMtNB433OpMu5O+FgXxOTvLmw9vfcnSzHu91Mat
9ldF5WB0ZgAEr6VV6PUZfUYjNusx43HccEslX3x9NxcfW4107YRlWv/JA3cqyhM0PwUnd4lS0/rm
ySWg/gas4lkXEcl9jvcIZDvVP38GncSdkcGn9nM1SKSanFmxOHNiTTECxkfTgzfdvyH3twoV7Uz9
ADRoNLnEwgwPsxFZSlhiaCxJMtfPnRNZYrYNkWqmta4zZCB2/BtFAUzDrRjYNs60XloxtzOac9E9
o81qE7ZtmE/nWRJMpbtIZMR734kEtxXizKrYHkCfz0T/TRT+X3+oJBDVMHwf87KMh82C4RrsYQT6
xcgHGaqGlSjC2IGb1iQkNPRHZ24ACiuhb0pHquIjAkRFYyTGWA0EhdLCOrMPOODPrbl4Cg2wa6kP
iA2uiCYtgWWIo+4Qz2D/PFgoVfLvJ6KqyCokCd76Da+mzKV/JzrhKh9NlQ4MQONJk6s8fqwbZi1n
Tp7diw1T0HNSn+dzHjbQ0leb2QBbVolp9sj0MnwQelJUlQeEDxDPwZG0o5tQd5hGA/EwvUnmJMfY
BDTyKlRvDcbqxD0mQzAhoaK3FY5XaD5DeVqZk/0d5GML8YLIv0i+GPYuzE75FkRZaHt3qKq+YO0H
Gdx4h1FVTq9aWJ2k4AYMQpe4YC66s4PDhmuKfiIz/GitQKHKw2KZIRxl8wGvskKBx4K+kPfd41wE
5+RV7AgZLai6K2/G01HBJA9oORrI+7S5YFYwQkVBBb7IJcK+FE2A4qah4fBF7Qk15/4ElzVnm9NL
HQuiFM5gHS9+twYogUeOgvL7OGutKiSis7lF+QkWfd7EnuxCmtA2O3np8wRw4GFwIOKVCOyUSqP4
Ch5i4k47EvBach+fzQuwJffb9y+cK2RKB/UoMh6c13TmcrhakXbsATKH4g94xsIlFGy2YjPa2bnP
wJRwIdU9HTnDZa7vBmZ3tK8uYeVqPIjbRpyWlBaAdaWvYgOafyI9ArMzfxtA1jdhF1mi5C7AcvZ/
6B1CZhjF0/tL3BYq7i39N+jhAQxdyZe8F4HH8Oe/PBrqmH47RTho7ID/OEMRrW8b3OZyYy2UHGWg
YSzp92xE5mdMs29yOPIpP5cU2ZG6aG4/CEbTY/mbtrZWUEovJW/X8Ie3yCk/kalc4YaBLDl2+j5s
/QraClJvq5yKxGV/lBXv6dqLRIcibxkXFMFDeaZaKlroxvot/3r/HE9ppzZQox5ovYCWk0SSeZQy
caUKEq1MWnH3yy2t6tlaSUs6Ewa36PCrlK6Vtk/rl4qAhj/VhMtNyREwFhw5qQw0juITnLrsqeXk
NSE+bKPUe3o9wP38VFwLmlZQHyXAuzO3KxlT/Wp3VsN91qSG0h+1UlppJPq3AdoF+dRG+NzvsD99
9iyB+e0uMbi6+2o1AvH6QIjSHrMPkf8bVK6hLMXqUB/tdtrljQPooKdEljjPoWgafBPyUF8v+JYI
s8nORs8VhDctzzusIFwzQ9kHKbiONakwuN+kUMBPBVZ9Xym/JmYg4EiYSJWU9uqwimiNMKJbIHlh
TOjmLlBLbA/LhedYsq2oG5sbGWjlnaU1IdxWsBwQrLWTGj2sdtWkTQ87MBOgUneNMgNbe0+g23gE
DomGfBycdGGyhDQqzeeK/uJGgD0W7w0w/LunRdHPmaNcTNLjXD0RGor/XV5S2D8PX7PPatHGNVkM
s5iq5nAIV+stuIVlKTF9FWKgXBfmZ3jSZ6AhsYEIWLMpE2W+VzjlVIDGNEOEjVBEELm00fdcgJ+e
h1y4O3xTdYCZV6MlpHIf9u72IuuWAn+yv2KqqLXvrrANlrOt9jXEywML6FFvzVMJlVk5VqoGiyfF
eHXAE3uORsthwVfuiAZolSiVcVQBaGpqBwFDIl01UANg92hPg2/K3Lj/6l2qfCLg6hGy805FxTTt
AFnPxqKztBKBil/o97FzWO8L8rxQAFDyTTkqN65F9bOUf7UfPxHcj++9Ei87YCFJ2Kkvhwv0r2EP
Wqv5pFnaix+tKN34fH57qPi9eYP24N1Rw5RaHlNZI7c41bw8yQ0xM3AuOXv0UYypR2kRW4r7QRnF
suZMz7zH8cSN9pQORBFc8lB/lZ4p35GUAfZE0n01If9SThnW4sXE2AkpTSoimw2yLKB7fhNUksu8
By1fRMia5FXrI0gCwEDVbfWCcQF0zqKL67hNDK6bvYJnQ/ns7AJqQP4biegYrhrTVz0q6O8dyuWC
bdL0Ibn3WAA5EYq2Rx8KU0BcXEfbnJcJcZ20WBc1lgQ7u574Yk2Ku/rH2vFtMT9rccQkKdd+QBiV
aMfaS7WrlybUYENlR43fIPNDMwopIzDEBA6Zd0l0q45Wc2zlEmMZtnve4dLbnIzbNCmKT1noIOUc
hijsI21e4BBn9/8cGXvJPPz9S5A5YlfSRAgogHv+tQHD+e5LCZTwwviFynzENug0aULzjMT19zTC
UQTstL389FCIS65JPiquyk7gadtImTFEhXuMNDpEn3fP2sWs6J0LAA5o9jioAFIfaqMIS4MSqZhH
dLEoYTg0rLNN0Eax0m2H75rE9UuQbuTCm0p6tpMCU52xuhrTFKeMi00SQJc5RQ4IZV+06+m+IjtC
gl4/EXdNzkQTrRG08Lr53CpaZfro1X1XTFgVuxQgdS/utcMy9Y2j4ZwIAPnDr3dMTs2KDs+MKTUy
6clg1EcrKrB3m2YrhvtXnPuIshjUoC57zwDbSLfLgPMutyo5fdLqsJYD/GH+QLOEWd5Xqnn35BWt
DdtF1IkPR1pPjaDz96m/iO2GE2IzGKMiWlyopZvV15YD67YW2LG9qIV1WG1VZw0159yh9YylIupj
bJYfETR47dDLLeVarfrMcTYbEMkrKLG15swmVzT0H60Fmt2wAzVKmZEh9Py1fLH+2YCnDGQaOhx9
Ymu2RZ82om17T6nuz0IYO/YiHLrAcl4QPvGAaaScRd9CyrMEojVvS6TFOG7ZRo+HSfnDq91mbPdw
pcWjfBNYESdT51hVlBDnJrBHwxM1f2mWAbcWV0sQdH49v5ScDJxZq+SL+uhR9EKcSIT3dt4HYR8+
aHMy4QJgD/VgHit83kXCFOFeahXjIBqun5mIcgdsTWvnwbNWTG8Hb/zTlpFWKTcODAliKKJNDrRo
nLItgHUoWnOjFLBWp1SzaXe8bdsvBFxGwjAZQBVaclZ0qP+d67VH7l+eNMq3THIvkumkjL3Z5lFk
uCciIKvtIwao8KeaOmOHtLfyUOoO/zE5ebqoJBxmjL0JjTPcgATZtbD8tvB5H4Ql3b+FAuVsVc80
mPU7WEJKuhlhoLApMHvIfGfJGjS/qadFXcDQuXF0Z0KEnJiCSKVbjVE1vXTi0/9ZOxcFfa8hd7gy
ylUjAgj70G4b9+BQTuQRXYYyJoV3/jw0WOUgqdr6Fzc8fsftyBvb61RgCrj+jubNG+uqdE9UQCuB
b10tXrwCQ7qWCTNJDOn5iszwj4x382Z6TTBFH+phCjDXMlLG65A+L36OAxnqA73mdeUuKNw+SoOQ
bUSdmvUbI3EkvtdrM6QXeYQIyRjblfA2CzqiO3bHXpsIN7xIV5bqKZtrhfHAieS7PXd94WiLKNfx
yVZ5JkUap3LXc+pcqdWhLjxpouQNBat+ALupqljvhEFIb35jmjjvPJfFziOuy50H5/cC1QX+aTvr
MidCq028mwQ/my9x3futvOuP5P2FJLQ7mfxjqRsZwMDRb2NJZ/6IPKOcFcRB5D3toiSNIvBXwyPc
EXzyHLk1DRy+XBilZgahzv1NZbDLeuWAwWhIituijSNm3e2bO3WWlzaQoj76DNRnhFoWTqF4j6Za
RnhzKDlACIs8thekcF4A9WMpGf6K1gcbm7rRGjATjKLohrBXpgL+X925e6hBEwoXnEQD+zW/UR3Z
7BveOkOWDqtSXOMjRYnYDHT6yhNeJyJMVtLEQ8Sc5mgEE8MAnBWP1WsKK1rdDctyyPfRGPpvUmIm
AB7uzKXGBZQxfwUtcZOAypv6LwlYx9xqcIFAE+XmW7T9edRsrzLSjPtgoNbGiClYJKAUJN/uG/NU
a4PPtQp5uPUruv0HrwO/9WEkZscqLUGXbLi0nexeYW18guwAWJ1bjPBOyQpGkGmEnyGCxhTLDbhQ
EetTTNg9e/RbjuL+6Ax8itsYkMRErUfITtMM+11k3GrCr2fd2f+u9l95jKBEHmphWWn4b/vEKh2W
1vLoptf/bEyooAjB1Tz3G87NRjMAQPXYjsJUpw1ifK2e2P1HeM8rRcAaq4Y8OaIxKN46R6xysSO2
hV7EmN8jMkWzFSuR61v6rZiLiPLHrTvaHCRs3Dp1i7rOWPctN6dqhM3b+ndMOjP7oIsMgwpZUng4
xqEIOy6C0MsfhVZlaAkU3hn4U4xkPIOW5cnI+BIUExLuVaXQoZVsfo9oSJl81y9u0vV9kKwYS6vU
129URNK4Na74N92qsX8Vk+a8M1rSsOxrdTlToijhB1gwgv35Lr+d0YuXrhE5ZKUSle6RK5JYN6E3
2rP/yTGneqCdG08XwSkeM5Z+NFwIlxVr41fFqtb1SMEqvU3eZTKsEFQmpawq1ppKSY2swXop8Bre
T/0ttI1y3fPskGT7pcyd5Njn4qMh0PDHlyIUcdM9CcFVi0OGL+hvZEhkXn1DiSyN5gOXszuiINBQ
6i+DusVpveET2oPLHiEczfbKE/82azpV2WtXj7bgAN/JtUshe+Wp/N5jIOTlR/3kUHTOnNE02EP/
MubXk+ZRVMhHbHqRBKsYNuG7qhbOfg7IspKYg49KKlswHd5k0L/xKFQRQe1At4PkcfwQLdSEkdCB
/cnVF2BXfB8rTVf0/DgGCZIYuQZI8uACa/9I/4e6+pj8/iMYaG16HhpUKYY51i53b26enIDZr4dA
JfOwNEqWH5kc2fBBjOXXpgzp3hZKV34SMqMZBdT8NQzcSz47L8YhjzrBYPIOw1yDN1bfUIQ0dRpw
sMQyAEEnHtJXKH6sNzXvaKtB9nKqVzq68oskyjjLQviqdU7fN/jedo0H61/JOOQNjT61NbDH3MTp
5rSbwPPojz+95MMdcm9hgP4oWlay5XAMZafywzx06IoR4g1aOjHdIbTjSgR9yHFf65gx+Fx177iL
aGGsHLU91ERhg4iNzQCIRhIWrbywqwysPItFhgVNAfS6CRoShFv91VyXz+aCSXr46wWilQYTgmrg
lJUSS3oK2QezNygFUz5AKljSJYJ7qFpTShOYwPKe5Aa4pQGiWPP/mLKP2OKIt8kUUMjg9ar0V+ur
smJakrJCIF+n+MKG81eDUempjRbudaO2b7cPwNw1Zci/r6lrtOYzAq1lifHvfavY8D1it3bJXqqX
Je2RwiL0iTTZYAN+xNCfDlsgJkdW/ieNpmVldv0x6o8rzq/9LVpT6mHiXe6v8WOP1Y3RJhy8w9JU
nqYKebNJxtAFrE5/4vLr5JuthlsaTVy7UqS+c97j9HnYtx0decxY6OvCQSvLv6c6g4L5aN3ilBiB
XuPwiAi8KKQuawE30cXy//zi2ew42KB+CyjD836Hzm4+bVPgxCISDRkqu98N2zJc/H0CURH7RI4m
p43kt+E1wk2HK2Jb5EYJtbCU/tLABQts8S6QiW+lgaQxlIiFuwMXmzU/WNpaNjc928PUtLlzO/DH
3ua7IvgLd5h2DXdmnAPhlL5TkYuSKvnl+BcUrVZeO6Aiy6r6mF29K6VOFQ+tUhMg63qy0p1wDGur
wOT8Ivmq2VKQ4AV3RwE1/dLm9VF9A04Y3DJ0BwR2s+pCR4IGtht8pPmzFXAIOOHnnjLiwaiy9Rpa
T7/3LFOLIYiFI+ZN8vM/Gwb7CJhPbuxLVltsvlBX1S0ogxagKzdZIZ3AQNrMObo03raoUTJ94DmY
zkxEB73qenwZ8smAJ3GpTHiPpa0AHO7+jWkgTRXUjB7SFuZ7RM1lHKQ2OlYgwTUk54YWXDoHP2lN
SUJpSwYwaTM2Oy614elF1Oi4tiDA2qFq70EDL9ApLr1lAA35vJkGelcagT/OlphuMAAnQV1iwXxQ
y3bBLBuAOtCzDCsjlaYAs3C0TODcJJ3FLSrch/sM5MtpZQbGINf/iU/cWUZjKr4YxUKOlo8e78kV
7TvT4Nqh7OJ95VL2ttxbifxpN9v2ipK6+kpGwyI7nkRSoyVvxVGi8Z+7hP+47D4ysP4f0YcGb5IF
36rUptAMfCe4PABHVje9NvBIUGvSXBwpXOOfkjUMNXIUq4fMdUovrDJRh2tNS6Agity6P1bh7GSB
xboZZ9XbUwsXft3qzOIMA25GC7Dx22bTd4wB/V8Br9fz3DMymxVMPYJbaKcPxQVqDPzZlz4TeFb3
xzJcnTfgO894JWHs1OggM70Q9NBIoX8lV5rhL5E1CTV2UCHf65xSoofyb42hA/EFgknB6gnMk8GD
aVhnr0Yw41uVW4EXbOD5l+2EhukTuwDe4wnJwshRKqn2mjSQXpvMwgCQENy/4Ui4a7weaDxn1Wte
b/I8Imc+1XYmJyBi2J3Mvsylf5OB1Xcp2vCppm1gpsP3cTGoPxZ3eETqXppNhXHV0HacybG73IXw
SH36Kwjc8nbg0eZty9vv3BVg9dcLqOhvRQzFZReXOoWDUovle3s4HAHYk0ThG1tl4VpPve5jFKWY
PUfT1tsctn4tnH4ZGf8bKQ1Rg8g/KfaXSvDB85po1T+Cty9kXBHuDB+Dyw95t5Uxw/TX0Q6ZCeZI
D4CaX9Pgyd2+ck8xPnwypkI78rvd/DNCufmkm3iolG3lgU1m6dHEzFLv01rjLHutRtyptz+ky1Ic
0M1mrrDWqrQziQ4j3mnyvxsdWApVT33vk1busvTmPB0mzXKhLy/4RSRwLgjMRVCvSOocskDIv+DG
JjwmmSzdlTeW2KClyZ9uUuu+QzRt9eX+kZ44VVk9opQISKUTiDtT+XCABZzmytAHHK1AMgr7AdVj
2ikyuagjC79nTktYS6J8cksrc1tWKO4oaccLWpVGZmczSjNN5HH0wXz41AYMgdvVLp8jYX7Y7NLQ
lZgd1OHfnlIudQxeVysZ70vO4/gT3L2oVeTgPDdESzdfktv6vgqlhG+H30Fh5jZQ3nl0uaYUgwKN
PkwEKHnWCbCWsE6hJ/tooa0FAWMwfALFHWeVRLRWpiydwuJM0kYaWO3+psEcLeeTt7l8XEPSNd0t
fjI3DDVcXGyOc9QfbDePojkxrpPtwlgaEIzJft9pnAOGWocz3DyLxc1FCCFiwlpcriFS2yjU8in6
fph53M5KKgbFse+cUYlf65N69K8jNy9CpcvtaANjp6PUG8jWvjiFPIS2DokEEOjk2zzkOESZhdX7
q8bI0AQCU/R8o9GnCgZ3u8cUAMK0pR+y7EVkWwjS74dozMs680LKikVHgnb2CJmD87x0uV+P7hc6
g6w6jV3KdkPneMOKO8RvvcpbdHFoIeo0ZvuexH14xHjPUfNoAFJtjTM4iwAHGhqt36AAAlyR0pRV
ZsXUuPR9MBZDeM2AqRixICmGiXoYX+DSL0ArXP8NsB+yQqfGXP5OPTwQbpgJqd4Evt2oSULMDUaJ
+q4o7ckoX3TgXUswh0WP+hIAgVxUhs8oBzoHq8P79bDWFO9ymczSX9X/Qn1Bky28K1yW6MhRsXyH
nwEo4b6q5NUqc4ey1paPSn60frWEBGJ5p6PbsT9+/K2jAjZnmo4uFd19DVEpz60SxDAjWh7WccLG
fGZmBM41XfbdrJFo926PEAGfh5lTB/ExupPHP1GiYxNvOpYrRXRFjrkgHP/8T2e81peXlNpXLnAe
W1lcdyY7E9WEl0CrEYzqVeEsSx+UANt+XlvtIqNrzXBZAvC1ETgXJfwEEt9gaxw+e9BkzEoJE4Xw
YU62lrXk27/4kPtkmxYXU4jRIPQQJsDSDDMfyCaZFp84BIm+hU2OYYeURkGLm9TRzds8bVIKvQci
VzuZiawgNryGPZQ8xn1IzmPbpF6WBUfSDXsbOCMs8swp9csNQJ902pnxDvt2DRLYGC6EK5gPKMxN
xogQl/4Z416t6PoBMXUcoosM4B8W7mggj2Bc3TkDk98KX6Ezc8p9N5NpuaZEnsF0Cp8h9KyDbeba
9ra77aiVX9luap6uCvXXJuMbYdDiyXj+JjFKzrzCGXoOytL7aTYhiVmfOP0DIZWoOSQum+yiXjY8
0WzYY1uibMovH7fYifGAlpa7U199c3qDsAyUeMjNKPS887BOsvlJz1m+hi6b0SQgqLDjgBlNkf1K
ach32P0eKinhJ8AVttczDeP1FVt3yqwDDt2114EJwQystCb3mhC+nj8enjnuV5M0sp+PR0gVn88c
/b0K4G9++J5ryLcLZ1cUemXnYJmNhas71qZdeDsFxpO0bc96WPElcqz04ajbXHYjHDlsEIwUy9Kl
pDCjuILvzHn093q3idjlhXAQx6lJHlIRu2SXGyTuCwb8v+6LZBRBY5rBqqObKTJHZ0YTpW8lB6Pa
99VRuLeJud04BAZI4Ly2+sGbbJUXY6KYrIBppIkSf++OuaJHaiXRXig/QPtApLBJfQkNfOx8oCQe
3wnE340ZTcBornjL1LTsFgBWa3DsDeOV4ptyB0DbciaF0njt1+5PFqQD7yIaRJQKKtRM0rhjhRkv
CH1zC6MV9hm6DvUtwiB1nUGvw7yIu8m0cJa40XpDI+t7oA2Ot39PNmhvDRTx232RA3duPUtRQoMF
IZkDwL577UOWPS+6gdyR74vi03DtvhvCyT2oc+prFpVrMVsOjQSGlqcyP+5JYjfHi36fH+vnGWBM
iXSUzMNw6tC9rP+iquDkJh++lOWVjFdhVTgoH3tvAN5GkotYGR/jegtgbh4IUJOZ+Rj/YzP3xkwM
yWJH+cNv1YH0kYX/vWtkrN+EPA6JUEHHnCcyLzM1Sp9ixCbP+cMraJ0xeej0FJulwyR/b8bO5BkU
Blc550Sb66jG0esL6vXPGhH1tz1Sy14jIFt8pD+jC72tIxsI3XyALnHIJNHWHuLYYYIPaNikCRs5
xt1fXDikytqAwc7dXhTn5wFJcsV/Kk65IMmFa4snKMyU6hkCTAd5OzCqrXR7Sy1q9CotRglAfqLL
xKTMQzbcZqTcHxx9ci3p54z/g8vCldnw9NaCRUuiUPrGBQQ/+7XRQKqKtnPvU18VT/3IxRP+KUPQ
2MTMOOfQ/yx6FHiOfxNeYYQHzlz91jlx6NnfYOFotPmXdCcJJE7xVy4BjQHCUS9gnnzc1vYsGOdq
dx6Q34DRI74ivi+CMu7fQM/gVFKuOf56wbhYybxlcBUCemBpP/6Byv7S+wi02Js4SSTqgO40hIsf
EArT06fWskcBpB/eXwgKBOMTacCJ6vyjHDZE5BlKoFLNY8TkaWCsdS/O0Rgzx37cJ9Sjy2a1/DjY
o9ZAUCM3FeUC9V7KYUutveJI7Ld1XtTQYRQ+mz3MmvPLp/SHHZkhD7cme8iTDDAWu9x65g9gmoZt
vg7ODWi0c4WrcZWQO6L1tUIWNmtjAQNsFh0PO1X/oclxNodHMI+WvGLLD4VVU4Ci6k7p+lCuBf4w
fb0mA9cdsb2q5GjJ08azYfsf+rDnpEfwkJ0nhfdTnIo4pJLKnP0yMtxoyS2Lv/ibDC87c7j8GH/P
S9YWJS2gP2jgpJe927Y0qRB79Jb7vZFLsS3waqJ2y8CWczICkzgpbLK8/mF0uOdPvenu7bxU/m0/
SvGIwdHj9LR00XfnzNpxhFzOikI8S6WJNgyynnQjbDOlKJY1T0X5qKpFmpDMb8S82rmm5ayQfMEe
1rVcqq6HNQo7PHU/gbO4SqCbWm+5tD/LD0AeJIytc3mG4UuTCqOtFK53943iQgYQ3YZk+7QtpAlA
flw2VQCPF5uZfGzRbb8+XNZaA/bLyexWUxx7uipp/QnIIG9W6Wj5qY06+iRiqvrJg/Wws6IMzx/A
v1UqwJu22KlktQDLFHfI2cRvmi1ihvNuTpumNMdwWaWBOKBnBWvSx+ppDOCOSkyTk2VgkeC35j8X
wiN2TrTTUehV03RcyUwlguyM5Quo8GxHlDrQ2FyZqJ8MQvopq6wgcXGZr7mdLopvnJCidHA5snSo
KCu+8XI5VOyVDWD/cEVmHjoqvlOi1pAqchNRyTs2TAwGtGI09cG65TkPeLqf4s0F3qWKuV0QMenw
ZVaoUz/8h3oGSg+hlwGuFqsu6V7bVgOpcj0N02h7MmcUo38WA4rxLyX73LpkI8nhg93b6X0xWp36
PceyFDffDDiEhQmWwj6fC0ds/hIJhGtVTwNZzyeycElishq4bg0eN5yeCH9x4eZLnhQuzWPflJy8
ZnSV3QjFQDSdOAJFPtBMnHqXsVKrDv12ugJBB6ZIjMNJ42hq3CXAttTfBVrZoDvvyNwklwxhzbCX
QhZ/k/R3mrnDindwKZM05AirBczE4ypfgyRr9njXkBLgb7G4jPC+xB+IOUDhZuG/c2ENpGUKUiqS
qoDx5EXXq7He2PJgdGIM8fnsrmZ9OdqMyt6V/DHUVQSgROG3dzscR4yuSzXRKk7sAA6zrYslPqzu
spAh7YfcTu7Wj3om12yuWF/+AbzVMi+MsIsYj5/f/EIz9lDH17vdfJADNgNT+w9aqdStDOKMFkYb
TwEp1NaBVT2z+wW2SEkuBhjw5dyMwYHeerwMQBdYkQVEfkE7HJhd9qNXx8s4jUvdlIPXlcjWVX/+
z+E8iomknXfLhYCB/upNvJB3Q76VuKLOojdkPUSnH8dC4OksL+d6/BxNJISywZBkl6LW7R5Kauui
PcM3IyFN2Hwzt2Vc6UhzwW+u3ErCnMEoczVbTx5sJ/VcPPUz/weJl26f+MSTwubfk/Vk3FsVIgLu
XVGdQIXPcGEHR1ZE2FYbTZYa6rdW2eJxkrlRApPOVesvnzEW/yG5AkElTQnq2FBpdkiNtwaXGyX9
TL6zVdBZcfEHOr7DzItKnXAiFd70neZar2ExMgBF9phnJhaH0+QBduepvwlEEArsWduWC6psYdjf
YkSt7kBbVPPbPO+501o5gXCVsmdUnH5VZISoBMzUEgMto6yWZ0N2D/FojyPflMz6vr+C1Mo4mLNv
oyIiu2ikA+3i8GUtEa0JyIFIg/KEybh9KKH1VYkGU/4FVGZpd0QLP6ZEUP2jXehshxvH1Cet/WNj
H10IJRg1rzJvpAHuColP4sByunNQ53cx8tn2Jb9y1PgE4k/K+eDn8ynryZjnrtgX10WwVSzYjVdO
d6ehU1GgjUFHcuPE5lZwX1IVC1OGpg++IqsquqYl27kx3GDELdTWAAPJYEGf2xMxCPX0IffCDuLt
FINlo2CCH55maQKNEf4sCxxJwf2QTlO1+pIhRdTZ/FhoDF46R54pH5elFZ5JHopHuOCygS0R4aC1
qzg4Quf7/cOR9rtZvjETst8MBFVmuziX4N9G71895yZZyrOCjO1xaLQqU5V4u2jHzxLA5BBLK5uA
pLcsDaY9MN0bgbrXWlffELYy+rG7O7kgrPMRYM8JA+RNuYJMG4Js5Z9AIor4+CSY75s5vrirSnTX
93xNRXcB/ics3ur0BHHSO0idxSDDqGrtyfoLRSWdKZ3YPo6xFvMHtYj75JLlKxMaOneBFa32h1Bb
SioSslEELmIsU7DihB3dTJ/ZxeG/RGsIL1BPJyW/uWPl0xCfX/7PTWtFtv83ROejFPa4VSsnaqQ0
7ZzTPwTSQmGDh9eqVotR4zNKCqUykRi88N3pzPpxz7w38q6wcY7Gs43pPMR5kSZOd4TlP/6rsFpU
vf60/n15nqxrCoXCsXKUeQielTtYlBFDpehndOy6okvtHB+8RIiJY7l9CZReK6G1ZD4MOpXKWEJ9
slR1xODxgj9HUHjWaWhr58O1JncVb8vY0zhZDWWDhRM+F10El2sBbvRD8H6j9v+IZbGSKOHXSnnC
5Xqdt/zo0JRRT+huzZp8SktuQB6jqAbPOtRcxqnI7450+zTRyFz0eAe5dBU1NEv+5cuGUP0FGZn/
+PSq2XGGNs3lQcTOZFH99Xgeq63VwZ8WjAY2a84IPAQfTa8jEufS1+EViBAjpjGK0wSZUlL2Tj6K
jMawVPIqniBUPc72mnTQr9ZrR8nTzywPao61GjHQvZJ3pOWysuIHFVE57qtSYSEaY6W9LQMdxCAu
mg9ZjAzpYU5fZgSBsI8kvU2cri5Z4MiJ+yCssuGqdCRa22vpChOffx8th+VxMuL12xwcaV0WZ1gk
HUJrzAFL3y9dyVAgnIqRoS6U3WTWi2qWUCceLqj1Nh9afE/ZLqdK58jazEKZ8zrTPdibGlpOavZo
U0776yfXdzJ1OPudUds4tGdC13ZZYEO/u+TMdM8dkIpF86LnF3qBahu4ZG7oN65LUQJtIa48o/oL
hk0qPT9Cqz7CPVWSP55rSv9ca6XYDxur1INc6Al0Nz1Dgf1fA6c34HtamGUv03xVwxGCRvh5bWOo
m6wjIueG5BoGNfG8Oci+rBStZKtdHBeVpNT5jGzdcpieabe+XzwSmNfNEYCYj+kVzMUXiT8zT/1J
pinCOhlKpb//yAcO7XtErwYhL8rcfXrzXiTrLcrqipSEwQUZCknZ5RLeNsmPcAB1yEOqt8fmHWM8
3EF7nRI27Qt9mwjVGeUjzWbu3vrKhDDdKEKST2G4tMbAe1kaj+AdMhCO1fjVnhCon0omw67w00E1
IKiu983MaS/b7dcRtTZoGldZ2YebY1LGeiOJa1gRg07bIRhSgUo4IRLghZqQJH8Z8R9zJys0AMxK
lPgtrhe4w2YFfVwOZRYTY9f2JtcabzPbaOrEMEUI10Vj37O6D9hJKAfVukANkvpnpaj9zwpFPRAq
f4Ei82H3eOFPojJVDIzvBZzkTrTS8Fi+wdRdQiepwKZIMMT4W4OhbypGRAeAg2U/bxi+XUxjg2up
Gg2UqNxyMZWtLgTg3FyAfTmeAZ3oG0FmUvYnwVs7E7KSxeg/XbUhvQxRbYta34I4IijAscUImPiQ
xNdAI6aZ3JIz6CXyCWQvOgWN0NzT2+Q8C0gz4M85rooSJljguNzN+ETfWBezk5Ic1A1Kc4VdPrhh
7x6K1WL54YH06cs0GfFQAHdzxCGltVazuCa2czm6BtKd9uO275uE+jvAPBTKS6e3tdctBrpxmBf/
1Q/YHFIhKEOxgpoVZMfF+4YDNlDn+AeO5YeSYe9CUVYFZQfXNk1O1Limhnn9KD8boVW8UKlJbT5z
2q6fw3yrvoE79oMRCTpfSOBBmc7QeklsdXOk4fWhmpMtzoycc/XW8cH/wXe0qPJ0Vo6SyofgHPkR
NdpxXcROIWPFuhS6CLn28NkXyk3lg7YJxzPu2evahQS8olFF+bG3uSvGS6NDU52WvJFkJhz96RNi
9ID3cN7odIdOWotQgkLml+zHvxOl9hkHDlZOGkQDeEmfifJqwljid5mnCET7a0tcHKNza5Xd/O7F
C2HfuC1WAbXs8ivWJ5XYLgFeKWqo5h7RrqNRtmY2XGN+ZTTLjoosKm6yb1l2Ge5+FYWO9tT5uROz
09rrjI/0mKm5lHY4j/eNMCux3pIrTkvVpgFWHSpcQa6yZs2UNj7PFIz7mO3cAk3vGJJbp30I8M/P
Z/9SaDMxVNsjwhDEOsKIeIlu+pz64O/n1ZdcoQ7Zm+P3w8SIYJUsPs1t7lhuLrnaIX5GcxIiKARr
vyl+rGLlKUwcbxHP6laRo/CjZBtccU+bkaZt2U8BJEOwT+sqza5iY4vW9NhntXM+dL9xOg+KPADQ
8PjzsvxKnVGJ4EO9pcxL406wwCut07pn1Jpgx0U8msr+8RDiLqJENSHJw7kr21LllY1PApdnzLiz
mCln8mIh87E9oEytg25C0PiSva6e6aWFQHLMgtStQplhYdsPMwcDVX8kqUmTNGXlD8hNbqKp1pH+
JAJpRG7xbYf/UKXbI9qQoe1HSKn4KErI66OVy/vuc2ugwKZyh3EhppfJPajOsvRjhmvrbzIUt0fm
t8ZwviUjtakHPZlQ0nZX5PNZrz2kkoIOhUE+4NgmGPcR5Ut/q7Zxh6F16St64IQxDbjTb/LNvPJv
0X4hkolwmdBXLHifsnIeOxS0Ijj3oV4Eaap/ihU9JQRVtWi2gHaeME73AtaQE52G2Rhlc5Kn2rCe
AU0simui2K7iQKvEZ7tLy00mBdGG1kaLXPMub9HlGxTHZsCVQga1t6LyVCI4YWh6xrKRwMHcIZSN
bV9i6gAT0pORWsOgpj1jQO5WC96NJS2IkVndSn15DHZIBSDEytEupSX6Cana2QUOjQVmwRL7yRPM
7yAH53bD/0GFg7LPP57asb1/RxL3OQTql2DNjg26opycIryhsOv9nX35IoXMJaZ1VSQ2ya/CwYIk
7liBURqSCsQ4czdeOWgj6rfUD+VYWvFZTAfWZ/3S1FiKMQ9cLLzD5+f0XtXfI5TEPJ7G6orKlQ8M
l2Dw2eLIHmq/x4uro/ZGXCZcc+pFnPSUkRjCIyLDNUGDb+/Jwy4ayZstou/G82yOO9XL+eOzBYxV
OL/qN2TAnj52dUesZlDohycwp39B+YaAZvaw4IZthqVMvwL2JjH3QAVDV5WmrXJmT8mTS5ksP5xS
TCL9abmXmyIf73KinfWVL2K3kkX0DoHIh7irgbAUY+hXj7ji8R7n4Vja091TLqbmncSeqLt+onWT
uxPtdUB2DL7vfFLyUh639kzEKvRdGF2aYSIA1+FB9oZveYNOIS860yspN1+oDNL8H+9IZqCCWNbc
JoNW4iRJW4Qp78wSUm16XIBOuJmGlsQGsqurXodT9C2px09w9CIvYytbSN14un4soFy7wt04KPgE
uBeeG0wuv5F0nRt2/WcAlS3GO7xrdGAsTTNkU1R4S/zJrgWxmXV0MQ+ANHFxoXbRIRse+JBUF3bO
FQu+RHbKLnvznJEWXpYWiXzL8ExzzQWNbdRzDGEJv1NseNTL/KwWRfkZYE4NqBeAAsu/TZn52yWQ
siEQ55r6B8byKcjkxgL7tqpHg45O9wy33XclQNNNdlVbUYY+TnGZtPI2KXW9GolqVYmx+Bz5z6Sk
wzOTnJrasF7A5cuVmMFDEZ0ijL+QETjHvHDDoJ5hC/hJZotG+4n+gizVLTaxDv7VxaoUDvsWlGqO
//duxbp1AMaDbaTNNGV9oYVA1xhgTiKvRDjPitbopsLHzTNntAeBrbOBiiqgK5A2GwyvUj8J6sUl
5a3KQon3L0T+rMD1EFoIPz5Aawy/IDNqzZdqP6i0hx0PFXr0oT/cmFk8A2KLtXeubUA5c/Uzor20
6a1TE1QsWDYvHz1ze+pq5aHWwkBkqJgpMSnzso/pmGVIyboEJ3G1qtwHAjgj68SIocae0EcI1pOR
YrWVHRFhxxjXkTlsOyEQLHx8ArwyGJaKiyWuheaOk3Ep395lv51hdfxaaqgJ2zYUN7tF63BaOti2
YBH749T73LcfydfFAiofvu1Nz8HB4Io6WDO7eTbdmS1VdReN4sgK2ETUwTV6Vipd0bHNuxn9hVtR
BDZwXRvf8d+tWsb1gFUBogFLQvUNdz8sVyJL8UWFBZGNEAdc6qOcvq61iMVvnIhbZj7/hqaK7YBb
de7PBIAdvrJTELJk5ZSQYMs/ELSg9o59c8h6UlFBI/OdjSSm129V99R1cwnt1X1NDx+qVScRZv4w
m+mWuZWkvHydpVkpNSQFmrZ+VBL38nly+eGWdnkTANwHIe4ck459N19+HCt4RXblJ7omIuJp2eOM
t+qYD6inajmrgQ78FAsMqA/jVYTYXZKD8WYDH2nwBqEWAgUZiSv9gy4jceczFDGo3zDQosMzBg0C
r9nPiPmy/XfIdQFufvvTBM2zRlddkHJyK7nb6TE/sjC77uukcfjI3C6Bx3YlDCBazq/RopcMVXcQ
Sg/095Gss2Iak+JTUUy8so6FYiAn53tssnMInzoiFMp2ZEyI5YEGKOS+mxCxuHiQ9D/Q8YuhmJNq
kqAWwkHNyreuKF1Ekvwc9aa7VfJSpE7SrGbGizkI5QzuxCgRcoDUFL4KCT2qkOEq+Gsrs82GBxF5
FtwReJjtWAecthrJT7GtcRYCMhg0ztL8tK1HY5lHLG+Km9xR0FuAA2Los0IVg64lr5YPPQXp2O+E
VxvUA/qfCfC2SmM0eQcVcwrpkMbmfwkp1GTceyZc3Yi1O6KM5kvv+ZFzpxLTdatQFDR34JFQC10w
u0Ouz6IgEbZ1zPy1pRN4V/U7SxyYBeRkG+mYKrxmi6VwJb5k8aRln/b3vkPSB1cz0GalA0a5rSWP
EXANbtS4//0YnmCfuOfj5cJlV5OJhO7KgL1Uw2uI81WnHAs5U31F8rVASjj7lEBnmrxr9qjjimLf
pAoFDqGFfDrMxNti+/DRCiyBDhLWmoiJCBA3U8SZGPED5NnXy+Dw1rjZ2cRa92Oe8c8R8pknmZwP
hitPEqAQzI7rlgNMGjQ5d9mDkP4aaW8AMhiRQXcSAUQ1T9QQbLTxEe0uIehD3DTKud36JM3uB3LD
VQrnX/mtyeipGWyHmNMyMG7vJRnZ9qDbK/4q5PEHJ4QEcCxekkP3/56wkvfkUT9wTZ+PErZ2zKQ0
iSpGSG1wpWnFPbK2lbIUsUk3crC4JkpQrd3KC/g40aro8EE5PbOXLvH4xPsb+i6BIj7oxNDVCkb3
6j2UEK0eCfVTzIegf+DaaCvp8uUIe3kPa7ifoAC5RZaA8bTdR2dMIBWAoLWFnN8ofHy/iLXw4Tvi
O53R13O1NlkQhkUMOgICDLMc86DANg5pKIDn0y61bZVHth4iaRT+uICLjkbpmCVEXRz0mIpUay7U
YusQ/grjIZT52oO/nEzCtuIPXkUFaUAIj33lRQrHeKlaKPK7j/E9ZaG7kggffq6MZXcGlarp7Jgo
Vi3RKpNWVgsbEH1n9pij4wlDZpwFRgL8JNzJ/FVdfPEEnueSr8/rjibxqjQcAZuHs0ldk2i/NhNM
98K3yJE5eaSvLjAO88e95KDyWC25YJhSAaHhGmruqtCvEerQl7+owaWza/zINFTAco3uaFI98oTC
G7wVVYkZ4IwlTiHcPWU030Gqp21+/Cyuhh6lZi3s37B03e/Fyc46KkHGD39ARtp2wfOnpbaeqrwW
3r7uD1N5nLel3nThXAYTlwq3vt+A0YfflFnSGiEduug2nwYyv2GEg/LS47NcYnsufbDTnL99eP78
kMiHypJqAIQ9IofMjGQm9+MQ1WkylJshusS6LGeTy+cpcLhBqpb4ggXB3tYf9vpuMeM4UQYBCRue
GXs2VMLUuR6QqIcY4FMh5lR2xeYD9xA3iEEJ2udNLsxHwFz3JGovbSl6zP4GEpjjQz5wgB9kTtIM
vFERrjr2yEBdf3rjc0wGBu1CuYpZh4GaH6OVPL8eI4S3mqAmZB2AvdjQ8V4ogPgwaVTCbM6uSxjN
cjeoCPHyJhw37Pu5U35mgGa6CNCQm0+jvGSSumv7wYVg+L8+W+gKyQML44HdLFAdKFU0VvJpcE/+
mCFj5KQ9+215KQvocsxjP5VTErut22STnFZiu5uysiIHwqxguWlx9Igg2pl+isr8RzEiO/e4RDAl
n8RzrfK7cN7zbASTf8BU2+uw3XablQJTyf2kF5r3z8W5rqLdihGgkUZ0ZVwy7Gj7+BMFJkIOp4rw
7z/QwaZBS05WDUGnjCitW8nmJhLMuoXuV4zNkJHOdVFRJzZtf+Lz3dkv1MaoIclxfQ5Z6KMwCwbz
4XeB9fJbVmXnHu41uRONaEL/dc9gzLr0RDWqaVmEbxWhXTmPCnK8UcefcKj0uJsHHiUcm69gEXfs
Ky8+XoZl789XwFHkS3pXSZjqcKK3USXPbfg4t2NYfMAnEgzNYOAEOalmWIzJ9snudrw/k7xO31G/
V5Wg+Aw0Au666WqL5Tt+Q94J22FVVhPnP8xcS7xPt0gXvu18aqJaiBlu8Eqc6GtYly9rdWG4DXAA
d5nLCxkY/JZJQ8JP8Ek13ppsGq00AnskwcazebUTwF9tS+uVz5CcQ/AwTyptIwRuCSSHUJx4Kv7h
kjjbQeQjXLDG+DdTqBnrOO5c7My8PTBqTny4UIKA/AXmTn26jCg5Fn9TT5ImhT6WPLWDhn5mT16c
2JDp5hRMFqzJ/TgyVnDFx2ORx76/WTHJ1QymkifzA2/0jVT8D1QeSEfCQ+w0xSJtPhBHfYI5fyR5
9Y+ULTZJ3YVz6jNykNuolGi8YFYnuNbrOp6Lt1bzVYz9APgZlfWvBUOuZqGirW2BLKCS244TkMaQ
LVTAOwWbdPSOHE1dnoqLLzdPmypsZw54XVNyZbTqbeVA5MeZt3gRMZEmZOXrgzFdFZ6A5dhMtfyu
9OuSZwSMbkNyBnE8d84+ChuJWa+mlu2riwmKgiHLdx2fq7qhDYPjjjf+J/+7QbzP1aUkLOSBSQle
g0vXocE0lwGpTmMx2WtZbSW7xR6WavaihOn8kUa40E1LNVcf8OIL8akkaagkwUbEiMsot1Vn4J4p
bWCUwznP++sGzJ7j2ul7XPihzViCTIVHY6fZ3qJycatRB2zP1mKWEGkBTBH0o0HkDNvCeHEXsqd7
K+Z+ILFuoLGs43enzcIuo/O8QlAf09DhaMpIo+SXBBzJCLORzFrXFbZHNv96dOPR3AxFMD41ZdYf
6M56+dYSh0C/hvXJxgewTHvabzaJoOGAeLPy8ZLRCOU1HU2/e0ICzGxoRfYzaGH8utN6sKdjLW1p
Wf2mtwzyeUhoh5vTOYhXW7zmLNLHmj03GfzfDLqiGRAROIhs38jdYRVXAQhdfPp/QiMGFvQCk5bq
MR0F8gDrtVpTeTuYbM4bVtJt6JuWg3ZDBpPZlfvHm/UIdfFgTGRl97S5nkEx6YClcrDHXDX9Mbl9
5sUEsKXVIcj4kfSZEvKcb4A8yh3EJ649hqWvVD80JLU+KeHg88Nav2+bNkm3aEuGoKuDU1w8nscu
RLl77q077eLeSztGlIwlHfLFMwHn4o0ONOL9N6ObYxok/V0ivRtxeyUw5G9Om/NH+XrVNPtcJ6vB
3RCAOUAZk4jfJTqSiIwBJEfF3+rbQZpvdjg407I/9HZSQvwrcAH0gknawNEj1XQi/KoqxdCvx3fo
RXF1TBe6ISIkVZYw/DfqJSs8OWavmdGLcgjVSIFqQxl5jEPppUFpZEOdRtG1qXloO9f+0qksANGm
79Cj5V/SGKRi4CczU+RCF9tqbvL9+KiiDsqwWll5G4ex5wHc4HXJZVgEpcBjFhVciBWz7VvtJSXV
cuEaq+JEexbVWGcPk6G+Q5QoIGP/UNouN4ETh8YwOvOyE7Cl2kBhFs9+MHKTTKDmf3q9ku6UvGqC
5d38zJo6Im7CwsULnWxTC1tp2F1bZWYC8g3Obzvy3K7xh4fDSoaqVE01EFVPX0In+7Q1RRcdS5s6
3EHQvth/+ITmoBHIB1FoCdovcoZYuIR9/2aN5wqniBeS4IbKAzvF8Yj0NhwsOO0XP89UU+lCaEiE
jvDkcw8M+ow5sWAGra+KCGV2oih6OdU0Eb7VMR51Iha0ZRPem+0XE9d2urDm0Y0lO6OSwctUoBK6
ImW9THjAIs1xyetmW2Y06yXEOUMfvoUsKqYhasPVulN0bJQkR0D4ghwW4RarPdgrt9JZjsRxYr3p
HaVTp0rfLHY+9qKZ7z+MJiw7rksJrd/TR6v7n5Cw7yAfEywRRRvUo/MTHE9Ey76nwAFIbrDcYfMy
O84ZAQw4UIJ52smBY643kW5q8RqK8Vd5UTX3a6bJ5kzG2DrhJ1qd6ZwKOzqmaTXHJdzzOAVBPVwg
0LbdV1F9bddWw7oDHwWHU2mGSjM3cBhJHqWDL2l3EPjxWMTciaLrNs+mRR4cn7wfKJPRuAZ0KX3U
sFyfErDzzrK+K9pSIQQwQrW4za2Hfs92vvs+jUErAwhEfpMLaaFqq45/VLossqmkaCnrZWQQs3TL
oqPHGHmkTb7IkuEztGyvzM9+ZuEQqYBYn2VTb/60YccM8zgEc68n5KzTrGxJVHJNY7O6Qr5YtcXE
n0hYOyCSI+7v7u0BIX7IwqcFZO8hEMY3Akb2dZ38idj29e9NYGcHpsroiObbI849EQ4diGrdxy2Y
jZosumDTbp1Gdu8rkyuM5wv1I7wTuOj0ZLdCQ5g8ytxeMpN3vdSPM7zx1bzQ8RAIeIvN/uikwUI6
b5Z3aqV+JAUD0wGF7te4TTFRKF5MbK68lP2n7bV+8IjtTSakOS9Ue7yXita7YaIzykE1rscsH5vO
JGRQl/vgmqt4DF+XBJkGNtEc9V9h7oM+BsLw/maE7apJOBNyS4UGuy09zOKlB2eWaij7IuwWPiFo
f3y/Yu8WmDFGbf6Yu5PHlJce7jJVFlDSZFW60VwTNgfVHbkQboHOQKhNh859zVS1AqYg6Q3SfQMs
miAv8t856MKhmCrfIwk4DC9U4gaXNtT5r1TCtNXNtcoxOfWuMdWbtGVZCntEPCGNtk/CjhDkqtwD
oZ0O0XVaSyJtYdLUgk2QPzjsEb6Z73agx0rzKfDVLV1a2Y88pbwNRZc8jV/O6FTCHYob9mkLDaJN
l2IhbbYYIDTtcSTZ4C6ZKbIGidbnAJagLttvX8abAJqEZKpUm3Xg5wIAJiYk7tcKOBLz/ZKlQYk3
GVjcJjwVIeJrCM4TgxygqfheJgbcdrlVJW6UeN92UoXihyo5vlBpqWM+820QGatKjWZjghXDALqb
8kXT+Nn5n1yV10be9nm6IOYMfjdoEAJfCJTLP0B5s1P+8qj1tJDPUXqnzANNx47FfKeBgqzLhfNo
3svVMCNPW50UqpiCniAadLqK4mmPiPFNROANdlzic/16ZfUwKOPpeNrPv/gon8eQR35OwTNKCSdE
yrXLgC2Nj1dwEdiKMtKhxINSxiZ1lxbKqkm8Krnr6hYOYZ5ClhJSXt7Iq/nucBgRFPOYlHHCAnEV
c0V+CHeLQtJW3e0KmwrJT0K+LpTIQb0JVhGU5alrjEx774cQeWsUNHohcRXicxFNFQnfKhOQ95DS
3eqseWc0wenzjWIHUyM2nzxZSJ0P7IWopazDrLe+qsCm2/XMfQGHCkDiIWerT8aLKZKb5IDQXlDW
OoR2ETj3ZPfsfZ/8xVK9o50G34rW3p1Kcv3V5eIh85qyB9TWamEjaT7x6sA35mhPYkYeNf5zMfYM
bVys2M1qQBaXOYCIT1RqicXWtjLAXY6kuM1/jwy1YHDYT+dQqo14zKJ1FKCOMsZPYIskzkc+GVd4
srz20y8ozTHnz04835SofCkbSJyNx3EKz/1pEVUISU+eE5r+suW9woRbu9zenm/vW2xwjZ4Mu9x7
Ga7BOk5KByNNykf0ZIMU0AwcUorFIDpPlK9gMaALtPGOryR426QJsDG0zMZWovuYdBE6x4zAMKnY
SGq1RN2hIunshd4cfgmBiF7PQbKiBsH6zbj+iYvQLi2mSX6577zuNGeYMZA9NJOMkYydtiljK5Ux
ywTwYaEDO6Fxrhh1aANWputvzY+M1+7Vay7kHhFpJPeLCL9J2npj3Ok4q1SY2rIlRQCWIdNxrZxt
sq+VZAX9RbrRj2m5TCT3sGfjN1BBC4PvGVo1Rv556cHKRQlpI4m0orjxH0KLFoAs4t4vjBYAFtZa
EDGzZ3HK36hhuiUxTaXqj388v3Ny4tDRKmWN3gCQ8tx7LNIda9AwZiqt9v9l+ZKhAeUTdMpt9DN9
b5HZP7pqCmuvWAFtxot/YvGDsfn2et3FKU1Vfnyp8+iCKb4F3XqZNq43ET57/C4hkvdi/S/tg9wf
x6o2vtqN/XbwZo0QVydijVNYMqZq7Z5waY19ooyVvYUdQCEMH14WmNabO1s9WI9v0kFiYi0DIjza
6SXuoT0XkN9a4112U3Tk4A+H4lst02A4vezNFCzwV6xZ2KNQVxp1+vcxb+eIdmxgxC6adg3erEF3
dilwtbge8exbjFuxqy11tFxFXpbv+MxH1WxJ00CqHkoDtemXxo5PQKMtZK5KrKadA7kKfeZ2x/5W
I/Cd+9OFJhHBeVXf2BEwUl4n3mpBRm/tS+KVPf1Fi2hCvhrs9eA8UYhv0/zhBVj5R3xiXcdvYcAs
23Q/H4XEYjQtHW7IDT9jlrZMhA1WgYZziDwIAIJipe55vV+1y/AO14vrJsW/nhJxYnTzK7+PlF19
/5RXXand/Qjdi4OUR89b79x3Zioly2PI7YDG9OVBJbQcy6FDB8/eLbHXrHcNZA2taT+npptv2Scf
0KT8P69gV531yRRcj83t3jo3+euY2bU+KF2bW6HNN2RHNLbC7iXua/MyMarVr2khUWuzL+8ZtnCS
4wLK3hSz0L2bkjBMEaQzUTn2reO/SyXZRhKsvIgOrlXeQtIxB1zUfZwoWZ3hXRX77ZwrSISWXTWU
siXau8lf8xKiV9gmQ8m3bnUweC2R6XUdBTDQJ/URs3qSVHzVuSzrq7/lliywz+gOnxijMKH8H0Qe
HYAJHtDNc+mdFSmEG/CcnwxzsA1QUorKehgWdimbkRNHR4cIkdQVoOBiVNzVjaIcPOkXWj1ysDey
1OgCdD2VOYesxhHo73sPh94ZR09C4A3rNcAXSnJVRNyvYMNoDwcObIhVaa2K5qikwbUHoCGR1PpM
vQv6/Xr3nW2oeJUFT1ACpwKdjDJQkFFAL1TKUxS22Cf5EGZjh0Q75o8jspGUA+lo62gWTaLZlrtS
x+KzIsrs+/z0gauu2XLTzaBKrNOGuHMu68zis56LSeqnfDrr3105E+nqTWpgJEuMwlKdoBUJH4v7
bEPG9wW3zLEZ36FNOX2nDpSliRG+Jxh+ayACSSEDeesz5BmsD/ospYQMQuj5XIBFqf2d2+DL3VtT
/sgiMDPau8+2/Dnqyjx4DCZWfrRj4BBkLdhdi+BNqt+auj/Y4PXYEZDdbOb/vnASNgmuqTHEvv/f
bk0BUgQais07nVv6rYfx8KbvNyn1vyek6bs406OgKWDENjTJ3E1C7y5bRbl+xiyFKLUDnc9NzeTD
FXmLTIBCYwchmstS1UJlWjiXVQ/S5pZGM5d1IX6b/9jvzl44/i47wBg2bA/6nlU5N9FWE9BfH0HB
8EyY6eMA6FmUbYANx2N7bG93xqS+t1MtU7+NNRwdvLaDKI1Ftz9PR2IV1UeQvMTwwBgyEUbn9EQ+
jXYqD8Kt5oiNQSwIX1fjqb9YrEb+XPIRbmkP8dF9FTtMRSjaWKJwalWdALAwcrmCC9HG6euBYOeD
xj6wVzVXN5ZbgWwm1xC2bVWFn9ZWrk1qvmulbYH/yATxC7aI92PaB1kZgdOkhftAiytT9JF9sg23
AMrUkbOfltcgfS6tObFyLIr/Vu0CVPytyJ094QnruRwg/LTj7UAnQwsOA89kZhY9q9csdXgk0/S5
nig+4a+3wvNbTyNu0le4mHhKw7MycR8GlcfWR7diGrzwFRjGyZfNsK2YlHG06mpf73hDQQBEsBan
IezWQYcyNCfhnk65fHO4oNJdGbfbCxaFMP+ZxNFYl1FyXuJQANIFKxd7bWrzwaP56l1PVb9fH4hK
Eh+5SlVGIamQkjxjI6GCqViezYDl7xRkTkBZrrwngirYsALCm5c6zNiuLI7kEMjaXtCsRtJZzONN
wyCKZ17GAnfqhmeaMdVwdrY6JVHK9MgbjXTKuwl/H93s0VjqW7sSS/lT3wI+hcW17WfXDx1eoUaX
/b5MyfrKeAe7Y9JrCApPdxv13+e1Ezu6DxrJfXvbhvHNolPxkXM61wwue82509N+i2DHFfmrvocq
Ubc1/RtPOpSXuXH5cyMn6rZUU+dr8Vtb/0iPX1ffUqcFk8aFwAMbAdg8i7HPK5MAQHnH4tiTHCGJ
6xS7brYoC0wRzcquu9h24IQLPGcoTDoi/fZ75Y2VYNYR2oWfPzVkrUcFWCZyIJJXgpeIOOqCiiUr
WTQYwUo+KpHGzKxSVRokJIPSUubSVzk7n9YrihL99a9iauv9dZBzmPhOCr7U4Cywoh3Cte2zKbxa
OFThpERgeIf8/d6U57iAE0qO5R4+U2evsy1QozgSqO6AE97R1QgPr+p+uOLoc63WfxrdvniMi6Ov
KdWQsdACrNrwG5PszV50vAFhKE6mOEgYZUQw5K0xcJTCADTaLiM62OujS8Nn4BCp8ogPZAjB5HAQ
Qyet1EKvUj1Gk4MGseflzuDlLSaXbaTVupCDLrq/FALHLejvgG4lheb8Eo5xKtXbGzvl+NVBJde/
911qFz+pejTl8hbptmQZncbL8d8FwdVkpMIxC81+Miy5eTMa7cJiu4aQDA/7D6hsYshyN0zlEyxW
XH1PjvlCB+kw4c0sef3FbU1k/o6J+NZDUfO1zxOQdXVTrkITqQ9uNfVXRXkBtsdoxYB4MEMzpCg+
1N4mCUfB8vRlWhklRFybD5lwmgtQ72XyXZ4H82CRcloiE6vffNkl/pCb/Wex1qEzC+gt3k7gxkl0
RYmQ0vczFWDeCzTmqRceQq5LC/cUN9TVY9BOcnG+loL3WV+Lq2diGb+2XZo+sYwx7OLAKnXWDyQC
XgxQSVYgIOJcmfQze9yzZ9Wc8xlTpNA7VlabYFtm7YFjzRTa3YQBzFFyE9Kqryn64cZ6B4c5kvdn
KMY+N2dHuxB9mNmTVFS3kH2Pmo7ngVlVyimYiNTDxCzD8tgrxW/+jN4Z6P5P4ZZ9DB5GPt/L6T5j
l4Rqvw7uUoC+TYXSJdOOrQOkQJ+PxD+2at0glpPLL/IobQuratYRaRYRdD9JJXiuuPGG/UQstllW
iG+dGJ6vxk53fBSzBOPLhc4mVswv2vca1W+BAaazjm+AGUlLK15Gm3aHbzfJmbQyMXXrlUMn9ji3
9C8R9eMK6AkEAGBylQ6nP3JN2Gpa5o75vJPG9fuDj6aSwnZ/xrPnNvGIiTiTD+fyneIL9mmEb1hG
LjXTpPvVh53PP31Thva8ds8WTrOmU+XnmOa3skNrD4QNilosCWvqvzAkcfiIa8JGAa2vu4H5FH/Z
8E47n+plg+GA5uvXt1IScmOnxpBpceM3X4M8kknwocKlKvUVuhDJWQY0FNGyPU2CkJxIBgoCcyl2
Lu11V/sOQlViR0wRdBGQSnKtW92Ibji64bVb7NwDK7YHUKITwAGcJF6zlr1Txau3fok2UKPSaUvf
WHUcztq3t6G7pUD79Hhea1RlzXwYzLYjG/452pf54oUyWWFW7x8Fy40JNFE/c4BbDCDzfnTeDzS9
rqobCm55a5jGnNTjC4j9DEpBPXq4+icyZFUnv/OKUANWbbxQgXevzxfjyReCWioY2CaZ6L7fEkFe
y7tPMHDajNY7U1ASd0wwLTWf91VRU4JguNICl0Y6o0z9LmTVjaPv8th654f7nmP8oTY992oWZW7u
A4xPYxDZp5WHg5zK807odJEzOJ317aKr3qvCs4QbNDEzpFpApE/iCAH1yn+NsytZBpPTtu8URdnW
LFkIE4pwLYBjUT9/JRLemqRrmume4w7dj5Gk46BpJYSqtdIuFo7T6Zpoy+mSbvb7mhHvFALQPz9O
GvrHW4qLu3V0Xux/3tupDbLTW4Fh0fWIvKtiGc1NO0Aqt33TjI1NmXjUmcuAjQAHKf9sHkRPlqnx
ZVKYmPDpEp/Lel3k/Igl6q7S9pZE37ZYXqnctQYyZT7oIlDKExXjRf0XllBl4XyH/1EvnXccKsop
ZJZzzqXYpWAEsR1BDVvT3AnMiWxgm2/i28gEf6b0lZ2aJ0TpcCGOfpibs1VAoYBLu53QAQNjp3CG
q2rkJVavGsq8PF2jksX7LHwZGOTWMLjG1NzaXZYZbNGXe/RuFbj9ILQgQaMVUPP7vdUmL8npydWJ
7dM9LFHa+X5lnmGAjg9UHFyPAsJp5n2mV06aRS/dEcTVP/fiIY79820qcE8DfGw70J1rfDDJmhNX
MTXUGrw/r95rM0c+9vGMxMXpq+p89579zjgR2uaLWvKbvHrJSPBxWcDxI2u4madW1/k1IPcz0h7J
FOW0RhRKWp9Px+aBv0o+BL09Fb5JYLbxaoiY0Wk7ah4YNkXtJu0aG5YEZ6AGN6HyyeRhyBJUHeE1
aLcFsMGSn8ZMJnkvin5vydo9jopQ0Ek5NMGjanr9fmM0BK3zfgWvhRaWyUSx4HJG2jMhjXEpiPWO
wjalQgjpzcwKkoiXGuCQvChmiaD9etlsoiNeHyCxAUADIiV8UlOo0//gxaBCsVey9DJXJjl70NRf
ach1LpSXCbv8fusYgfJVEBJmkPyuTN1IMRp39hGIuGCFmIY2Y4zA6SFhTwfckhRRZ3dcFuzJIy42
DDIJgaVmElaTYmEGDT5AYaFa7bxR3LEalKZhmYJwHC5Kltu21U7Sk+7n6AGpX4hWC7nOsZw6QbrX
W5urbXlw8mr9gsVWzvBYtYlsmsevEYtEBbSDH7IF0kFfT6PZi0lQbROUTgRQ4QU2DHPaKp9//yz+
1F94CVSCTCwJhRLfZ6b1UhDyUqD4Yj5ybayOabFZB3rV5bQbK4g03a4OOZGMVfkEIDewdOC/lYLa
sRen4p6jVIzWBG9ECcFPyz6fxJYg9yJe7z5mTZLsNKCsL0mdjO7xoRM0B3HsBnsliluqYXGNYG73
Cl8orL7ddL0IiBKZCr3gqMDLuhrjqN1qdKOHX7Is0WxIUKIuHtXI1+8q/kXQMU8f3fWQQaFyhW6q
43c251vo9r8zz8Fxo3tF4DI3h3a+bQPY9M56XiLXl6CyD4JmHEoUGK8EvxDemRhto7MX/8uIJsI4
gXwXXKAsrJQGwYer636qm6eORLte3b/foDt/N2OSoEtF02HYnpBsEqj6QXP2ciyvuU0hmWnuTpLK
SQcLLqgb0k0joMZXZBDXrLfyAL80oemt4tQWRt3aCQ5hMI+dRt+HNVSocGdEu9k9fKVNTSzQLYlW
kSezmYOHBKghK+QJfbrsz7AArDEUwxTS2tQRjkBxc9Fj+kJ6g+DeMhmRgC24+ak/NIhsoCA+YrWd
tDqCJOSkq7wBCasFMpOB7BVXlBHBb+lCyQkBwf8w/z6PuJhbV7PLVJB1+0Hm1cw1Fk9zQAM1xSWC
C8LZkHJEpT3XqDPnnCZj/X8evt10nOhShvNdoBOuXiZVR9Cku9aXkGrNPEgxo5q+bioLl7U9lRjm
66zwBHF4qJmBRraZ7ebZ0dCqYsYdG1RC4Fm+IdCBoFb5XAapDvjr5AhoH+W+TzIFjOXaRelrSBI1
bdUniyhWS5ZFaDz9esRN8JryrXAPt75CpNaAv1677Wvdxqs9PmMoAWGrYYDmYjHjkhaMVCFaWSbC
zhCxZsGUzt87SEjCge5U5mzy0fyopnfrL6CCHePrvc5SfnPh23JWtD2PUufrl6qLHjvnZfxfmxvp
ICyy/jQGxJ8PD4w7ZNRPBaRHOAx+h8Zfgha+gs8TdL/WX9DiplJuirzvw+PysZcjpMnSLStTK6JA
um8VVWkfy7xb1coN05i0qdZLAftHFFUdim/NZZR/4B3A1iiuV5ivaFjH40Qc9kcpMVsqh2vQe2Bi
AVH9Wrq4MpdQ2yY9HlNtYwSonshItbT4BGV9ipq1Q9EIBgWJWumf35md9AdZ/94ZVSccT94wG3qF
yMHmlGTuGLwPjoTSk7kw1g5i4HdESt+HEHEBWTTshOURY5HGFFlGMr4z3lH3gQfwpIZ2J12srPkG
BpsBG4QRen2O70e14BZ82+DNJrTn9XS3gmme2n3U+5G6mtPZb6hpR4lqjowUIXIqDgGVAH28EQ/S
/DNJsmIBRouzBp9kFAwg7JVstFrFQz2XEzSXChSwbN512W5LUAr/rZ8AoTRbcQOQE1durV4W75uo
uwdCpU//FapP7v5YrFz7NWHkilO1pZ9eBd4k0Dsd8je/WBLflm8SFD5MoH0GtGHVdY+z/fvTPlem
r2jkR3XZbiT43lw2+v4L+bfS2uZB7R8D638s7EYr89tStidHG5k8v3fJ0Ws2shmAi20Bz4Q3NV93
cWM3K6oU6TinXo+dz0cwBbZUfWo70brhFMS6ginpMIkjnJteXvVtJ9Fehz4pAuDkK+cfcDpz890H
1Yot1LwUJ1olP2O3L+Ti3nuj2jTUd7psTml2UzvZRYFZGuR9E3I2MiNK1Wnzr7hd5oKYl4ZgY09r
OB5Qv5mWKX6RqXizm2Hp+junqVfUcHWTfN3svqEUP6bcHrgJq62zm4aZL/bhbguoox8sTFtRSEsn
YZ5SgXFH6FthlHLunPUEj+/D8CtCLlr6mvohNT7P65X20mGJXtxY+2TE0OIO+yoHGKDLZWAp6Ta8
1dEUzKpsrGab57EZIq141WtpcmZ9RaqpNP+2SmeHlXatpCvSrtS/EicjKklsteBCDLdmYRK81jLD
JHugVo5cGgE1E+g6//di4Kf9oVHC7YVJhAGLHOAzvBlq9oP5HuuUPEqhGYvEbyR3H/yq8t5LD6ol
SNmtdjeYMIJkgtbXXdKDJn5L1CcfxH54/EZqZZopq7IVAFwV1eCv3bUS4M1nZnTn/i5mrp5wkjIv
W6IAKRqFpg1xfN/DAB67m+0x4CmhU+Ip/q2mTAwHzvhI5A7d+0MdYENpeisFSEQ5XUV/BKEoLJaE
dLQVHmWqBKbix1FHNBdGnYVlBf+8WX8rZYaJ9Dpt9sfamtnK+lwXqI58VL4tbe5Jzsa6uEi9fxFh
EJDp9gYJlJ1OZ14BTLZrPWamZaXcb8+i6j4kzQLNkUI8FdPGVO7Up1+BxS3QYohJG8ywccW+2Uxs
Mgo4sSqMegMh0uWYyj3UjUqUmsytDLB2Putc2ajy3Dii0maJajj2JviOOH8QImOZ50ANTwUpM25B
oP0LGpL8DGAH2y6gtemfqTAuvUN/5SJwnremNUJaU/LYCbCVZc82zqJ0QQN64wcTseFbj44P9SRG
mwPcJTfCLrnZovihzZtM3gMSFWFAWAWFoyKfYuQ9G0FfHPwPS5mgo6zrXToYp4z137VTwHAcmCcp
g4j9/mRlN1SaZUWhrJy4EGtlbHqfW+KuAIsiIBtjQBq9Y2RmP3ifhBsOpUh8PHEOyb/90xFjOIuf
0mnCGpf6TFt2C/+nEgQsOfGYqp5XqeiRsmo1mEFobGY8Kkkftu9cANYMej9yFw/HajHL28Xutt8T
vY7AJkRxbKeDAVn6UVJv+McS79COUVurgYD730WDAMuQQ9gWHd2MQrLcyUGOwTz4nIyWAPWX4abm
X0bAgPL2KslRixe6ERPQm2sFzTcuHBsf5iwnViiUQ/XaJSPZgrpeb1SnVSaIDBF2UZqgfaAP2n7X
lnUSP+b798U2uBKzZU6pBtJjNXPMl5l5oqE6/iozNX/f1fwnR/lRIh1isXuHcmsxt4//Vv4blvsa
Cb/8YFAoOpd0cRB5sj78/GkRMHD4llrjPNrS3MUi3U0Jf1Qx/bFtlJySuu77Zw/ljjhRekTzYxMQ
vNZmQ//XmCHJf7F+OnpQa3jewfWElUKuG2BGajW+grQLHDcRhr2wkL0DjDi7m11CES+oFYGraeRU
ryFhAjR9FHfK1F5k5MhptP5L9v4jxWqvxjGOxMFjco8JTuOM5W0NSfST+wpW9ZrvxxSfdQqc36Dy
6z6S7RVheKl1cw7GZ8bVrvnfSrGnhH06UMWfsS6GJM25FQ5FK2tSOE8zyink5l+p0obzSERq8lyS
Vz5LMdCplY/J9FclzIOMcB5TMp3gBRzGvP8pSVAscxTUG5za09se8eGtvbWPZw0avQTORhCqt5eo
806v466VfYqpnrheH8C/tPa4POqRF8Ifn6vRu92oyAW1BTjVKDo9OBRWQDPWYcy5wbMNEqIX97sz
UEQGs8mAaExuRGP2fm7yRV67J/w03OZNqzkyDw3VILC+EePKQtpZvpUKJrtbWWqIO1hLpBfBIVOI
SLavppgAoD/KqllDDvbb3X9FkgBAQ58RqZlU4WRYXsLtkg1YehEk07yDojP6vwQ17reiOBwXfukR
w351/qQwMSeZB9K+ukxUkICFeANgWP3OAGqztXRaTFloNs0Jx9L9hcDyIWTQyYf7fu/FNNQE01dv
5+7ZBmmeRmwoQnVHb0FWLKqpCtr9UZHJNuca11wscyEl3LGedj2Sg+h3SzTUPXMlN8kHp07Q8Ow6
BletbZb8VFz9xQ6yxyR0rqSvAPyhzymlK/GgdEuUESAiesCx8qAWCrvm/R+Sqsx2QdJKCwN8Z0jG
QEZmp5cCwadwOnuLsRoNDiITifEzqEBHTOwVYZT0mvc27k96+5jwTjBNBBCSiz+uARgFwf0k1ysB
uzY33MY8MMBtSQWoEqbeZJ+zZujIIsc2Zt1LCc3EfJUN9w2cOc7VsLMR2A0ni4T++mvxFDWg/60g
6It0JnAOptHYqDGdradw0hLD9mDM/3He5nFVxDqSbxIAmijflDBIsi90SPv2J9Dxy3wSKCmoVyZ8
cDH69pxYKJT7Xv+tIzqz/6B5LglzhV7dFL3GsyuXLO+as+Pd10HNdkE1+tR3FuIK1Jr3dcI/ivdK
rCTjf7bzWXumYqBgNOlhfvIaw/VXJ1NpVoDSoGCEo3eB5MMD6jjVWuKfhlBLC+hiOT+BKwZBnZSY
SwooyKcv8ReRnWGxqo57532RfQH6vn3F1pIbWWSXDRfZPHDoz6LadglVOKE4Pz2L7j1H1zpEmwYz
D94MFZ5e0fujxnXqlSXcsquLKCNKRH7inXUII3sezoCsksClqOttW0518G0tZrsi/7/Hu31iHBfT
zu1cqIw81t9hDY22ZOVJW0fMpqMIOwd1HMBFETHr7KiejgL4sKJGpUWuC/12S1BXOs7QX+5mS3A0
qSfENhFF6FbvUV6woK/97875ykL5vbY8PYBz/UkRmX1oQhJ/jt+H663bfZ07bGB1pLdFzfJkItj6
uz7L2MbFnnv8I0o+9vRC8J1GkusQjRb3hU66vT8PAKsz2z/RXFsvEYdsVdDRTSNVhcpfC9kD/qZM
jKqfQk+5oqaLmgXsdo9MYer1u0173Se/eFJnDRRzUbi3fteuvGnKmQwTSHJe6Ju/oOnRN1csmEJO
Doj96/2bphuJi5UnMUWk5KpsPP/5vYOLGe9oPGQr2HWE5a7YI0NZxB4KdiwlHwEtRou3w0mMAdXR
Fc9IUnIh8SuZYuZEd9OH416OIZEBUac7GcETIe2nOyJ8Vh7yqc4GxYMt3pkCFA1jisFagqX1/+0s
wvlcFcyJ45hyfQtB4CNNQgynYTT/8Mv764Ymu6LfeE448T2JmDpbAkTbdCPIdDXrvA4/KoOrK1ck
ZDklb1smryHz8eGNs6j5+y1y+QPan35weum5UiKYi2DBKnF0aUZ6F/nYz78z2jB2SczgDnORYOYW
lGb+Aa2jo6Nui7paZPyUajvpxl2n/T/PoCA2DJJ4oXjgNg2vdAAtFkWfF/xU1r9P63YCgFfqjnpH
Mui0r0/cgjpBHWWM5N6aL0AOVy4j02rOi2D89+2d8bsKqp/86EQ42cCjbntNYW5ytybkP3kqnUJN
QVEjJxRIOpjPxTJ7PFNqkO52M1M073OO8cVrrPC+tzFaUcyZ+HjEY/V7H6zmcpfYn1IIxq8YZeb0
sc2Zi0iJDOHsPVhKds8yFs0Lfa8MeqB/WqPcl1b+L1ceyYq13C7Qu/CKsKzBntcHQP5Z5gKs4Yfc
QBVpkSH5fYgS/myqlcNjgqkavaRMBcfhwGcmbHS30VJeUstOlZuyxIkgAdppAv+s/X3tH6c9mx6h
KvHqjoH4nE7AmpgExd2btGkwZVbTgJgGnvdRiE1FT0WWjZ4ypUURjP+tieG7QCY9mUSWxATmjANi
lgjLcayAx77dXDLLmfhZTDlpIDCs0uWBVUYTgD0x5w8njPk+H9kwZObOJF2ho/N8ZOEsyMAzTTRo
65F8uMHqEAqwNkJ+xUDT6w8T4gGpakvGDcKVnpAsqrsvc/wyWJFdgaTERbhfWr0K7ql7PO5sEZ6/
0ier/AA7d/kJIj72wo3uHEiqFzT5PDlZrT2Y7R8eAo7qSjm+mwjR3O4mXp4M3ROSEJzNuekgdCYk
mdsketnTFUOeGvzoiS2c9QdaDKlR3ipDHQgEnjAhHtp5sUXP/u2KvJtCNNv87Z1aRdl7INsofo0C
0V5GiscAW6drGMx4zELXlmoCe7iIloId7GnmRmc381lokpyxML5NUyNOYscDIbb4K+5FLfdTdjQ9
ZmoL2ioVn7rguOx+hGOEtOf+gob1Cecyx09ygu5lvV/156EDpq97cwFn8VYslMIby6GAuIP5qMBV
pX9PSj2bica7AHqkqcmAbaDTMlAYguPxFhacQn6NZx9A94qOQCoSadFlAzu32GrYW1sVnZsoye38
7YrPsYr0uRYJ1t26mYEaHPR2YLyGNdc00FJSlj5t93s/OLiF4hGxijjokJDszVIawLdTmNx2aTii
iblZEp0WzQZYK6RatzwbWpY2fBw9fdSFFyO23Nha0n2jljPHQO/TNLpTeZZYCXADuPoyzpxwcA6e
slQ2bWqJUqLgi5nVjXUN+9Qn9duoWUnvq3vknWdzkloFzi+LCC63PCFTIOQdgPVYpcrI/yr7WJHI
OTJnVs4eJu9TIoBUsZwckAKyiTvRASFLiEkOa7hD0TKZqbW47pDM4BvkyENsJm+ntuOmcA/iUaw1
EL/79Vf4w9LMPaI9fUr9845d1bCHnBv5olxZ0lStrqdHRuV8mus4qArGXZ3dBQ3R9LxCD5wddUoR
id6RD9UBCA9Elyuq/voHvyVZ5NHQNFmJ2BRab4jGNMTxJRrp+gCKyAgXGA0/kxgMSX9VYyGOEpkZ
b3sJ2UWGDUTu0c4A97wqdz5EOJPJHdqjGTeRgmtM/n3fSGEdONjEscy03pOFK6lk2N5Xw/BCIufm
4eXzLGsi2NXzNgv3mCTVDobRvHG60Qd08vOPbGKJIpwy+kliP+olOBCmsdrAPvlgK7tmoFgh7ZWX
DK7NXnYIGM3h0si+gATOK5RzHs4pGXrBfJliyPADGAdOJAGGJ7AUzdBYT1GfLOllbbRkfHi5ebgS
v947cPtbXYvXUUCm8Yc3ZhA7pWL9R1f5SJ0sAuLl2FKo7CcYD8CLONsvTkcZqvdyCnn11cQpZzY6
2yT6lf4u4eUK9kHWPQyAtn5PQSQiqL3gqv4GoyHRxsf/jdkvGfy2ZGSu38Ykd5vLLuS2Vck/Azvy
XVvYMlSr1Wz5B3zjoPiv7rrDSfpBN1f7lluJNGMuWCeSeuQ9JpFi8KKmopHFPMUqKSjlQoXbJHtH
FlZvubJPLNW4sV0CN/W8lVVYSmT3Hpdx8kcemH0NfND338RbWEN5Hx3HOCA3oWPV+fNKL9Q2J74e
Hy7VGTyIPD5aiBbJBnj+gpS/FiApK2d5xbd56jfIHNEq/Xui6V8zeKvWpxXM6T6GtGtx3E1NufLz
U5SOv5+6XADPPowWZo3+hS69rDKKzrtKs8SzOG5TvZB5w+cVW4soyly2QEUat9WxL7DBoLbd8dMa
nXaaQT6qNfjANfy3aCcM0CnzKZ10XqbiMTOTb+jpY8LwJvzyE1M3Aal/TDq/FgDUBdwPpBzbNDO4
ckXb9b2PrsoVC4Y8xA5qmXh4HosSmr7PimrjusFM1Ubfc7jj5s8iYoLUJDS5CODBwzjXkK9lgcHK
d0uc0GsARM8I12yIXbXLaS2S/742npIs7WpX9xdJD+8LOWyAYhHJFUF+dkJxy8pGOUj4g4/Zuw64
CcVdjCS098Ijw34L6u4kNn+98GCcYR7e4AHxazn0TOFHyf1/aLHI6Lk4Y+MtOzngTuNzNx1f1w5p
V1pe++kxaEWm8nSze3NMeCNAYXknT6gwkynLL0SDemV5Ze5qBJXAkDhShgWQi3+XgIEp9zzKXzRX
xesbsGobnVSbdnqqPBOrdMlwAyNkF1fm4K52CCwG7tQtz0CfTKQWxxS5GeJfeXRCnpKzGHziMJpW
9728b7kUncbAN8m0xCroaeq05qkZXP3BQtGyeJapKuZdTAb9ySD0JJuWt1O6NpAd6V2l0C5Zwo84
SBsgDtJLz+/imi+XTe+/3JRv6N6Pi7aFyyVi/bKyHVRl5dhZiDpCkTEzl/om/CRUL+LA+oFYRLZq
ibiBbKlKsFkFZqwLNF7czfVaVFiuBDtohUaJ+HXzMWL8H/DNCZJBCOzKbVNaT6/Alx6K4XPcRZDS
9i+X3nvJgaCw8aKGv5b6dwxO3efB9xGqCfvCL+hbSHWdn5PcLsnouzfEFS9+CChws+cAmeTL15As
Ymxcc5kV/bA/YGP8OxVPpvhLWSYyz7Fq3SJ4Cn1NkSZ+t9HuKNEu8STt2BWrq7Bdbk0vZJ5+czNh
E3JvMLFAksMkys6eZ9dy6ylc/nIkiXmxDPO3UPkxEHMdjxybRMx8zLgBTrEHtstmA8HfmoyeM2/A
GmIiA7+xqvrJfPOUbND7Tf6sG53STWzS5wGm2jUjfqG7cQzxmCabty853+Ot0DnAx7JsiVbDsVTj
lNzLqI4MJc6f+3yqrWqsXUpKhB8/4yG8Zm262pjslTiHveqclqu+Bhc6L0GRo8QDUobuslm/9iqM
/1TUPHhccN0vrU8OiK0ZL0yTcj2knIeSFmgsqqs7LSB4A6yQpvM5bQVOdbBLQaBcjGqyMKF9g7Vq
CIfSEgvRzVTX0ER5KzUqpTBdS7Iw+HeUPIeumHOTgmqNeeRzZ2eY6uKjbX3CUsPQfo6hUVusC1VT
88SeZJeGQxzw/SzYlcfEeP+DaEQRd9c+pdQc5QSGRlztGO1IEDde25CFu3HUy3PnOxTSDoMHU4pq
N3KCe8ZVDhWVWCfykiv9Syf4OOFc4lljN0Eq5HUo+ELKruk2Zhvp0iu/d9eib25HiGhoe9TuHW4W
N2H63QfG2crFOeC71PtDuGFoNUUGQkumXTNCqDj2n6GVZKgDTT6DTJDVN7pYE8bM3fHX+v+qdSGW
SMqYRA9lNb+Ojagu1CrfvkDtEjgcBiBH8wjRGivt7i8qY4H26XF/BWWOEFfWm7Kuukpva+VhNLhD
ntP/IqR5uhnThmQJHjujWUwFK3WtxNYmqLORXKcvVpTJ0HTq6kD1mB+XWwWN9zuL50g0s3w1Jsxo
El5U3FF3K91qxlH6xAef17M7gohiW9GgoTNKIZLcsVssYEAlZvLA/8PjWK13ITa0S27jtU1ygi1U
Dt4QJ2Q0GM8UZy/NevB8EG0rm8sb65CfKqMaCYCQdMsM+fSVKVlikgsixBBzhfx0lt14bRqYNmoT
tw/cDH0QFQ6GuBn/lmFtomN+SUFlnBlpfYZpp6ujcLsD21zvA2tOEi+cdEGblHw1zr2jwKoS6qOa
Ze2+bWD5kV3rRJjV/bKSvMNHTxxX5enqOUWRTNpeFiPPPXk59hoppALTnf04O2q9WNAHNC5vSdP9
AUrp36Cyi/OfNX+SQUrT4a2fYQEZIIg7fBp1fwRzLDVhVLlOHTm0NEn9rKlRMnpqXv12Uz+grnA1
VqXcY4VkZEozaBoxWChEGZ+lEYTEnW6J+zOk5roxXRIrVonPDVmns5573O9ZiaBj4DeFx4x5YJBb
94aivTcOizNnyNvnINrUOx/teGztbFBALHEncE5jRCgrtyaB6Qw58fmXBDJHLehYUqIdiobpl7Cl
tfbKtGXuPv1PiBWU/l60vQGXwAPW3qFSC1UasqAQL5cFNCjhbe2Oeod86v1cAaaBcs6S4maT1A2d
kHu3nB6ScreT2pl2twv3LJ6GJusPl/NZpGC7FO1SE4/OfCDsMZqZU1aLJVRr1JNHxc/zf5uB90ub
sJRcvTUP1ffKjjbCLpmRHh4nGMKDwlOoZOSvHZFRKMzvyg+7K3hVtOIy3m+jJ2E1GOi6mN/EQ1p4
KAak9eqjyVuvc7F4sPrz86O10Zf0q8rXEpiYip7/sSAtfbX5vD5CG1B5qraMn7RyoyM9fH3BaJJA
fL1RJiYVpDkRv63f+uGhMEszKQNUoTym7J1FDFqQpihbT0oJrW6LU44oFYT7Oq2vBW0P0z2pADo4
SSrN85xSYPkY94aSNQgtMKd1sPFvGX1hYz/mjSQmRfxeOIRzy72nlv1cTCHNb4cCkziv0ZlN1FDK
aK//t7ELL18IiRskRfApp8WFBLMNDpvl/6iqvZADnKKJnnMhC0YWc/oAOnwHNSr2K3U4fuIk3UsN
ZbnYEfQCtr1St4PMohLMfebimOKMoNIAOfQEVH+UpaYDxb9TXX44jFeD3NpmsksQ4vLDTpx/pbor
uLEPZdvGfHm0Z23IxkvwIdh76+T+AICErOMONQq5koQAPHQ1O/LqIoDbGn8D3ZlRcVYuiifNrSJx
QQ9ix04LRuoTWffmrEbw1ptz1mvKoPbWfw+33LN4Eq6pJdwgZuBKzSP9aCtyyhrJXec/Y0GJnx+a
kifWF86ZFR8gdJ5TgxnhnYuSy5mWCX76Faw6oIth8Uc/1X3AZoF9LJFghGapW84bMQcfQEEx4LeW
qDLUm4KNHyZvJTyXuQpBQ19qIQLt+GJYRv7zZceB0JH8k+kCEDN/QD9iaA0WHXKH9OgJIr+UQIuB
oQ2KDhrL0e8IPA6MOyPpukjRK4ptmzzoworCgKIS49dhEyDW9sYMUSksiKjoC3ujno8K1vYD4pN1
8DB5JgOvNMDYZsl+i0uzyJ3wQ4232P8VV1UgQl6/ijWwYhbcZT8iw10AdLpEyOGA0cEGJ2zkAyto
xS4B5tDykEKxcNRj7yZsFcT7+JwNoaosu6OXNJZnXvWzKNHComo3hqKDhSqQ/mzb6i/FLv6/6YkW
g5CdShvL/XdC7ZFrF2gjsLsYA5mNx5Gp1KJo10H0c0N/BwGIsAwJmgSP+qYWUoHQ/HWu5GOdDPeM
8rrXJDKV1Dg23TbAcEBpqiL1VUNosAeghIrQTjFcwXWSe2AIHfzCfPcoLKlmWEp30QhOo222sGrI
WuP1RKxu1qWXeQxLlncr9pwpPmmtMBT95pbWfef07E/ESdYBj6mxP8xH+g/1lMd77u/xTR26p2SE
QpqObf7UWEtb6/ArWtdm++PyYPdZfe/GKe/VdeiWBzej+wi8zts+12V8ZepFkTGIZ2LY1XSEW2zN
w/7TXeRCHngDjAjKZmxAuN9qoyPiJ21jYcVQrIPlcEWFIrZuAFPEN6FXpmM00w4+UcBb2I/vhjod
MVfcznLYiGjK53pmk76f28QLI85wfWAm6LCqhmOLCKz+EWitmyo17g6YriwIPuvfHXfzhT7haXKv
w2+ADlKFwk3jg9a4xdGkYBfpfLHW3BdLuHtIWkPB7t97bxcV1HcCTR+x10TFViACJqM5IxtJEXm4
52iwO1pc4TOmUxTZpObu7upxecrbDaPI7NgoFD1vs1B4MQfKdXRsqDOGkjni3KFR7w75QbKfykE2
JuIsjXCNZyQOCjy9SmdpgyPbTzLZ9+Th+OzHWhz+vRsadXKsijDjjlwiMEcfLOXdyB82NN7hoWnb
pp7pYvUVGLvHlExQsFgUYaV105xeOG4avxZokih2Dd4jwZQNHjsYz4rTJu9quNEmX+fqdxcS8poB
ZmkVrjrEM2qASJCgoTnRdIrK/kV+egqXLPxlmaC/LkDO7PMK3tWc34OOzm4OB5t7McfLUPs+Fqzb
+S7Owi9lQ1BXynmRDgkBWXOeTQggJCqcpNHZPmMVhAPcaim/Zt5H37HJBN6OW8ISk+wakZBKr0yG
VMksyLAGlIgIpIqqBYngLfILxn9SunyJ31y43uli+uiB6sbMGiF6jkV8G1SrzpVVMsOoutWljtXa
+JHFmatuoH3c8HPn3lhH/ltgerz2/wJWNa7j48KaMafv5rimM1Auhcy63ZZgXjnwnvTbDXCM72lD
tNcaO81APRAe8QPe7dnEmwzg21kiQGVJww2gbSVtpguOTK1UUuN6pSFJHO6ALaNwv2OixutR/38a
9ls5IADBIrAHy0L5OLxzFWXBpaLFDsyImqXYLgqRoggeZ2uPwhKlqZZ7MB1LcNF4eA+mMm+mj0UW
Qh6KuZIXcly0nPbrSU6csUGyvvYQK2uXYXM98DaT2pByg28l7m+FB/D4lhG5LNoxQIeXLXs4rzM6
Idzqa8TxGhaYtEPu7N7+HobQJu8IlFtfL+q0wWEQr/+jMgQJd8CmE+Zba//02SvZq9n2d4knMAR0
yOqzj/yRVbQ/zw2L5hPb4SAKH7xM34Ocjsqtt3EGJDADiBKRa4YgZQ8r3QYzvrl3XoNwu2m7ApnH
37+4sqOzT85/JV+Lt+an0itPesu9k6tbAH6vSmkwBSc/VCR6BJ+RFjq/Mq59Cr6OI3zJqE2JoNh8
K39cJskP8rpxqzpb30HeCk8lr9BTcSAfQFUzNzM2MjQItfT5SMawcMnq9UwojI0FCaMBDMiX+3Nk
ydGLruF3qZcPBBKgjhi8dGfCNTc8xQQZXdyjp59tc00/otdLbB3MqM/9Y/2dkn0idzr7f91gus16
l0VBwbEJj9NAza5iFkR+EXTQWXFmgMULlS8BWh/Cswe2lsyXPW2tfNRJp5kur6N9nriQlFWp6Rc/
gr1Cw4+1zJ9K7OpggLuPGAyWOFLYXFCjXqKaCNHStHo1/HbJDMU2IBDr8MrXvre4SUb57nCpBiNk
86ARQqR5t9CZH/kl2LERr+Uv2szswKaOFrosI6IkxaMNNSP61XFr2S2WojnfGfl0fdfr/KBeFYuY
6WrI2ENP73NLJp9WwtNbPoNlCbVXoAUb7WPZ+6lOxwMSszbYf9DFMyIhP0OuboOInhrBHVHWZZLH
V4mrOwbuKez7Igcm7/6QGGt26OO+sTNpoDC2/A8dM5IMyOPKCUzsO2rU4O30bZRt5qZqS3ghUk0c
Hkuufl067ePSFIQk9Xg3m0ykkOFU0o/NKY7GH87VKQ0g+zqufwoMDtqGMQYuPUB+5fTpndtlmOlO
ZCTgGVZPft7uw/KAoCv3VB72A2p2nk8kF0yVBWRCJ1KeHv9PE9wRlNCecn0GhPxHjUue3D7f2Xw9
990Gncj+POcw3UvK04r9O+bxsCKmnmvbhOHAzFaMO3z3GXFUX0asTi7nP73TeLLk5iHT4xLqW2ra
M4CXw6k/+V2tWdTMYdG88lC1LrPbMcKeSAkO4C5PBdJPPawCXm+v2DHeZrK7/CC2aCj1FTZ3Lj8U
hHOGdxUnm7A/+kNzsAvERYoP+dtAm58jftbwQTI3HSJBBj45eHXtKX5NpFFDqtLwNBP1hsu8IEbG
m12pz/BZk4haURaQMvdtPjfA5o5RDGO6J2+HWdFbDMpIE/4qKg+D5+M7+fxiV0Ura2xX6wqz9sr8
TAwyiFFAV7m+jQnxqP0pGu6My0+XzbHL1kTy+tBOCeuOigj04giEnf2EWsMgcCOAeeyu9PGr0kRj
yXnurmZLYDl1TjItHLPX2x/35+8QTX+gE+DaLLiNG0bvinFlfr/rKAUMmcsKpZiQUBEZ9JiDlhOp
IQeSF+NuuLa/mM4vOiOhx2Vb6wXPUxQqFm9syWkQ9/JBkPz/1rV5clSRSd1jCGkOAlHffeSZpAnl
84YQnDi5pLw8MwU37ODHKJP1+ANG1kEvJGSvPqKKJBO/fqEapkJe4OFtXeMWNF73lpx/7ioz3lxo
KMtPO6vKNN1pN2jQRjp/1r9OVphsKMAtsiDNmg3LipjzEoO7ZP6JI3of26OkenbLQgCXD0R6pTNR
ALN9v0CaRJmB7XnW3oLeqWo1GmeJ3PgElfA0JYoh6Wuvf7/o/enIB4BIjCrNNISY4XreS8NzgYnN
+9han91hvdHQddsJEckE72leq5JQDOudX94H954vDc0ENL3XWBtxgBnaM1Nsl7tWxxlWAtyfML48
LhbcnGKoJZwCTIfbnH6YGLZZ8jZCji5CmwkPebMm6b8HgFRz4zfyeB+556CKpanClAWQUjpq+I+Y
/DQ2MVzEskq8Ml6v28AleML9wKQPte0UD65jO4RwViZFZJZMKTCgK4WDDjlN6CFirXKCG6RD3G4s
9dRSYDX47xjJQyPu+I4Da6xmWWBh5Y39/IKljBdNiOwims9a8sxJJKz/T0n0Svss+eqv8P1FoeWH
ja8PnGXlBfTcSB6ajGxrMz7F0x/5HB9FB6ViCJ8BPIYG4c+Gz/p/HSxabJYE1wB3ljaw0Q17sKHs
oSdZ+JbuaaReocgZkcPKfaPRLD/Z4cHzZN6mC6OsCw3j8fbBFHUDCvLKXCAx5PC6WFKMXX47Hs2a
5PRzxAyG+6xvtKi0hmQ2amvKq4EU9IeMCdZSqzMYYp7r6wZLh+hL5FIQ+1RoEslD1CR3+8SDRTMv
XKWdcRK2Too0NF9zFWs9aCYhA80a+HC8fh1dd+m58xvf6ezvoDdgrsV3F2Mah8dcxZKD7wzXriY9
4h7LwMNmSJ9WzFcl5f8K5QZ/uj/p+DtmtbGxpoXTmX6AOzlWuSt5sWzpFb/49khHL4OxyOzOjgv3
jtyJjPXRUHodppraWHDFOGbDgs4hHpFuM9wqZyAs4iIkKUZdei/9zyUps72HBa4sf3anhuFDp1F+
e2ZVNwOvMJaGbsrH6hoB/D7lL4nRXUUNYiq9fJT9PR9MHJXLvkr9zKn8tQZrQ0siVoZaAe4QRU02
VG4hFnlGqdceToVhDR2O191pai3Du7o4IOyq0MddZ/c6Up1zXwVDy3wrEPinr6kpNs36dykG69m1
d3ZbyDFLpEUXcvvx+MCq6UmnT3cqrFbEvyUISaAoWc/hhIEK7frXXACPHwhxlxQEeZVHZgQhXvsa
tV3OcJDgAQ2bLbdSEcZNgWwoiCxhHRMx/cIM18YpF4VnE3HO+BYM1XJsqdXbK3RJYefJKBwyFreh
dExkH51JgAJxEbFtK3MCGgF4v6kSQRDBKJ+1wBPvajHanwYbzqJKdA3v3wYE0p0uNNQd5xI5G4qH
Mp9cYzl9xS6a6VwTa7AIuUVQSmV+MGhbifd8bW+fyKi81x0UbXutkIM+q5ee2HdUMnOCs6gOwlRJ
oZ3QXydNAUGEFz5EityFal3iEt4f2xTlzO4Q1vULDURShyTAc5l4kLpkV6ikteKoGV7+tIfTX+Cj
4wmTgOtYykJDR6hpeBHShAzFOKEsL6AeaQCfUtj+39DhU8+oaJ/CHDNNQs+svZKItgk90Q24GoG/
CJKy58sA7JObqonljB4FjLxsaslM7u9JF7/4yyGB+TeuREX5iHnS1URuof8LFlmNkx9JUwfkPmr4
lYJmt5rZDT3WKgt5ozg3OmIIYb/Bqv3VsKQZsuAgFCSaUuIVFd7jdlqgrCkQSzqx4tz/ROm1pIIr
098vj24SKuOitc4Cfw6oLL08FGUtOzwvLLRVs9AteMFyrZJJv5DGdOI4B04yB9qYQQmszK1vFOgQ
iYeHf5E00Ah6n2hslc/2pgul0yTlR8QKrY2DMAKSC+sLYQBZkHRxoaYN8u4Id6C5XgxPNGdXATCn
Pld0+nc0CoiK5Uz2u7xuotaax4t88oG9YDV8u1Wozqx47kNg+xUR+UBdCu/3SM+PFTL4/CB8W4os
fYsv+wRX6k+t7fa2TqF8teSnTRz1Epydtvqn/Ypc8/KKRf0hPqxozeBZRBBarSKbAHIQ1HL7nmZY
be5RNgXwxjHt+MevP7lr4AWhqmVngn/yyqGck7uCrRwwfujIk6449k1l863ghy1Qb2M7sUXTi5tw
GHnRe53cOHQmtXw5xolic6dJRT0hPhlGfSF9fhXZdoUhfGAWqG7WxHITrKUW5AeHDOT5wDJjzSow
XfCsr1gr32gCtjRulGOPrg1hCEPldekZCb6UKC7DVID+V/iCy/43ftano4t3S1kzaC97NedHiccv
MMC4S51pvClAgm21gmvReHwgGnpUFrwfXSkTAkAee/La+Fehiy8hRxfQyQPFAAH/8oCztx5wKbht
g0PPU1r3D/EoTF9Qp0/B/Z2dY5cw+Cfs9mVivb5voR1tFjTJUlrklvzSjsKlCWn1BWFt4rXc2M/g
RFkCItvTVHgayuS65+v4xM6oF1gLxPo1w4RYp66on1wRZ1BFABeeuP1nzEq/IrLzbs9pm1N4lDNm
sgoYtODj+pxVuI79APE8ptjAIMGl0+yX8Z/vDHhRlDoyq3j/c1ZAJ1O2xlC+a36iLJTs6Sqbcs+j
Ttmp+GJYqNMENpnGKV7XV8Ui4yC46PS0auj73l5ojKPAX3ln/mQ+hWUBZ1DQGT5IEMsF0Eu2H0LM
QlilwlaX+2ZZbNF7eltA4ova652zxbsot0pIjY9/fyiW+l3+INkEzR6BLM9EwCXMnmgc0wLsLVDk
Cz5p6Lyo+FFECUMH1ZNaAs3yP/USFXGl9EK/dhSPl0W8xmD8D4Lpzs6OmC4WH+NXLyz3EkohDetp
1441aVVmRDyHFBvWA0gHsSfttS+N0a07lTjVXOH6nxVtc3WgVBpeg+RY0A2IiR3sxFKzeMxd5Edj
x5DZaanh1TA7c0pAN+Y6ZUlgjcFeC5HuariIQ/Rrz2hChrWvrCdmlXZmGVEWbT6cntfUZ7L/PtnA
1gqtwrHdvhKtsuDZaNkF9zEFtD1jpGV/15cZavRHKj/9UJo6gQz8ktioln/i1hN7QEUngnJJPlAJ
fyZO/3zJRETxD7+j0p9nSLGgJX8utHIo1WP8wo6V+7RZnUSLB0EVo/PVe+APvSw8aUoi8s5rALjT
O+EcY1kGGdk5PYHPtKm/rCsrCvaddLxztbRpkjwFHW+UF0RiLi56GJssow3r24sb34iVHer04MKO
oEoUGCSLM9zxHNLkVbLUfmAxVWBgJa0T7g2eQc1ALedYB+Qp/YZMaxE5Ys1jDuH1nnTteUV8X1KL
9jOc2TuBzATyoXmxpvaOgc1XwI321s/KjRGGjh+CEgybWI+sCRoQd2j9o3CUzrK6hayJ4BLs8/Gz
5CtGSNu/KSlzLT1K3qdtJFbkroxKMvMnahr+D+xLZxFyPf0pTE6l7ResP+fZLYBtgVvABtg6zhDs
JSFsdEFOlcPC6uo4WJwEHWUKJHjuGUV+lBkXmHKXScsc9JNQop1ukG59lUPewmWhcNZ1dikZf3cc
8cyiwVpTd2XcfLAJWbZr7gVU52h88eMPusjRs4+tUXmKI5L6tbExXfWItmnLYFaBAMZ2dp2rA1jv
uFjPCWdoehLMHivYRTSKYmurdJvtpxm1+vSsnA0jXc6FAiiCZP/8gae0VjEr4cKhAHQ+fVJBq+bz
84uiAlqN2f5I2nDypCfFYpURJSAq8jC+VSNNuCJRCpFi487N2zwycsPvnrew87hNp9iA9Yp2vFdH
sawaJO0GQtZjxCbhxrh42+BH/f1rhE6xF733x1kTryraYZZxbRJC7fPs/Hi3Z02JKjL+UQKfOGz4
DnljCn8DXKNFo2D4ISiuzKYXSRnib+izAI9YT8oNa6UeYALRbeG9ZW96QB4T4t0KoveUGayHP+8j
68C9sDgD7x8FCpAQ696jJdDCOzCqXiin1CM9tt7CxEIv1owesr3NhuPRsRslJI1FDIOrppjBLxcJ
BRDWVCKlhZTJWv7arwqG3qNf+KxtsP4DE5UXpcJIzmXO5mIrCNzhUAIqUnkbsnoY/t5ASUS227Qd
F6HtlS/76tXqKm7mjXMeJlJQXEPaCvTT1ZwMgeKcl3ivY+u7sCpCVupsHAm3Y5+hKYTbb4jqkd3+
hv7+tEl18amgd4v62q+ZRTKujKNuuG0WgQs6i5dHuM4hsFf1o4rhE/37C+4AzPzvYwi8NEDbb9pG
n9mOKmknNx3gPTJNfl6B3jQg4AW2fUdn2g4XiEHQJMPoYWt4VKaldxUjZZNAYcrfZEKBVKK6DOYr
d3PgKfICMbgj/c0nUn2aESzjdao1r8hYZcV5crcA9oKeYbv7u0FoxyNQ3aR1t+Pu4F30ewVHfGZq
Un9erkQbcmqBD0LCyzWgOIwTPTh6aMShT8kmamviX33OOUyS259I6mcpDxRDyM142sNbsYWf3Glo
x0q2qv7G/bIaGsYfmMwrX8Vcjiad676PJUNptxwPQoYUZ0nStu1oEVgp6OZctyiyniqapHf0/HnD
Mrehu7p4R4zts1L9y8a2USaXnxPpBzCVskeP06CJ0PyesEFUo7YKOR0pdmJ7VJJEPDDqJQPY0rMu
ytMRBkL6CGU0rA6RikPufkQTWYaRE99qLOlONvKOU46fotSOSl9FOwD6OVVBWjKHnW/KB0IajuQ1
j8MBbSeX9Va6XYrkMRvzZO9lhKxWi5Tjsoahrt3FLnZ5UwuJ8ytsiVlX12RQt/q9qHrpNu9sSJ7Y
KWQHxkJgtMmASKlPwBT7JpR/e2nezozSv5ggQOeqAQx4zBgYOjPjAV/oqhTW2GVB9PXKe6+CZlPM
y8Exm+q47UrCIfUnaRgcVPFohHsRaE5PNZ0x12NQfKjT2dbeGErkpakdv6nXvnRpGvbVv3mGRoAI
Yn6cZVG9tODi4hKwYm4hqhJrDhpqbNihF7vvfM4hngdUuhXO1j9UhLARg4vn9a7rIPD0LWlM8bCF
FaSXYUMQ+EAFNoF/0VX3ae+5xhZ7X7glUeBnE7nBbWSwY//qjC+AAD2S4j2gfyoux3cIzhly2y2W
woyBVPOD3C5hrnDJoB9mMuZasvq26XbqzVZ1RWx4JMjQe7SfdrjLt3egcZCnz8+jR5KlbBAZUD7V
arPCGtXsFQ2s7VoV9EORS0Rys1cMj3PI11MiuIEFKyD8klGsbLZa4fQJ+36hfoh+C6MF3h5IjgaB
s0XAimUTE+3O5X7gG3hrkmGBOXx8tAUt2R8hSiL4xkmXxnYHMriWxV4qjXYVsak9zU98YxN/xs2P
3PAJr1pqQNKJXHZEBn8BW2I6nzdYZzBopm9o83IiJ6j+1VeSDRFrJbbDmRMyfmxS6sairmRhQJ4U
hrv61xfefLqgHTBwXsPYU6NeomDgtgIOV8yY7SCFmVx2ceOjnfeQqTUXKBNYlrjJT5Eu6wj11FRW
tlKjQECpTAU/pG9m/FWio8sx4gPLlKGAbdQzf65igA8vHP5yYyMGoXHSFt59eCWh6RHmVcMwkDiw
6km0K7JFIAYoc4fY8107mk2CA/Mvsvwivg924foeHTicKAq03E/jiUGSgUO2EfuD/vBoW5V0kawp
5En5Eg12Tg59CKX9QdwV67banVzUCgX00s5D615Rykn25WGUVuMGRoA8uLXl1Izjy70GpvgOBAKI
g+5VUEmxaSnvMvHt1XqTXppZArDWgPp2i8NCxBS96cxY+6cQpaMdFdrIBE7I+s9cVn96zSW0S3Nb
HXNrjaml4Tc2xoqWbSBDk33Lg+Q5lDzz6gIzCMm0mYmsZfKcqEfK9pLh+onIc2PRg7j8K5LMxPoM
60J7MIXUyAJdADohGXjWmu2Tl8e1ihxeMVlNtcTaPEelrZIPpJHH9Pu7l/lCIVvLLaO1gy6HvXYD
uZwYbzUl3BU4A1hIAC+dshlfD3tGgC8kgZUILmQbW5Bb4NExm7amJMxL+E6sTGNjUpn3hpnwtHMc
sL3DTstmB7hO7ZtuKdjncoTv7VgLCGymJWrhPinK7Cs95FWZLgY3VO3jGxps0c+SfB79yBfx+Sgo
1pckKhjk5CHEBhQC1Rt8mi9Tg4rWJaQqKAQWPvcpuZR48F36fmxPRYYjVFez+owkuvWLzkrxYYAB
KcNmdABowaFXTrF0SQwyipy/pt5bSysIImQgCHltu5F08mwuJENxm1L9cU5tzRavoZe8mLV9Y4Mr
/3fO0dpPbxYxjs91ffnxnGab3CWrd/tbPzcVH7lmEgtZ83wIvHr07PPTN43pMk90E19b9b7dCKAd
38Ui4Bz1uejjN5T2MSUkjx5g7Nnq+T69W47Np8SbZv/m6XeoSxn9ha2JoCqycQwsKesqxSMW3fn3
yo7Cry6IajF3Z8IBkcbmcv+mEkQRP3SLLmU2SRBvdhQ/2oEgNtAqc+aGBZM4veCMXusxJVb2b0HU
hGJPDnRTp5cMvoNa2Pv2Qs/PPaTpm/GfoF7n840DrdoQ1XZNLPphSUqE+HNUJp7Nv+P/LXA5Psni
aSbU0UdSeYoqkYTaOq53HM57RYWxzGpdLTlWHnpyGo3DWw3pEI0nbx70khLOuMFQN0MXckEsidvC
zgbbgsyY53IMBJAv61al1akXzidArA1lpad8YpwM/D2PHJAb7t8JR3aHb4KTHoeF3eec+fAtvsNN
hGrDAPfMEQ1tF7ytXJx2B8iOMQVb1yfkcyjtuGHdxkrBWVLtePNC4Z0cxTHPDvFcwAJYgGhLIgP0
MEsi8weUWyjeSN7jUwSB5kOzIwg5qvTWFDesGNaWaq3DPMSawjjg21aZ/tIGslZDmQu7QWN6F4v4
linmzZ8Y5esNOMjtaUhaA7K5tLGe693kr231ipcmxg+rDXJpkl24C/fZTNjd2GBYNFiLKEkqOWJ1
4AgGo+LhyENccTZ8txw4BlkY2x/BSAzs6AullMU3CQdNUMMxIBkEmWfzpMwcmmyoPkFTz0OhcOHp
Dby5cW72JHa01KArjkUI2XfY3u66pa6+kZsaoDJo+51B7W0yiUQHOtZLwBt1IYbJ0WgZXBCagB2x
awYhT9ikPanl+WWmv6nw7qK6BqrHElVzDnBGqWfdRyfLiCoOfOQzPE3cYienxZer+i5/ilBIlD5W
3JR41yf7jVvqsQgu36GYfTJc9PwZl7czacktZgyw/U6c/jtKGH5iISKwo7jogW2ln2Pprc9xDzA1
KozzifyakhRa5O5OtBBoBLAVXsNRJnPSVSF9eNEi53r2NIW7cZ44iDh6OQxdCh91PfTn6fL9ADcL
Q1oMkopAjBY36ovLgkwKoc1/aT/GAl75WpTA416hgg9eYMGY9kSYninb5RkjfVBVjejmtScb3+5S
FpoG9d7X4z8b2TfGNiEhc2w7IYIQmsAdL5rKLguQedSDNFRbq59l3czAYoMldxN1D/9gKf4DFLMH
KG+7tEjDIxU+tJn3+CdDjx83kYpEPfwAFQeAVZ/mHMBq7RRATwwxb+y80J7f4ZaYQjs6oeVanUiR
K0LIB+3HmECqXlr1QoHV//gobyc60yMkUcCfyEpf684szce3FEHFT9bulNt3MD4XYyT7UWaGWY6H
NvsF3ov7VHdhkAsubV03xWyrF1oefE699xTxFm0BvEvF6V8nAQ7X2lVA+bRa0TaL7mC5nXvzO7s1
G5V1md0hI2WVhqX4Ff7uyhDaxt8ZX05ga0AYYpFwL1NdDqUnX6DFmsJk4ur9/i8r64jbyxl2UCqw
vXh2cFWqX1nKCmZxk4AEv4E0edttnwvF1SYI7ScWdY/AXF23e03e77DFnhum2KswizUI2kT/E9wC
lSt0ZzC61/pSsm9fzflm1pOYi+t/lqGwttPNxJkGB/F0K2T3mYtym25TRa1uKgIyahMsDvwWcDuJ
ThRsiICi2kVJihCmkMi5M5PKe8iwdsyUvdy6tBagiKgecjmU6BveGcTS+ufr2dcdS1iXLLr2nxP7
8nhuDzvkpUu1Az0rxqMhwycnO8SwfEJNCHCJfVfHSFS6ybst0hP1mbfoMNDS4//t6lkUQYflwy+r
i9TXRd5ZIqxfQvBffFE2wiC5FN3jEYl1zGES2doVXHY19v96kLC5sLL1QlhJa6qNAg0tEfLsI2OM
rSLqHD8xR5FjQek+/kuPFJqJ867UhYIuR/tAPZtftv2qPo5xZceNzFDwfQUT/wB44hSepxvBxveu
JPCE2eRgEN61UhZoy/J07+b9TYcJtB0Cefrk6R/FSeR3N+GJcDM9LYfiw6Eh6FKS5UWE7H/35XGo
htcsPXTMBTUlYJEpO5F7NYOUd3hVA4WFTuAFiXkxoP5IpRcJIBBFsTNY/xLhtycKMIz1ttNY4GCG
pYb4G2ibLEbeni7+VmxmCJnxrSE5hK7TfrWqtZ6nJY0w3xRIT7GrUMS5S7WAxZYX/xMOhcRJ/m1W
RYM8dtr9T0vWLja6ye7MeEV72d8mSZJQLieTUmBVVxAVvF3mwG+aIPthPWqCxFlm+/NCvBEjXMpE
vQ2j0M2yXyqOaNr90Wm3Ew1jEHikzMVg7S/91BXgYxV4oZnyq4iY4U3hd2YNOOK+MzM5nhF8+JGK
BbeKk5fgFKkbJX85XUZ0c0NUeTtamCwckqqpVityAoedyltrYZfBKu+MaT+U9TkvLLMUS9QSNvRR
tOa/xCvVE+v9ThrsvEgO6RiwnuphpKgLTZIdmv5LZa5igQVG5Ma6MQ8L2MGrFrS7gMFsTO8Tr1et
lYjJ66H8VcQK1FNIQgbSr5vP4QKcVwCReu/GP1FpsEz5ggHDb26XhrXnswhLi0nEgMeeD631w3zK
qsC0CWBqbrnotiyZq08FEfFvwPxVZxS5LC04Ox9TzxSb/XbtjLVogzf2xUgzFa9OdR700v3OBYyV
eod3ZBxgFng3eqQqAf7c2oWLvizVRrUHE99X+2nriWJ6Cn7XWHJvZ++zSM8/EaFsALD2Gq6SUX+9
et3d8C+5YSahVKPpW1YYD+A7tl8bC02vAOw/v4thhRF6F4eHtMe7EWK4R463Rj06kyLGGJ9uqxV3
iTJ4bcfLdl2W6y0e9B+A4kaQE92mequLljiLnyRAxhSUlNy2Tmw/Zdc2BC7sgVBXJIKJf6uOSNbX
AlzvvokGBA/3VEgxDInN9FOjHOToSCBun2FpyqXkN4i5JaFS4sactFOiXqfd80RDRSSs6fSvVJnR
zoiwlD4sIscKPw9YiWhk9rn0GYINMixM11A2fKY1+mU7NJw7lqwT4YH/FPTFKgtEAXU6NslS1T2V
2gQKN+BBRx0evN7lRETjFA55aoLSh0ECOxDrjytiVrfKz98kHcQ08QJiBlKaT+WQ5i1/MFI/2hKK
+3K6DGEkAJ169Ye4lvi5j2nBcfkRzWOFBg7rln4/NsbScGV0+JN6YQclM7b0s1aITCsUZw/PJdOk
vJ3XY+AfKBvB8vG5L+7ipjm0AoBEbcnmjJZPaOs64KFM5GzvfpKSLWFOtwVbh+8OSa7zAehKMSMV
sXF7eqD/OsktJ8g3KhFl0z02mpM7B7o8k/f0sR0bYiHQzKOHK327HgFz90yQ0JPOufMk+tUg3w6V
QXjm+uGyLvXYPyCzjTzRbIZ2QhEnPV6k+t1y5Q1CWn33CKiB6XRMfMdFTRKBWBflev3AnzFDQhn3
4gvcXrVPHlO8e6O74zaySgP+VnAdXqGODGTqw3h+OW/oPf4SZDpx2rAu7XXkTUxl1NTE2t9lkmo+
g897ZZ2URO5egEA+RahFnHbSlKMOV/B2LEUTy6OBgMinmUYjCKI/XpOa1fAZKYHy4x4LAFDQEuFv
IfMS0fUcddLXH5C65ZQmlKDDGUJM7ksrXUTYtqN0fBHdTVlOayotZqNLEm2xRJ1pnJVUUwwiii9K
n/gS1FoxJC5d5o0qPufQaIIc+m0vo0jxfuP3vUsJnFkThGvpbuNh0u2o7/ltkiZWLfTQFYZb/Pdk
O/WiBlIFxu7zXpz2ZS0zPuX6qQ3pRXW8p7WKIdTpVtxV2GWp51eoSRTznWHyeIdUHZeFQ4qcYNQg
H8ql4IQSNKYKTrB4k09cGeJu4oKBJqDRJ0oOR6xuxvEniYRYtRJ6x497YXJj8BJF8NycvcGsB9Tj
bBotbJqkFto6hUphexRMksGWFdDZ9iIr6HwZc7pA9/GF2ZiUnUj/34AxvCGwP4dLgALYu5B+IrqH
O9XKyq34l3l5TmFtYAHuC+Tk6LsEHMZyHN3QrBmHYgvvoNqlqng4f4r+6uowe5vVhmxFzfTQqpQ3
PHWa0vP0zXFRa/Vo5VFx+72xTNfetOoHCVUBK66AKCmoC4DL1YZ6r3Ap0+IollXRlt+79I13oip7
/yJougEmVjchckmbv7ub0WqobZZMA6Myf4tbftCfGgp4IfKr9GNl0VdpIkUSSKXvC02FDQv6kyY+
j0wnUmrh8msX1fR2RjnB1pYk2ZeJa6nu2k6WincPWXfYlasKZH+MbSq3yIZhpJqib/UbpJAf63Az
0w5NgTYS+bVg1F6wsyQ9O2awwkf0Zfg6NNENPQYqqxBKsF/92Xzd6eg5rxMH57j/zlIt1UJiaZ5l
T6pigh+5LAWAQ+FqHWpHEIR+rUD9RZCLnAWyEzvyjxLunugwN7McaG37LKdj4oov/zItYIL9EI5M
pbtuA3JOYoTOR+8GLNU4Al+Zr3fEZwFXb90N79zo8vrNl/JsyFnVPygcNMyvY2OqeumjAEIJ4wUx
eF7z86QaqKFHPau5VqePVEcJQ8hHO8cgQ3nh51bR8hbkAFxac6uSbrLH72y3ZPar6BzaN3EWzQDM
F4PQ5wp+3+3xofHVEoAWWhSv8xlKF+zk/5m66s7yKQYygpwVxoS401Axre+7M8XBiBXZBmmlSk+6
eXe1My4xiVQBLMTunk/kcbRXefaSZY+RFFn9zzxkIyYYm1n6amY3Ec/MsfahOfNUmxNfR9ept+JG
Aazjr9u8+C2mJaBALHzA9lYOlV4uPtnQ8ytrVlOs2wjwlM318k56WOccYBNCP/EE6vG6jUs7JDSC
AkPQ5av6THGf+glbktmz9/Vn0qis09BSknT011FzX32p4pmw4ZPoha92afLUdGsVG3N1R1DhgNBx
BCgDe0cCtH0D5Zzv8Ckc51foR80u71TM1sYLaX3/HrHRMXCla1tj1zxVJ1KHxOBZ0aYeHgKOVAmr
Xvvq3zgr8ZWtzEoGs1L+X/I8V4xg53qAPnaaDba8tzsNta1PPCPcmjSYQrAjYhViY0kDMzGjSIKN
paSbF4bu+oSWSeMGJf0WJALD0+9MQOpmSiGY/lUpN4XROK5697tZaeMkm3la4e7Pw6F5/yNAVSC+
WamhUv9wFv4y8/WWQS6xzAAg0mxhb3KRBrTaQuM3HRIwt9BhSx46bgr2/+fudMLvIRLF+iDBeGVh
YPqKrd5ILw/0pkvOeIEDZJe880BPEnGxoIKY7pzCkAFaRBgjVbx3pmk5x+MNMX/nSEo6AKi+FMva
NYHRlpIqhBOLtnF6DGcBti3ENvtWZ0zWM2gAxq2JIytT3MnC9dsZmhjuwykR7iE4YUExAQHKPJxk
zqFG6Lh+HClKDv8mxmu8kG7+MopTiFvCAgY5BPWiHOynixn0GyOLowhCEbdnh3WUzFvRUUzWH/+O
b1rMiMVuRv6ztiCjTH4EtAmyS9iVlKjtszRuGzr4FNHTglhJcCl3oPRwrQOGpcktFqMradfOfoF3
4A88A+J5nSbIdnF0CoxJ9xGxneW46bpHhn78Fn+XA4qZtdiEsPJSXDSvenu9S3TyXBbrtekS/hQG
+lJAfDnGetETpYOmL7+yukliDQKZ1HDP82TqQj+UX+0Qh/nE5zjaSOBUhXdcHynhtEmDqkg3c8Z2
ufT4fw7JvWMCJ2wQTRLu19SzgM8Yd96A75J5VZ2NbU/m5GEhmk9mUwG4KhQ3wTwQnVrbEdL+46h/
vas32BiijRsiVkSVHsv0c39egovNYwWq1Y88zt6et8NANi2D+LudE65YLQxZYwTSb1o2mgGH7xEQ
9P0hy2lHLv9/N4EAsq0oI92gJ6PPStfmuRu3TZ4RZ6+OX7sbln5MWG57aXCsaASa/iJ/sZZWdf/w
yccAZBWHPC0zl3mONrPFo27x8uKnp0dCHDk5dMYKArGTAUIF6HQh8hgifQ9/lzap43xfQFd9nWc4
L+7hlmtBV0W7OHAEozbeFDss9xTBYxDAb09Ho1I6GKhpcho4svoZOb7vPA7qBXOeEhF+uQrgf0Q3
fAx9ViIM1vyEhJ6aUbok7+VQXXpcU/jpjgjbPjA7ZXFKLGZ3YvR31KIOJRsjJulNmTXUBa75O7nx
9ORpvf9WqNzfS6DpWcR4NM8vUtLHM9/uJi+HXvHNC1b0vXNTwarRyPqiXifGSDIFQWsmff2QS72K
na4EAxjKRpe31RRAeDHyAZVXTApAhSW3RQv49Ig6qNiWlQ/ZluPpYvM0djxWBtx+LgPOHSvEtVF6
kRq24MS6hD3StklpUNoO1PzItxyCM4xogkYvn4MHDTJ5hMtCwLt8BTPqChuVF18kbrfUbs7RsRlJ
GuN6CtBlnE63g/G3qRHwXMjQDRZBYha5UqhXhwS/Qm4Nu7/o9KtoTsEaR20KKIuIrUt0s8+pBKmI
nJmjCqTF4IQKmdvl79cmVU8Uvl15OY/izogdBo74zhkcgsac9q29Yxdwaqs/5x4jp6xKYmpsC1/Y
/CFu8X+r7QrdSLRHQFE/XWctyfxPisMZc2rAyzyhH6/XZ1RuLTTi66b9zrxTLA4bJDA/EF9F4APS
gOSyFSyc0fNI/LotvQLGOkAsjVI1S3y1mLjhm1V5wIc/Ivtypl9GaR3H7MrWVNGV5sBSfWhtaD8i
188TQNJVnIF280WJiYYsxSBHffoDxY3UfpBxoand3BmobaXUQSWd3ijauAM5wMSGQyDg/PF1Q88p
i/kOvRUKsxvWeHcURFt04pVkdruH7mVKtGPyplAfawFijbjjirca41sGoKKmToqwbzect3loULkH
nBcaAbMotTN1uUV1Day6Z8RZgGMD5dix4XzTIJjwp+6/6qcob4UeJvhEhquR4yBMe0wC4vtmagqZ
UDhLlr7782gAZRxJz9zeuyIvdwPgWsMj5SldKqYroJXsrxfU6vmvCyOs/BFan5utxUGe6z3QOt2B
PAZrBsnb4+/jiRuGP0aF4x0sIfilKnyysWd1Se7a1DT2r3K/iWaZuL8mPwJh5NdkkdvReO6cmkKo
6f1e4nKA+ILjP10h2w2mwWj/wk6WVl6dD6+IoPAlxpvJKADfiEDnfuTnPEDy8KPXNIjia2bk/2LL
6Nh4WopY9jqpRJD6h0V4yi/pxjTxwRakFSpaZpZ07axXOf31LOI/x7P5YKb4iT5nJWjKXvHN+0zz
CBYO8XGGWocjb0ZSPTEi7ZMoA0LE40rgfxW6Wv03UE0nUEc2DIOrEjmB0FIyR/JalYUwTw2Gplvq
UaRTGJic8qzYLxDy098oXKzzq/V7iqyclsKL7xr7kllxD84rUna/U6iEvmVNQLgiVvwI9pKOhwv6
xp8TF/oJg9eaKAsEg8Qnyw/nSa/153t3d8QBFIXkG3z8+Jsqc1pcEc3jmw/GAaohJflay59vNWG1
4Nj6gjIPoHsQNiautugDjDdey4cPIuDOdRZDlGmMel9c9/y4hPsltACK67/tYH88W6cyLW54uuSa
Om0RP2pb9kPyT5RCiivB4PMOYV7BKwdgr9xJBsBNxQO6xAzAZnZH3ZiG8+ydaJMdgK1YBsxcYkYk
n3UhN7+AzJbhzq+yvPNrlujuZoF7NaOPvXUIFsdi4OdF9mhc5CqF0MMy4FZyyoUQdHo5xaie1B4h
nKef0QuFqstEfON4fBywLnrK1cVLPslmRZ9vZxdhuBNaGG9UjeXZ1nOzxca47h8sucl26kXplovl
unxmM5GcFTy9xcPY4SaKnDlR8d5LvE1jlty8hz5sc0dhgtCCDHrJTdLS5yk51fVDgYDFFd1Rr3eL
arJpp8AyJjD4AaXPF6opp9u/mnTS4kNXaoiQW58oSfuTEwpN5Dc5xdGUW52H/ogvyw5nU0dnNI22
5znEBg6ZQpfQvPcf9MYa4L7NcgeFO46Co6Khz7hddmXpLTHaKIAQDrAYSx1/O9hdVS54nEY0bMHk
IrRdXQiZZZJv0ePsU6P5rIGBioamUguiG9b0TpbPqbg9HNmFqxTGuDYrSJPMsK1mMCrz2Pxfs70W
pdej6jyB2tiPbvKXdey2BGanU5D/CATZJsRh+UmaYVr67uEjAzHoJUsD1C+74e3XwTBbv+AUsh3Q
5CktmGD0Q2kjLYVu52vFFwGCtIlPetD6QLX7IpsI5AUFYjEAgwYYJ3bkUEZHtBIDCQqgWKwjMEIV
i5yFJgQnM15GPNN4zg9qz1OawvanXtI5r1PFyQNJhja3NBFdrpkYb9sSZ5kbvIsugyxrMhmIppmE
8I/kkIUo76KAJJGjufo8sk1feDEqcLxIzpn5bP0NBSPoTsFrEEXNVBWG/uu5nLWY5mPpiHPsjhWo
NHXhXqUasJ4xd5KMX3lolonKOnAbHOG8mOWaYCPBNwcsBBqjmSqs7HUx9J2LuR2wRQZdtBGr6V2P
0BGXEzesjntvmaFcmle+zIWVYEvS7UeXrRYZDN/LXOnvQYmtXFwAFpm3k0c4W7zb33mRbQpuFO7P
ZoRnU43Ac16DDAFzPtL7D9WdTpQYheFLqz/nZqBu3qFPSc/zXuIoMp55P5HTe5ZWMCUYBJ9gFJSh
kLLDxGb9S49NphgXuhBNu9HGybuY2+xsNRviee5dIq6dPqBVy9swTNfnRtV+Vt4CF9NFbuB22c67
biosuF4lTmGCg7ArJ3UBWGsvf1xug0kA6/IEM0WZ6XHGmucgfh3QQVsvI+OBmhyaGgtQX/BcHwNc
3c8LpDsXAJnq778YXmBNvq798kFrzzc0TuL1jX/G1Hl4B8p3D5f2tvS3BsMQGKd95FWFvNiLv1Zt
oDaO4YupIIwMDcZPtGCXTaS70sDIUdOjqteooT05IP7N9lKmUit8x/ImqBYcAXIrCeJYIfZlh5db
9oUy8m/MyUSMwHPx+t6H6Qp4v8QSyQgPLguMnS4MRR5nx/AaDVWVcvPrrqey0LCUEpCcj83HhkWm
KRRrfo7qday44suyfCXkgt0EpNwfjvGyC8BLNtNnGc1HMGEkHOkmbYCXskFqjMR5akV2q7R9rIrn
CFSSVGY80/aviUjh+vZTCE4I9Al5Ws1XDptll7ZhMnKLrNQUAgAxpEiGQFm4xNIRyZra+o+kUcOO
9XItxpBkqbQ3gz/piOSQyEoITdnXiLkhR+/+WJF5z0FvZSMr8a8/QMKcQCnBWICA/Cet7kd1g173
xvF5BLAFxDlov970UiSqjpDy8bXBjlcUly8f+E4+Fw8D0xvumELFG3Aly3PAN/DchTJYRi6SOvAx
CO3HAapgMGpPspTiPHXTQDbyC6ovxBxuV2dbRAFIcUfoDi/HWVhBgl8vn7m124ydBpMOszJSuJBt
ukWn06wpaF+ZPdNGxOjoQEAT1Ee0KNUhXT4tjhKDlad+6W/uU/QeJol/iir7zKTi+KlZSfgitrVJ
kSXxwxgMBgphhjHcu4uN/UUBQQGiAbA+YzrK6gzKsMQHN8Dzvn99ghi5uJE4dzCxMVLOSyXXKt8n
TQXpv2zkZlS6oLwWxEfeAYBO9Jk7OI2QXAL/n5JnV5X1IFELbT7oGEy15/PX85AMOlCjpebxx49z
F93kYyJoh5FAu0NtLpK5STtRDXS+pivcv58jFUO+7HRJBwz4ODTDuXn8iLpwjIAbcKaPjyy3rkk1
8/8b8vJApfmkSv1TF7DezHKuk87HPtUN3HT25CsHVganiauTKDkVKOOwGXosJ2zYxl+I6Gh89Yt3
PhWWgbrwgbFppYp6BgP+/o8igw9T31WTY1K3qfes5QifebziqSSJU2Q7YftlQ9bL1wi3+emJ9M6T
M32PC8h9zr6liPKq0JtMIm93ErNa8rRg2taOY6I8bDQ95NLlw0Zulu/BmCydCWhgJ0xE/6HVOrVz
mMANo9pxW/7Jo4KHPLqprLrWnm0E8rfvZF1+FxmAhtSeYjHVlNQinBDouPuFr47FQ+DMyyqCNr25
vxRJyPKHRUmgr7YT7jQxiALW0VPxGrZATxu6DsuFFGPgNVj6kL6/jaA/2IwSsqJMLWs7gXNeFW2M
NyFSmbdagdGH5X4ecw/8hy7fFrIEWuGgbr4di3orF2cKUMRAXpflnutHjr9pyQ9dhAEHpEIfVp6/
t6T36j5hJ8BuPgFK+lYQhAhbeIwQPUtO0nh/uUE5hjwJ6j50JJY2FBNJGclYALJQAPXvhhzH1M/F
7X6r5bl+txfBSd9Wl117PbjMVgDgX5D22h/lfdSsizKvBEy2nOSm3b8J8Hez9yD1wZO7nIKFSoSb
s4yp6Jbijhfhv5Rpn3HE74eELPf9lnkk8PxPXaJ+4rqttky4mt3KNoIBqXbMqKNTloUBDogsQ8Yn
jTho/DCk24HvcZyhDMT3JTQAGrgL79wV4Fvz17N0ddslvWDHo9Ds/OVnyWHNvmbBQTkseMU6b3YW
0HJJ+vgqui9HN7gqqxqw8PtlyCW85pxqP9USU/KB2jgMxZOl7hud4VkvJ3oauT0bxCXTAHYRT/OO
XGWdPqkkhAHIHh6duiN1s4v1umVQNfAmVe9mrh0PgjvY4XguvjAY8iUhjre8tEgE+sxJri78OILu
BHXq48TJQo7RFYO4jlIGiyQZU8ZpxpnGq4Bn0XM7F/sjCItaos63szG8Sfbby89lVQ5ZE2aCh/g1
sMHW6kL+tJYFiPARahclkOQXTG6ApaorA28Jfs2mO7bOpslanR1moB2fJYyLdCGghtDGillYAIPR
xDLelZRD3tY8qOY8cvT807dpA8SIoPzpQ+569Ii6mRX1J6ZhXfjqccTlZdmOiOqvdYbtSsn34WW6
wZlm/BSwduqTJk/vJ2tgBIh56dQnV3tFhDAMAoJ7c4ckfnr6GCH2VSb4PGga+qwAfZY1KsuK5PPc
kwDPY/ebUsv4vRUjkCDb1Tj8jXakrDg6ei4aAfNvHTbcEeL+X0r6XxVYxlvE3Bd06FrV+2EH4wKe
GOv+jzsbFQIT1g6yfGPv2kCc+rQ5Q9DFdzGH2gXxiK3Ga2OAjtGZl5D1juSsdO72MNo5hiqscBcG
c3mPptdO6o5aii5/SFlS749mfwX7CVMy0k8ePkMzvK7KVXMDZV1xREbuMBajASKyTDAxwnyekph8
axuvK/wcZhxPTgCXS52U0aZgXwwQUXFiRjTsomYuS0+MFv4ZW+Lnwbgdv8nBO0besEshpsVCxWhq
DuOtIVCdZaZTwVH1mGiHQm1C5QFLL5uO8HL0Jlg2LkbVm5bwN9G8iz5+/3N380T62aU6evb1tLqK
1DG3iMptrWl/cNIPd58vS5lUV9yl1prk0OsKwhgy7aq4+MrRV/ZVBj0i6TwhlrcbvQkroctpa7Q2
b0AF85AwhzSgX+035NecbSp1dPH8Ytdnri0Zh+mxu8xKKQZpLpRGNklpQBPkWh7F3Nh5i/b2BA1k
VFsvMLV9+3g2D4KPMu/VqjzOndfT92EJK1vI/MJQQ8+VCnSiZMb5TTuNsInyhDD6zH02FwthjQvb
Y3UU4GVFP3KDJqWR4DAwu1rApmFJ5BlKF0FK4wbOy23fHy5ef44y+0QnyEeOKPdsLX3UBFPKndWk
T3RW4/mT9qPlL17d7JYNK/3LyJr7u+talO4coNAioYuzYczpwf8/H1MA+C82Zqm96l5H0MYLhPn7
nUteqYNZZ7oHi+hVMS/hb3/B0vw48Nbln3MfvUC3Alws0iGAB7bvG89NXFDgNyKdLTIFL4QdXiQo
13apOHYszXBzJ8bzoh9R37WyKWxmYV9a2AE8ZVo/yd7sFrxZ0RV3yKACXY5GU1RnqfFJsBSjX2Cb
RxN9QD1Hb5P/GYOPM7qYJmmPr2MreDxVCTTdK9G0tXv2IDHHlz1EVBr5DJmjyDgxiCRHvclP1Ab7
89BR/Zp621Cfrww9R7HfvyA2XTyVD5EAyd/SER4c7WWjN8SBDsjN2vXh5oiCI/IBOcg1hDhlqdpb
mmubKznqgC8rb9GAmuf+BxXOHV4hw/POFb1+DJ0FU+HSZ9M3hFPsKm5JAyDrlZbrvowIiJIfBANC
diBcuHTvGL2J0DmN4K9RYNcCVQoilN+mMK1C093j0oJKIKWEWJwolV1DKGRTygHOsKp6bqnSMlIG
pcajJyuAChHor4Y7cbcxkbhtpBgYYxezFxHdHuYQzkWJUA21f2jaeWs+2O+pVYW3n88SVZQl9T30
ajzYIHIHSJJNVyqZlQGDQTAp4EZ6x4xFEngjpWvXj3QmXvuAeWGrygp7wffq8ZxaeTfCPCNAXGZi
Se1I2Rz2fgrPWI9fdL4gSutUrs4tO0ZMTew0i8FsYINrgQugM/bSQQ5B6tqz8nnnNNjAlsEGzJzO
oMmtOb42L3luYQaxj9anrwmEmElPrdeKgI8nGW2EgI2urAh5uKg3nVZzfW3FEl/G1CCqFAJZn4gL
wOpf6HZ3dhNK2FnZhI7KumLDVPFf2I6/wbfivg7XpiS4LIoIv8mvOwhDTH71TV3JCGyUOH34NeyX
jssgrHav9lUwCGbpKv1CYniTo/MWtvnDLgmHwZOXl8xOFtqZxTzxx1uAuxQyHoPzwpqEt1Ks1VBr
bJ2kgHaeHW9KMBUgRymvrmeDVGINZTrFuM8rY7/2YXnIJKAT2eOTbiVhvP2knuiVJC5TJ5p7DDmN
ZPC1YUbxhzWc3RfdSa0i3QMHmHBZnUWebqPkmPBhaWw4Sx+7EP4BwVGhHEfziE5v50UZVdO5LjT7
aWFcrPRDcLpUuec6Uzt6E13hOJcoYuB12t6XJpRnVT4gNz4dwW94U65pfL2e97FP7R8ZsT6QdN5f
lzzUW+t5DZwJLDCm4ezeul7Rw8Fvu0JyvYAY4n/lbhsSKRK9+l3+QgAJwV++rQKH4I5SOI1ZusNa
W+BPpye5ko5lUwS9J4cux1HORU5bHB9rnF/4oFnEokdF16gwKuq2jmAaIs7dGiHbzjziie0SRqWV
x/ea4phARkcQQxtLHsYkfcbmYQxBGr1o6zK6q/1oSVk01wxfLXK6g8FFgQM9RwhqSGRiQcdr61SA
Yb8+ueOP8/ekOd7lhhhZqlBvWkGQyR/D8q1pDtxl/0gf2uHafotklnnInnxN4/rfOipUaORdogHR
rWJGlwGyWBrf2Lg8OifnGK7VhzKXi4XgYTnwFmO29RrAxcy2hsuinthMOhA+hw/2tI9KbdqHvv46
3+11Dzv/35SfCWPbvJZJgqmyEcJeQoStD1g0VBxG7ZTT/Et0cW8ZO6KKpm9Yc0B6NLXA5hmfTLkL
GuCX+9ma4m9ffsn8ngK78gxa8tcdo16uwD2TiuJD5PcWj6fBSNyM6sz7KZYV2IVFKhRFW53D67Bd
QFSppAZpdF+DtE+yNk/lO0Oh0BzCAVE+xvpMSENSWaOB6bmecr1C15IQcrE7NdI1zWmzq7L0eVBT
vTXwa+GeZxMte09KwBo1rUnOUA5qkONXitKDkPhl6MvbK87S/cO8YuoxSDLsNzdjTcig2FYUPNf+
XjRfiMJWVzxwOenojbCE/xAoYpd+pu4OPn6pypchx6zFHSb8UlLj9N+iB+3HnFtHn7I3LvXoMuGo
j/McV4hK4s9tJ7JEZmnljk4uP6IiwJ0pBlLhT9fZ109Qvbyy2B6AVdQ5kM8C4PIeGLILgR1oZnaX
oKxlYjUKrTsXCBRVquqCW6dLUjr05rLTLuYNoB/7uOfRYNK+rvorR28eOaVyEFPyvH4Sz0Eg38jr
ogpugJdiGG7Ykoeh2WmS8Dt7qJnQEkw0sH/Gr+9jthL+hpnWNJ7tlnbRTx5cvy3OZxn80aKoOWyH
0FeVxhQze3hmqm6TeUL+Vej2IaN0FPypxqkBHrGEb9zr2u4ThB+A1SHrgRidywykEBqqzYYV/s0O
/LnE2WNsHEdczK7HL77BczgnkxXZn2KRS59F5CeVviF1BLwq3Ayz2t622fqzYjiTyBV6XENQS3+B
vjW86TpicpOQwjs4ysU0At0OVPoCcIh9I2SDN1JqgkZstJXqYnTd1U93Z9gyjaeB1u2rzfhUp8FN
VcWXCDI4j8gB50Belg6KYpym5aKPFlQ7oCJFKGgziZJBnFGV+F+c/m3HcgEX6nUBguB++OZi4iMV
kRavfy96zIt05c+UhbSDGhy2CqDocEORXtXIOMBbPIRANO2edq4Ad4waguiQEYDRRbbZZlCEcRq3
yZ9itv+dUPwiheekuYvbzC+LjFDMi9Sl6lyNaRHI1ZBScHpx6OD7i3D26Q4bdm1dzogDFwv8IXvI
2yeyDJdpuaCYNCSSMXAWMjKD5+tvUDzontekrrPILW3a/jgLvPeCWuGLPIj4hGNjNxY1dODe/Ktq
byTnGr/130s4GFl5xkzdfiIvgB9pRjqdfaTwMwYRTbTRercmYBJRQ7gZT9Fw2HHJIv+pUQnvYPdd
UPZMgxSO6FCsYvyIMPNhWFw6FRnHA0OqtdQ8o1OWhmw5JgiN9KvbEEMMZwL9+lC/C0HFGpFz2ZEP
gCk1LtKqHSeC8k+1U9GsL6dBDiFpJJsf4jGAY8P0hP6hTbHTbOlqQP3+aKU5I/6SkUMNp2Y3oEeX
u7n9ZoSyLIjeTdSrEv76/4EMnozxLYCmxorPuXl685ImXq2Gyb9pjVslDJmwcK/IG5SGDGH9OIuY
UgPSzWD9SohAT+YF8B3NSH9LjNVLqftzj+CbZ+GC4eXJBKj5S8+P0Dgvyg5cPzr4u3vLlp4j8LLk
0TSHAsd+NP03gc1F3LdPiqgUwhzBRCq9xa0y37fxleI59Egxq7DANkoFUlUxH826LuHXCqZ/xERq
5Z/1fjkKMrsWpGbtZ2kiFz1amZfYlFDCHFpWPGXc8gw3NkOCS/meSm5WNx1Cf3VMBmQqIxgff04t
K+Q27sBc2UV5WY/hpO8FyXFJxsMd8pHTU2GyXUqyD5FjXQ2UUwIOIV4NsJowgybBtuMgA8anXoIk
ttwCDcv2vmzfHClie1uXYv/JUpwPQMK0TYGFNyLBGhETETDMWIMXG+mTxOWedEJRZWSUh3xRk5yI
fDVHVhm5ffWXLGDBSfoyKKZ5y7l+qjcTtILqLuAp7POwhmE08TgE8uie3hGuI7jbGgs2vumZqc5k
QnRyC9nn+ZseW0CSRd5p7zI+uxnd5eYDjyCU8/uB2giHrGOwHU8o64rWxGCzMBdBEqC2Hoj9faVh
2sJ2NQJ6H3DiVX2/+jYehhKNuJ+3cjxGFKQArWHlJx6ifMxRAp30zm/jY/vW0dipsHTrj2eXwSEG
xfHbz7SdI8IPNVe05FB52s+Dgf4nR6rfQ3tWc60nB8ynzHO0f/kW3XuG5n4JIzGvtHbgOcSN2uAR
iXZxRTr08llnH8DGCJA7SML2KOvWMNkmSMCzZwEvv8U6hsgZ7749T+hXpmiAmrp/imfsc4VGP8rO
RMuzibNJKByPXYEQHK0uOzhRkKwcCLPZIE9AAB1fnhYUpgcn+Wn6G80FLmHMzvbKzv1vfA84jX2G
/hNu9JF2JLe1m0x8fMI7WMtYTdpZ/fe4w3kWoXwnz57+yo80Ez6tp2bgG2rOuVQEefgM1R4aQgHN
r51Y7WBvmlyENp6wPRwJbWPs1qWf2HssR38vDpWIhebQdsY9m1acA7WnxZCRJDl7Ag+RatFnEM23
Zh36EXwJ/W5diVEzx6Blx6FDrzsr1b7SiUfN9pORDjwys5KrkaoEu7m1VqRS8szXHa0hKoMfPfH1
A/lBjVKPtjthsCT/iO311VfuLvlB61ofiWbE9GhDDBUpKA01Y5rzzvMPFTCIXvXxXgow4V8PeUrK
DCbnLtMYS0zaTze6p4lvtXsz/PlWFSO/3dnckEo5cGExet5nwJtiTcPNLYH7yOYA9UI8W9PwRKuH
iIkZixEf61yQkcKA43uO9Pk5r7N4CCObG+0r/xQMLWaxh7OYMa4qEbbksMOQa3cvFtPjaweHbw6K
NxJ7BTIuu+P1WGzs77xA+DFQ/HnQRrn5/aA5SILbnAW1nBEam/YFSFI+3Bd+ENvAPgdWm+n/erQV
Ok930bji5wh/LvXp68uumakCi9u1hxcofxWbMo+InNqVtvSdedmrgVLCKDR08qXEy/re2esHL7Sx
iU3RRxuOJH9F4OX235oKkN5M9rp44rtXtjYEb+gMb7f9eZW9gbiPYI+jQqEWYGy08gWX/ZRTtfbG
AN6PV4bDudiRatVxM4b7Pn0hfMiit7+zln9Tmv/fcORdtrRiCt1tAN85/cpA2sv1hLrXYD7GHGtj
t1i/a0ttlecU9C39Na/ZyYb/GFhQTw9qLrSkWwscqf/uaDVRajOnvH15ot7RtRsXnoq9p/y1sjbA
g98VXdKvW3yTe8YPoKkoOPNwvpdMTrxOdHyJTv4W+E9Glq2fqSRWj4WcuYep1byfOpo4AGsd1znF
Br8Ebrde5eKcRzcEaLy/bGHCLX1vTuM1s+7c8QDh1xdFVw+ty2mNRRhYM+kfo7XEipfAO5mWdCnK
gAWrzHC6zP+LeVNDMvcpTLSlFTe7rxzfENvch3ZBtP2KhD2kzvFL9Wj9QGtX7AfbTcbvYTifgwcq
G65QnaBeI94JqusRsN3Y7wFVFp4Gzr1jkBPty+rrh0WnIECRngI7nD1yh+NqP9C357m43/TRhlsy
mcH6iTc4wHKmJafmtcODA/BA+uLuTy9l7fkHOI9Sp/IDazKB9oF2MkRZ4BEMMsHoz9+pRTRkgYnP
vPtx970BD3IKOyeW4QQFT8TNAdL0V9JCysvmJA4faOqvd2zxyMGfNS1aORYDA/0qMVLnoSjmHI5e
ZjlM4KSZgMqDDN/w24QTA/uxxel/DjCu+n5XCpibdx2nYCZfdw98CZK7D+MfVwfxsIJROAmI+mSG
xg6zLJ+nKbSvBsDftBMlxCe0m33O8PbnOdTnLZ3MJv6EgW+3i8KBUMZOPxKZKzwAxKKlICQmkWnS
2IVvKY0ey4w6CYZUohP+LOctnD9hS0EoTId3QslRC5Ab+xHNozcaLg6nEeUm6JkI6sjl+Kk4sAXU
MAotEWDF2qixVWma7zeAkHMvThfAESSNIr5+sdSb6nsRiJsmitv8f1JU5+iZ3WlUxANpPf6AFpd+
qhHoSoSYEFRxMayKJUNhWmP42dzV+G+eaBkvI/DtohZfPObkSbYuHpCJVZRaiHSoTmO0jZHGBYu8
qp+LUYuocrFxBJ6MpXdZ98gLxbhDjYTibilLnjuwFhBGj5pmUSIl5bt+5rO57QPuTl6X19JUmfwE
PDAFKybPsfNi6+j/C6UCa53j3EPCBhq5zk+DuZyOswBCRrBWmxO/bjO8AGjynW/RS6Sx8m7Dmjpl
7gOGGa1Z4cv5UwPtqxePT1qqMwdpXTFn6UxZasyam4nFMlGoQ7fpM3HGGG0Suods0Y+QEttfxW3r
okVdLu7ANtZ/P69U4XaBMj6RYg78uY7Q92i/yqlIhrEoCp/mdNk91P1OEseXpUqxQ0O7fwIJrZ2t
mQN+o8zG/SheYP7nLh4yOumPzY1N8jj785HNsSFBCc8+v3stWaqF5FCymS6qqMpASUBw0K5BSm68
uYGeKucxeBr1Ty1A1H4ASNoQi067XfMSQgp7iYaiQA+toMzcjjn5VENvH9KnZg4prlVSpm6Kqb8e
9pW8WNLRdvqiP51R5tV1RYAnz/GVOIls0ElL+nFxUc9NIadPJ7Ip9JW8rrH19R9/rrFnmqf926Kv
xMDJWwEEPOci9GW9nA08wQf/2sEOPR/WFFNtLB3J2xodheGNTf1Q7R60Ry1v8/H3J26tkOpSb+0W
sBNYTVvKt+AlnHmZpCbRnU6g8XtkMPJWCbb371eli0Okpc1yywY66o+ZmaQJEqzPMM+wjiNfUsY/
cqTDxRTQB2EyEBDNsOQNLqy2bm0un16sSecdtOhoWXT2+VwJUJ9cgpPTTXLMGsnlA9Ag84AMyr8F
H8G1bH3ozr/IYh5WCbTXN68xgX7xvJuF9rUo3zPUrmactUZd/oc+xLzGGjCtFqVxWgIjZ+bouHG/
Qw628zjSoFoRjusCQWOVJ4DTlIauOrMoWZ75CJBSkHcVj6wtbbysx03vy5ZzNcuGq/fguzIoHb1T
e/CbpRV026RB+Q/W43WxuDg36z8h56FHyHiCznxOL2x/mcXBcKQmJRikrNyS3dWwRbm5gYWLKljY
Zk0WLSXrnIkUgBoA6gGnwAUp1RsB48NcmrNA2znGJkn3G53D713WSB8HRKVCgbDWBw10s++WIx/b
mzOKHMyMWROWgjNPG/D3jTrSvYNHutUdrG9t20OnqGu4QVp3HVRURFP545pHIVj7vv8pFrE140cR
wG5z7kCfvtbQn3v1dEcItjsdvlgf/8D/KAieasxdc6seDgT/1lXEjuHyVQ1AiYRk508MyZSgMLx/
jJe/Wikeiq3hbH/U+MiJeWzECx8GNcU28i4Lt+UOkIhe79PXHA/slAQeLrBXb6aRRrec5hO104h6
NqPbdfWjZZmt05iFXCu78d/cTfWQGLupe8A0GrzyLG4O4EU6sok9IHXtlmUEWhcisJTJjcxVw6FP
Ftl8syU1+Jq1uBW0gWeruXZXGiTcx2M6MojI131/JqOEWVlTOt/oMCYVhh0Z5OXHJjt7nRb3uwSW
G7Tdkdjy/gstMm45v372IA7/HpxWIKU755SZgdFan32Tqzpbjj2WUjOtkwewCb+dOolRWGpJrnqL
9AkZuiXKdxDTYk+jk8DmZFl5T2HyV8YWtjSmdM5WUcBuxgv4ytbIiBACotHbLE990WusioJtpqZ9
aOQGtgkMOqKgYQbBK9aViALeUhO9bJUheBn8Rbn6c6GcYqvWl6HPyVqUVvUq44l6SZ/YTDRk3mxj
0LYxANx3QAkS71mtZBMgon98Dp60rl9XMUWuTfvmVmje2jHLfvOJ7flzzKQN9NdnBuM6e2i0Nywn
2nweL/BJBpTp0DHXlFQFTJ/0NJcvWmIDvmsdibUy2TDBW5F/aJ+lPwt5hrzUJCD8arJHgFHj44ay
SmA1F8hBac1PCsKLk4RgbhfnL5devaZ9xtmTUOPtXHsjPFZamPfe3VESWCdwHmgLkAKcEBlBD6t2
EFFgWFipUdT5MYUgqRbTXXP83dCTu4xeyVElEcSwETgdHPuz9vjztU0u4Hz4x/x6eUVf6n/7WRMC
+ViMOaDYKcYh9NubnmNokDlj07tO4agZLao6VCY9ef9B2wcBY5RHT5UVUOEqSdpunTUEqchQQlKU
j73u35v65SpZSwf6303FkFomqUS4bsywpvCwsQdJf/1m3+Z7okshqcTAJngp3vc0ofDBLrK2S1OH
dhenkJOierFuAYPl38e+/eX1HqJ7ssD6t/g2j6Oqc7HjeA0u+IbkwkGOx0JZivuXFI98o3J18sdy
lIwRV5oB6YW5jrHuqnNppJw0JoWImTVBAmlILTCw9E91aK+rNLPDfQdCVYZJzK0Kx97zcoe0ytyj
tcfdAEQapCWSFpXK4LRQeW2JyN5YCXfFDwAqiIHaQj5ixGFdNhNDhQM+FTBkBkazvXNKPMIyPdIt
x12Dgi9xd0fr4eVdtPFYDxuf0COPGW9JPyg9ZGxaXxemk/Gv06fPnEP2PKswjw2SxdnlNTBxWCup
jtEv8eeoDXSWaUGiX/ApeyoiKFq/leYLz0rwO6uLsB/DGbPKzfPjPc9ikukMjtCi9iYg3sGCpq0a
dBHbFqNVvsYtZHNiUA7/6MI6UhyRddpc+8Dr4OCviCZV62LGeKmwv9OLO/tZFYIAGqDQZC2cGUMt
VVu4XQFE2Cs9XI4hLT/X2jpR2r6nowwp+b4l17uCtY+AMYYwWNtgDqnH32dGDHtoxSQIeufRgyEK
wsFZQs8LbLxu5cGiZywj0NH/5qdvUgL1MbW5mSvxUtvG1qYrznRw+LYfjoDFOJbA6lG9Fu7WLsF1
LqcconGOktGhuqZe0Mqzl7z8sIAjwjHQmLHxib178fbWiR0GPWLS0jjO5i44aGe1Ip9NlRhWi1et
5hDG+izEgIs+cFB8JFvoVv/rxKi/pQFSNtMVWRtdvXj/ktTgRdXJ+asA3JaLFyccjXqCa8ibSnpE
QIPRStkdAbH2W9gfcxMSdGWh77+LMQUUO1xhbY9L4nG2NtIx3xpo61aCQXjiwPuzJ8hrTm591CQk
LppAd/6bIdYRAah+/gjTOJFOAX0OfSZheC24VCJcI/ffvwKmRP9aaO2ni3dt8blcVcY8nBRQoZQw
RFK4DhYjATfbWfZnuqqI6N8LS1Y39cPErHCTF8lFgLUscFcbQVKErh+w0m/aypSIZDOqHNxeNyyq
ly4tYxLtBTKlgEzV/7KrtZpuw8FKoe6SUgt7ez5+t+5+sXjCwD2utKpVdCq5JTgy6UBVedKsOR12
tmPJI9lGMzJS+gdtl1MsvBChqnFW5s/NgKtHsK/Idp4WgV+06RWiAgqyq18Rg/pBhH8tf8cnAhkY
rIhXN4Kxq2Of6QR3eUQUMFJMQh+wRUKglDVVpPxy+TPw4PH2vmqaBQG7nypKFPMDl/XFsUwgfs0A
ejb9zSveCXMgT3+4qcX6OjTH6rZ5dRtbkyXUCwjSncM8gP9di9ZZnM+SqAyE52K8g7GPrwO2sxNn
El1fxMRsnyCETn2giR34BVGTpBlQ9nHN/9q88vNeAqp32xlsCFNitovEh73uMu1mBGvfejthq1M9
2EW+/KxBtnZpZ4+w3sNvy/D8HIsx6fQyPLNMt3MJ6TbLYrbHe2jYaYpszyj1Xs8nzW0l1XkZAvM/
EdPI10YVwYdVTDq2O5hHDOfzE8hePG/853mbPUWtJIsJddoFehlPqJOm8WJavfn/QGElq4Sx/JRb
ds4IE/Oa7mZEn9pk9iGcSriYZJa7+gVO1QHXRoPf+1hfL8vjzqHky5L6+8EaSZKFP7SWlA+xzbUY
hBFinvVYRGxRH+XwH9ycVjyQCOWcAkDWFkWpuRwPZFBErGPQ1MUPealmoLQqMcNbpb2UPG2Oc+3i
tgBJohweQ/5JwHcc5fTRy7FRB1YdjquvXrB+6bTGRkLQeYbxDW7GfI6ujlnMZBEH8hic2q10ByvS
pTH16pkxYVZ1P0b+sXSKXxN+GtdLEuIiX02BdYjwY43DlCjIqLoFR/LdyKeL2BhyjPz4hqYQgvU7
y9LKQfcDsCvu6nWkwkIi1snVNM/DYq+0f0aNWIrAkn6PQIGPySsvMzy12GyBX8Hz/3PocDc1qVsg
ucGto8ol/7RUG0DxI1lf6eK690d7tkkS6iTR5Sk8PUmC6Dp/PjDT7EV2zNUerkq6pNfoK5JR7ey7
dGZAa7YbpH6DmBq9qfuHc0JcTDK+As0dDT0UIy8Yd/UffH/e0MOkadkgpC4uxhonEVcsW6lYr5tF
lt6jR6DG6noWXTpRNBdtOpC4nwe05ObougFIRJuNtdCuybaJT3No4+y3CqhFZ78UryLxIeKerhtI
BvOL9fEEAfVlxxbdbco6g+BNpLUwchWhS+E2UDQMjhglTJsDQ5eOD1pZNCjlPg840E9+IsctObs3
4ZF0FTomx/6gpRGgNYE0q/UIQm8hqlNe1RnpweTTK8pjCY06fqRHx640v8X0E//2qFO3i+Jcw2kk
xZ1rsQ70ClVhu3Yrn/p/wDbFFxVcYyFlgqVoeWFGkfU8GTXzKCUypQDFRhDFBbqkicHWbp3GjiV6
Rk6Upy13dP0Y4AATioJqnD7hpPrM8EvyiqcHUL+JouqtAmtnt2wfVAFsY2UX05EZSAu1FuP/9wd+
FeVE8VLoZCKSxRguzsuohjAW5sKRRl4fkfJIS5UCT0d62OV4gR/LUeq4WvEcV6r32iUUSrqMRmj2
g5NlftrGGXOHyjaijoofXWDIFXf/CF5rtL9x1OgppSOxZoRvVCdPlt7XCQPcA7dm0U5Th3Bc9qTg
VeU/Gaz6iV7fUKXIoD5NSADpu49aIuAPF4Q+c3D0b8y/pmGpwF1qwBs+fz1UxmuJd2x6TMkCIjSt
Qf6RsoBl1SWXSYl5K6j0sihISdOhayLLsdNyq8pcQPSxROdxKdGUYEfaqDF+kwFsCbUmzlBf/17d
kWVUgLcXvr8wjh9P80pVYsZShwR8eKNQyjdwWDYlnIyz2u8hcp7kc1Rwo+C1cvCbJ+sHfjXDig0S
YBg3sXztb+cCqnCYpKNOAUf7qn+K5GS8KVUHb1F1xD3p9o2T9P/VT5ERh5Vmtw8VDK5AceV636Is
fQdlYbqacXNDTC8OhqNGXQJrHR9g0xY54RMYwABtVMfiD5YYuS9mrJT/nCSYzG15SCtHtvLLyFG3
lDzMpEKAWFarf3sB5mmxMXcccMBoza8HEpN0Hk0m0ymiZQjK39pBokyXDdBfiHKmyPNHH2zMqVYp
ehptRL/q+2XbFtt7pJbAwC3oH3PKSPRX5qfmNCI494lc9Vm4f5qvBWRviSnHgT/iN1dxcr0EncZF
uR4UbMy7zy9f4eDW4lwMsdLFux3XAqgZbYf/aQQcw5PX3E8EN25TVrPkMjkahNQiYTZE4uZKgimh
Gq7Ul72eeBZpZVsUy9BvK839utS5kyr4aXsT6ctxS5mcRZrmZkQdh3aIhWzzl6cGhAmp1x85mzoH
PAnK7GH1I2R4+oREod0yV7lfxHagqONRzRhZuwI3tdPlW7dzuv/nLelO1ixjufnC0mplcp+fQXRV
ucYKF0CGEiPjuxZGNJ0WOkRHY64DjrVRqiiipu2jLvAUwtorA3q7eGrfMSDvyVdzab1AC23YLvK2
2wOIvUo+E+HLR0skdXGVj4VKGvHn+ry/8rek0OTZGL1KQCozoDUllFYqriD2TNdL1RdhOCsHWMrv
Lu9DpGDNSL7+xuAF6GvOqX0IGlmbVa6nKQInMrt8YKN1YmdUNMQUnPeTa6j0eTMG0ea9pcDfGrCO
galjoiXB4F5W44OXummeihyZqT00On4pN2wDk1ln+7Piam9cl52tHzpOnurw/uppVBm/yFNkLN9X
gfJCWbVmDBOGFVYV6I1gChMEtGLC7A9Gn2TXIYQo4RH0rbXIN2yAePpE+sy5o6dyeyhSBAmFFM9c
zOpyhyyvzpOIH5GV58kPpN9zeUdSXfZepInbMpVtctgh2g7KlSlXeDS2mVChFlbUR6/kOGWtEpf6
6di/RGaVkkIrzD0SdLlsdvqxpYG/L3g/p1Meo1z9VaV2RlDg2HNp2rWlpCAVSt4ztmhYDxGKKWfr
G+AnkBLbiZIm5zZCQ63Vs5bHq4Jhh1nXBsH74/rTF75BOVqiAWdWd35rZTcW7vYlRS+OfT1Iycl4
VJHkgzi0+ttVgQTNmHrPmu66i+TB8fizTbWdfbA97b7ichq6hl1mT6aY+gEo3j2M1oQietNYB7Cx
ZYmcleTBd5/a4HRGMMRip8XtfE+N1xgLNfOlO4l0cw2kMSYGW2/Xq/JyiiihU10jTk31GvKCEDJO
uB7u4c3yNeF1Nl9zHvUufpe0jFcAdTqZxIIZCUo70GAT126PBwdtdKHPS4XtvVOUmk7DnHVaoZvb
fnkaHHZY1TohAHPzlZ8zz2JaSufOcuJRMkFM7SH7dOKEoHWYkdUreCifVgib03f7+GogY6dof7Wv
rMAfkxTtR+04W7jx2pEjyFzjzB7hLPNOU3xP6LrVSLdcMBALyjbpXiCZy/WzvreLfL98tfAwTIQp
K3H4XIIXNGM4+NwBQ5Cj/7ZPR2j0N5SN6+Nk1Ha0JyphdC1kCiLGwRa8IH+xF6woxhLWqiI3+axT
LWnVxfaPBW1/YJGqJJMU8y9ysuLB4RWz31j13XKMXiSWmk25kWlyUUUDxwwFmMgFBSZjIXIGUtUq
mu4km8+st8Jr9Ej8p/MnnOixO1Ve/P828d/ENIasiHAeBO+8NVogYUsYXtXr+ZcDlTmh6MHiPaTE
APXdCLz7UW9ttH75hT8r+eIqUcA0/A8baY7nxWh9zb/8BlIX9NcLC6rTNYB42Uie4vR3AWCAhkXw
I42ROiNm2OOvhJu/ygHDyT1Elr9C97InJioI3dvvJbbgZmbzHMkv43ckyGlHDTeNVqfEjzsiY/cn
LIiqERM6THP8/LIPG6jn1zyjDyuwXZUEgS5IZk4bWM8TcjwETeSoHilWvKTqm6CnmwuFMJ0pQjc+
iXnB2xHIGyEmRTCexHQ250pGy9RpGGHfP2UT1vOBRtIGRwsAyKx5cscZweiEt5NGv7XsiQbCVBwl
RPpJXbKGCjUQZ/wfTA1n6oZvvylOpmO72B2tfBQDWn0y7cRb9zUR5tXR/6roVt51qymLYAtpPb4G
Gpdo2hN53tIrcrqDc98k376aahV5rN7Js+RZ9Th/a6yHQEhf6qYeDK2zVH6BTTf11MkT2mN4Q0y/
GWmpnHN3yc6AZisoixDsyqsNxRnnEF4wYKI58Cl3n4UFPiXdIjaoYF5ej0Cx5mVNoLw7rHyosZpM
heOsE/mXRPaG1V0GDEMDhF8fDTZey3H9KJYso98puiL1gBxjwTiozRarJh7is+bBTIcon/xh51+x
P3hmeFfoVeok60FO9XfgY/as6Ksd2dWKkBTeuSmyhZXVvyOuKPbncfA0LHP3nKqrZ7/Rap1fzEkh
M0DmBvTTCPEEQ5hub/HPA4jdAdhoarCYSjJUXXnrT5/JxbvzDd3f+Zmn+9fsrX27p/L4Dku5L5rz
n32RW2M4/AdP/KKviY4fT6BpVe8XVJtHn1Nnjk4EKlJb+uT1gUNRGlaBOymbFKYVQdHo+wmAWnoo
hsZx5Eu9HouKa325TSTyB9yKJccMAume3ou1Py34Wk0RccxcqyS0CXe+fpLoOHSAQC2exGFw1Ag1
4957121mmfKWfjdf0z6GRrRD6sF0eLGQjyNif6C5OWPQ3TW2CvHH60XkT3RPzpxFJQfrEgiwEvIz
tEHKFaxRJV/WjbmguzsIsoHLyQCLsjKHxEUUMSC20XyQqb8rbrN7r5y8DT7JBK9RbDhSOJbNcZyF
OBaHqWgRKEB3lC7iEOywb3k7rkTid1sBYJEfbt8xGr3bo/3tzQRnvwJP7FwZT0orKOPmVvOn0Kr2
lsoMwdktWqT/+b28uBnvgFHVFeXm5pobthz+PtPXks48zOiI96mJ0G6m/YCno+REq822wYIfIk7C
l/ePex8Wi9i4pQbgvBMEIeG6mYZZJxBQz7Lf/ulWD0FLFXe/5p0apUvs2xnEhFudzmTxCjkh1fCp
6MQgcn+yp4eRD8p6BAEFn6XbkpZD7Z9cUXymtvEs4ktOSxgtC5a93evz10U9CJjIDXAs6wzAr2Ny
s7pqXuBpoB6NZTjjw02SpIQ9KcSCCSAJ44ry/Gc/ri5NUG0p6jZ8QKjHaIZK6kC9s7iuzUCOWcT4
0sCHa+JhPfSLZHo5AxYbfEaOy8PuNbLAEVx2tnPf5FZ7FPM5g7BNNPCcoV72yz8paEJd4bQcIfXP
MygvcJVvBEAbMBdt1+9f20xjCY4+IdkGL4xaut9BJym2G2MxFDUJKVdEjgDxHIf7vXWqCmLPi8js
97sPtCvlppelTXlyi6PeRTGCKVQYozke9RMO8bcKS1L2Y+r5OBlwk+PjAXSdzmCtxo9us5tdnZo1
RTr4/SNUo7+E27QiK4z/2lS7z/BxMJGI21ZLxNFG036mHEOvqSgZFPyTPm6TVRXqPNgjaQMy/t3l
Pt/WO2d4L64z5Oeud6YaXHfACPsDPau7uEYnXB3v1FIYhORRPEpcKay5YfZ6eMkxKOFoGtFYUwjD
FgRbEgn0yfLifaP3NvoqouN5A6JPKmHTCyDr1du+hJ/uIUGiDk795lya1V2XwKkXOJJjd6tvvHlN
UFe+2YYEjvKVeuivxVP4S4fTQbrDplxgUokyfCZRqwsfkYzeny/tj4jDA9S03UEXobxr8iipg2jd
YVxG6zd6dGtihFh7F3uIMaxBTNgLeUoOBOPQ0V1Ya/DbRur/t3kp7qVvaESqs8mdAlzi/ABoYLWK
nDZL967J/LHf9zmEDeZKFUejeY5/UZ6p4BlfScK39K3qOwSri0XLYWGiJiB+L4V3/tZGvmKakrY1
vkeffegALl1VnUYnxxbuFqtuMJbDcOQrc35qtRXwkivnCStiekcYZZ7H8OpA1+brhGkGZTtirBDd
IztA9zcH3J+TmVZJj7XZZaSbncPa+LITM2VrhaJmyPLcz0lyEtle6CywMETrSGRolDk5XZsTlgan
/w3SeurAa6HsQihvJp1+2BOnUfnxH3ZRriXBRnV81TRD5oa8rdrHWocDY9LZeG/Y7RlLfX0IKoVl
+9nxxG5QOc+B3NP5eB+671rxEIsFKK4TMy3cU1b99Mb1aHPGfu2gZEA+AFF4izH+VCD59gHrgJ64
nsMpNT7bSmxr+tn+EPM57UjYdFjuTM1AwodsrM1rgRsZYUjC0AKmV3VkGeqKNKhvE/tLSEMEKdDg
pgWJkTr+6sL/WHRarnX0sYpDd5EayeZofiwzcTP3QkzGzkpKv9B5Kj7xQnA4R46RXovBKDD4Ngcj
6Vooet5icRLfa5n9+jY8bYEnT3oG6kymZMFfJmN8WwqqIh59TSMdkPZs6BxlbwTfcNR68xUTVsY8
84qUAIbFEtINc0fkDFn3c40HEyVlir44ewe2jK0xzYp2s8pHUJobOyLOstjiP3rn8I8nAnpKFiXo
T+LYrhsD6YD9KYiTW3bF5waJXozo7od8zauNHmHRrDFsBgKMQhD/j26LorTqt9gU/c5y6gp1wlMe
NBLGc/VNuMaHv+u9+RpCj+MTVAKohX8e0KYJuiWHdSk8Z4KjXuO8jcQYFPJfldCe9Tfkadm/v/7W
DZxQQzaz5XwCk75N6207p1MVRs2c2e5p+fTR7qU9dLtWnizC/6o6mimjA3CF6ZEMt+yg2YmwDF/k
og0C/fYIq7TZ735Or4iqL2cv3AeTCpeb5CyJkbTaxUifmc9YKdvfh2vR02QXhLdHq7GGup+5Mp+v
dZl3A4TRs4F088IMEHjlq21r2STd8LQVSdnQ5u/+qAp9/cU5OXGAMNg25o/GEVLCzt50P3Y7ORGc
MvN8X2CKvpBPgJ52SzeEMBume182RGdr2hRL6S6pHWuzRpmcY0ilNL+wQAxO+MrMxLel9uThMG14
RP52fbmZt7Runc7CZR6NZ0M3xsFCjpy+3KuGrsnqLQKI12CtNSVafZGyPEthxJHpEjeajKwTmP48
fe4IpiaPpuGl5F0sHNpppiAJz0aT0fI8IokxroJD7Aya/PFI8KxuAooL0a82zHSYerthWC5aAUwG
3pDpw0uvsg9nVEAsehZKgbChK18ep0mZOub+xx5d8b18FbIMPYsI6vEtgsUWslVTnQoXvwOl8xBk
+EiaueX8ggGq8IQ10/6CF+6sgNkV4teN8FgIsfpleTKRppQBgXSGZWDdx5YH65jd8j2sjsfxosP7
MpE50v6wcF94cOQzn7SygONHkkNnJ8paB4HuuskJGim7XZHQr2PYRBhsX2rMJWV8l8UPa9hq6Q1O
yCFnHOcexOCegptUZuCVQSFxPhLnlDbF4fjgzyTvpahvepwvFielQ1Mh7bNKTQO0oh6EdWTPKJiB
eHevMjtPULoGzHYPrajF603cAhKv79EF2SeqLhlX2+lHde72cqQm7PrGeOTR/P33RY31Txzn+Ef0
vSb1O8KDmYN4MhLPxlAK4nrDbv+/Xbk33MczepBfiG7ERJ3EzDcS+P4YzSrid46MKDpoIUBEFDvr
P1I1w7Bo3XqD5tu7O19XhjlgQzbwigIXsYZuwGMOw+10aSSOLuQcNSLTsiFDjq+jhFO53UxT7szr
3CkqdmrQD3jhKP9JU3GFaPce8TMs0s7gRk0J+XnT1s81G6eK9wGf1eJPYuBz/wXagMdbYnW1B30y
TmmMhaTFlD3OeGZv9bHnChfRTxT4Fng69P0Gd7Cb3hXb8DJhqigTKzUUzA1tUwOup0e3j9P4vUVq
hu3RXGWrdNtLynhpbWSzrwCrNRy8PhHyaoxVZEQN58DqMKRl6bDHJtcZppNsHjkHrGzI6D3Y5rZX
hPSzk6qEljXsybjhazKkpxl30bVH86NbQZx/WhYGrWsSl9jcUHvQiUdUWzkQPVpsxPZ03YMgTQ+R
bTPSdTuc5jx0NBx8r4JAu0/IihpRzewwrnbxN53K6q/3wXrHECVfrdMioUoc9hMw17zB8vLJ98mS
m31h8+/tMJ4+J/Q7jaP8DWqGlprJbUvido2Ds41qJ/1nQs3bkmRw3WSC9q0qQ6JT4CTkdSytmHww
lmD9n2ObKpoQBBalYzaAsr6EDUCOnmvYKQ3hExPi5321VYPE6rRNqageAdvf5dBdjrJTG0mXnDV1
+xI6EDHJuED4OJNvX81hq0OBNit2Phl/KD9w/xSZAChwNWLKIEyaQJdPSKf16/7ai+zARRRQgBDQ
WfG3DP06BhldQ4mV19bvC9HJHn77KPXwgDEyZumRl/pvxJpqHbY9oPSPVcggCRfMjiB1xfMcx6yt
J/cE3BWx0WVD5qV1pVSmB4jm6amj/f+JLKZ/i1lXUI5/pDqxGRNTEHxxRdlW5H+7AIm6UQhG9e1M
IgXOUgdqvbjSPBgD2GNET/39HD1uFFAUM+D3CEu/L+OsJo+veGaH59HQJ8QccgAxo4ylgcLgm9bQ
swiKLCvMBSB5Flyg5/4vqHRmy6K/3n1WOMZgvhAOxF0bmPXKhepOabM1a8oQW05EnqNQJ/CV0xzd
wTtqUkz9kT18mtJ8l274lPNXtHppx6EYMdAQY3p+ee8QDrXNraQBQVpk4ReX3lT2CSnXRV/76vKQ
BkM0XD3moeWDOVKwOc9pKnVQV0lmUnCp7UV61V9Yq7rfLms6zMDAbRf3R2BpGhjif996vpx6B5NT
rqIOiothrfw85DArp+3ak4hcb8PH3QA8VvM2ruRXxqTjR9lnnb5TzktPwXqe1rVm4NULPHlDo53S
lYUTHDFZp6aEuwMUihbCi9JLrbjDWfcL5GzXp2WCZUzSzblKcvipqNYRRo6NBkL9IPUspL05tOrR
wAbfLadl2SCs5YPngCDHQbvtbYcWVnL9nRQwaY/dG6vof8FJX6k87uXkdRYzZfuMQlxaj47dgTFu
OiSOKbXJISrlFtQML4U8Zw/r91aqL5U57nkFyNHGu6cneIgiZwoXg7uoB3CRgkywRqYS2DTlZLBi
x4kBpghdXD7duViLgC/AS83xrcouq3IAl2SAFhVG91exHL0ZKHRHkvZBVO5ohyfYPnDI1Qy3XKTc
PXbtyl9Gfw/J7mDzvtrbkH57xDTCZo28Gf/UcFZFxT4DFs/N8rzCHp/6FspSe7qdcchR3fiuqCmA
OGlDN2ugk5MwPXo+qbxZYl/w87NNWBIzujhvClOJ6TMrb4RxxTO5BVc/T1J8cS9mFQ6GRL19iiXF
q5aPkDcRb5Fn+Hg6jTxgfvKmTlPsD3ZQUOi/7KCycGdgLV5G4WDHhWt2NcDk3pvpLNQ+71R8EbFE
Cf0bpFtnVTHrfg5buUG1KaB8KIr/AixjLF6Y2MwlBRxt362RwHDSF5R+1sfSFfO3h4QBMlEpBKuW
LikhlmyaVutwVMsDD0xc3ggiIUZ3uZSVWwcauTeIf+HXDrRmJ0JJJC9j/EjkUZ6z6eSnEWhyuNcP
KqJeD+yyBRk6+ddIcJb1jI1xYOujrcVvMpXfT7/rzLAOSwe0snp9sRHVtCSjs2aEiNKElljv8B7M
pjT/d8rb04aU10ka8KFAXwFdid9wkB/SlnE9NtDlcsBDjM20F7A8fgXa5pCQv4+q9K+c1b0p6L0g
Bo2Czc2D+cKj3H9UE6ciRikKS+EXvz5R1dQepRvPhg/secNaC+bdOKhA9PE8LmV4smHAjs3veErr
+zlL6n3OmDYAoNpBzvRly4kHct3A/vbNPCdbMr+GCrrISeJr3yntVxc0lNkjef5fY+EblTKVcCLK
ZlUDbAUkMeSFiMMqvh1mtmDqN4C/CjXljmvw+WKirSbhgVoYHfTuK+LyZ37ECJtVU05R034JKxrx
EUFPd7TDT2m603b6XMUaeIJ9aaNrt0vauf/T2l8eiu4sCz5uAesz7rqqK1uK71lhuJg3kQNOwgkS
uH0vP5tvWP7jq/ZdmGGLYiqPjBUS0aMXbKUBOPm8tOrV18q11SirAXXqxmK2SDFQIM0XgPhH/5cL
dr8ULu1iboMA1LyRQ0EO7saqf2JvWavtzIqrht38Tcj0q0f1TL1wV1GF6KWMT7Zu6lpaimbn6ojT
1cglCm++M21gG6kOoDG+mOv3rINJNKOa+XFAQDMN/+I6BEowzRAS6mizcX2nsU4kEeENV0J6zfvX
g4bqAx1E41Aw/XDePITYzr6yBjaT9830Lckeyx+xdOeWSSucg0/DSstcu2o3v92X0JmD/XD2Y6w6
oHlQNlizVRGlPGExM1qdblbx2PAz8dESUPm/COUvxoxCOiis2XrhNSS/8SeAOiUURi3j62Yub9Ci
Wd4vnQ8qmNNY11r7TqQ5N4onL3dmuH43He3wALGLxNrmvWeZLWkiHbO3phfZEYJ01hxDwS8fBMKH
wT/92g+NIIWK91F7xnBLXHuNe5s5nCGfmFWKj9wxxfnnTVc16pKLCamPu+1QzifozRPv2lWGq6Q0
DsmWO6TpWrmI78nYNaCnxP+uhUGTyg29tbXsUAuEGpnHrN28boNZJQ6y5C40a+1t0WLrk0tFA94l
meO4TqWFXQkKxThiWwfkATh0TKI0T9In9ejEixJk10GeNpaPO3QqIgDiBnJ8/Hy26BWDTtd6q5wq
DS1JZfJc5877a4X+ERI/fV387TTL0KHw5gMztPZPJh6hcy/p3dOqyzXLG5GPGwahXu7XWXyMt/3F
PijbFeEvzDs/ESKUi8HwDtsV/U5bvUcbvvJ8nGqO8zB06seuQiHiaCmNWxUWH3OIdH9EsJW3fumg
Li65kcy5HLrCsr/XbkacyR3nVURs5DSK+sOYr59OdnXewkPqddJHxl79ThL+OA+sY9R3XuqGQkWt
x84zsyvou/qUxdsFLEG1WP9gnbkirPrJaZ52sqVh+dLldKWyM8rkc7I+ei2rV4Heop/2zwJvX0tq
cGyyp6VLBiNllUz/B5f6xhGtWvRmObA1I1GP14G/sSgMKgSLXyI0oOd4s4PlnVyNPwb8aZtGKwMD
csmf9w2BZVGbFDZ+R74iq00/wF6QxaFSFR4NibvigcEV4zb0wCUasto4X7sMQl3YUckWhe1ZZhh2
C4QMOyxJ0dMo0Oq1Bszj3SBXK+jrHzqTPYYQballUyMeVvj6u1cW70iFDDQEl8C+mivsztxxEnHF
ORFhkIPqvA9kZ6tz0Veo2axpMWsMkf1z9OceF0jMPFt/0CKGDUP24LogGTTCDBpuIqeL3mbPAvx8
Sr7gETbKEs75B0lAjmPUVpFOKeOJKTn2Ih4ODFNPYcenYxoG14KBbTs+B01tLKjvNJo+K81szXTo
taIet9PhSxP4tCDUrB6Yxz7DMDKMaB6FY6muwJUFfGoO7XKRfwZ5O0biVt0bpJuovxA5nVEmP2li
GiCD3Pcpmjf1zM9PE2vxGFoGkv7eDtwaeJEIudVBMqm5mzuy6xVEZscmEm0LbdCbEbz7JblfquLd
G5OYxXYZ4hDI+ejz+DZEGcxuFdKy36icHpLltR3gXFGj4nxvIpDHeiV4sc0aEauvAkOQHEQ8Pr3e
iDIx/7S3+bps3wVMOSHFChsTUYvqRKQ2x9u8lHrGDuwrese++H3q6ToI+4sUZmgQR3Vb0x8KDrXc
GpVnQJNK4gblRj7uonlURZqXGdQTpA9Af7G1FQY2451cMB9sRaNLQvagjm6anJ7ylzXOAbBtUQ/U
UTcM7SGzfwl9e1Wdc+TaHdIR3A99ktSZ+yK49ebGr5Rgb7JF0tvkwGiBYF5ezP3ccrVPRL+n1MTO
8UoekqwFMiUgYiS9kBVxAUOtdYFqBSADcobfy2QstuTFH/KCM+10GgoTdeFmjHIhwQ2837Mk3YSY
YShzlH5boxDuWoSX/UDipkA1jt5/w/Mm0GUnlNver260rwvooAMRGTanYllysp2lz0mjc2G0Lqc2
VjySI/y7rpZJ6wV13nfGywRkpLLVb2fch9FtunriF0vTifneFjXuOns4hIZWiKkRPcILoKqbii6v
1myEy0PnzTR2qdMrlpicK98h+0bKYJ54sCUcAnyLxGnZeuO7J98tyWNHNQnl0/pU5tWtafzZwQnb
Tpz2YhIIwLHlxJhnZ7RwzwGQ3H1acxO5XoPuGWaqj5SbjNxLiJYTUp7BuHSPE0czZC619urTadFW
DDcv3Q1RZqJk1TfcIgcyAQebzSB/N7S4tOL2imPT5Fk4NmerSbhcSRGFxvDC0elLkGL3b/6cephH
B+rygbr2nfq786Fwxy+nqfPDYu1U7J3tKWJtL3yR5jwTvy+ZnI/q5TEjEs5botoNwLZhv5hTh7Zz
IX4YnfjybgTIZNqOeiyYhZbvFOcpFmNcTIKieYyhxfMxbObA1FNoZjhGi8WZXUPEWDTm4ISnej8C
enbMrN8NJXbDAtmoQHC6sUXxpTfowiouuTDuhIQzMPyLntTALV/zStMQMGyl+ic9mjPGm43SD2jq
d+bn7NMncZVAbrEqAh1VuMdmdKy10RtwF/Zb8hR6QBXEVXsZFwr49VtYRa8PaHTVmMR8EZLcW9Vb
mIvxLdoAUeNGacCWPPrES6+0E0ZSNfIo9QOJeB0yJnsLNbXJUpNi5pYp7wy7+ctj1EyE795Stlgk
GdWsteZhmb9gYaXE65+R8dBPhMA9yvpFWHT6jPm0dMlqRWnBtmshOjrV+/syxE9ewwFKILLDpZ5m
jx1DVnM/p9Boiun0LucMDufhzBGUYAwuK/ra/2FvEU5ZkCCv6uyOc1Gw5ByYGp/gE1DySUUFNcDq
JO3EyfmW0IFZIlmjxkx9vflCdByCBHpu02x0zE5rWYFtl4UUD7KK9pFy/Y5pbZqnHhiRR7YChtWo
ZbQcr7Gscu7GBWHxPFFKXfpaQAWNhQhEDIRRbq2tq7nWstYJHeHPr9iZraSkpsevhwY6TZdXVLPt
f3F8oq4L64+dKzUBJOMGUKC/mNjKIzjH+r85KGpsUbvaJH9i9xU49bXot8rVg7CXxEr6E9XrzgDQ
Qm7Mvu+5t62LzF7egB+v/gXjXRFedAHLd+igFFGyBgmXSm/+bmc72uod4Yi1TzmxTu/ytFyrWAK/
owoI9rEEBPWdenlLIeiJePOXBBre5PegKo0FG2CG5nn3butZTKaYBzkWljd//PRvwtr6VYWwa1s+
zCarfYDXPCQfiB3VA+qNn1IhdjzSmO0uk526rJfHqztKKsvZTzll+4TpX6FuOb+3BYD7C7gO46rI
yBq+xeDVj20KQj9jJuN+Ka19mcxt5X34RhoBI2JVp0sderjj2kaaOsDnZIjupRty7PYzknpbYe+k
kQVHH44Gp6r93qdGo7L5cEMdASyA7yh4eJLmLHyPpkk+6fmyxC+GIf1m8cQdN/2zxye+74BsXz+u
0TJeTyUiUDCJoHas46SyWM4CC4Uy+GahrMOvi6JDt9Gi3LKfPyVs1EVvOyPobUdd98E1eNiL/bgk
r1169kWqrSWd8v57WrJjvsbszLaPVB2u/FCafvrsw1+k2es/ltKmNNrFK7XMLDjPOpwxD5lREoV6
l8zO77Ho81PSLUUTpMhl/3choPISWAWi26Qv+xvePbIACouBOTO538Q4W84uqAR/CIzsKp14vpCp
U3hyj/WnBJ0FiJtME3tUpS3EP/eHVrWtBvR+lr53CykJvp7gCWnkPFL3viPksmIgGFORb9zcTlrG
c4WXE15bjLNjLoLIDP2OodJR/JIAM/vJV6BTa6bCNBHLipxkRxARuVSdttI2BbKJ9K+2TyGo46fc
1KnvFAtHkeKgmD2JjMvrV5TD7gxu00dfr/Gl3YbwyJi5rBMUZER5YDzjPtE2CblhLJ2IGYDCRsLg
Mo/D45MDNCG+IBn9UcPxqibPmbtI2+vDD4+XZG4Q7hqWUQMvTIPufNPV2lGUK9sIPPFwTj9svBGq
EOc2c3lw9A4IhPHJtQFVUkxbi+9eR/B0Imh4noHFOLFxIdMTBy9J12i4cQfqg1pvFsvqPA7JI9cf
kHFhqU2fUUx6MnYgCki79i99Plf9M5YSMnUbAUTabjHYMVaUvoDSKVpaRr7IxwpjtZpPasdOCdgi
+Xto+xy4Q9lmKIVPnSC9KSdzAerklwr2tWEfz6eHxwCl8CwdgxCJutAgPqWZlNjg9oy+PtOpRzDT
iX1IqWHiJ1vM4m+TPomTeUSuH+iInmkCcxkvXII7EnjM5z3LFsM/MbZUeFs+uIU3ErWdXOc2wgoD
Za62GzwFoCxOTPrb4Izij86B1li5mrvfVaC1GijSj2uuKqC6HyQFubX03eIUrLtbOvCXpv+DuFQb
6ZvhEkbSLp2dQEtZFouNRCWPWVydo+titHNTCHatOJO77Vt3Fg6zrkTHKkF/VQo7nfTWJgxSCeSL
R1yUrzJGKIBMV6SYqDB/mb4Om5DzfTU4AkePcITPCDLb83yxBvZ3D9slK97LDoQofrHIv7wQN6Om
DIiCp7yDq9E0jjsqHx84Su195Dy6tkgwsDdK+Qi7yMqxw2D70MqxNzkGHjN0cyVwsscAITglzEw+
aCl2Oap7QVT42Pm5NqhZR1w5KzLn9mimeySEje2qkSumwLTfpRH60dJTz4kL6WIRj0qLmjVJ1LKu
s9YOy1jeE16DTQlo6YPwh3Dhub1x5Z3IU/j3LexHHn1PEI9HPAGTAW/qgW3yqiszMvEpUjgcnN78
AIXPIOth+2dorlkaBt2EYYIG1tO/DYZ09W+Qt9QngsDtbed/Z4rQGbotQC0hDIOshgkAxBToKuso
NASQVXRtOENT9pxPOiiOk2Xg5R2qQD/aweFoU+x1+9F0iy1gf8X7tZkBKTvdiS2hp9hAGmlSBnr1
TOtB1jNN7pzIHm3ElOcQrRe1ODGpDBpO/do1XVG8LbeGxx3wfqwBmNhVe2a8nbszIpmT/c0P3hy8
Yav6TMCH9I2Gd5brpkp+tHev795iFr09yJFZ0EGxdQnivnGXEfoH9nK3RlcxdKLddvDXRMfyLgsS
BIR/oMfB7gXBUnDzcWVK2vLKKgs74qTmHayPpQ8eyu85o6zwN0koKlwfwP7Y+yhj64UpTR1vNQgz
7KUtVCmnCtGYxDkggmH+Wgxkv4K8D35NvYtjyweO5g0bGqG/Litmsg2/bRqy47m2SUjrQgZYy/6b
LBjJZmXjC3xvqkL0TayDFgcmNzfXXhfw+C5rnedoq5RjH1zrgjg3obv7q5V/Rj6VcE9S6u+Dd5bc
3hEI3CjLSatR5Rf8CwryjM3o/NUed+YQCib2NFU4bKs3sPW7NWOSMSmBDv6qIXawJuL7bnFkxopQ
liGU8HuQ5zEC9a6I8O4mmDgUaMmx+xI9jhG0nKWEO7hGJI/vTT25vwocV6hii60ZjtNxtTUPhx88
bCLjx6Gsoxt118aJ39Yn4fzyVqZMaEbJqUY0ENJs00WTanGBpjSwY7J2vWxhCwm181Szs7SKk+Y/
B5jmPHOrP/NhOHIDAESSrZe4e8IExEsLrxF0jrcWfTgwBiqu6UrC33k5wUDWGpGTDZzo5/+n4L5H
rC/Rvli0lWiYcToj/I3VucIPRE75NBVr5wiUyHgTZMz4pY1eQtg1FNvBRhSNKtT+JEZZXnCm4JSW
wpVotC1osC2vH/XSQPRkwXBjlmYbEt1I+DZNYHW6GemM8yDxWHxwrv/MADuf3fI63viTBce3qLgk
h+XyRCquZWqhNm0b97o/XnsEsMV93Mar3RmPeCF9gvRgWuG36lmfM/0cfMjYw62Kfilb9b7eMUR/
Zlh89W0f6+TmkyHFl4mwjJhQkdOQGiiBvv41RxXj+MujvbqoI9r2iI1D/FxIK9p6zTJLgB03KvfQ
rFeO84eKgYtZ+mSaa+wSt4vnTzF5L9yCW+hWyR9buJvWROCQ9QEIct1hbcK7dZJOvJdudc+WgwY8
vVrjbQJ4Rs9C3cVW/wKUU0Ml7oCHRr1U8XIbO3v2ZIEMjZoEknrZBvP9+h+1nAwepe5/FxWNnX+L
7SkDNb92GkDGJ8ZA9l46ttpdzyAemrquQbDHCPbhJtifMlAVg5P7I5uvyXtXlraxPMQX9VFIHaT0
057z6Nng5VwSt97m4Yryu3xYsuaM2N1zEM87MDgu41YO+QgDWcG4o33nLuCr0+qSHKXFUBaPT+tn
u2E8ArE6FW1mDnZaC0myxyi0sQHaXaoWRhXwf80CY/vLkWE7A2CA1N8NB/CDWmtZOcd3tf/mEg7C
X3xSS5v2FxCpKv32VWsL7MiaZyq+VHu96k8+I4jNKLpGUzVKrIj2JG4fsp1aUfC7Lb6clXgl3ast
FenAGCFl+2F2lxVXjTO6BP3O877mfOUrevM2MwwuVH4Lk4T5qOb/I1IPiCye2aQNAaQJJQdEN6LO
TIt1lVT/1a83yD8X0B/j0z3gjblvYJmUHakBpl4TtBbXsaPG1QVJ2ZufrTuv/rigqYWySI3sTlBG
cV3Fm7BtzLwaKvC0NmePe+sYCsAWDVaSFdnVGj/m3BOUEYgRcg1IsvcCWysUbTazaMpQvrW4sOOo
Bt4tBeFAWaGBUk+ut0aBq1I+UDBMYd4EzC9ZZUiiAg32uVbAAsLu7NHuscgZbnS0b183RSR3yRg6
2Lz27vXTdVtFPsotL9Xril6FP3Ti0EwrDGoRGvD7etmG4jc7UXvwUM85xjv74R7o2RNGHqj/mONI
JDeZ7wZnuFwVO2x3gQrVsWP9NEahnMjH71oCqvw7s+bcps2Di8aLap5nlZ3/lYr/KUuW4zRm1gZs
4ZKGVKCvRhgALWecOR0yu7yoSnTtsJTYP1rBd1yr+21SWB1lOojobr39QKvGnNegwuxtmsTv0Ins
RFXuydtD447HuO74fVDCKMpeZdiNQMWyTH2Xx1ijRC1MlUHz9Lh0hpci4Dn/KoC91u6lCdWdy6qN
57moA1etqaqwwDQj+nQ3010YAa2k3zKa4Lz0suZ7MXFKIQc6SUZMlFdxDj771ccJTF0NNs01oUOf
AwTXuw39zCRios0QwSUs92jkgpjdeRMZZ3nU5lfu9Yxp7eHYx54Kunw2Qr79Nc5X4UIUt4VNJG8k
FYX70MXXXAvNIoQj4U1eFfBLBTWL9Eqi5XVw4PT+vZjdc+PPCtD5LxfJraeH3OULgamXUiU0HLka
sh4XcrWxYEYB4FiYqzk53Dyo1+1BNpStz9XjLyJFdaRKVHDdH6bUlgdKzv5hFh+h1LX/Z3yta3CA
/EX2OcnQf+l+srdntxB8kXgjl1xrPFNXfCyVjBDlZCdpZMRilIHkf1GPpGuaWqsel98WHK+LV3ZA
AKMi+JQl9CvKyKOUEsLmfvPjurvq7JJGMjpsnDTruXffF9cKEuuRf+AP+X0YfE5xJz7kGyVVn1KD
cxdV6qKH8pEmAKnsf0hFUFnIOilut+i91/34+gDo/5p6Wac10SCuC8O+Yao1BiUPMU+hXVllJKu4
p+TVebkYYxQ68AfOVhq7/IwmV9fNYJ/6hSGmNyyW/7IYaDmfmEpLxohvm0p+cxFvLiJc/4r3yHW2
DLWwXKIxtHdr4ij6eGmQ3KT6Tg0rvZhMgVNyXEcY3dWqAoXxcZTFO1exUl/PgvF/4Z1FFJ/dE4t6
6gOex1F+nvWK+XQbZ5KhM8vShARciuduNLHjWcwvtLc3WpCKcg0xCwUvu0qNXgSjUoyyHo00v9ix
+0WhA/sNrLNrppxEH2muc9k12LeXY/N751SbGBeqSkIzgnlH+gACkdbzoAdN8nvrTwO6GRCmOJ9o
BCBfvtbPRPWQeW2umJTaNGT+Fm/Ur+G+7WUjGk/FPSrsJ+Yhf2w40em4Iot4lAHVx3SLJ8KML5W2
hDwcyNiwBGKzTfwjM+bNnFJupYMJ9bJa34Umv63XcH8WSYarMS6QS1GSJ3rkEwqRANJ0mUOP/lW4
wFPII9FsCCYX3ovc5eA9JAooRq9qaw1liGWTgaW5xwNDGEIZkBQi3gGNeN74HlWhr5fAoybjcTeT
2cygZm7njuXW3094FhsctLrMXzV/Oe/ISmRh+ZXI3FDmuH/WHsRG2ZYDcM8X+y8lGGdSg8Es810W
UuX9hKb5mTT+DOewXgtV7lEhqwgi1dHH8EXMcoO0j+uWjxbtNJe+4x+40PcKN97qNblPj7LeSkSG
VLM6KTjAGf+U7kCleY/TtSIyYF0kM1KrydUtQrSdY0d78JIDZeO39PQQ6v/+fVdxWjAuxY8yieLF
gA2bZqVhkpJx6LqhT1LEnSgdfJ1qc1RScnwNAAuvmJPd7LfrS+mEYLyw8ez9vfbDMQhUCmFnx/va
pTkSGzYl028iP/YyNxOIG4l50adJKG6ufwT9ZXld71025kVgmtoTz9Glpv6IA5dNBglsSbyop+U+
4JKNpO/EbjYWnigTfK5BKu7vwtRoHtRlJv6KGCO6oUq7/yPluIuEeFbP5VD6Pti4fFVIot3ctvHg
Hzp08U8IS9rC6NzjgNmTZ+qUy55WmwnVMdho/AGvzySuqusj2RTc3QRop5UCuFv0oaxJzumaqOVg
oKZBr4kx8QMohiPix8elouK7aDLGXz6NZpZSDdIDw3FcKl3bcumHl6Sgi3BJRdHUKaBFwT5jLYGv
hVdiKFH1mPjRQYrv8yxlYffMGFvEl81/TjcWpv8RLGqQ8N6SCML01za6RnKDbzeeivURON9sANQ3
3T4rnDIi4tDUpL07PDXS30MCiXv+TvGVy49iqMuq8xL4R/Nl9y2EsWn6aPvawjEUIV2IJyIUMN1r
x64R0G2s+vecbZbmgxqgoTtAqnagcflQicp6ijn109Jp+AfVOrwkzg0GI6wX44bz8DSFXKBdH6TD
XOn0zt3OeMzkt80p2nMxgwZpo98OzAu6k8dTi6tJBQ5SUTYBEczA7DhmNzvgL1n5EmUI9KclYnRP
wMYr0GQC9pHFjDIJtP9G1ufxoNlOfFreuAcJv4g+qeEjDA0cXxDz2t4mF0+dg90eEavobNymIsje
B505gOlpp8r4u/xA9BjosCFF/umQ5Lvi/U71heJiN7lNpeeUtlkyB2HUFxf25NB3X9MwHacVb4VZ
SMS0TWyMq34dlyNkiJgcCs0Kouz0kxiZq0Si/5E1kY7ZzJli7OSYCkRRxjSdFfwDkTAN9o51kPYv
2NrpMoQhHn0eRDBkNmaVMYQQEvIKpgVFgpaYLAhuJ7M1xKxXx3K7Nhz+lgfZep+oLyXM8gcRoag2
N/Lh+MgUIAx5TsFH5pCFinCdHLU7DiTRSNmYwdK2oFSgCpYDRfvFoBzBefro3En+MZA/6xSirj5F
Kyp3STSH+s/CQhdRfYzmBSkQPsFuz/y+vkyXqZPLDGAKmyfvAYIoctfT47wGevPd44LFTAQ//cQD
4VMZTthx3cnysnBhbesS0JGlSD33BUcB0jzLzdBFK4dg/u98u8samaLUdi39mJn1cQ5z8rrAafG0
+CMsKHpeRKrgvgnQVOO1OxgtvG+By4E1tpZE/+RfVD1k6Z8RE0pNGH8vHvPPY9TR9INXAI7w2uOL
m2CU0mWtug4rIqSvde52kQN8cNWslbSTrufLSOqNQIJWzNNHlO6CcgJHYPivswyxcarcESF6bxEa
7kgmqATzLEGNXpJR9PBnrpXmi9o5Q6R33BOLy6RXSK0dUtMStbD/iPHWGZ1tYcaT+gOvaL8YNrWx
dtCFcEOZPYITNH5lrS6nUBbtzLBNVt6NLeIbFApft8lZidSk1HYu4PWQcuGTjw3iTXMdoX9si2dt
uprXKW5sFZI6lWPYLqEseUYrpYVMKGpCLeLDW5JC87zh0TJrqSrYG8gyWYZMoCXdlODPXQVia9dS
E2jEmNGtUrJsTHQp1rNCpNkWyEzh5MmhW0wKSm7+RY9m/XpBGwwVG5N2gakub5IkPR2LCeecV4ih
rGuFCxt2oMy2BSIr20LA0UT3D9YwIrzOgY15+75eAtTrfIdVjYtBP4URebVLJLul4rqntut12/mU
IpKVcpyDf844b6uBoGAKDIvyuse7Ca+uiZa/onH+6KoVCEW/FUOgryP21skN7yhDi9Hy0mSorYwC
YrJZ4AcvTuP+R9vj22eYvPafIhFeK9n0rXrIvOdaYYNVV/pImYEXu7vQVJPi/dljvSkVlb1cf81C
xzIValiheSG+ddXsy4RYXJCs1ga6JGYGfTr/O/PeoQhzKq0+Q48SKw+OO4EqCUTqNbrnfqJIyvKg
XxImpx4XTwQIbWtPgIF2viX9UO1wAX1oMdBG+VnSQQdP3B2U6c/Qy4Pq5xmaf/tH89SmDezbUOPw
cYH43wz9PNOhmSKKvGTq5qFd78mdHD/J4qjPQkbyHowfdgh9ZqWlVYkOsW0MgLPO5BSw+pvVZFDi
xFYj0b1h1nRKPA1sHB2ticsP4uUddnhDTRia/x8yjarOBx+63GoFJIJEY0W6uP6/btmrwJnmH8MF
tzQ8OpO5TsMTqSf0OUSPhpUrqNTbNraRGMlhV2fDyn2R6dudm+BLaG2xRQ4Z9kDapYzD6vY/ocTx
8WG9zP/FsC7CGMcB/n99/bwew0zf34kOWEluoHVBIivhw5FSQ1d4R5nt4z4wLB1mbAwPaXpjZtZb
ESVHFV5kiRGhmW5tmZJlJdCzMxea1ps7ddRue1XMWcD/fa9+c5Ur27odTwKlq7grxaOyL/hBtKEP
nJTfhFeqFyIMGmwvKBL3uW8oJqKY00iVFyX6x9wOvgqyC9liBWV11X7i2zHZx+RUSb9HQ6DHAXiY
bQhgzPf0hl2bzv4r/s7bGOtkK6OqKum1FG5NCmVTkCWQBjo0+45ErYK9Ki1Agu6YxkkKEJ3T1WK/
C3JqGz40O/EZuurmEyfdJR8f4WXO7/L/V/h7fJizjwZ8ajoFx1yqJeXzfEbAE4T0zPjd/T/2sZ+D
X1dsPEJw63cvW76oMv0rTB+jMaT4Sw7SCuVtaperOsTILHRMqXFgE1Ayd6v5gHKXzbyFlSQjk7Bj
WFa4zSO8krlv3gB80EbSWjgOrIChwP+mfk0/2ExrJwBXQUIsmCWp/e0FuqqCKFzwWgn8GPRE3PGi
jWGNK/FeyRBktOJbVyqz2xGscjMzEIqF8i6FvHHBeEYLKPPDMImXr/yBHdXPDTNINyigh4CQltui
SFLjdiW0HGy4DwF9DWKuHblE4ojmdanlipIOd10p0qTkwDWd3xhA7jMp8Bt1lH2mFowi0J7ky28B
h0C+ZYeqHvSPGWHyTh++iT2AXzN9OvXzgOWzi5lTs0RUDVR/lZDWDnF2KFGLloev1RSFMKBbhTIe
RHv6J71L8MHCy1WXcMo/6Rzb3t2qyzvfmqwChohDRdrmxdFhO/+iRWlyJyY5ukD1i9W/IXrSVcef
8ZnqPw36ozLhQj0J+B3t0Fw8b9KAIiECAAmBhLZ/Tpb842KtY6poJ4l4lfuRngvMbyJzHCm7fXsa
OrpzhY9ELPcElkfm5DBs5LEYY43jG0jkq3m9ccA5b+uLsMxBxT6XWGOPPg9zBd+n09srYH99bMRa
LZ74nkL2UmvgSEPuLsh7a/eMp6/q8dD0jiyWPK5OScIMERFuZanJBlZBvUcreE2Sx+ayNNQgZakx
8t8oSZvyh23pqnTnad5o4xDuUvxnP4+484VpGAFs0tI8S/6gSDCCz0eMQpqVIy3JD0YSWJp9Sx4E
38YDZl3qrtqljO0fOYkrorK2Uy7AIMrnU/OymSNPSm+QYAX3pb6ewWsfydIWRZ0h/o2SrgOe6ZoA
FdgnRG3xoCdhB1qmqUe9/X4x38o8vj4GdlAEgcmfwCjto1teSn5N2Mv/Qd64eMY433vNGw4bd+5v
07+dP9QNXRNGICX0bozmNcD1I5dsQnnDbffb5LcE/Y0lPIWzBHi/jQRwUi5z5Q0wPK5HuqPMYvqy
F3sofDjhKUswhERbn9x/3AJBrgrTcc8DAD0Rrn4Hgb0Lp/smEGgllFyYiM0HoDhhlBEia+P8nelh
iniy9U1qgzl1sRIx1w9adSN5bcz1BCejPxaxsd/BfCdLxjh+Wg7CFBGvl3LHe5o7m0Eaapv41ub1
GTzTwDhwGbXBbdnaWhqtcnZAVaoTwNbT5KF8+S2GePtgG4iVzNYAF/uX2smj2n/2v7i5ve86RT16
QSRuqMp8bqz9t3sjmy/IG5BsFCZf1FhuJJ8R95TgdvCAeBP5foEJuV+uQsPRQ82kdfsmaltO+onj
phY5W3rCSvIvsmB8viITaqFit7hE95Q7wdJ4XJEPPjHVwIEOkT+jifCPJdyZrcwL/ELuQ7Dj8RvB
8vkcirNEHnRcAXQd+XI1aEr9Rno2BzTDEoO4PmVoyZ7xYGr6CPEwY9+hllIoDzKO9hxVdvFeiXeJ
oEyAXFJFD426yssvLLlX0H/QP4n89t3sTX8BZW4p3hTKUqE7vj3AzBtHsofAr/MBjvYEHNATlY94
NQxTy0fjJKR7OhY/IdEae2U1HlfY5nkeuJXoaxyVnAjrVY14lFu6syWI1uZO4q44b/WCWoPGyi1f
a4KCXuAZYxIPuLfB5m3mvKCj21qtGOQKA4Ecjlc8eUnE3vbhY+Kt5LhsbM6ukFftom1PflNdNljE
q+U4IUp6JzhxJOIH4FWuW8oulesWUrrIOa+266DoqAprdXpfLXyXUq70yc5eTunEc3nNO3zjvKX7
jM1O/OcWpyotQYMKV0NNOlkqRzzA0YxZOXFuGHrIZyWyRf8oFY6lecYT6cZTHpR22XWyNp1qoteo
lvE/fK7U7EmuIx7hiljIOP+udoVzJBVsNMEQ1CBnNFhMy1BlsQlc1y3d6P4uNY2fFvWAzfP93EX5
UNY5n5xDZGF5Xr6X5cu3PofippFOzLG6bnOx+qC/RjTX6qGbKvQACJ87kvQFAz37N3Q9PK9fhs5t
E9EGJo+aUwb9Xtdme5S9BcEd5Cdd6Hsg0nv5tK0G8tqO4yxh97R+t9hpms/b4V5Tws8vlo7o4+rA
57wBIMJnzRnjuHDNy5+HRYkk//4SAMJhOujmOpeQ0tLISJn+HzzDz1WvcaOHg3rWN38HvGD1b/Du
uxrAiPWER7GhFfmTGQqr+LNK5IbweEe1OWVHirbgPc2iNGfEIaFw+vmxofMt9FsFw0+0U78LkeHQ
3wt5npiJg1MF54KSpqdFRM79y8elxAeXYjWnie4jSgAs8aF//MXHQt6iSmIhprLdkIDHTJzejuK3
DYzOPX4V6OjCQNt5p/fD8iNLls2lmlCTYYHGOzZkvpcndTLsJBmYRZEe/6EALXSE4QsdXzNyHEc4
SJ+rSWLBJ3EAZJ6rfyFVtPIwYTEK7A5gm6E4jwOHkhMTPsP3brv1BX5ChkOdPwO7pcxXtWTPa6Iw
cCfhTUgZ+OZyEi5Eh/+Zz1aXFu1isXQ8Z5xrTrLxRrCV5jrfX4HvwVDSmM6wDjkBlvY8DDRJOpqU
r76kpqModYj+VWJxSz5mhSvI/6MtucKE8TRjrLYbv4Z8wh+iapo69nRb6Ay4u973Brs0OjV+moSW
KexKpOUMttwATMIvAj/tg+Mu5nzLx0vUvDMg3PwvOo3YgmfENv/TvZ8cnZvN/iXSwNPiizTgbNEC
Ukn8VeLvUD6pSbUJahCwXDVPOJBJpjDzp19o/6mAIDhdGKoPWS+VUeLoT7zT4TckW6bwx+2d6do8
MdtbRh1biGpntIfQrQcKglSgMyxEFyTXFlgKr6mKcA3KYIqRUecumXxbeNBPcmsMRN1M240uDJ41
tUq4nNoF6e5gte76n7LGhvtZI4aIJ24CogF6Tc/No3j3oAdoElmCSViWYzzOWygsQfzHsZBrmO4G
8LU9s3wMb6aDNUUWzdpUZlba5bzBOJZjPx7DkcAqqSz5fsNA5UeR2U6YZFldEWNP6mlRZ+4r6Nbs
rP0mGwnRKQcPngFf7jDAZ00uvhLl6O4z1FRLo9bl3aG7kbeEWFaCkXP5txe3YieUHgN0/EWpGTbK
YCv0hqw82JERdz5Z9HVGhrnNBq7bNZbGdmMNXU8ykGqZ9eA7NECk2uW+TVd8bOV/u5cgIQn2svZ9
RKlEoWairmzW/sgrc+wNYKgo0fUSZQiYDALP7tpG4ljSpGnU25k9heJuEHv4tYx6M2Ju5Q4d6ER7
94+TrbD85lGuFafxXEUafZoiBCx3XtSAcyTSh0+5M1GPIofzbOMMsTCdAj8REHX72m0qoHt8LV/Q
MelXfkQyGSREB7wzASkScHae9B0+tdh2vt77NsSkRv6Hb+fcKYUK71hL9waLMQ6hNbm8qlpJvLsB
cDdJbE9qQ3o81gPZb/K5tqGbNw1DcXOjRYbjrHoLQbygNAxTzEmXFY7hBb/uwzGeKSD01BW9J3QF
72nW2E8MMi7gpW+u2MV6IOilYuzWoZ01WkTNyTb8org4pyQFvYwIE6k4a8eq5C5JEjOkL/lkhv22
Y+uaHRZQXdrSP4pURTzwuqm90qjzr/xoN+W74RptjzvCuHMS+KTrvNe1AuOWtafT+Wzu/6B5zv1o
1fkMSN3cuzCnkCubKUCEZVCQMkxHx9ZbBbFKWY/7RLwnZMQ/L8waOUEHTw+unofErGvzbG5SlnKv
ySPU0MGD62J2WBdrrpnMNNBHZDx4G7uzyV/SXVAmLEeUFP2W6e2dS1lF4xT93znNlCFXGLORHxXU
7jEDGc192+gIwhBvE0TxexDkgFSp4E+yZvKnixP7LgsstN1R8OgISxGkrOjF7li5lCZDf8lQFc1Z
JQv2nBYvtxotOpikm5uZjHBhVWkv/khQlBZ+9uDd+78fRycgnCTo7O+x3BHaFzYy4zK7mlWGJgJ8
9e+ASFLy36rMGBcf2rXhFLcA68L9FLJ43uWKRAJC7ylGGDlAnt85ONjL85/UV5QO2SfiZAC4fIPF
qIQaxEG3EKBBxNeUHYqGz+c9S0RjIqrt8YsPNjmd5PfBD8uVaGJj1yYW4N3nNuHoDpNyR7MnYGt8
5nozmePIhpUZdSuUYm1F5XkwzGmkudS8RjFpj+CTJu/m6u7j/n3wmGQRSRICUV7OQo5//0CnJV8/
VEO79CnmbiLq385iVGdqyokpPcJM9gJvM6Hu+S4A+KQ677uM8epb+WteOzMLZFSRKVWjyvFzuUbB
yTY14d9/bTrXuTPvdJm/WU/a5FVvGTj9/miyMnzUohBSrv0+gKxdtoB1jbtABo5SY0JZrlU/nUl6
jRA1WkgyJuSpGWkrmGlBwFe1WaJFbk2ZoTgkSewxQO6HdwjHZPV4IPNMA8Js8Xz0bdM+cLQ5paez
uQIxNGGk399UXfpvHyehIJPQLqWBYhXxPjqSXLytEB+vucW83sR6snc/GNm6uUvyamHMxAQhvsKD
56JKPq+iJsym4g4HDBn+6UADBhVeLq/HS/FOCg4KRQRJWTaPV/wvp1tIx8LTzw73EMxzxRg9iqgI
H0RCALWpu3U0K15Gql1B9BirIggwiztLQWSTdy+uD839lIG14LhOiNLm8KFU/Ku1GaH5LzaKq44e
mHgpaEiK7Wn7YDxl1yo80xjiV99tp3OqF6YWaOKY+XsclwhyMR5UxTB4Y905eXn3JYVo3awSZFyV
4hE0cmBAvB7DTDUvdcKyf4cvgS+tDNHpj8dXwl2iEVwbfKf6nhHAqkr/IgC7YG7Gkj1+ijew9nTf
qFtLlTc+vI/+wzfAfuta7sVBOQW78r1toTYGNz/5szbPcifS7jcyNXrwpShMWEqx5pX8XuMR0Ewn
lXN/qP+PgyHkshviuNJqUowgfUaXn3hSFfSE20lb475ltN5NGBlDTkj6E8uEvbNWBB8ReE9ZtcmQ
kK0bJkpXAK3cRB2i15ouuYKYvto0SlPhUIPmcGGqI4iAA5fZc0AgGv1pIuhVPLSD3kSrbyFqDmVF
MCStzBTXJgAH2ZPIb+xxdgTwHcXMzjqlvEy0hkwt/kq3ygXhkoWUXZziFWmGMQ4FPQ9ZNjsJumYa
+q3e04Xf5Gjjisduu/XL31O3Ip3ELqmBj0UsuZMJVWAPkampnm8sy6/rak8z150Ke2hdUynKwLyi
DJ/xEkpIOeQIIs3qAf1TKytNTfulsKyhZAyN3W010ZIpl5Hud0jW2MNcqIeMDuwaBouzfs1j1an1
1bIOLQ7itsdzN5g29NCSnfBPfndB6lUBLLc7WP7NARV86cVvk0mLkHBxvVlKS47Xsn1/GO4zaqkY
bMI8+EDTCwKC9XV70IHMSQy0jnMWgSs5D4j3tRnnq7ET5G/TjbUZLa4n85KPJmjYGqMLn+2Bwv6t
bVqBSSkbgwrkf6tI6dQW0l/kSqqYfAR4XbmVjoNWBo/zSsOm8/YX3oovAtYrsK8rhTfhe7gr0c/8
3s6JsUSo8aN7lIML7xKlZh0xJDPrsI0mos2AoL9KsFavjgS7zEuy8FoS1Ty+WE1iM9YfB46X/a/u
EUMJBc6zVgnfsX2y5dukOO1mWgsENdjY2Kyfc5l2cFbNpWiPkxtXKSOwri0r7NAN/zngtd13rd7s
pF98m8Y1UKbeM5jKefDi37675ZlEHONGbIsAtcy+E2IbRs5cUBHAWFmpuQZUnyqUHBxErSHKP9zJ
vnwbtMDnD9q8RrBoQ8CiieHST4Fyu31vU+2CnnilqjeEV7BEpgJ+MmCizSElH9bz5fDU01PLtXD7
XXou+7ogEkNUl4hW80rJJiOxCuIyXXi8EGAS2X4fGO3o0+yzjGnAhPeRG7gAbglPhWYgIieCbr4/
Dk9l5L+kV8J1TzEOKCpI54BsiOvxJPz9YEg0TCiJTrIjF7iKSy/GmxrsBCo+LCSFRpUvVCwFMUxU
zJ8waNnEY9ANe8BfW0CfPA+xGIwlew3NaiQdsxoL6+6+jEpfdTU3KWHyCzTRIwQ9EhEFKd4Xije0
5/wYB+nlHbMte1XtMN+e0v2nkGmymXH4zlENO7ju+aFOgir+EnvHKsHMWVF3xZCMdI8i1JCKJaJ6
/eusl61lVHH9iRaDfTnaEd3w0YW1UPETvOp0i3He7l5gQlbtxRWOIahS6MhH4aWJpg27Aq5K60oK
+KzSfHuR7l2SJe6dflmxbW8mmL60Jp6cweQqCAEvxMRnqQmO8VwEwsexmmaYic+Ox0A81X2keyWe
FyyrN9sdoqHGjka0kKOvKYLXeTwtXdE+y8veMoQi4dAPmfezZ/L8Tj7FW84LaitxUddeUcEHIIjZ
MH6ZP26t2SoxADSvpaYLJ2r53lpVyaOS6cmUyayv14uw3PqmmeDjAhBBq8vkOBgCh0+ftTyUaZZ0
On2a/lakc3sEKNWJ6fQZZlHLTQQ4Q3R2n8oQuQHBJQRRcmryj2CFPZ9f1iuxN0OUtP0CNsvvSXwC
64t4Ga1Et7r/xRwOMFXVkMODgNSf8eWxRcg0gakE7HxS+xQVxeApz29YNqMWD/QUm1W8XgmlGM0S
spycYQ6p3p2+myx916Vt6JnNTey4wwo6KwLQ5mxZm660x4UJN7Q1SgnnUmQZ/VfZe6EqwpcblmHD
M+Z3RyAGnucm4LZ6qw/e4FZAvtgk5m+uDePNzuegwk3ZAcgR04Yq+K+i18Cuu1i3QtrOzMfiv4TG
b62KOa5P6UsRSZlrGtsGlHi6tVBddtg+9Hs6nMTj11zyAlaMtwqgvrpbY1aq0AHFpPieYbpwSNPx
uEE7YvUmowwODELeDqcHItPzr9k/ygtw3iMOxUP+4PuVmHiOGRRlKWb0xImF7IHr1UkJiaWrNmn4
BC072rMz+E/MdeL+l/cmJsHAIjGPEoYH3I+jiGBlKvEuu+lwoMrbaoN5nXbQG13NvNTpxeOt0POF
ubgbqWJ+vwEtepplkD6dPc9bnZ3Og0KuQ6IBZWbJKqPPY7NEZfyRQUSQkw075HN24vlUvhsjXvsv
TJxR6NnhXmvduOS1O7A99OuP5FdblVamnYQaLUrfXMI69fF8r7JOgUvRgYXsqNbXBW9+7tEaHusw
3NRxBMmpz3EUG0E0EQbyXuhifzc26IexvqhMKcEP5mIo16P+8rREpO0kcsD6+t9Yajv/cPagytc1
5PNvahvTnIO4yjry3M5C+a0ePSiTIn95ItvO7iFTURFjfaRFFTuFTV7cQIbhNZtaQF0FJwqfcKh1
tT5JnkjOmUBl+iXqCP+y+ZPWaeHF6EyXLViMWistJbnjmsX+ntZSYKEJbl/XNPHrqOOND0t/dXUc
RVs9PoAmgYLyQOvQj8sO+7lmMpwGuVvlATHX1qUsK5hR7VoecS+EET2l/Y6P+LIxVsHOkAcS6vbJ
BopS93rohevJJqxe0h5BWtQ5j3XpaqWzkwAm2P+3alnehCH9TozbbXzI/fMyggLpgFtbjHnSGr6H
TMlHcHu6TmUK4JbKr4VneR5EA/qravDoGNl+E/GlzNkI0g/h9bsBi6ZqH2nCjkKiC8EZXJhQ0CJ2
fzXilr2c7jP64Q5bKjU7toNYvLgAPIHlYpFPham91yQhVdW+FQQsua3ziZQVbEEOV6RlYPrQwwmH
vP9p2X24CTAUpJZpAhx6onFJHAnWclZGcrYOO8D+5uPxLMHYcZWrlZOXw8xFCJAH2qzs6ZRqI98K
nwEzBzZ66j/OmZ8RrePPh7wPl8NSKdszPmTaS931PX+GieXApTI7m4HEzbZJzdxyvkSEH9P7nBGO
Q3shLXzVmhQP24RyScqUe895JdYZOSKfsLz0s2MV6cvfVH18w2vw/3mcGHuHSXUNn00iyre0cdup
dRNthuehl7EdUUcPhZF8UQpclVfkc3j4P4a8hzVMT2B6nhOiay/qgPB2VIhBw67Dq6YIz7vtj8fk
tWFqc4XeDkfvRaRNAQP+/CPl5kkiXv5VPBvpXtgyR2ZnMqdevxZmmAiM5fPtgNuK2amtL2/fe9gS
IJ7OhBnRiq2zoiqN5sDd/aVOhJYgHrqyZAaXn4biBTmn7pr/QuDNGzayyMgDcuwY3qBLDtR6iDz1
at32QPllN80dQ5/NGBgOgdacfIz5mqJsRuU2YsrxVnw1k5hwieSjs3XbvfT1Xd9qr0letYG9sCs8
jqkl1oPrYvtoKDSwiO2v4+l97uQ4PNtayZj5DzqJ997bT6d7xoPj/f0GAVIagFiLPVZeltu2q7MK
QgvqunXhTpbwSmSB89o6NLojR4ZyGD6QMX/j3SMITPnWa8XRk/dNijPTzE86Ugy6TpeEgqBL8dJI
9CuDzyu09HFd4e3LBRBOi5RRpn45JmjmO88EtiNbaG41kKcbziacv1DqpD/+Fm9b3l3wEK8ROY+7
ZNIiQOWPf3r8R/QOQxFetUfrfRyy7E/lV/9di9mGa2DHW9WG3JtJXQs/NgGnRBuftseWV5/pb8TC
tSW/G5Tma/68FeSlhF/6x/F03F/2NlKPD5LJlrK+ZcPnTtrICWCf+YirFyaKwYd0ZMIZjMaVCg4L
JWKIgggkTeeoBdXnOuNgPlYSip/wmBW3dTRyg2oue+mbwZcxEMFKRc81WQV0JvsguKj0Zkq+2UEO
1beUjnwVdi/wZCLbv3YQVclwwHh3hmH64Df0sBl05Lj2n1A4kEjVxJuL+7815H0PBVSYKSroJvfv
QstKnqSOPH1JXqtwHnHSaKP4I1Ip1PQpO28UCJRih6KqQGe2aSfVembc1aH0Lt5A5zfltXb++cyn
MIVteHYF7pPBliKuyM3QxFCx88d9MNRcGewIxsF/7YMMukUtRBQKaYlge8cg1DmsLJF8G+S8a2ZZ
3Ouffr0AOwjKRjC+QtdQIl+I6bVVs3NWqi+wwZ9K28XjzRXhMtuOawsAiRbKGThyhA72H5yfaN5Q
xBSSQq5ApMNyKfA8s7PCFx2J/kS+I+zfn8+P7NhCvmBe5aXM/zTCbr3uIv9ND/zJJs9n4YYNXBUP
9zlSeU7aop5Prc6sbuSHB1TEZAyX+AosgSxetWNipy198Wr3ne62XMNrrO3TmEGD1I5NJFkueyPF
KE2dngXo/1NKjmr/BItaDwSL/u0F2FxXnV7usw0ziTVZtCIX5DlTczlBdbqZCnZgVzuxNYgMZjCJ
eDBKFfvZX1nLYO+SRJi76IyTtFNAmQ4aDN+JihSjDk221tsPGPT4FvceoXI7YErsNoUAFi8MzTXi
LRHJhEgZFSk+a2Mu+n1lCjW+xerOjHEZW2gP7ILa/ZFs/0wOgokQScfSzaT/EXiDIkxPVoEbAQ72
QFjIcATp8s0yU9UfI2McBVWlbC/ETIq4PFntgEnrZBL1EmK6jP1Ik2xFnVDOKJ+pSN1iKjX0R1d7
kn8FfGivUopBeoGb8OriMjEWSnDELhyKqo5/BuHhuKMQkJ3fhhRH++1h4DgNkvumHYG11mwFoLvK
2LEQqOwffPMcuajGzRjEokHQAO/mxrBUbsnoWX4mYvvmRLBz6RDe/BV9huiFIn6MjAMGAph2A9ow
dz+WUrvLSQNNpdlAGeQ+M696+Q3mlcBMkdyxH/DxGEGDfT31OI0XiyBSVq8Kze6zB0p/TOB6kIPW
Gt1zjgVobTlT89cj0eXXxaMPdF9Wz8mqhNV2DqMciNaxr6AOABYeE5nvRy2UKWRRti0vi3Purnus
KeEuUQ8hHZ8TOfXL+90P4G2VLBr1WYV1Rh1DRAApaV1OjaeuijvtZDA4xOymuQVB6k4AoYPp6/kr
oGE+pF0FNPhu1NhzxbMT50eJ8s3Eev+dmFd0x3kvGrC/QmiRxRyDG22PTeYWIX0iYaZlh6Ifn3LN
7kq624DxVG/QBmwFgGV29GM4EONf0FK4H7Wj/BTl3qKqXzw+gSgTHTn1UitgbBNNSlBJvCOkm/Pv
u+FwFCwHyyxvnfvdKoIUJjP2y4c6VRvfE9lE7uvXcK31aOOklM7jgSbWDLR4rX71CwEIUjYj17Z+
vFXtMH+n6Gdy512VO+GldjbW6Wls4zI3Wv4u4itxr05MTZ+/RsBRngBoDYJrPS/6lYoEithAJzKv
HjGsMwG48tAJuV/aq1fRqdh2wcEvyjGnV1G17Kcw/AmGAce73v/rZu0ejQWRpFT878TCRbfsxI+B
cwHPb0G2TmlSPST/DbeD8Eq2Nk7FqLqNYZq7U839viOtijgXoexXVvLWqfKxPe/GzSqTQTSDJSUt
MxnhwDoy7s3efnmDh4WvYYQCj2C4r2+MOYEPmVUtJL1ua/zlfjNfvwIpGb5ALEFnvBtrzBK5L5ZP
NfxWkndh3BA2GYUpk+SmrW/oug9/7c63mMs7h7Y3lnjKDzCdcQYsNgI6ojNmgevgdXtt69L218Hq
QLlVU5psA/Ha8Igw2EldhP9stMAlvTPY/CKR7nFKaKkiiEzymdghlVn5TvaEHk95/TvHdr/aYFuE
VJGx/OblG1RvuFDEXnPqzvuRN17V1EJQVXWf4rlpwVsbgLyXi8NANVpB5scpWOeep50OCtZOzu66
COm14HLvoIx8n/JoVDN4CL5YS5Il4jq4O/u0ySJFYHsKbCJUpjRYEoV9ZCrZGtpftRR2ZFGCKtPc
xSFKX2+Z25H7pMv7lgSglI8Pfq9AwH2TcHWCxlMUFXtWyb5WSRwRJDtgIMqOVfQB/pixyqYIj5Ie
fagF05moCYijY5FrbL6sPcDiID2Q7AfJMQHytZAIOQhtdi2Db6IAmguNlzBXyOo8Bjcmw06t3qBV
MIciMsLBh1rvr1OJQfZ9BcUnfFdvln3IFdvah1hNGjNcZCjqtExYqc5VPPfs9moG61nSXXqumhJm
2kZ9Stf5HZivKD6UTFk2ZXfG2khU4LvC8iPiWSYhpcnJcgR+Gxv3rijwQv0ccS27Ni2BFhv+W1Xp
0A14unAOEtL+6V5HRh+eqoaSfdLSx5C2VzcD8iS4JeCGGU39GopPejrGuiDmnAhy9ZPA1C5ri0dM
R7E8yzf7rnFKLels1cUsb6tPh7QlLuyeSB8Lq7AonVnE+Uvp9ndwObQQ4cmOmFY6dg8VuOvvUMqH
plxkKgn696OtZG2ZW40ct79YOj+bQAuE50+qYqdfkQuaMyzdLdNxYf8t2H28sn3C3OXqGxf5ov/Y
dS4hJVgtwSKH8uPpkw6bjp5QUmA7x3Wso4xd4c9hkhrglmU/GoHinvpxMK1xlc0PdGYcMwGDq91k
MT87gCS64VKWrMaW6ZMfsZPwLglhn6k5psQxYsTlmEsBacEe5+dzDtFmWQJofaZZgKRvr2+q/raf
sseEapBUjHHreC2aPU7EtscbUzBDywrI0uFl4TCQadPZNu8h0YvDcZZl87smj/W4Fx3vhH8Jqaqh
GldKpPBwJ+Cy+MX9qcbrypSKpeVX8G15KmugUzLtSVeVSOGWRn1qH0mzSaQbeybBVavtNXHjsoAc
XQgGyzaHoblGQBfJzZWwu9ByapFfmU0K6Uwv8NuZD8ZSEQGdVEfw1dGLY90GpS9CI9rPkxRW+16E
yw+hwonCqXUh5cXuguY5eOkVs4iVRvEH6oJFmmu1OsUwQviWQc0Iu1TUUjCe8TMU3yBynJU3BoUl
Zb7e9xrJHX0B5C1GCpEDiqaE/FvS7EqElJQ9hbTpMd31skPAkXMlOH9TDF0Rt53TcFDKlLejd1yi
NTgou0qz1cogFvTSfYr5bPUCTIY5XBRStUEvRteK/HxtlcWTchilKbcPuYc6hicXFXUBO/Irqyeo
HCVw9VsPkEmkC9+JMRGmO9gIF/UkO8/9EbqGEql0dU+lLlXy/HEJBNGF+uajjHQQgufiUns4R8dL
JTMFDtTwLmUQavysNawYfQacSmeLhlBRVJMCArDueHZYAwuDDMCPWHss/dAFd6W62aGPVBEIQYi+
+32ODgRUrouJP1CB27lwjaoattS9BKfMXmWa/RIlyMJwnIOzEyh3m1wZ13oGaxZP/ESbmGzfosPB
2PHDaybWHoct3z6WQufLqwXc7bgWT507lsm9hLtxb6zXCiqbK6sV/Tzabv7LU6L3UWzuw3wnXb9Z
SLPf3+IGMK5zcNX4/6DviP19HKoXciDPXqQArRmSSCs0Gubwh5Yld32APYl/4l7Ya7SSlbteRKoE
7Rbk1s5+yCkTZ71CXQ+EQrLgLlO2DPb+miO0hv5oryeHuzZcx6kCHDfOx//2GKwwDjhFdh+sIVCb
FIcc8hbZ+BkPfo04CHs85NQYAJ4yAQCB8pI+QEVX81jtZ/EQXEdBen2R2C9zaAe42CzwV5lM+LrI
W+tVRX3qFen0GAy1t1S2XdOR7HmXtxAKWEoQlie5P40XaLV7Ie1Jqi/8aYK3CPHueVFD5sXbX+/A
CYDkiYSy5JTDraG1G733O1IR3tLnje97YyJ6n1twrCHZTw0K1Rd83B8Y76PgDtTeq5Iha1a++W+X
HYHV4fYq668hQqyXU0aBURssWosw9CrgVgZ/Q3M3MnsZb3dkkuM5GlYpYFkX0bcx/e6/6muvCp2B
gjFc9Ldw8jz+LXpE67XceTyuTBUx7T5t3DE3WLCXRXRdU/9Jo/giDoJvW5AwKdJeYhmRa+s9R6XF
IVeG9Ejc3kq3tCrJ842lK1UUd1c721q9Mcpm8SDzHC4sf004qFG8tW27e8rpNlwHoGL6NL0dleRm
oaaVe9DZrYJgYcRhTwwbEzaiHDeQvABeYwv0vPz6R+ljQH2CIKY9Y/3JtxO40LERZyh5FOI1OqTC
pC+hbXNkoV/hx2pLSgNtgyLE5I8m5W4pYMc5PWEnqWPGmK9DIjVhRYYhoMjWTRAE9NNQyUvKUeHN
eXl6iogJ5XriVqQrK8zGy2s2ikKVTQ54f8+atXL6BMqez9slx5fiMM0cwKYXG+Yb6vIpSznx5gwW
+8bqIMShhlkruAeCe0uqgUipyxygBDZmgzEHD5qCEodBCdzJ6W6Slk9dLKzPOs/7hmH4PuGx/+U0
qecXzre3RCb7as4zimUjTpuBFuEjkgW23Me0yT1mMaPWqZ6CVBvlHftcYum7KVou2Q4+IkFPpAE9
k5elqSA79ag3D5jNHtzSxF32YMd22Bu1ORdR3NeT2O7VhjXa4Zo0CPAKZ7OyTIWuWTv4MeuwhUio
o7NFOZX1NhuvrgFbSX97NzAFHO0i3UtXIMjlwpaexShdR+/aJN8uzAajgwbi1J+axUcali1ZPlMz
O3pLX5KOLjriorRiqmv8Hso39KIICfRsV4KAV0PRRRyGsLAe/CWzo1NPhWjhxcJDK0qDgKUfToc6
H44pvrbBnWiLj44sG/HToUMkoZV8ehSuTACSDGCkjrTFNdnAWUwxVkZ+QgKNGdNaxnVvQ+rWUlX6
eNHTY54sQYBPaSRPR6YIEYh+BQs1ssgqSHwJqnn3h77P3tsyGKGxifYLNCpXUaQDLG3bsVmmplHF
s9pEOw7vuMCTcrDI5TEVjxXfdU3sGx2BJQqqmwoOML5tqI65g24xa7yKuJ8tQ0Mfi1GnWZ54QdIc
VOSqLV88rziCCh3GKJVkoAJM2kDBlA61SgorGVkqbFxp5dRbsaq7ZaNs2e0XsUH3RD4kIqlzZIr6
CGJS/ZcZLaZLM2W2psSWPqlK/7ZJ4Sor8dgtkXKMP91La9mDpyiQEHHivTzwi8pCgMhznAu1HJ1q
Nymko4QqPDjlljg2PQAbMFIOPfdtzyaNWqTSNOshQK4szbROyy1PvmZi0uxMQsAMi5ITekVkzXJ0
ZX1rkr39ZMriD8F1kg7lKxGYMkMisyjIzqLDQjLZKKLtDg0gbwJLe8HSoJpGSZC5bnAXGiBufaKv
TWl4eMCl62m78RQbkbijRBMlHBfPRNUalI2jV7xdM9XXppwREGQpyvcdOaFBTpP0JlKR4PNQHjUb
X1X/ZR4XvCDakFJHl2iStcoG7Jnf2lMWK1UaFf1vCc1hQVnUoWoVhMEzsfpOrmn9LtXTeut1VYn3
KAxhw4eRMZVK4SU5SzUK1XbE59pOubkEW+qeBkFC7uJ7JPiiLDZI2U00o2SRdZ+TeWSy0n4Q9pts
c17ABc75uRe1BbG3iQyeopYkjZnSAp7DCfrsDQ6H6LooL8/c4+qBn/HzvsMArV8TzJEYhV3LLzJB
WpgDFrC7/IvbO95sXXGFPZ+INGN1Qxqk+SDktWp+cqz/+M2UlesGtAdfAxHVYuYdG/bCpUEEbOtP
Ifq5tpRtMRR+a6ddvFj5CmxpIy87hYvCbvTiwPtdeyFQET/oYx3RUZy0DX8aYg1UPPE/2C7IbhxL
J3yzWn6v54ta2X5aAziKuYSm6OnNKhe8ap4+nSa20GqwfEouUBjjc8WdOL70S7QW8AWHT1xiLnjd
q4c4glrmQm5ivhM080a1nKncz4VVUpi3ITg55TnHHLtzC1xQxWLdB9tawimIZvUkny0GaQp12xR9
5ImIlipFwh/gfS7MyZGPyjXpgGTcEJlIkcS4Rqa1tiR4AkV8HYL0pmxFyplk1DYdBRGYGgQtp0Wx
vJrni7PVXO558EQVFm1xnsm82HDaZwYHj2Op0yZDABPjaPn6Dwjbiw/KRLZgb5Xr/D+OcHzn4dqQ
JrrxHUIgrGcuzhV7nK6oR23S/tDAcdlAMZMIZCc0G8BYztkkWQjOkamJSBgKd912xbUcsWwyfy9W
QFBrjc7z8HI6if05NvU380Lr9Z5QlcsIraa8hsw0ylbFsHfTT05HUa2cC56a8nsLl0DQNzu0uKdm
v3qdvRBbHqf4Rfv9hwGa9jUndvOgkR9tXTxAgGv/hrmoLJG8NxjIFnHb7de+x18bbBjmlhzIkHg1
jwfqLlVTUZAQlTg1LZj+qpuouBZmyotHBbZ84rD0Nt7rhEzsCJfX/R18ITObETMML3oO485BavTD
E3tjCbRRi8gXJUwF9F4Xj7IxMGLWKSu0ewnbgG3/pehn6U0Xda/6KHbgNYOg4vlK1DLB0I8+bz18
2zvQ1hIOSQK5gc7kTjYhmj0CU8GsmY00TCyzTR+2r7YmT6DXgWZ2EEOETnrZE5jrVgkI5gFl8SDy
krlc4xgDi87TFfTYgYzw+12C89fyHKoxvNNfbxoDLHLjYyBAz5iYh8hQBGuW5lz7Og2nY2QluA1N
h6KWl/tshF+hQd1lj1fa8pYPrHI249ScP9S30+RxfE5iwvdDpXD5jDCnTEvfcmqFX2GeIoDVOpkJ
2hy6uroY0R1EielzTRwrqPDVBPOJz3XT6YB/5TRPDYtFU3xGIUHBXbiceO4XL4al/OgmlYJIFQ5+
7J0ZTPo6o3I72ITs6AS4FDzx9kGkme/yqBP1Az0SHf4JDWjbareZXDP0rZKPFScQ1w8KlGVTcMPj
Cc5ChpOnCs41WoB3TAW9YihNZKBJ6gZYpiJsSES8UM26XbDAZxyT9/bLffSEtPpTd5DvOdh/j0Nr
u5TeMAMfb0bO9sTDk25Sv/W9RTdoeHqL7/iWnqxXX1MwttybA3foqbpnvoTbTI8uVAfCTsNmva/h
nlGGEshdVpwzAH7YSmP4h+F3Rc3eu7i0f2BjboVLpj75IT3iXbcDNd2JW4dsxtkmAXykhjNqRKCr
hfZFJyIql+2JESw4rDNuyiakBalv0KqjUkQuTnbMriWw71q3Sxpe5XNqvKfbpri+m9SFrTndOzNg
toLTwMrUonmhHGbOts+SXzkp30AIVIxtVNnD1GXw7u5sufiDPtUuj6PQuU8Hr9LgIWGIeTuZC/AZ
pjJpYsj5y4hk4aDMywUhDGItjAf66x+84/xll9ziu52SPEfytvBIRIIbZVFajR4KV3mnbZMCHz8m
Evlk4ZbVlTZ+NTQresWo7iPl7vKfNgvDV6g9U92sM4STUNQd93au3q7soI8HclE3korSyMy6Jr27
zint5qoY6d+CUqGvzYobP+/hJ5V4o2bKaDVU/809x3etuR8xZW1dMixFalG+VXkd0C2TA4Ym3Ray
R/Rxsk07HlVWYuO/GW+r3zDjX36z0ruOFZW88nenkyr6Pk9Lb13DIvn6DBTPnH6YOg8/tvy04FMe
ddCE2OxNS8h8Z7SwBO9QzmJOXxJIXxEXtNkspWS8/VQuJye5+NdtMbq5c05Lk3gNhAbGoelG1iwr
B5+Tn8ubTf6rJ3hQcX7W6435+KrUCpvnENHHojBmSu4qWeGzHScHgn/1TwDY7X5X+weLrMcaG3Z4
AHlYCAjDMelrufg5MVFJjHapeAMEe8KA5RdDL7RgJaoc0T2BrjxwRCA4xHTtskeMdYzAYF/l3++l
JvL00VEKyz1DcF/OWVMZu1CJWAG0Rry5usmSisRoLsfqWosYlgNBL2DzjTOs4X5+scFH4lL8CZzG
eIDoUlamjmuti2jfpCFpLVk0pjGojmhxyQ4DTZpBwmyDpOwmWLxoPDIuM0VM0c7b2fC3SH0rpLWB
TFEV9PY1HO+1a7qDbqgi5w/6nBXp73bvE/2a2lxu59GYo2zMOYgLfeHy0K9sNUeirI6EiBfsTuXq
Tuuu1ePPC3XCh5qdNMm67Xesnh45mk3+JQoSsZ8YigOH4g1plY0jDwXJp5fqdoPoWTfLWv3OR3KR
XuKcYxZczUa4M6M4d9TB4hDsY/YM0luH2CfnOcQrQU5ZvHrkyO+BuqQKE82yJX2q/i5HovmI/w9J
kwiUr60mwAr/rhrxDIieb4HRi08S5kG6YPslceic1OOoXSezBnvMvFnXvwFpQT2IAnKl/Ch7th8/
wSycqU7wo+BepJqiRCzLAggAbUgsRflbyBcFD8zYZFPxP9lLXshIyNLsw5RdZeHiXDMt2DASb3wG
ZL4jtL+7Jxo+5ZEzoCyMJkyKw4mbb/lxnXPIfZV3HK/nxZQ1aZvlPNU6P+0AZBKuf2jmli/HEplz
Dk3wj1ohd7Fj2iMXqi1cMdUjD34yr3lcTKDZ5IwTzJfdQ18122kXz8xVP9avQZBV8rQsATGW+X0y
jwjzRAP+na32YobVKPqpIfFhAGW5o9wv/SvOWVe4r4xOY+2rb0f9WP/bd5FCZ7zpiShXaeVODiMu
96LE7we+w3mCpkwOuhGsblLPQJ0WIU+nEOcjWTp6uULBlsskLk774jiK2S1OkPwccu4OxY8P1T18
SHip9Zc9r9KKH5AQ72qDD1WGW1w1GW0Z1rWTqPsm/Nae3heOVRRxHJkqPdY6QnrGANc9nfg5FHCD
SCKAiACmzh5YaRDglb2qxNjKr2s23Q9GMtyJIWoV4+Ki7CRcTAaTdvYsADtUz2O7LW2ucqpMsOPg
geFOunp6I0Fu9i5X1zYZDU42OSO8bHkhMgl3yXfCrDhG/iG/o/LSKKPxw5PAaVpVqQd+5aOlXUdg
MkX6rmXCFEdjhTrBSZEfD9g7d2/6JDF5xt4A7OflVj7xlKlOvF5EOJL+dd+HodU3wpL+58Rf/jO6
q0hl0tgaJFsSM0q3GWCb0Aob17mhtjoBPeddjtJqQGSoqUSsW2lJUnhiupUfl/UUez/HuyiJMw5q
WrHzGN9Ap1Fxr3JKDrJpAve15Vp2vRJuTnZgI/IO01Rirri208NRavXh/FxnrU/2JeqsWB+PsTOa
PzHd+g5Dz94kgH4VvbVCKUjXoxhpzuTC4SXE6HC8cFyuy76YfekSJtFzFjGnm9rIbUNl/TOxArKA
Rp0BpfuA7bBfbuROmgcn5944a2CuNHSbXx5WXL1C3RHF6A9qdDavJHmjN6lyAci0frKZMYxwDtiQ
api+NPNMChev+c79hF5fLf/KPX5y0Qnik+YUUVL4GMRV6k/jibFS5fW96YpqEYFo+3JRHu9qDh0o
SmduxZiaPS/SfnVlW65G+KDFQlfugBjUi93dlptWPypKRVrDnCWPsJ099OIK/XI6e7mtzJU88SNp
UjKtvmalmher98F/7NN1V0Uy5BQjHAGmLXHAPpW7o+knaU0xU2awGimgVctP7XqFrPkYbUw/DF5R
bVKYEbM98sdJnnxIz8axMh2wBQ1m8M2BJFgWmlFK+wEO9Q/EQHYpuhjvWp8l/4iAOBd9A0aXTHM9
GUmiYJko7qkVaCShBSHo4a6ttIfrKMNIP+iTF3KTp4sHj+ig0wS5Ja8HmEovXAzZUMF/8jc9d7Js
y7f+J+GNnbbaNJ1y3NwBtyZJffoyyxSlGTas08BVYD6X2+zPSnqlXpM42g0zaktQHcRBihB/i4q+
ZmF3Es5t2UxLeCO20O5xohrw7s9gtGDpr2qDjlGisFnEoKY2ETEjKJdH54B6r+tkXkP+qlImwsv7
k1ZWLl/6QHzMYOKRdqT8tXmJM2hkojqf/88czUbWcDj7W+3380XBXckqQ8oHeNvwRA3S+vXiSUG/
QfEHa3rKeyrHDQnRE+TGqQoAvVOnT3Sy8Eimaci2/9Qochw7TdoFrrTW0Fx09EFtsOjO2AGzvE0U
s5NNrIpDpxwxDifjcXU9XkX3xiFjrLO4B5/9KB8VjJUDXpCIh88RLxAczKl1ZZBudc9xsHhJTfdk
/zDaI0gu2QiVcAarBHiejUrkU2wm08UWUwZhAjI1s8zNRfboSh38wtiibqXevoPFAeIlyceEusWf
f6Wsc2s+nfjME1Pg2wu9Y6bM/lLud9DLw+oWc7CFsTeW2ytWkOPEvBauCLNIBOkebKdBsFc4A7Yd
BZ/sPMG8A2Jhwn9RCshDe8D61KNJjKEHpxFNwdhYjsVkGqyNivdIy4V80b4poPTU8zTmcfTxJcgN
jtBuH3qOCavdroNrneScJj48WTa7n52O6AClWhP7sEXPqjN4GSOTnxSR/V0b+oolEXbSEjNT5xZN
y/n+Qz8W1CbnPHVAHx4PUUqvc85vmvhc3L7x0VIgT4yV5unLxTIPa0sDDXgjBlg72g3hsiypLnqe
d6RwM4rs3ChQRQgoT1s0ofZ7c8DixIOAlclhhjC32UHZiJy1FLNJnMN/IKCqJtIi9QAb8u+/38Vg
HwVA7lZkuJ3cWixJTX8J6RDeB3MSL+X7SvJUpGVwwJ3nVMbgluyZGJU3MpW/cD5/7TkeYRDMzFaT
xoxbAGfCAOrCtvlrCT11eyli+OHEB88oNuxghwPqWis/kbrt4vGmE+2C7Yf1kLt3E6jIU3/4SANW
QcNO8JXMPBKq6AYBj4IWNExNEjJEsc9nP9tHUdDDcjE+fp/tBjNAK9iBdZcyGROWyiJ2Y2GsxEmg
knrp+EJzjRktthqb6BlO+FEdhU7xdCaNAQMOjCcevsSwxfNbPXS6brd5eYGJol6Yo7sKYjHUPunO
XEYVgWPg9lTc6+mjH2D3tVJ3/eShyOXW5yL7jP0ppCTQXHNBnKw3G7BS8vZftKT0JwjKmLpaZ1SG
QR9KAmOLiMnjhlzIDsCiwSPbK65CgZsG3+qE6s04I/egN2LT869la0K5zhiekvrtmqQfOGRQji13
GsRA6uobbgP7EcC7FXcDYjEx2Mg1m+6YyI4infsnaZ7+NFPtAh6qwX10jXzxyMiDd6UVUZixgiiB
M3J6+8D9ZZpNLx5Sdlg5gACuxyf1vp7pu2zOcYUpcvf9Z7QooiqSYkW+qsHCwcrgY/LzbwAg7x1S
s72cAADFnpzmseaT2ZW8BBxHRPxhXKe6wpBvzgmbY/qiuHj4HqBmpp0An6rn28f9Gqi/hbYntFF2
VLbbdJUW2BccfZYrQ/YN7IupRzhkaXh9UDPzgFW6m3AFoIkFUTBacDXf5hCRkdhcm0k6eJanuGcE
jffR3EPBm6B1b7w3W94CsFiSTjDH5J3QTCHnsvPTGS4H9IyQ0813td+3RzuyFhL+hGBGS4gOcLaV
lV5tgq1wmWwVQynwCjFWM3I9RafXvKN63s/P1NSpsquFjfUuY9MAsYJ2iahE+gsPMAc6teSgURtS
/Dq5gGQSKLEgTnlNBwoS6YZYwj3lY0ZW8f3nBBO03ry988M0duT34tVWuchKp3it6vGf9NlCpaVV
1PmPXtRl8Be2L+XTsxOn54D19P1YQwGV8sh/FdArGmeVcp9d9T29tfqW/VcIw845lozgFtHv9RR/
NaJq5QL2YOA+jK+FBjXSByzUxE85mXi6MY60AQM8y0oCGfKBDquw7NAJlptkTsRUx8gzz05nPv60
93Fo4csu/6T/qBkNfa+cP8vUzhIr8xuqD27FIqhQBjCRN6+eKU5p/G/BkSDOfQ39YOMUWu1aam6L
eN5rU0H30G2Rf8tnq56Mf8vFdiwy7BkuMvt5ZMortHCJQQhxSSZ9WRK/Mepv5eA6awMBkihteij4
+Ge/wK297c/gLgAeVrSFj5kewXMyoLGDg3Fa/a/eUT7lrzJ2KlFjJjk2pnczrlXnrbEGGQg/65eV
W5ohE6RVOY/74RnBNdqC0bR7a6TpTxL99BerOdOEhpTEE5MyGTQ3LyixfRaeUvWtgadmHEsDQjMl
sgVsnObAOh2TgbrRTFESinKfLlShGGLsKnkWp8euryaI31XQfVo89iUTMWfhImK6/yk/UKmiSCFU
4qpHoE2IxSf062Ha2BXJXR5o1SjZyUbtPi4AWMGLyz7jiisvlXZw5SEgtjdPDB7c82dSfVc23or2
XWD127o3BNGd2LPzA/S5iWfah+cURoN5tk5WLyhV+zwPDNiTlrrIjTlgSfhGZ8CP2W7jcxNgDUE9
ZuLl/RSkLLdGNyw50Y554a9wYhcmjcXdU85mBo/nTJuv4o9x2pMPHR/xh+Rcl32z3R41Fl1Pfgm/
Hpjc+0eWnQn2NfkSeFddRwBsvRCJ4InPJ6lrWYY1RI0XEsUuo+ZvMuOJxPvA72PPdbCdqwnnq8e7
1lWfyN1uhrUuvlPkgI0ojCi+aEI44tDX2D7SMu8P8pvebV2ITxLLTF+mVw+SluNfaNRck4LLEkfJ
3Du6Vsb8dT14p3X6n/nXpYd8qGYmKGKcC0SKYFQ057jVc896u19KGtj/NsNMl+njx88Rk9A6l3Kc
5Db1YdWNlbOYW0cmoxBpOPW1Er0gb3LqaewvRwrBuRjWFcPc7dYznYsA7Y4+4Hf3fq/JdAKMvd8U
8Y20AZ76f+sj83xeamwTGUuOIo6tougL4Wh+FKYZtBaLsZqLUnS0FLxFLGkPft3G8DqLYlbshndv
h8yRleEuh43GgWyuEt0K6jFMPH1lP6y/i4Y/3BasExx+GpWFE+Ztjf5TpDRGpgbNx+vtuIp0S3ii
m4S2ACgAB/7c4xQwjM+ttlK526cVJhPSCOeRYF7w1vY2vKeuvggK5uf8YwevQSyraHVtv0vNaFr2
H+8uqAjWlKLhaiR8DbVTwtrtJ6dh6rtWtoUG4PiCz8cc0htwXVIrRpN05wKxq3yrHonrkEPx/Xbd
UoHa8bbNaNmAoybtbzzKp8M7yxXlebx5ec1N2PdRpVPQQ663zfCxUJWJIE1vzsu1MjUd7cKxgUai
IFo0X6prgqTMFrP6alMu8rSgWNtwqmIisT+w+n9B+DLz2X4ZAShyy7CZSHNNwmiJtZ6m1zH4Cgf6
ecjnuB1vyltpkRhppN7yy9b5JX220SnvtoRclDjGT/H2Ki5BupHG8BCMs2l65Al7r4UQ8WnSzZrC
hwoQ1nRwkBmgXuq9Ss35XGPyPDWAJ9e7gb8h7Gqxot946JEkuzJes9h2gbkP1N6+iS2iXn2F2cea
Gw/dOksDS5Ppc9SVbbnZ9J+ruySVobnNnIqbQYmlpDcDbDlyM1ym5TU4sQDFnHe4/GeDL0VmcKgH
jgMaImJ0/GwJCaEZ89KPbIPOXPkoD2gXlelb87TaGaJCzxh3qVPzMxRDXCdeWS573AlSfpKMOfpU
WZjfsPXO8qVsLkt6Ih1IfyVa0ppkY4NmsGay8LOj3OZ/b4gP6HR1lrjk+OF4Re9ePz4IAO/VE8/w
VqMcBV41Bpo3JeEuV9vzgwm1Jw0nzbdA8g77SuUKSSeRu+QmQDJHwk/9KxlZkrMVGA40ORSo5QwJ
oSISvv4zoTRaKmo+ztSqAzkzOMkexGIZ7tvUOufuH/9ylFvKzW4CdZVlMjsWv0oSgFe7aiASy2dS
Ej8zpzBnuwBs/bCNnoSDNNVH7yhLeel4019lO3UivW4S5FPROqK7kmxdsJAfFppj1sfb+NCXieyR
MRTbT5F2RmqQ7vXMGQLi1GnhhIdV2J1uzQZIyFLqHsUbFMHgej82u0eP6llDVgxq3sy5nkPieSAi
OkZQ0rhG9IvEEp8L1LAXAXJItn8D+1zoU3Oc2W7P5WrjYY8e7J393EXfmpAq8a+a0YFEEDHysGSO
I45Piy5hibNBAAC8NT8UL57AEbDkDGY45HsHIcwBaT7urdybD0VSzfHGdL4lIFcczqGxdj4iiDEs
CZGt/M0Ayz+QSDoObYvxYIdScsusUG8NyYNywZtMfMucW/4Hx6J34RgqKvvDZo+uzi+c1e6+rVoi
nmP8OEEsdP1vsGW2NPC9Spe66xT8FINRM6v9TMksy2kWEG2U/FH8NWWgSIY88hXs+8sWrwcajaLd
85VLUR+bNGR5xp/803gk+FwEX1sQHcxr86nlK3bh9xNJkh3IMJP1EiFCIdq7xPjFBbitnno4WR56
SodjBR/RDFVmJJpUFfVmBlBR47/+AzV1HBL/DHzG1LkBuWlJhTjM600G2VqzQ8Eod9zxdFs/0jQm
dtXecPeBtxHz2YniT60/xJyMoOfzvVfdasfPqgswr32sX7va6eFsicp6nekFs87Y1kKbi8tSzuKO
K6R0XKVrA0h7+3murALgydh4PArssrS3M0HhOMxQZOtHwSlC0NdRiPrc8QTxrRGQKFlq/a0O7Dp8
/DNvusig2VE3FfIB4bY+BzuswFLwQfsVjqqcfjraju41WMy7XVkCmUfSezQgoSDsocEeYfhOteKc
rUvN5HUDkwZIRUU25Rdi9ozBFVjUeUEmokTuFLgow7Ik8qJ+Yd+LZ4HvO9+P/y53MJJJ7K9rmVW1
UBO7p8Re3xl8895m4W+VL+2IqnDjJU17QmruT8D7HFt0/a5vwP9OgY2nWUSgFKzMRUCgo+/HkvCw
44UNUMnmDbO2d7yS3K72rr9ejF5+0XW+zYSJcyXhzvROkv+Jc9JP9uB4X50EuJouHNC8u/P68awy
1nsJ7E+6BgXmRL+vNmU/RoUVj3SVzcpb6hKjQwkpqj2BKVRM2Tw4SN1VIsfdI8xdBGTrUUXKq9Ll
fiFrcjoFZxGeWsIbcuX3vf6bsNIwvETAP6A5Na+FDctn2BgcG+Z8Zan9HgJhp1AtuLDdWfB4yYUO
FTx6ef8EhOXswr27ZmcqrAvZygOUgzZZiE+NNy3x2eAgxnTxxlNMslbe6PrX9o9nWyMHnieC0cwi
VwEgJ22Ds0m6j3+yZ9fdIRQuxRP3fNf8LNt9L2EiUpmW/4KM2SvTyvL3QGjwCZjnzFJsqRjN5E93
GT+GeWfczoQG95orp1N5Rlu+E/J78lTa44W2qyEjTGQ53oU8hK59K9VDKftUmLsvjJaIFXVoXndv
7Jw1+ddhd2BHL6AGh/yJOaFWUHmjoMJ9aBtUN2B05sWtmBUpkF7lPqcDwMiM1MtcLnbKYildrBME
4bqZ1WqwsarfhanVvcOS3yGYFKn2BORkgVg2UKwvBgJSrgM+VGGU4+u7nRaHu+nTHctawxwCHfuc
4nf9J+tSkCc5TV+f3cCJP17ptC/HwqLeOrvvQvr+fH51+qWWkbRXgNDQVBNZnLRdNELm1zqtVfKQ
zLAZRMf26AMle3lSlDq6MytGcP7DhuoMdTWdlhlkD0mAaJiwS/4vJndeXWtL1FCBxfuY/xS2GFnw
biCesqTVat7H2mwtoNXzxhCy13UJM4HaxPa0YWhtL5G+LELnPCOc3zCnmu3WYetfdleJyPKK3bT/
0mGwCqPYRO6vM1aXEzVZOSqEFRNsSdL7AYmHLIZBOfNDEMzyS8VZkJWi+SFqrLdYKyO+00GoXZGu
lt+Aa8cpfLFCW8dQXEKRJTctzK5uMG5ibhEvqr2ixlDZ1Tw3PlQDFh9zfgZ1fvRlejtYqvs7qMjA
w3Py0Jx7cc8uSI1vJUae6vl+BwrPICqKxsoIFMEceT6ZzbJ6QAfjKeptUmGJK2Xh7s9V5A5Pr32o
4/1WFqfHWZ3b0iw94c+pNA7pouvluiSEAgbivfQaE3tLFs2ywLrcnSIFKyXEeDuox+GQ8Fk8SwUK
5OueD15IIv5FVS/hTGR3o0jdG6A9A/b3HCfbsehXg/rVVjOD+U+gpu7qXAqwmbbp2Mgnt7hykNKC
Zk6lCg6O4VpjDUo1tRlxwdzkMIv6Aue3aSqinNkX+a817dFlb8VsPj/DloK7YNDTKafpMlGocek4
0StOXiaWCIK475aLh/27bJPFTfykfjC3yIjQeayvECDID5WRTdEl+yhJEoha3YRQlfMipF95ZS8U
0JeKZaaaMQr2+CBwoCgaqm2A0Qn1kC4J7xyr0dbEUJWkK7MkVDXvqO/FuXfDZEtERLvGAk5szpkR
lS6MvqNAeMMh9ZW52qkf7gnDrCClIJvJcZ0LxPY2zQp7/+Y75lSqiVOp4WanvuAjQuTwynvQgeJZ
ZKLmwthDRsNatjruiaHUq02d7e0GLrRX1Qh7bquStfdlm6jLEmH1hJjFctuUM90yFozfNgT2lsji
jGT5sNguRWnW9j2cnT8cL4FRYpY9HmV5glWO+aLgWlGwjB4+2YDReMOiCVY2ZQCWMOSJo/lNcg3V
OtGcgtfkN9xSFF7p8etq38tj9Wrni4AmDCV18xRNv5PtNtgz3OCXVOjWCX42GGhWla1q7UtYm6wM
Hg087d0JEPqacQSw4OXG3/OuthscKa3WifHJ8JEuhaFnXFwPnqlUOU2Ct6JpxoPszmsZGIZUlCiV
k+J/FSDHQKfu/4IfTku+N5LhXPMVExo+fBqw0Wv0LHu347Qa89SigHh7r6uhl3UvZtr9puc/sbyB
2mykdV3Fp6uWS1wPJdB6WCALAEeKfEiVnkAZ3aOD5Tme1VFrUDZ6Xpow9/n92o1/mlK9m/2+dUAb
qvia4lYNqP9zNOXd6FwHVDjyUy7ofIefpJQZMSdS3QmJ5BlIL7J1utLlwPnYz39qpbqMY5ez0YFL
+VGM/rf+U/6BjeZp8PR1H8eNhFmE5DdlowYyPgs5a1SK6mFTK0ND/siqwPTAt9vIXUWoiU8VOqGs
aQOncx5LsqVfLWuIgay3SqvzGuzHF0lSKa1vQXm50Chr5gvIUP2RUYKs12xuJDEamCFMfIagqRrY
BLHzqC71HGO17pjzi7YzqjOirAZx4LOTysUzxLkiG5xwimlJREcX9G0aes5B/PCwbOOgBZKWQNGN
ER27rVcQLGGQ2N6aIiN+9C0rvt5efRTTBQ4I6EQpw/S/1qcTR40RjgdVgvQvSuHuORw48ZRJ2V5N
blwGou7rMgpyE7kl4Y6/6k5NDfJHJJJlg1wv6X3jEI8EMYa1J9aIrlMZmVm8c2q/Ina6Et5igyxL
0ZD+4YiOOqHRUKQ5k36kygOVyGDwlzx/TIkyOH9eafNYAnjhnNBYVc5SAHagZs7JB1x4vaIOFgrg
u94wSzQMqcEADZ7a/EQ/6ZLWB/RBBQXVAI+0m3fQABraeL/Hs+b1X2ZW4Q6GSMNeSUU99iGO/IgY
fnnMZgVndGk9V5xqOP42Y5LYka1bRlA8cnL0/4SWvg39lzk1AI7L+AaR5SUvBM5YC0BZhk3jIpUy
AzMF+lbY0OitDPr1MiC+uB0bcgCuLmxl7odrz/PGs8QTj/I8NMlnCm/xbnutRAd1Pi3fiZYQ3iEj
KyBbLVOvUBg8Ozs0y3MH9kxXDaGXqayMZFPv4s+OrmQAib94FwjLb5hqjZnOnu4RErO+XEMJHPKm
B2tWFB5nrK6wo3YR7mJXq+0W8nHiJmmxdox6fTNf4S0suwMrVZoT1ndkJxQm88REWxnUXb1r20Ko
cwcKMrZgAHHGH0XBOomRtNKOCt4tm4bCE7WSkI27k2bgZ+XzcjOrVJdMddsNQIQ4sHxEKg1VFdv+
vorEjBJ0z3OXBPbc0tURUyLkgFObUaG3elPn5RDQSMHYjpIlOL0aj5gyuXRqMS8/lNSqygEcvtDo
jAZzk/1KcbZhBZ4ic451KAn4dGjLFEnidNdotoCpEZAi76jc/bHF8Hhz1tbMJpOG8VjB+esXn1Pu
nPIhhejWrYxjm5hSjlGpSdw2ba9JUaroPO/z+WU0sms7FJbjlfTzM0jKtaY8BwelKQ8VLQl5EL4y
vWZNt3hAF8LufjNVd337dUYsXW9TacEVsyOLMPwquOB98nbw9XQLi/roKFgKSqm2TqgwiBV+e5XS
puuNj7iGo/hh4w7wjTLZr+bAOIguEXvellmmXnEBWUIqAft3ALPPIJCu46pc3nYHv645B6BxgRVt
AlM2RCo71hd+jY6jICTOHKL3qjNXPV+cnDFg5rTYP+bqlx94QF/0rCtrvxmOZJX/Tr71me7Ayyju
TYyOsmwl54iO43Ol0vZuAePLtiJJ0GnRJAJv2J9FSocrpOiRB3vBm8x4zy0k6hn6L2rBmDuex7TK
jJND1YY9lzq7afVmDcHgxl4hP/WNhLTTfVwfbO3QpiBi4sPn0dScrfWyWBD3v2OERCVkXwgMiLMZ
QLv1Zn3ze1FDrw1jPnedPg0+nWPjlVIfcxyLzvCzRcQ0cV24AD+DgjcMB2n9Xz3QTRyxq6vK/+NQ
qfJSqlMO0OGjJCBAEVTSvRFxABgphUcH6OhOd+jLTLYUHoKrCEukqXB2LLr+Pv0kqBkjoSsaQlqT
WKZ9Yz9GVwR1nO+WrXlpOMWdTjuzEWGuth75XwoYS0NnIMVnjAYhTFfN8rce4Cnyz8kmBeDkp5jZ
jVM7YE/B4kvUjfvYE7iGY8lT2ol0QpBC7L1ikuPRUBLFyl4kylf9Pn66KGjjbTgVaY/kOZQJjKSu
G5P4emwN/tGnCTEir7tvfBFfEPXeuQNgj6K/igvUwA6DjT4nFUS6ogUhfyFKp7iKAhZTpVkDcTAs
GEsOlXJk2A/7XzbKO9MoUyakqVg2Jfx8RFGiAXckOo/IagtXQLi6NSoEcnZCSGjncC2Alq18MYVo
bXrNLSJz5bKXwG10PIw0kfsIpU5tYfsZ/mcyAYycpKppBlfTBDxHyy4dTuHQ4/mmCH8ZL40ARb7D
lpSMJ8TZj2w+bX5zBQqW14Ub+ozNWjSdDwxpPcAvYWREgS8PH43YQFddpIHD9tjuUNatw4Y+KEN/
GSkatfMyc9q3yb4iCM+4RuysbmWaNvZbj4l+bqK5ttqfIx7m6s87hj4ZyRxEVqhsbHDWmnnWeXjS
bqF6MEeNAaqgjAmJU8dJOCqI4WRdKnaEX4/h+38pVtIYgCj4HoBVoIh/x6s+M/Xt7/Eyzrb3fDoQ
c0LoV8JZIj/U7MeqVBwhUENxn37zuaLyLuUGG6pWj7UkWW2KfpRqpW3D+ilj2/IhRAPW/xpOo6nu
HUAsiCYtkGyxXtTv6a6/UjoctBobMXtMmLAWjYMOnTPYvdMPa4d+DWJ/9NO7ff44vMrYYoe7GOoQ
uS1S56vVCXQrWwG5DflJiNmTuKWwORMLumW1upWZ1E7phzfONoWWbGuW2wmHffyYhwPVY+6PHMb0
GeewD5VPYge4LZ1Vru4hppmtQeUNKJJnPBvFgAXtrqgdRrlNTmrGgWWpuJmEcqmdCuoHxznfuKar
eRn1dNOvLABFjhK4r9HJAIcz/5GW/bWOjj1/uA7p33SheAOSpf2OyTBdALoSa9rEmCBHeY+4Ougt
qIjiqscMo4sFx09O/RMF7yXoYu3W4Kf8Rlj0EHDXz280ka+MhPbRVTsX5oAE/T3uDtrGOiJRgu+i
erL7hFTDkK4OQShJsSl/bajMlwbCLpNm2NGC1N/mi3gy9wTv2T9O9I0RwiqWUDb5rYfdAz+2Ij1Z
ute5YoVQo+/akPVE7x1Eg91PpmdZkUR7bBNHYWEegiCGjiOjqIEiL8SRsRDHEPaiO5gwVC3gDrEy
EyvvyWBBjLT4faiVfpUCX2VxhMQnDCbfcp72IKkd/9BWqaO0lPGuGxkm6FaO5RiMgGzsYz0XGQGP
83Id0Irjs4pVcaSnuOHU9n6cqMfHY431chvBr6usp2yaEGnIm+KgI5KS6N1RVNpIopIiigYg4MYc
aPJt9CKPCnTyQq2iNR3BnxhpakP6q8tc/E+Fuu+DodTllfx0NwQQnTreA4/HKNFwrAWrPcVvxVTh
B8QI7aCHu+Nu+xFNbMW3r37Ha1IXo42/GiuzbgHXZb7AYJXmbV1sQL56ols5FQTDv6ElKap9LbQb
+fYTCKhciHubCkVlh7LQrg0DgaYHSCER4ept8Yea5lY2GFZV5SBO14TLFJl5yGo3nus/bsx8fDSV
ZEj7dhzcExQLHLklKK1xBrWJOk2YFVmfHHEvqklGt+vGnhDuyv2IwhqY+MZqiKzr++qTmDjYX2/R
aC0oxqvmTGX2wjmJ+XWlOWAWBVB2lsVa9io5DH+0vjxjHVTUs+PgLG9FkgIia67/l+XieeLR+7sO
XVAZ7imlEwEosDnUllO6iZAb8PInMKWv4slSGFKLLCoRPc3jFByahu6cYUSS+qlgEEn5/RDsChZJ
v4iEdI5vXllvt1ruGw1SEIs0e/gww7j6l2601e7MNwBHl+3PdtyG4/mdUydUahXdahgBpqQ1XqEd
S1ZiRgL/Jg2E0EY0hk25Dto6q6PmgUO0MSOBP+H36ywbrufoQDxOTaCqPrewNhjX6plXkNzV3PIG
Ow2k+A8Q1E0n1h69a72J4jNwVAdqUOKOLlSfB4ZL+DaIxdMvyH8KwvlVC435eFXRguXQrYj3fvyK
IIN0f0vstJQtVXEK1SOjU98J0AG1P5IUp5/t55OVAx51N4eess0jFiNKnMH2ognkU19YlF/cbb1n
RVx8cWBh5/mNdeGNRVGKzf6gyRnrrcNHG5tSo8YKfaMaQ3wYR7BuAJ0IKY41P3eTF/rDae685FYo
7jTmmQBS8Hwj76hdzWsAXwALxz36SF/KZT5xC4w7/qHhhqSo2MFeP640dtEDgtXnRlyQ4ue3gv2Y
Xic5Y0+8FDoRrRPKHuk2jJBlPepmVVEFGbjV9h9v/q+xrfXJINsJUEiJlo/peInRXgAYhxjAWSfg
sIdUCy6qehYhwFEhwiboO04bK/GVprf3Ot4zEJWYMkNHQiRJK3bsc8LlffECTC+syEx0K60mM6ZD
eLrZ2t+7VbAjAiAXrxrWLjFdfeLNyum8rmN9qFc01tbsejvKY7Ai1KEVmDdi5paYk9Q1anSyIxF7
cuC0wMa19JESwkBoWvKwptlfV0B2xubo32vrprqbHu49iMSVTU0S9zYojXvyYvgwKaUqcR6mNZFT
uDzT46OFYskGZ/bzJajrMce8luBO/VMl/gmTsUYMWHoFFchX+WfznU6jSWkrslOoJvUAERurHohS
4luOH05ATWmumU+2uzQZd5IL4p3nAMaeUzOGFsmhfxDPIKMCuuIEdvc8nL7Mwj+lbL0F4rCibWiS
txdMohJpmlavdS3oIp09D5Mw5vKwcOczUrIhLdz90tgq6RhTkSaUZ9u0FiwOq+UzRqidEOfjsQqa
HlAyXphxe/+UoXTycrI10avyJaCJsDlkwJXB6f1cGQ/lCi9afgaf0eb4ZM37s5KG2pIeG9ARWi/2
qOsI49ftQxjJKdqoCLFlDR7VBbVLnDIh17H+qXxH6OIZKO2gXu7+S0JyRrhKSCE0jJWYsPupZmNV
yxdCvemnqLUB9OCyP3jnIQDyC4PgI+8fHGy3Y0kYsLnozulXUpiDnWcT0GxN8abgzbOP4TIvDQSg
I7QPswwRDOrOQwsX8a9BAGUBje5kFKixXjcnpcfs+7hyMbhjLcEsAnRKAK/ZqVggL2mXk3os78wU
n7+2/6fgwHpoWEih1aFVUFyiGw5v13FA5Osd3L8909sC9PjIv0vSYsIkv+2Us9bprMkcEFNeVNso
nlJmf+zgfadhB0Kh0dJLKKCsJjADMARzqKZmZLS5J52AnMBhSOepRd8Vg0J1dKnY0lyirWFjqrRV
LaHdFbSCbaCt1rFEY0U2c0m2rDKA8FM4fm18sA3EFL99oy5jTLnuORm99l2zYVRM8udOa6PGiWNE
3JgCJH1EsQ26oVn1GJ/Ar/A8J0eVC1t3LLigYDYLAJDQWNnrxn2aV3R6cMCIgh8wga/8mH7iNsR2
ndTPkz1QF1WN2b0UYbg3b1nZc3BYkln9jxDzYSrIijMwKlU2rKRwSG/KJg7BuyIrRNhABNm/FoRd
XRcCaevMfc4IUumh4BSwp+2m6uIluqRqDonWsSsqJoNftL+Gxkqh999yqoetf1YZAXlOJGvhfMzm
TC9IHT9eA7AzPPaYF+LI5QMyeGHrTqSuqDtMdiOXdyjX01nLWbkJ/ozQEa7q4J+rD2LhvhdcuKvJ
fHBWdnamppN+ZlyB0hmqysMsz2rk+AKK0SOqMr0Uu+nwmlgxRvUMMFKMcGjAP7KwN0mPQUfE6/Yw
OJP1ZjWR3aAhtTmha7wutb+wp0roNMvn/ZG0dA4s8wm2XoITpnjejXVD3BTcM0fBEHD6LnlJAHkv
3dtNfsFDUqsNWeScn8kIuowDst2u3+6pW+BFX0oV56s8Vzu4wp0pTJEq6AOyiFaaXAV4bH7rLIwD
JLuN0/SSRrJD8W272KewVmwJbuxDNM7HXzHo2mN9OWBM7kjFi7tDSIeUZvkt/bpvzCGv5+aMti7b
y7NNwFhk27N8DAEAcqax9x5Y1BXmxwxmBF6QVno2vTVd28mEwr0zJrUokcgW1+axHnDtgQw9S+7e
r7gVERZ8IfQLSgHwKUE+UkH+SG3Oauxk2L6eeEY2+l0scJgvawqIxLc3qVS2NiXpMdffzT1Z+t+T
/lhtjS3HmnhEnm1JGk3u9lpmQtfCNrzoAYZX9irbwi5+wtXqJd1G+7oLelwLURA9y2ZlAFoQ+piq
elzZp5vXV/QIzsM56+AYBtk4mqI1F5v+1S2z3GYGN/VwoB+f1kyNKnlyUZObbtDVfTtLrd14T8JA
arCoOKn5rzKJoCAhf2EIrNcuekt0hj4BkDP3HGFS4+8dCOY0pVctPDc8NkVPIEd4QiXQrDMVg/cH
mq/kk25MgHK2Nhwmh320p+0TJuOQrrt6D+sn8H8e1IJ97qOuEvpld+lMB21T2hXZUKZUjs0nQUcw
dY7nwfWqAsIYt5vnSKJUlOj8fTNY56NkNq6PwDV8uj5GVTC4Eg/JZtBfAU0NYz/HFbULq+4268Ft
9BWblG2+R2mqZW+rmpa/vFj2rTvNIr+5naMwckBMYwf547Oxpq7WzWD9zmeTjOpwNx6ZoQ70kOR2
wk/bfpEt8ffEUezlfvWzjEdrKY04So/n9Hax5rXcfjChzeHVlaeussstUmlJYCj3my7u4APdkWfO
SFF35qllv26Uv07pIi362WIBVvD/mIsGlmMXltmEaEWfvGkbhTHLCQQuTHrB5QMOKN0ehWSmNmG1
UXe3L8R1FiS7BgOGCSCwTLLi1IOeoMc052eaYUsl9sjt6F2sFJymLBTJmKlVinGKPPF4F4Xe8TDL
/ahU7mF5lXH7N426ZBtpvWr1GuTEKXpesol/1C3KKvJs2f9JEtjoskoGRKfxJWiRK5INsiptSOwp
aTo6hQ41enj+QwaGuSl3K1Ozbwis52fO1jESWq2qO+nk03chfEg9JwPryV68C3KVc3BzIXRRmjt0
WJTcTztCh5b+3BF4v4wHHoIzq5/L6PYBNiT0vdf2yGGjUHkFgZI5AU8f287DHH3GbbR11rp8ire8
8vp6syx0Piv+rBTILu3gYw1mLIAG3uCwckdTHcHgC1cHa3KXmQ5x49rOW4CjCrhvj4APbZOzTcag
KDqZC4Ap4qZX2KYUmRwTPXxKTfBL3PyquEMw9by1S2sTT3GhR6TqicJhNOnO/HHyPnAefhj5us/A
WqPtLwmQEcjh9nyjHh9Fw32ppEuav+f8xh/sgoEg+fTl4qlf3r9+s6kKo6b68Oc33zEOe8r5v6Aw
4UPpkPdzHW0UFwMaCp+ogWOBvISZOg6HXSB1fKRrnzHdpmtmmDhPJ5HXYz/rRlW6QGHzktIUjcOd
Vjxky2CUSP1n9j8qdZL/m/XtrfnAuytXLabauQy1dULYRtKsNBVxL7Y8CImC8vedjtM3cxgSGxaz
ZiVFcuhaHtnwEvA/7mqHpjtw8121W8V/stYG/3/P5ppOCX2K+fa9QcE8BHx6nKxV4b+4/7AdWIKr
AKLUfpjZtC0dMtiDuCpEp41TKBKIK9k9FZ1lCfdLsens410mDff1afcGlBgmXXMWnmN4iLz9ZEAq
4xksmukrLzBdnPo6/YQ/msBSlGJo+Rol7MYvPnpBD/KeOPWofnODWHAGDwqkpsko1caDaPHb1qwn
KZvAlsLNzQvO5/JWYsubFIdOlzl9nYzQDvpszS5u5BOu0RYD+d/NKziRIIO8EwtamH+8qqZbGfLh
xIt6JAbwUCtq8CiGc4VArDduMb7DL95vI7/jnwZL/zAwMG3p8xKcpK0NvcRjQ65Xt/eay/D8Whtr
ojzaNNTOi8opafoxKy9UiUUBFZ3lOZDcG2LJ5tYwrK3AjANpqRiVj+NqaW6UF/yMdBcmeVX5C1er
cSHtMCAF4PwCrkwuweIiyYPgU4xIy5mU76yFTNW2ZJLoXHCaTTgKYwJge/ZYoU02/2zRR61TTdZ+
cxbT0k8kP0C7/l/XFDd2eTm0fuXyILuHUAwRaVS37JS7KZr0G8cdOyB7vyTDD+uDJip9/1JnMR3Z
4EDwlIseTdeVodX19sO3bfGCnhrL+jzf9KTwbiBprnMlBxwbP0FSVyz+bJoCfEcwWXaEBsPkY1GV
LwAfFbqaCCoEu9X2bwRtOui4H76DNAqAJNC4/7ChwA7KkJH+gAEgLK+lt4PGtK/0qYwRKtMlnGp4
wD1u3ecuUTlnn/12sI8ofGRKGEVpUl5wol19ui5Vq6C9W8U7FKr+lJDhOaHhVNGqBT2EIIfyGLyS
+cQ2WIDWO5f7jyM8eZ96Oqrl+kmgdwaz5xtLN5G31X4AV0yuf8/RKQiY9EWsO1WjwPHn3iaJH49b
8SuOQL06bny0cWVFEe4bFiF95FtfL4vbqF+34QyyUErwN+a1GPFpg20ahgEoD1LeXwJBNyuYM/wn
0j8ma8X+64/3v44WhPUjAYYGju6Gk9TWi5p9xq4pIHY2dJatHjjUMkf1pwZi9OaCT++Ofk/Cd8Sc
WhN0Aw0FP3KPOTBxwXoPhnu4XacOrfinFTIIpkwkMvbBwvQBEHDJcA7n0rjgCH/7zQ+MwqOLveZA
fLqQe9Amionh87qbxgP3YjfqR5UIUwalLSQovlN5u/Fg7EsYuccbVL9hG8/1Xi9qe2/MZVI2gZPU
3Nv6DdoPKvReY5cQxq/+Bz9aKwHxJnblSHzU53us7HlVk0OPqJej1TfstB86PIYzHj0bJP+Igoz6
WDrVi0i/IPWJ1yzWx5a84JtELYFE43zTrbencmkZY18Z+we3xvJafjaqZNqtRHMOWXbAZsRWS8eV
+UgFZH8ORAoA0eGcUrwDUThoKwGrUrSWH1qCeg8istGEx40HhSEwsCA5gkxZIWWRCPsUfdobKq55
W6OJlNNkhaTYEFkcRfBsSj3noRkcq1L5lWf9SHyHXBnX3hCDPajtBrOj3d+9NWaSGAhGA3MZJkdq
PVy45bK13KiGup3wQ/dps5PkbERNj5/A5hPJhmkujy/IEvQTmQeJ+hey8UzvJdi4KewUPz5yQd7u
jk3jsvOYWa149wBzWB9jF23bkDgKg53EfaMTyJ8KwK92ElfBBq9dOna+jE9/ZgDdStOeL0Jl9tj4
0koV67q6C1SsIDedR0Q9lSlOxhAaHia9cTRju/ULqstPFNpzNrySX8BXC8ytYKcim2vQ3xtx1zME
2PdHpeqkEG5ujs5itlCzeyaHho8PjOTX0E2rQ0UVE84y8xb+fYUW7Dfsu0tSd2qQwX7vs0Yf5ZyY
GNR6GuBhM5BqY0CYq0v3M9vZaYA2DsNAXsvCm28BP2M9LY0iGbT4jF13+qvSiyaNvwgiH/amgqYe
iL+q6v/rXfPP+hrK4bGBwliefse3nIhzPRotQH76ZTpOsUN3y+wDh1HVNV/HMKcwdAZLJTzGeqJA
fmbLAz+ahwXiWh28haor0JQxMWGqjDgedd/hlvBDubD5dSCceuwGrwDPgS9DRu0Bu8pifpxIrMYF
EQ44rgGe/ixqVqjQ1wmemdr9rMQGbwjQBPiapbxZuwczXUh/8XVdiWwvZFdbv5Cpx1te+UmZw9GI
+3hiXicD66lEciWb+Tvun6DrAxRbhtiDejgNdL21OcjHMV2ULgBo7jNxloWOBEPCeYpDgMddzIG9
7yzgd/vcPrCbc+W8SeBONAWxcNSz6SGf5rL5PJqTThkoWauAFVcAKXWk7pf+y+WuMjsM+OfU0K2b
ARfHLbjrs/tO02tPk8Gzk2mYKT4Nb+G8Qo/3rFZKYlaiH5wUgJ9sKMRRB4ncfdF0RshCpRVobuPI
hS2b5r1uli+LExKUmTJwy7Ul9y7wnbWIL2LmxvF9ZCpS6U8H/jyCBJG3sQkTC6+F8AyTkdlADhJc
Bx3v1jRAx+0adO/OBQTPs3JZ5RRSyhd5UD+BG2u7kctKzgIMjdrGH2FDHpT5pjT3LU2h5QSb8EQT
gy5xM4jGhiz56PsIXVinIV8R1Nr0zk+GTOXNVQwMMEvK7d++8z5L25T3EhtQa+uvn5ooJFI4KtwO
JtpQRti7zQdPbLez9uahi/+zVUdWQ+mhG0tBt1Oish4Q6PChGqP4Qk6dzBuRRC5HE9Z+G7xYHPlM
NDBJDD2Yz4nGzpUTlICzCd3WFQLMiIEz8CdtdwPbmNTEw6DEWd+7djvrby01/K7Uh/BEObOSU7GD
Xxq6KRHGuep6CcFUR1pOjn2EcT/kJ3cdLrvdyy0K+e5Y6oHiBC/92b6HbTHlyxTzsemxcHTKuLuO
ZowCPHSbAPxHehGxEKmpaaNasfzrTatxuNwr7lPH7O6PNRgO1Eq4OX+wqQbOwCoE0yBRol3qIClx
RxLqZfQ7rPeOIszFVle7OKLWHXBbxcQygooepOkliUlYMlPLEEbxemBnPsCzGcnrYRMJlt6WGeuv
rchRB4bcdy1iEo6OMWcRkWFp5Zty20Zf/1njP0IrKLOOWTguzGiLrwfSyeaP/NnRu49YKSoGIOYW
I2uxdX3qyiyRlm9uiUEMnnMvqgOMJpAX4C8HJ7agNDPUn8UDEolanbJUwlctzpDDh9BUuYrN4QPO
01mPn35Mnq5t60HRqlHK/P07jsQxch6k3sA6/tqbFVdSHu03AiBqs4hKoKh1aMFanK6k0+xpcjk9
sTU+4PxbxOAymQnUB2/soCbI0fiDAwqvx0DZrgKdIWSlUaXhfm+P3sf8Knc659ieUD3AexzbwyRt
5NUMgh3ugmGCwwgIi4URTsrVLgr+ebB5FJ8JfUmq0V4iuTLb/OlSWL1r3uXOpZW0b6KLOIT2xxzR
p6fUEKVrTHhuk8PKdp1UHZAjfofk3Ge/NHsQvyCNA6Y5PnDOfuvwcRaR9R0jmZNezv89y0C1bxYb
zmxD993Wur7lRbRiRG4Ksc/okQYriaaICOJxJkMqQULcnf/UsEAF6Wg6WxFZSkJYJkoDSFqWNnWa
/ulq4HRKfYEdUy9HE8oJU7K6YcBGZT97t1ARRpmfYvuYT6pKl+RKDBAwsLtJHgBydjdlCclW+WyK
IeKnlt/sy6qgAdqB/iMYZ0trp7y3vjzTSgLuW0VQMh5G3TC1swddaJw8kwb1MILhF8p+BnKJmsQK
wwG3VACf+DlI4lWOzYtpf6MWn3kJTFhCSI49G/BxivBrxt9kQRWyQ3qaOFydFYvSWt4yPalutinK
c1F84O/qDVXp2BH82k/NkXtwCiZelkllUeMU+zGVQZKCblX5vIkrGMpRRtTfn/+2tUk9zyIhAh3z
bcsEP7IQMVI84JmWTPyJru6+HSaM7g6JPUdWVddS/UYVg6BzBXl7UHDy+k0U4WWx+0zXH6lsF88E
T1sVbkdPrwfDmauee5DX6UQhgf+W0qQ1QPRxME32ZJY8jteOSv+UBd3krZ5nR6pccOZrOEzgCfll
hvKDuwhBrMes7ICdC0LZ9PqP1eFo3OM8mFOExj69chcS/DePFtFLMnve/BHHufLlPb/HDMWLEpU5
bOzbW0v9uZ3jASYI0kacfAIDv9C+t+wNf1Lfgk1V6NRwakQ+QQCui1Y/xTlNBV4dv/M4Pa4mGG2i
xtUOplvRP3MhOcMKkMFyIPRa6YEm16cAXDdb4Wd4Plts75yzCL66GgIudoTCel5eRkmwtgr5vBQq
Z9ZSdXjDmaStMwHyLAUeDoSgZ++5A4NsL66CWbOFx2gwe/WCQ1/CH2R9d6XG7J80w0l3RN4elHJu
H6oR1HHCRVrwCdPzaZwHn49u5bZexfHKnlj+OndxagKIk9QC2ekakQValok0YGuOp7yHXpFqkA/Y
k+EXYCS44udH235n4EslqY8pPjVMB/9w3Y3Jr4TRJ0GBoymaXDamAHuZP1CiHkKPYQTHQt4LIFKr
kvITQ3aoyIR7u48ROQk0oFdnCZaHbLg5wOu0RZWZtcwIZJRm6UvkPk3ITJtGc11n85vcdXsUG1Kx
AXGOpgjGf20Am2QQV6MJD6ywEsvANNd0DCtBQ43pHTv14LohWYfbs0FwadOwVeIS+xN6fgsMrDI4
cany9AY6eDDIG0/n7bq7Ul+yNDmhQsekL0pdgoktpVi4yMbCmcmZlrH5jNR/I304mDOVYvi0JXIC
DiD2gpIwNKhtjtqdvE/rd18GNhcRVPSuUGxitFhf4RQnyu8EgdS16n4Ht3FD0c3qzP0JMsoUtVjQ
Tz6g17edbax7UlMtWDxpbUVDLaWalilg8uBVjA+Eee2xNNd/QEM/ULF+bQctYD/8vd5WsWC4D30f
vtsNotX4Cikrx4LO/K0t9kPwrwAalJUq8LISD3tWr8sxvsVlNhFVPbKvZsVIV9p4TWCLqvxdVueW
+KQ/ZO7aSeIr+HlHbta0eidpjTG7xzk3ruLUqWerhO2aKUqFUGxyyzyDe3bBa0T9vs1k5P9vkIxl
JtBv9AwD2LwU9IjVWUVL976unmhluLVV49oKzHoZF0F6BE2FQxlRBwn6nX3PZ1LVtm7abp40x6gM
eQewJBT3Uu2OCN90vJ1EHDL2vL+pAk764hJCulqHj0MspCnKmqu636k0UvYy7dfOUFh2QATS2Aj0
JpcymECDsOT89qYjHbGlKNzQAz67v31a1WD7nkk+sed1z0i/ub1pGkf60ArfRn6MdXhQeTtF+T/s
0SwcvcZbFBRdjulLEm70iXb8Ap1DIUt4UWmNAo2e8Jho2T3CchOsQolFF/dICkZmZShOLOBziSVC
fpxlVJNRakrqqjhgc9NJAL5pkj7e/RovagQMUd7ZwYVId7izmopik7VjIDqxCJxZlYHQe6dtpnAe
69Ws6ITpFhTFFt6o+l1zefGm0NTyweWpaaSLXW5+zC9u4iNm0CM6GYMIGRxYk12fEzPH6SO6hDzX
IqCXGtJQdevPpS5YNMTMhC5ErWYC15tuX/u7Ae5TTN94sJdtVTT+bxDLZrljrcizDBCrUn9qiQFk
hfszddR16U0Ny9tKGNCN/DTmKp6Mdi1XGZEX0Rp4XJ1cF+BuVvPCnuwqklpSwk6cSuqOjKD5R/e2
fcTn+d3LZEG462ltvIBlrfwqNI6FCJUr+3VfimFl0EN6qWjNTG/8ox4vS3oBP0wKdlXeGBi+/6St
OVixLtx2JQpFx3H5E4b5PV0CQlRgR5mCkit1cyyCCXK7GnRDP/tXn0yQ7PvxMswqozvlaZ1Ppqum
QcFcJKwpFOMqYcN8peWEvqz0+sBCnP8PlGFGyAGgGc3c7viza1wagjTrb2cQSgIDyhmcwB2RPp4t
NnrX69ZgOjQKjk0aQ0/x+GzB0CbPOmOpZxBg0+zvxdcRXR3Cy1WJVdwQBcDv4xa+IY1FeawjNqwV
0ByB0y2bbxKri14sfdqQrH1m8sjUgP796RhULn3rEBsPDwreM8g4mu8opn+yj+7enyCaI5jpgMGh
MFwoEYHv+qtZma83Km71+5Njr4uaEOzBuQzDofr4JRAFduDYPqJKc4Ez7H8bcWikPRajxtnunqJX
CBawJp1WKt0VEUx4om7KS6mEIG+k2LZ1aSCVKawPXxzK3fMfzyCH/D1sk6M+HqZ5dvYZNW2r5WCQ
kGHZcb2TOCmW7/Eo9hgDPzWho3cRQSjJhWBVc5Fr2zve6WD0Tc7jkfGxnfObJi2epr++n69oHWax
0HUKq+3+dJLkZg01MYiXlo0M0tzUU/uWsk6DNboKQU1NBb+0S5xMl0o2w2HBE28vbY7XAN6Y/YSA
oVTOVOGGRsqg4AzBFFLj9PgOb8P0ZRXJr8Bo5kR/JbHYV3ecsrwwKAKM1ZgBCHsnKxhJhCE7BpJA
UPxcgk9QdZdTl9pSdtSoSbWzGvKOsC8uhOFSVCTAREhDCo2PI6iUHyCMR8fzt0toUDoa9Y2y3KyC
R2Fb+lJkYWIN+pXvFzN6E21JFbPblwDhiYuT1756DsGMh3+HCY+QpF/OJann6xkHeARQmnWKI1TF
FXpmnw9lx47pYbs5aVACFwbW1IUbZm5B3XCh4vqNjbxcjLbOcMimmej3DSqtUwvzSRbZxNfppUIO
8/9P5iVc7KN02KCR1flyvnUg/CgM1yzGov0sT3K67HlJmYQZq++AAM4GH3YlRrC4VDiv7oc3qPQq
keFztQ5xxIHbaHmBKs4BidPlkNka9qAXoe/C9Gm++xxEKE5Q7/hDxy0EnjuhecgwvR6HSJn0CZLV
L2SaBM1EW/R0jz1Mr09JntohK44TjUPrg8OUJtJ5kgaBCxyXuGwCN9N29DgkHiBMlQc9iNUv36gU
SXyJ4uIoaSmlghTnAUX8WLTrF9GEykR0+NF/H3p5mZ5hZW1kwIC5DafhI8WyY9/blo+6LX0ql0rO
psuVamNxi0dSXfoKsfwcmipB0b2YGm4fNiLQlONRB0DYjVudHfw7lthdtH8ZzcLv3O88w/JW7UXI
mYcYWG9lEhW9psbV3CbRaQZKzg9cEOf04jF5PUHzu1maBtZ8B4Dq+jp3HiWO4AAwF58/i+aQ4Aq3
sRl0jr38DP9Jo4n09Mpzg3OMCDwkvEgDgciEm1Ly+oTSq7kiY4uiCF6Rk+joQccYd3sE2SB6uVEQ
xb6K6hmWbkwBTFfkLBXrTQaajAR2OIZ8+7uQOw9Q7xgBkCc1ootsF6f4jhsKlHZgOQCd8HE/1CgH
uqiPGZBzqjdrduV/D6WyEHI5aFovs4glF+hb0sACR/a4u3kpEk+OTnMbOxtqIavggNJofV2xTiLN
TOrXDRirte0QFeYgkiLdqrNNU2+as24bsd/F07DrVkPGPOiYRsYbdPclQ9wGhwNb6fMlswenkAsr
riJ0QumLo29lsKMlQGmwLVSpWV967ucIbRy1JvgNFSomh/vvq0iokHEie5iahFVkg2wY0CTNWZn2
X5EZpNTvsVM+0G3KuyJCYd2ugbdn4OQWR4AoEAusnHVIFlVHuWLsptpaRVOyMAJWTjFrcHxZ/RhY
M/NZvHMDPV29Ukh+RyBP2vswuxUZPcfTUc59GDVS7J02RNynpaBBUE2wuHdwOhyZee/a5LK94ltM
MDOJcLthbAHOjmjNP3Za0T0nMunrY+6CGfpcMeYr0q6asxw3yw/SqW23gP23sSvo3wglTPvzNdCu
RN2P/BKbpuLjZltI1+e35g9mIQHb7z8t8cO0IpCMnfnzq0qwUxyjN6+bLqwjAuda+pi0JqrB0Ydr
KYG7Qv5+9MmCAjDUVeoQTNDpARmXLcumVmMhRE8oeB8A2Dybv3wgw/qgj2bzQtNBAmnPUDEamnu8
BWsAHj/taGgQnMQGMnGR6PbnxI010ibteqgXhR+lGepIg4uJ3ULhEm20rZqhgTNxG+phjGnHvzEv
qKWGvVgfK21NNhv5oz8nCDtpM6ciCYVNEamftd0IcRNfui9giF2aK7FOIOSop+3poJmQPPK+GG+j
71u8wdekB20YwLAFhq15ARPAWZW+HafToVfP92TP2tEeI1KvYF0ShC68Z31p4rKCYUFxuRKNqOWO
/BRBdq2ja4M2EUyhGRpmwMykYrtVoGCuQBddIgx5SVKS4v/nExEpXxSMSezEE/2LJHZkTBp2x7P0
NV9rMfvJpQeYYgCaePOJyYGbo3NdVq8guQav0wj8rFyQqXTLlWgumI0z6I8zUi6Fj1Bhn0KJF2Td
jOzwISc4wPSjerB0RDQVpPE+qHMeH41uVjuGJlr67g4mRHxSSnAMLOM2qweeKS3HnvKb56iwbMi7
Cg4B7Ggqd2Bhofg6ePmut3wJ4WDo9DYqLOxTSRWQGUQyKDnycn7en5CRXDgKP9oB221wAm/kjmX3
85Pd+Z9jwLllIfSb0yryCfxz5njf8iaF+rK3Gfb5FOkJJJnbBqJTCSbU1YeRHupTXcPGnXsSk4AK
DSwbU7uU3ZuY6NddVJiuEMSD5ZFRFQXz01ZX1ZBqVuAid9WvIze+jzZqyBTJI7BI+ZmGb2BIvlzC
cpiBAelwMJqcDEpMUxpD/bLr16VbDK2shUon1A8jDTXJezD7AC2JjBJ9qyLjfSMwOIEGMsGiBIFZ
Dpfz48/KUBNMqGZq3HNOpYlaLj+tRqbpJ1xGF4sp+Ndm8vIG6a8ce8sURDtgYygy8p2T9qX41s6s
maoyHEtqCs3IfkaN0R/UUKFnNPbQXZt3c5TuuWr9Ow0UeTTchihQy6x1OfqpfjKIZl+V2T3Fdbgv
etyyRaX7m0Uov0mLnuosBCoR5e971E/uP8TuSLLxk/z48uPsNhd6hhGXoLRe7mQQTHK4+2bVHjKD
+vEGDUlHgtiidzcGfQ1MUZchyqxaEqCfcA5z/knh62I0kgPChLGu3uV/h1YVeFbRo+UUJfv6+8kD
pOFU21dqXZrtSIHBsQWNC4uC4/mjz2meBxnlNctIzWqlnxE1PReOPfm41LXhw62BJnFbhzZaC6qa
N2Ziwf/Y5gtuMnLvZHv9pUwt4/PpIUBvgCRPpUrKy4YOAe7wtrLUiVJmfVQy4LpM7T50Fz263mkX
braTw1Fql8SqWVtfU1O4VuFZV0Qvpct2jlySKbPYTXH/VD2pfazvu5oJGP6cMnglb49UJENYN71Q
4ZM4Nebxs0rIrbxM6WZlAAl/5/zCZEwseRCOb4uMm9EXHqISZuRWI/aFha23HCrEWCnKIDQlIPi/
f6DIrNnIvY5xFOWxPmpwc/rsA7Z7qiq/nrgfe/v5yT5E+fnK1KAbYre0PzxnwICO3Fu+HW0SNfBE
wmG2QUMAms+VJGUhSJjIIXElvICcJ+z04ZLWTlqAb4Zl8brUqSRNOcn1cQnyyNCtnbsH7Tki6te0
mJ+4f6XWeXlfsUcEGovE3reGzIA6H3+IJRBNMKBebHNUnSEPVNJqUUfH+wWWYxX8UtEBDBs4b832
YhS4S2DQxIAytJpVJybZu2PPJv0q9+NQ4rBn6Nfm5j/CKvaNUSlxgVS48n0VZIAZyBw2UIivwkC9
+TgLLn1Zv6IqiXJk5m3baVQ+pDGcD/GEylmmqAKp/M3MXDtJ0vBq6o1auTG0znV06oqWRBS95+yN
0v1sbbNf2neSJQ1+gaevAWf6/rrm1t2rb0ndqRIfhvWuN7S0pTJsAUmlNBoKFhV73cJNKhziMIFy
hxJartq030NC5c320xfRlTqIdcTCUcYFUP3NX+4VzuktAnrX+/8rmISiSdDnQ1+5Um7DXzmWfLfO
0hEFJhVrbsXR3EYG8VBU7XV/GEQ+je2thZ0evmCkMdU8lVdtL+bFzJ0bnxF7mhBkZAK5rZ9zRpbq
1bMSnuBIkElTHEhnqSnX/P+65VkDxAeI7vbL3+A/f27dFXhh0ZH26uJQ2SIl/nBxPnX5gG8hTq4h
xQgNrDqLwFTi06yxqyEcfKj90Z3HbAFtM7Xvq5PsLDT20hiyA2/B0169rViV4Qu9akX9UBashQY8
LHALKRAXDecGdV8p678Y6whL977xzf7TI9jiSA+dtsA61K5wQJb95XE+CMpn+hJTchlKYqXlk1hz
UokyER8FmlQloBbg1BJ16j1ElJCaF3s4JhlUllvRBF+tM0ADPbI5UM/rb0IvuXUucCn6pR0GB3d+
BIMaO8Waj7CqmV71EhZme3VRxZzKSrTadlnBMTAwU9GpCc+ANbE+NHN3IcAC7PEOQjrhRGF3nq2c
13NMpqjY4z3/1MIViXKq2U/O4i/OJ8kcxKARjqGtov0twdhSfJ/1DxYDEu0LSLi20Q/POEAeGGCU
NpWngTKicagNtl9/Uw4aDEdAdMJgT1jHR3ifSHaUF+XQ0e/GB4L9uEJK185u+Rhd93RrGyAkjBj3
x+3tJiOS/D5fnzeOAfkszBR+n1BiTulzf34m+Ao/3fIzwjbIOpHFlxD4oEAZMvPxnWevFgd3Vj/D
u61TbH7XB+yfwtvXT4mW9z5zNtScYnj0Qm1/BbeNYNinPDqY9zm4kBb5PgcZiuvtrSYKgM7O4/WW
+G4iWBJynrC7fLwfQt7bgHqcLLWA6cYgD+yxJ2ReeX+4aZ9HA7rp6Qku1aRPPoJaeRenU2EOe6Zw
YYWBKiPdljpQvoWtXB7Pgr5lA41z3cyOqCCJtxr/z+OO+efolc9LUW+/GyUkXkcAD8h27oq1p3Pk
7l/6Sn1vi3xImLmKqHsTDtTLNp98F3DL3rDSBme9/co280JkC6WH/PuMljY1unxJtIsvVqbj0DMN
XtdRi8INESJ+IbeC+n/QeQV7Tv797nGkCqHnj8G6RL0tOThEKAykbGscOhP6U7Gx3bAvJCS3/WNr
pySXUWGLIOfWyHfkHRctWpvFRVZ83OLW27W/mVL9Qm2oT3NQ+rKh75g3noLUB9v6wfdTFb0KDWL7
RHISlVi8ksGzbdWdoy9RyQdMnozX/1U15ByoL5IQvrGrTSVhaGVQ2FwV0bRBVwzD6j7Ii/SZ5xi2
7AtbSMzfu1d8FpigwZNuqLqKZ4j7Z28WulMOPBKrrB8Q7SYQjO5g6sYJ4dXCJAV83hsSB31SLJW5
G5x8g1RK2rTv2NO+KcnlLPRSi4nMfzjJ+y+h5jX//gaFGSIuq6wlykPb+JLoy/AH81oqCFkYSf0C
/TZQz20bnwf4DQBN+AjXSUGq3edMqbNiPHCw4gtwMO1mPGP4kJFS3K0NzlfSbS4jWch0T0GdzYpD
uN4l+eC3xyeOIFhJSRoSm28/2iurfJG95Gjazd1uNNWG7CfT7W4HikARD5AZDx7OjsCS2m/ABVtE
eW2dn4vMiTpOXGyU6FJ178BRY+z9DZvxCGCDqgkC/OCgOXLsXDLhTOtnVG6v1xiib+dYFaj2hLBz
qL4iO0g/CTzZW9ZlCARl3+Sdq0qEu0WbLHZ0mv2ZDGK7heZDfjJDPCkgFS5Bsv10ree/NhWeve8s
Q6oj3j/jQJ8s8r/RqeEPQSRhPeMd2NGqBIv0ZGYNwmJjKD1T04KDXITG6I7OTj2qHBjxnbaiohtU
ISX8m4O1xowLLILY/o0v1+15z9GVmm0CJ4Z7uI9cBAbRv7RzNsMNHcv3uWlXa2DnPZUwV+AbGbk7
VyckkjiuxT7hht7XuRJqwvebLLO+3vk7rknGYkmBpuZLa8bFtoKYfuP1mLP/XDzgMXrTMeDL9qGf
dS+nTYZUTrssZ2z6njomcR7kYT6T0ABdlM5ssYlmq869RT1oBiumEEz+BmYGpyaacZ1HJvbPks3R
Alcs4zz/01kg5V3KXqC06eD7USlNZcFAvqey7mr+3lP1rd3CYuQyyOa5SuGtVMi1QZ98J0cOnvt6
8mBZboZba4M1a58hNtUW2KU/YhZeW5sRWDA5PmxTXINhoAvYLK3Gt+g9nOeT/ckuJ3qhK4/A6QWx
xnhnQOSlvwqb68Y/RPfiPBgZo7qedj1Dgko/9i5n/phdnpVFQCG55fSUuaD+s9BmoGZ8ywzS8mU/
DwVdNvMAkCj1LP+H4uHMlw5D4asYaYOVqWvSoRBUJ7Bv3vTVIsT1D2ijMwbVK/+9k1QcLbQgtRqm
xkTduf12MOinOAHCAqDVAVao9309oEQKDbGWW8+/UWZK9D1n27VE9Sp+lfolYot/Pa3jHnn11nfu
+loG0Z2aX7M79+L++89RemV+Ze050ClghTPNrDowv1u2/dy+d/n6DDBI/Eab8rodpILbBQca2CpG
s0A8q6uOC6sOwvQiaf7YREoE+iDUmetd1oYgUxjSOAYw2lSZlzKMwKyE7NNu8e54fdmgxxaYeqhl
yHvAHRulvEMbuyLu0FwUiIZXzrGtLWbOPC58k/cH6n1Jb9CRokLWVp4D+MnESz1V/mt50e+Zm3gh
YYhs8rMR/6Av7Mzt/uGfny1STXFo+rEeGVG5fKMB2BQg7RHp3dRLICuwff/32kpdcWyFhUnjViri
ynyiXwoOe4u+QMyXdL9Nu+P+ln8Cx78tgD6H6lyzmKb9+2srOrOSRIoB2a2rrq7u9gzK18aI80un
FDGNBMPRIPpTWPuFSCTYMgjvg1zLv54bhWx9A71tmmwDrUuxNgDv+WXZndcoU3GdCU2LWet+gNTI
aPgeT7lRtiOaC8jiZAY8KJCh2jPE6VA+ALg9qcuYwf4vzm9aiUn3PuF2MZqp2ijPeHpUS5vvB0nz
NJSIsreTgagaLAE2mt29FcXX7gDjMGuTkR9ruZKR+TamT/rc+dc/R/wRimigAcBTg5M2xKl1/H/O
ffChEZWABMc3JcFEZSY8MFYakAaKFohcGyGfwWvIU4AOO13aA+LXvomYptDhPth8lne/E/4DWrot
Flgs6osf2YRmBx9UXsunTmB2ibLOxC7stsAnevbVp57tJ4RVoI1EuZLcUTGAdsyIn6In0W0xtPmU
xiQ+uHU0RSsTSY8wq4S6yTi+P+3vIby+QsEU2VLIUf/JOgeG668dyOGDHIozo8kKorecs/KQrUKY
k5HWfNd5a6/2fkugR5gi8drNempJ3QlP/4uZ7kR8KHpJwXVe7bYD7mZFqUFNfSYJIx2xHfKPZJMe
mOacysGh4pRfLF4f8d1yxSLdTM4eYV9frVfddDyCnu/DeJxRPNUoWc/cpD8/rGUMKGyeoqj2j50J
fZ0etLdFkyZn+s2qleGJ2hy34yid6801n2x4RGRWuQ8NTEex1FIsqHLcm0c1n7B+9dAvsYNkftvb
Iie6dtLC1CT6IL0mtxPyC6dVZ27dysyBXMDgWFcYuIj2K8NnXVDbrhfJawTkbtUc3Mc1cK5blN3k
JpneI6/hkEr3NmN8z6OrW1P7ZCsuMAkTBBT5odxhgCb7qaHXRmnaEBHkB+3J/kGE2OczTYGJtESH
saqxThaDWs/AfWyguZ5nPd9qz0WwAMFXp8WAMn59BKMH/TojfuJV3WQx9dqCdWUyu+6mRb1uyFK1
+//6maoKNQhzh47DG6FdS44HX9d92PBm2aX8ZVUVCS5Z8KgnFAuINkXwXs4XcYitNXWiUXQXHnSY
vJ8TrDZy4mzukVGwZRuvYfQ/KMObXtNFrJIp3JKBeZ0bWLlu3PNYTS9WBe9Biqj/8jvhqLTf6hBh
9tH08WyRL8OsWRUgiLlNo6XADzewg01KfZFqKSLVFlcQq4rKiVH/0e2HHEcuRHXP1WnJFTZuhhjb
zdXRyxaubwJIQZDcL+RTZoTOvalDqxwSZ0lxmvTj2Hn+5zu8g9PD5LE2zutGKcuHnmC4w56eGj9t
jg0qxNGQWcX+9k9vcSMUZ7BCFsAO4sHo/tkCh4vD5HJ9l48orj0e82Snue0+/Gphl+3GGBHA4lcB
xbDxW2esbT00X5Fo5HtN8EWt66W6STBuNv1mfc1sJB+t5TV1CHcJGtC9JD6bGZl99I/wWiWzRqtF
n2o4slz3W1N5Su1Fv7W24EgPoGFuV7Ic1PrEdXS+Zt0QLXHw9K/a/4K76mKLuUG/l7cMcJzpcrpy
efrqlKsOF9t/pqUcqGdNa2K0N1CRDaLwLZwSgYEYKO+2xUY+aUyYQsE8T5Pbze/FKXPcCsvvVujt
R4iWgp/poAFACv1I281FFSEBpoD0qHBuxgAAMqC8VS1dUfXFFxk6rlDbMUOwGE/bOFo41Y8fvvuU
/JaADufX75KI54CtyM+sjU+yj6j117A6Om87jLKlHwqMXaUOBo0pmc4k/kDk9ubz9iNWkuP4pQZG
U2Bnl1pJ3epC7viofeLT0FdzimeRZK3ZFxPRbJCxf950ULElD8WAOaLFQy7QZLZiV4M0Rm49yhaL
/iXG7zSlQlfc4fju9yNm6d1QFwR5iy9aJYNpi5dEDABefz/fAwP8zCg84htbQJAdf0psLxQOvHVC
/82x6atU8bxdgxDx3daoAM21qGUUscVnaEgOLuiKHpgvrYLMfgLVlj+SmJj78fA2mivkqQb8wMMM
qD3zS1IyMVM3xNB7UaUXWjGRo+xKVLCgbZx+I38jEgpQRBZ1/KCRMNtELCcOAIU7rNv0F56qfZVg
wszxJZ6eGZOysmKEXAF7wcOW5ZQybW5KDOLK2nNCKkTJdX7ePD7A5Ls6TM1ocHoXNRmSY6uwAEm6
eSsz8YM+bO9N4Og/wsy25Bt/jtZFpXKOT3CsEDwY7IGCSaYAyv3vC7pAmy3GgnZD6tG1+pzF2T6X
Ccy3BDYG+g0FqZMSmVS/WTGvBvGfgbvRMau7ZOQniWAnBI0N2TRN5+Qv2FHyvCa7KyOc+49a7Y36
3Avrn6RB/ZVttaxmwqa/FSHQzLsYKHROkXXyA+wcdsJuLGieMo+6HQTPsDh03XPDUjwGmX/Jirlg
IUIOrOU834PxOYAJeEg439+0gc+EVvDnEouPZ/mbm/o4bzx2U5mSAXWfYZ94/Uap3HvKSptn4VKo
hgzq94SrznN6ScZIwdrUmSC3I2Xaz+1JMMSr61jM8J0A7QQn1SatVMahhy95FGv/1M+5F4MV2RXM
A84Iei7Rr6cDfuCaGcdwGr8xH+ETPLaFVAHYx83rQ+hrNdHApqn5MJpQGxTyXCKoQz8tyyTxcVYw
pME28x9KAJge7RAnQQ67ZzIKQvGHsLlj+b5Q8fd56kkVjM/TsLo/W383x8ciQrHSng8fpFmJFjTN
PhO8DAd0UhntRwAVcL9s+C/zr0oW+qEXQfC5rJ5hGbOphU76TkZuUkOyntppCKCXxxAKUYcnKoS8
1EA4QMMNneCuCFQ0zElsmAApd9Lqhz1pbMmi3/WlPo/ZgIG6bIlveuGRHPWYCd1vFxp/oZHxN1fQ
UqsCUNp4Isj26t8PxgCZWMbiE9uQSaeFCpA6JyLbbqdO66KcFSfIvMwcK1Y1krVVWxkvEGx4ANFe
RB+5x8dcDTAjmJ29okLVDRf8xyY11GoYb8Woxz+Hti9LlWapzPyxAlf3Vz6EvpbcRxwJ3qXNvkup
tZMLUed06UixIfXUvmZjFg4TbkS6rOF6zXxXta6p3Xy63+tYBimhdx8tISgGlTemV3W0eVkT8HAA
4nUqMLNhZ7KfIHgUneDFbtgNmbtRMs3UyAIaePoTQHJzuR0pseW3ANeN6XKZ9Bn48O+O9uuCO5XG
FpdBcjgeAgd1uYmZLqLwnZUNyqK4EJlpwuygl6MAsazpjLAXlAY1OISDLNgUAadwGxCwt8f0jUva
IB+S2SQuoNLEpJeG2xE/8FDd59ww8CgU2tCkaVxk3eo0thcO2ztljaEEI2dl1TUCoz7ToHUaycxs
aYvVX0aKBa9R9cMGSSzLMAD2jk64rnp18vAbjqIIcT2sGWQeyfM8h400jyzb5uxCl196SMiPcaH/
fcJxG67rvQKuuFgMJvTcftIzGrDQm5xWm3H+NXVb+apUd0ur4Ou7JteWexI1FXA4wYK7SftRUerK
+4FPuW/kbNTSBcAxrBC4qvkgh5X9FjHREDgAlvuAyNIfNKbJWMYx2IlOZGhjTJJnpggbikH7P0yS
PudkVer3qTEPnXQXvMS4wjJPPko1W6aAbg6XJDqdGis9hZEiXXRB/+ibJbK8Ibt8i9moy8zLiN4U
nvvgKtStF5XAdsyvZyUQPwRnSB76jSpFC53UPBL0eKvHr+JjZH/O01Ffu+Nkl019kjRccJdDggAJ
W0mvQUiCHS7icGsfEGS2E87qp51+ln02OZqOyL/wDwQ7Ww8kBVQDz6g1NlUrfd++4hC9zjHtr6FK
iP0xNH2Sq/voBOw8PeXb8XqfdViWTMRkppFVE9NNME0pKWrLPWeBG9880Ccm9DN8ScYXeJj+bpVc
SurF1D773ZWNCBUXooeREojcFKDRYjcmZe/yLGrVbRzUHX6UDTL6mgENYvYozrOSHuihKnkd+fBL
qkfWhY5JArey+b2Wm0ehtnqrpe3uQZr+/WlAAGS/FIrs56GnKNLmykgqLmpmJnVOBcaQQZgQqFpP
DE0PPzUxmUiQxGiYLVQ5rl/V4tRYEznUc/sIRXBXw/u5F82twukdIDET6Ck83D2u7kLsgPYiGTbT
WV9bREtfiSBYUnzDDF0cngICiIH79Aw7zjviUU8igxa/NFp7nakj4gppghAYrczIUTB02PuCti91
WwIs0jqGF+V+fFfR0M+rewA5qvN0hhwAv8hI+8Ob39U4IZAosSkK8lG+sc5BSv3XdcZOOa200td8
0NIjyDGKCCub2i1hN7uW+H7ZGPwLra+8IrEI3/cwJzBQ4IonZILivtqsjmVOMMX8VzyS7MOK5syn
MEbcWQ+TdxJNAaNlPEI9DGmeQEZEN38qNRbozol7XMlKUUjgW747TNE5riAi48VXreqoPFujtiMU
6W/BQ3hqF4bJpYs4JdibqVfPcOa69z1qz1LtHyshwzUtsBc2yuu6ATv3gtih+gMwFQ/2TUYBAHXy
MPjsAN7NWRpB7bzLSNfdJ8Nql6BpZLDn2dw0PGYXC6HcMy0WVpuTPvXQ4aqzIu4L6apB6PaOR+l+
tNV2KCo9itP3vT63DDdWmA4/1NbN5OfNEHLPN1LuxW4mLEmF6h/lxKLNZ7JNnLdh9VGjowSDTOSd
R3JzQO3g2xUAsWZC/ewkzKu3HhluEXenAC9q3bW2AQRCsmcTXOfYITP9cOnoSCQmnLgVk6d+vbrF
pCC7OYeiVRnJJA+eG2Pbe8Bvr7QgzvTkC337YbLosGbuSqt2tTSl5hNhCRIy93mdnv1oNANXE+65
YGqdacnXgDwR6S/pVl23IWSa70f7Cm3oHCwDPgv8KCg2BS0wVHkPwoSmAGlZNX92GC/cs754edpB
6uEr7Kuv/LErE09Rvl2lcJY4LneFYRysByJKn0lVryOBAqogIUUXdKr3yiw9tNH+GdboBrIQ6ZVm
4gxuzWLy6qis9m0E5LliCIetetQRd8Rz3kowXIVvIxA89Yo9M1LV4HHYb8tzXhwUuo1pSJPE1LCv
ysgkp1m/xJp2ihfeJRC3wFFr/EZg2oUID3ybse/s7K/Kr2HZPFp8P6pm3V0Qvl9OwpglvzUdu5V6
rMhhkQSq7AvBuy4dd/b1LvsLjcQfDr45uURHO5KKpMHskwAhtmVkk5IBV3TYdHClPXThPGu2T569
EPwQ0F6rOYEQpWmVeIv6w6zDHennP1ckF1pg+5tpQbzHXxypzSpf3LK20rBaHHTPQVbD71/pst65
le1QAM+thGX3vi7MHnu0n7NmxnNqwNo/EQ6MjibXabzUX200kCxk73kQ29YAlRsKCBHkDh62Oll4
OaMZwD3nCvj3p0KUjycT9hJi1ioHO6fOIbRnlrjFCelaoeq0F/fVq6TVH+A8hgZqQK7lI6Y41+XM
OrvGYwzjD+2+YrWT79cejQThmiZQcY3nEimCn+4sqrQkzuK/Sw4XMaatrtSxH9wlckZLQZyDGerf
ANVMCEp4S6c5IGi0C9pqbV3yuC1G0WnW+IQ7V/kivLDbgAkSmPTalOQJ7ab8OCq1KuTPTMKxsYR+
Z4w+ZTX8neSntcZcaLD4ANbKgKNV+TpITNhelIGtUQs49Vxamy/IE+AFjuS7ASVJHdo2ps4E+bNk
bDIc6h8U4nXy6OHMEiJp2y6Dl0u4f7pY0ukp/DpVBdruXFSt2khkxUYyXpyh3KiQNbl86C1bC6/G
n5YB1pp5xyvR1UmZ50PKSrBZsIQVbQTxUNf7iKgCgu8ZYmHraPzW/RfjOrbhA26tvSiDt8yJMGwW
oOSwqhqfHxvgJTqm52RW1+8Gf2lAtgJ04ZAh1Ubpf1WzJy8suyq1wNvdp/keeYm0KCCVT8V6n7FI
bn5hWG/XC+wY+5dPVbHEHY/LrY+1Bx6xQ1sLnWRzPRoOH3KMdDFd0YXtz84Heb7znLii54u11mxF
o8xXgBlWJ9pqB3tgxpJ+fciTjm6x2DE0x/IQS2vjPY5Jh4+iVbWWHTIqU4aIsBXSDss6zFKISY08
zWFBbEgfBIBnENL+nWcTa1oftIyfnQ7MEH9dvuL2vKv1Yl97ohU1Y5qAujRwqPg8+oOBgcfiDx9s
OJHv63rvj/umFRI3/ON9NJ9r+UYMup9HXm3bHzpSJsnKfzdGpQJNLVuIS/HWY+06EBFJwsO1Nxxt
fUMG7iPoernznQhNgLEne64g2GyzSj7CpZnwv2izUrS2FQTHzbVZ0IIsMyaUVFhuQkMmSYu9qMUZ
0eG497Upffays/mT8frHuc1my8pumy1XgiaEzpUqeuq1/R9GloGQnYqyY8Ly+XfdTu/MciOuzNxh
W665C+cLPDpXRlGtiF0VrecXEUXlaB3O8+k2ykKSHIU4wOOJaJFHcEtEhHPK0P1CuBftqVbCG2sb
PH4bp9yntJetslRaES3nKaQzomm0oXZ7Sh2DnqXYMyWox9HotxYn7xbByTUbkKcO3pwXpfcR572V
+AmmeTqJkpsaGfI5ZqQm+JiDR4/BezkSwDRTodjFGSwrUuflsPsz9vQxcpnzNASUqppoQH3+rORX
ZpAD7WX2BfcyK0mGdtc0NFQpFQHIlxSURcydAxcmjjNzQzG7t6ihIySWWS/q9449HYi/V8TY8D/g
AFCwetNC3v5H3ChwdjXxfyrU689AJKn89CG0DN+plAgqKPbDe6XlAhDAgfaxH8iatvgjTuLowDPc
5gzhTQZPzYARf0b2uOhuXkyR4yZeFGF1SjXer1eHjbKoG7VlgU4ZbK7zzztFk7SVPz6ndn8qSzAP
nwMIdK+Z72UtCJR8xO8qyeCCWlJijZ5p38LKY1iI1B0rPTRwrQZ/Hy7grqwKU4pOXd3GfXMP1Xt5
kCkAH6OpHcOz3cE3twBFSr3VAK5RU9GBXXTZ+bpyYu8sARtN7kzSInzKT2E+oj8FqcGWx4uiS/Al
MzIvZaC0qwBo3SMxgiI7ZztR9kjUM6gm7l/ZvopbttjEc6IQNl2Yx/u6+WmQDiglxltqY3MjB0b5
pG7n9B1I7DLhm8K7kgFmqKrWNHihspYw/yR36e6Y9wRZ4o4mvhCfCMcQUCMomucJ3mLZCAHC85V4
A69cQHCaga9WNkqxsk8CQc6c4Ou+5koj9gK5Q3zXA13K/tPWtyvG7dN1HQcfhBmRv5HnMvX2s+Zp
HOuO46YxFN+gwRslYAcPcae7JxEitKpn3NaObqZV5dmEFlXtM5S4/oSCHADw9CO3mA7enWYEPfSj
wMsD6nqeZg5eWcTNNrVtbs8Na04+wLRokctywZljx4vZWGypB8cfzlFvVFmS2m7uScsUQN1fUXvi
iC6SZgd2MT7K/ci8fUCiKinDEdsyEfB6cYPq2sQyQoOQZSJyJI/uXwjWaNN87/GonQx4gqHZlqIu
g8iL5/hAT+2jly6u22bGTrDHS4MQNT3xIa7FzknZIO1oa7Bp8BvBIH9lApnRqoiO5ZsA5PVWN+xC
DLMptnV280zYv+XQ7HwlJouW74DnuKyyoq9CzctFbS3ng5ZCxhTdGzbgTfvXas588kytIne7Y1nO
tZvKMPFBGK3Jg3Onzy/PuqnVcFW6pjtjMQRoCyH0JWpKb6ty5wIqLxP5dziG9Mxbi4C741nEPmCM
VX7IfLYETdkFSKT5Hbnxh61mTvHs08AmkLykcup4vjm/k5s1gEOADokrsScuggfi90VUfjExNraC
ZyG1Xhz+aU9nuHc/cIDIkZuEw7fzVu047ELq5Kadu4lixvvfpnQKWyShO3g83GJAlMlF+SJzRsZ7
OEomsuMlXu0Ok7N2b1H2t9i0jn6G34m/LncysNWcg6nC/98slF/BsRVpDvugdet+RrTLtDh8eX/0
0cp3vfZms+yJgZ1/cl5a+BDa24oAIraPYhFwZ57FeOYUgSd4h2m6Z4XfAcRzDobzoHsFd8Cdy8Mf
DKjFVayqBZcEJBoX6RhFkvzOY/H9ImainLiSQCHV6hhwrPW/aTwPwNB+RcLuE2bQ1DsozPLdKFwS
Rckx//SAo95QK5r5N0wZsVK+aCVIa4KL4J75vMkIM0y+LNWg6C848wN0q9NiYM1S4p4AIee6lQVa
Q3cGDwUXRSuEyDE1QX/1uMIPTmVF2iR63VTo1x5fe0rx848C4W1U5xTS3D0W6Jvp1XgFgAPOzo7z
9t3irInkHaKSoHQr/lyh0TSv0jhphElMQZzcsN4zmYYHFVd+TNTQkZdh4l7OFm8ZWIbvmgOV++ic
GotAm/hMlKUnOdcGxe7KIKOfPStAn59xVk9vzNrDQja4NdSr5Uvw0AQnYj1hd6mgKzQOiSAwnJmb
nXF6GaMFzie9o1za/s0GpzM77Uzdf9qVN8wtEJ7FY6FAI2Imhc+2LTPkyKDi5+DLDejpRmcnUcDn
yF/IvHPbpeTJFtKv57z22j9UnzLPOBveoxZkwtvjoGxCpRM305SidJRdFMFtBCkOV94/azW+V3v6
Xebcsw1sOqfwCB7S0rbWj61Eib47SUXF1HJ6ou+YuHKAd+0sbTp/ufz/e0hdQIGjVD/gBVUlNtoX
b92OVT2cj9IWc4QJNHgaNqi2sDjpaDU5aAqRGvJBmytrnMZ1YmwGLYO8neMZqqooo6t/XY37yIXH
OsDW9YAyHyT6N9ALfmzi18KAtNgz8L4qb9pdHRqU7hVqAn1ESGfoWC6oleeqY7LB1ykRgzLOGSgI
Bho81vTbSO6y1I1PSGuUjZ4+8td22FzlK0w7aMKKz2J9NHkkvrOs0KgLcNtGfJDZ8+eeqNiuezkZ
BZIwwWlagjJPpp4dHvMjhBjqj//FI4pbDc5yukMIqrb25Xuxu4VZyQcm81pnDKfiRnSDgadL4oRP
I+tFn5Gty1l3sfVlujBb1Dl6k7aLc+7804Hsrv+PBHmK/OYS98FBZYF6xz1hCWDEvZke4F/K2agO
7htgJSCxFbCBkaT1ClX3OGswk1VQAxMPbCL3xQAreRcy34ObAUksECB1T5xIulRqah4dGu+fbRsQ
4z1UB23xvrjTF2JuJ/sCX4eGSvx/SZsuwXE5aN0R0fZPSw0kqUAWYL9X0p7wzVhiVrY/Kr6/InDo
3r+rauZqsBCd3+yyJ/P0RkF7sJutFgnbL+CqURZ750JbWd3wHtcQCXrYENNDGNgTYTiAS5bSfH6d
PtfYmKVaKmCtnrD2YngbzSJeEiRWTldvHxLPQ98Alo/Ga7RdVVG2mTV1epOYdeDTCOqMXQ7JJFKh
TfEfzBAGbAoEhh43cLnpDgiuu2OWAZvBY7UlYSl0wJYdISQxsM8RWUuinAr8GOxXG+LA55Rs74rZ
LR06dNXQmqePjU5TwpUHpQuzT07h+I2vBeiP2j/xGuuzfYsherqRjdY5EOJAnVSkzj/HNZeAbiE6
pkKnsys2F2HofRIQux9xv7BM6QcN1+aRBi7Cgs0VL2DFrgVkZGQ+WxadKHFeLUI7yOPKcNR/SjaL
qfz8P/QISDeKJQy7JPKm7Fow1mEx4rjJKCXlz6V2gzpK+eOlSBDqvS5EKEGzmb/jg+vQ2wB2o/Lu
yD0ApKpoe9KglKcup8C6sBJ6xUvUYYLA1/X3o/7n05gx+hdrfVB8lnreQrMsCqlMt/vPfEyHrUzG
mRuJFF/IGwCf9TqPBt4K3wPHhkmTTzOjatI+VJhgs6LZzXdwDLHaajgeLgrXjbHQdqUeIX8QwmZr
7wI0SuY6mMBG+eg5qMdSpiSDvM97935/9/gzFewagKEp3Q8BKkcPiXYBp7lrSncn4ylI3zFQI5Ao
uWFDrCoRwU1fc/9sOBHpABPbpQvsECqArpaslYHVwV7tX8dZeqVb/bgswzVH+vMd9/ipZTdYSlMs
6Fm/f2vPVEMzOLYxA7FkRRR0hLh2l/PbgrJ2RWgpsx8Q/6zshFORR3GaSwr9pHg8VsHVjRBfFRng
SKBbig1zAXJ6ixiSFmxisJCT0uz8eXUNDQLshWYhpBc2cake49x9tD94feN9Del12WOylMUAB95W
YST3lXIbeUB12LOUFuy6LjdzsZm92QjrhbXuRWwPLYVUb9RT8rS1Rpn4w5L0526Jq5d04A3lUOD4
uGmOEAVd4sL0ojMRjY/ICze50VDMaRNPRtSsdlfiqcTk8OTCMdX0r/zpPiI1rgLGzDMAF3OV6Uud
B/qGviTo3U/72uDD33ardkTD2lKvEwZxBLvPxfHRidMBmgqebjvdvzMjkH1VeRVqrsK4Z6S3gtf+
C9JYF9N1CVn2VmUaCWr9O+YrQp28cpez7eninnlRt+1dFV1BYZwR9354QLx1WPBB3imZD4VapnD0
ERqrmZ6LE6AtpYcrXwz/1VnRrTcL5mLl25ccaNourbX7ZNhEvNqNrv+xnGikHLFJNvj3T+etM4+S
vXG2qPPWgZwEoZ7Aecd98w7AxhSguZjQ7d9OtAXpjomFo6Rn0suENCYGVCygkCGwX3iJNTEdTkYL
Sdd3Vz7zYw1hbb/o2e3njXvH+J+wSmQJpPoKPPc30DjSuMVq/czOMKV2PhJYE8rKM421v0NEA62b
8Ml0D8xn3JpbMZeG7dN0W2HDbVuzYk+xoUrwY+wX4844CWM604SBuzmDLdShp2HR/R16UhEW1hmt
uoDTT4zrWReHYaBaA+3eUQPANb0BtDt90ox5VOz0MjQFV3hyeEPPkz6hM+ITT4SPLJVbkR5IkXGl
OdkEW8/EBQOK2cLT9lEw17CMGP85PSf2BeXds8h7qt9ZCy/YtMxAhBDUb7ej3wnE6QE8rooVHxS0
1FTgQgrE9ftHP0YqBGwt5hEoXN0AvyAup/njSCW6SDJU9bfPiwzqdopMRZxrgsLA7lsUXs2f+SFI
zjScCyDAsCWRYQysJs7ObyauHlwZbYGCc+LAT4GHnseC65mDr7aVp3F1oWOdqmHcl/6xFwFMZtSX
6+q6NYtEaeB4aAmHqHdo0BVtt/zuzcOZPiLBIpJKDc1vccXwo+GfoG6fT12KVDtmkB719iVCzOjh
TOlY5Rl7aVUaECEVu9pet7QLwvj3WmnNVMIzvAAqrwK7CJYdCUawrXY8f22lcmTnXyu2YnJQ5lM3
Lc+II48JkFDZWhsKDGTYwdk9NgxpNAF/p6d0Khx4c9EklnZtQXC43fS8MvHHIFeVzlv4f1r3V7pF
qlDYIrEe4bUmHt7dK0Aii5kH+wHnkkKEhwU21GamKGGWgMV/BOa3vb4JfVK76b2Dx3nZ4NjsTvpg
lgxfFpgfkKRu32Z/GF6LsPtLdmaFqLy8R6/TzPWEYGT37L5Py5+KTffjHII3N3dHJ3GJ1zIF08Yi
/CNT16AuZqqpwxAX4YboeelM/lbugnoIZZ6EnCDN9nYuo9kfloOhBhAiHS2yzuGPqs1vMG78z/NK
jvN9FY/UJsnGZzLlpY81ECgaQ2Cp1dTtmgkkhtzcsrG0+aOYBrNloSs7NnCbxhXbBSWiMrKC4e+Z
CPFx/PFu5H/MhxOPZpsLgh0qV4Q0Gs1X9ZH2Ytzs/rsV9CyGt8z/3kGIs26XsodmQ82ysI1uf1vD
eM0/XGe/YpFmNIh0fGWKCwbGQ0amajEVnwIzmdCmVWuTioPmmV4zbY0X4h6GHNDOlBzyeJi63s9X
u4bes6iWrMfIL4kAidVrzXUgVmQspzlQahTF72/Ews0wXLEkRmD/B0Z3kuONLVJKa5n3olcnfwrj
XiJiLs7qsOYtI8BH/B3Ah4AhvWgFl+JPcrvGKbDw6aE2hUsGaDxufZWcag9o1qmuRNQUM1yfi6Gt
3Dvj5wC+eWF4xciPIKLB37PwD+AV2D800QqTYuE5Jt9pwp71WC53lQCo9iNabAZ3lU2mBQyZM45B
0AKlZywr+ZN8xbLvRoQ8/a0yNOJDUzszcajlcACTLQsE0ALmZ7BrBdVFxLvaIO1Dln0h1PPdThdq
5ay/wGy+aaxYLpu6tE5Y0WO7ncGPsVZfyKxliIGK5/5R7mCo+zW7sdIMYqERUcayF6ipLKiyosB2
CYjXdykrH8lxjvHjq+4tlWECejCKRr7dy712uEW0ey34lGbqEc2TCQBVjTYWJzFLaKa/NqZ4ZDCH
PE9C6NsLXqBe2FsxE6/w6WNw5SqwHV4L9PtckJeUCszI+ID8SSJkSF8vawFmsA9j5pTbtiKoCdMu
ls7JVMxkCN+LGxtJhH+R/lRz6Wn3aIWaoyZ1AX1g0SxJqT3BUIfBlVDJqe8w2SCMyrRaR2IF5SeL
lKFKWB3nnQXPHf2PNxADwO/MQLznGxdTNnA54IkGq8ibh2YZTotazQmHHJ9CYn3ajchlomE4RE1F
hg4/2rVk2qAwn/J9Y+Q33xAk5894I+0S1hiMHe4bv7JJGDSdT2duLHh/adjIRuyQI1Mfdwdc5LoE
dKnWL2gocrBL8NSJSeRHQPD/7FIYXPXnO5J4rg9T523tJVPxDy4BZWou8I9NYLqkBSuw/WLfxjly
wnb9EhfMgGZs80zaxle3UTxZn+lMEADdzD2nxNEbOuwRmBxYm2SacJg64l5PmDKdmBi+7rGyvpkd
C4gyMRIx4ML6GRu4sxNp9rqBfcfFfLMwyO1rWU68sKT2tTnrQg733+iGoQ8mx30J8W+wPYB0baOV
ybqmo5Qiy/bxaALrxCSpT3QG60fV25DjE1CJ33Ap70gXENef3LoTHk1oDTuaSk5doxbqxLz0A8Ru
HKTQzBhVIMwEqrxv+/QsYL7C15kasWePpTt1EXQDEp62akD5hWnPJdmxSvA0160ODHH6cArCBtl/
/27yyJmY8/NewR7mG8LH/O/jbhc4yp0M3ALp95EVHmo0Q86sN+pfXR649ntKkuT4ai0gTjhLHW1B
zU7xMq8wgj0mGfVoW3fV+NSSlLdo6W04H1wvnvc/DtqZ6NxqqwqEexm5gJP4g3+4tE72x0394Clj
zYYKvrEbbJBTsSSnFMJVZ07JCyo3IqlHXUItrpGF1peeF1slKE8MCoUmqDaJ2qU9+nQP2LMnI6gt
fk348mdrQuc1MLIR2Kkik/sRAqMTtjFIPMepJRseT0ZQbt2iB0SC98ABmxtKPp/GgmaVPkaQqiiC
CPfKEUKayfynIqwJ/OxhvM3uEKeCH61ADbwEficx988NNUYV3vOSsNeYEdloz7B8Kw2t7eL6L5jb
NyIZRYALsD8PuPMKaig5QRw8sQ3nnq3nT9nYKcOqbQ8j/+X3Rfr9mYNUujNCyP9SCWIHfsTM7xMo
u+CpCnCIdWYVJYyKETqhJUzfoRBobvPbsajrX6jThS/MXsx+S9lwpAlf9vzEU3V2gNaTX6fpYuRM
BMfMhJQuKQpxrtIiDgbizvUn1KrZ3yw0ehfk7pIsiSA8YTC9x+viL41hsEmWdDy2jRr8JvDJ1K83
noIrbMO7doACtlDoe+IipIlKc0S36pAUiJpciruFwV9C6jYl/IdFNaKzaW0XNoNa2iLffBJHHsrg
nIPSjp8G+5T4dppYCB//9MvpXnLBl3ywrRr5DJSwj2oZfGADi9PUgD84Bis9G1HaEmSVINRrS9EY
ccnri/vHS4ZQkNW6dJSSrvTKMocYsjQVZoZCszUSA0I3veUI/w70Vw39Ew1Zr3zLJHVaDJozcyAt
s8wDH5VbN6o5V5K5Nv54z6yiL3Rdk4AegYUxf2d2RX0vLJYeoaO6O3inZ+aMtJr4X6UmObj8O59i
g0GYMg04i4RFb1ts9VM2s8VQXGruyfQhGsy8qDv3Y6wGpiWxFU5PIyQ8VUsjqZYqyKzwft3oD+Xf
DAGe8WRbF0EGmMC70e3Mes/p7p9BnEiYtr/zI/dhBwSr6zkRHrjGDQtNh8aChVpx+OZoXRbLgi1Z
CMGy7S5bS89zS7gaCzfWrozqAdmYnUykqEmK/Ivy25C3g5CG5d9JRQFPK5keSQxaUn1lRljAOnB/
haZbVMT+825teW3w9q75GLR9iB5sLY3cLekHi/CcLBQnjcjlKh4zj1CJpqaXt91qQf/xEjfTPU/I
RBuGETrG5h76dkwVXnJCpt3uFSuUjXhtdddqKbtwJCmHSoLYhR110ulIH94gjFK9/7d1hP00fnIp
P4+TuWRWMXhP0EpE4G2ZiQD6D8xsBeaR4tnF6/nZ/dJ6+jeFf0FIijr5ZcqCMOhPuC6JdspgA1j+
RsPg7Sf7bOFlksVhefwcmYwdZS3QauNOLEHLiccJDPE0iOORoXqxSEAA0X6HZt1cc3apRKNljXs2
+oTxSKJzyUFhQaQH9MHnURYSAgtsfOmY1mLU4e1wuGvj0Ww272m61OLRW9f7dYe4A2r7p75ptK7+
3X9ogNorcB45qFTq09Pay+Z3LX0jYjJ4+2I/ThJyXNn6YjBrHhLI2t02ckjJzKsZaCFHE5JSGAYt
y5Anvp9xtJVPuggKOvaAL5TwL3WHPIWGkEuBk+yCOwbN5Zku/XnyR7PeFJ5PFncOpaQz23cxnFyc
SWyOD7mzZZ+zNlLaVhoSlNIOfRXWQsuL7fzyScZ7ER6sUyq7cR0RBmCG+Vck4a27VcnHZhBmuXxY
IDrFttHWcVZ0Jjrt72BvTiXfBvGyTjSD7sp2LfGx3zauDH4oiaHlwAVrZL/UA0hqLj0LX9EB7TLr
5qmMI0et1ULL1YRErk+KQpgzF2+A36hEvko5CTDdjCn8cjppFrYuC+Hv3heV6LBdJo9tlgwWRZQ2
W85fKSTN7Gtan0DBhFqLZYHA/e0Nga/7Lo7ZbCpNhT81FFNjLa8TdBEMkglMk7FerPA0I6DGEpev
R5LhI12mn81pZM1a0ZcaeStpRtYWi27B45NGQRG1V2mmNO45YgNBmLzZK/3mXYvMcwjdEu6yv6kv
3XsNmLfZVfcu4nwWY3m68ANg9rSkJBsSrf/Q4Qt8COW5nHtrcF0Szg3OT3vqqbr8JoZ+vVR8fSqT
86vkNQXYfsYvMB7+eF1MbRcKMO+zgADPrzYC3zA/40zrFPjeKjVAy+tcc3KeISD7ilzyBHoXVepy
yq+13bhoUklBA0YHloTy4mznXVi7XQ6vO+2FlB+DFyp8oJh0HTcZzRyijTATSMg5J90vI6YUaVaw
eiws3vogfd9FTGmNRqFilWF1mu+gZcODE56xbabO85I6rqMtGltO1W+nGq6AED2H6/Tp+/lNZDZG
zRMv6QGxF8cmR92CfEP8GZoj19aWBHqqFV/wQXpffg4YkItqYQap60oTp+xhueX87ykgAFBbTNXW
666LDtT5QncuOKcEJP7twgAKOxExeI6eqgb7ULGyOOI9kKuJjtlpYMx2aUEqCke4RQ5flE8mM2jr
1NibhQ4Bp26Z2ojhTvgjZLtqnbRSXegik9tCX9GBJLA6mvOnqQnf4zk7dTVMYRj9vYxLtcUpdaD8
Uv4Gw2wuIWZk3law94+ME8l4FFIdyPBXXldgUBlgrbAG4GSwyYpc0litT35KfUCYEqL+LtGFR3sG
TCWziWcgkD3OESZ8Zm2KYLshvjOuZc9yjGYSfbWCp7sJ+lGdUNnLBHP7kykUieinwGJEagmqId5n
4V3eJo6rk3VmfqlQOZdTajXsFpUoTdC05WwYpR4rpDmdo6cVq9//mh9vW83w1rJZ1jHid1d6uNJi
yVP4SZYego5scCgl+Kfv47+WR9J31ynwVgd07iaX35AJgnhIatTHgCy+DCKP51UwvAA4tlLswtoC
P9srnmUvSCL2E3Y+oa5BZ4AQo+PMSJKglXOb2Te4m117o/3PKUR2Ry+QUfvP7bnQGPKl3ILKm/i1
v83eKYkJ4vJaDT1C/Zre3thmk0Cg4m5t41qe9rZvTFvU2cPK/SZriwjh51jARGMigU+uT1OKI+sD
iyGloMuLSGmKAh6koGMD6nqUsmbBQ7HzlGJg7Zwm5lm2R3+2sNKoL0LhYTtNCPYuOzXT03Oa3Afw
pfNl3mPIiqtlE+2exM7TUpQt8c3mxCUTvNJzcTipjOhU80WbyOoytev7ewik7KAEHWyOO6/+mi9v
yqWILGtUuwaopBOJe5TGcrP0TNLPScUMDFsaxYBY/rvhDDMTmBTfGN6+QtmI/Xf7w9hih7vBsNBL
snWViVEOK9DFMcXLocTUEHWygz1pzOM1tC/tG7vneXtqtybxQyd+pm0EZJZucKEbs52wjFb3fGbd
DZW3YsnMqx4YOk2yKAJIwt2tUYSnmSrY40eii27ITWhz/QTEqU5l0/8fHkxJEXK4u5caakoL5csH
VUi7T+26kN5yzDhod35piDKzb+RB8FmSZ6VQFSBWRPJMStV7Sp8rnEhy2cD7DAfHJezJmfXCyUWo
aDwcEntzIUjR/A18SdWj/jfEd1WUO0zwlJ+OF42+JnFTl4zy6VjXIRZ8wxgaUahIzDLh+k2XjyeT
FxZRMeuFMGQCDQ0Jt6NfRARDEWPogo+5Ia3ixwvctVZTMV93aEgfavOk6hyWPoHhP9FSnwRVyWkS
sJbG7btRR/GUlxi0r7HOAJI/IXiGXNSqzwYpHw/mFJVi9D3zTwJ3HaS/WOD5zfcIilfiTT3HE309
IiMxbgmQ4zSJlMVF/QbGG/e1CUIzhiDZcmjdht5RhBMDh//qRemT9GoI3MotPW6xcudyncKzpLvQ
Y6GgJewNVJdND7pp3XeVUdtrJHesnNh0cMEXaR7ObbsFO96hDuY6en0Gp5M53vdL3u6egVHM4Ysu
dpF3+RGnIwoZZzuNvwomPOAQSbGxcUqQTkpHK/8WqZ1jVrc+jloYM6q5qd8MRNggg7D4CfzP/EP/
LNzu6zyc9MdwU9M+NHinipVI9s3I2m63za1wTPf9W8RG+RhgX6JD0QDeWdp/gatmO1otMoBAl779
CRlPFjnBTodNJR1eZ0OfX4Lw97/PJt8Is/Bb6Um2VqeW9Mc/0/5/Rof0gIr6kynQHq2cUE417r+O
JZJmbUcTwpQGJbE7Ua8ZlMwpQKGFEaKDmnKrV9fbNG/cZUuZPKRvjx+6Q+6EGTiK2jN68QPGmt99
I9JTRFqmzra18bHy1mOYJhsgzAJpmuysD9fuOD9QtX7qJroMxmRy3BWuWax0ebj/G1sqWwfTKwup
uZezWJ+r3t7dX99PesxElwGf7cap2hTfrsrO6SD5zd43TV+9YemuWXRubAJD99Vxu3LL/o818Jrp
xVz7E1ynm1NkAc6j38vcHBy7jJ0L/0xP1Uu0mCI6vMpHYlfUpcIpgPMyt12pDjkRQSEtUoE4BG8I
BbQjWPU+yZWePUqWhemtzYEb7AN8MMQFwBekR8ZqIZkZNjJz8MKwHowiIi8GpApSVCV1gz2sr8BA
eipJHlYzR03xTSCTQ1vGtkAPGW3nw8cwLtuVIfqHV0zGO2AbkfGOv5++LVhP4p2d2HjBEtqKEioO
F/14abokJhQqGGZKgMFCjb5jdJDyOFiesbebG00gSegxuzj5bCvTOLRZWFwZObGcMU2UxIPYj7Wd
srUtODxlWGYY8lVVyC0IhBpwUCB5OrFXbSu/BKJMuaj9tsr9x0hz3jMdYdGTuKoKcZo0jPQL5JLV
5BvqKrV9vfsNe/UXdCh63PKidXZQrdjECUrTP1gzpy5ETNINO92WqPo+r9/n4WeOKOssj11XO8us
ETFrHqKJ2wsFk/hwHMguUOqkhWbAQY9mZwy8Q7S8UPbtVas3pC9jFR+//nqg6bLgm8HcJs4rEfHe
2tXC1wN+eHnbXZgmk+CVya53K8txaOm5mS4O/4oz40aCB6KvCyQpSkJqYA1G9MFGHQU8h2otG/KE
nAY0kZ4YWeMwdp3IIcBlmeQEe7Htzv/vZspikXhSJ4HLDQDxY8pBQGCqgqDx8zTOTUnUtZwwwoRv
vc9eceD00PwzXRZf+5kq2zsLb1T/UoJkoz7BdqTHzE4AXqSrXBOUSmonl/zjEqBkLmP+il+RcZrv
rLnlZMo+JEOmFmBPdfFTZ3Hn1RZne6WGJsN84jX/l1cRzeN8nUN2+fgI0aEXhBu7Chn25ue0qVyH
KwuxMg8ThhxITOplBLZwOKNxgUtz4QmfuAJKvqoCGh2CTgGS9kOUQIjj4UjG3zCSlH8PaTpKUYHo
20yXw9Qatn6cDD4zU/S3wvsBkZnnJGEvtMIu334j8/sEO5vSDRUWFXEXPQ9ZUWwxcrWIv1X0gL8B
Eh3i7ox00SMjujfzCfeB6JTeGOUP6E05ebSqtZaho8OO/uGCnF9lrGGX+g89At8VYjLKbYu1vc6v
ADpgPVTWo1vlZ0d7FUNXelxXnPz08612v43+XCDQWNDTUmB46r9cEYTVg269UG7EJVRDsSX28TE1
AuP769A5b2DFTB8oW3pKDRaKcFEgbzMZKi99nRtT4nfJk7yfLycjK535j40zId+0xug5YVDUyXYN
e9B1iJD4cr5uME7Azln3JzGg41KWHuA2G96FM7DYW8A439iNSG7IqpWKadat15d+dhXXtO++d0kE
ZVzpuZBLh0VIg5evL1BQ9FkrDKGlXvs1qyCjjDNc61/TdPoLbehRedGL6u9jz9id0yGuOEyi1rVB
3OY8tQBwgeSwr1VOhulGqI32P+evZa0EENXJF+gGBqD4nMHhWVPT6+P+ingk8DHPWj8JcXyyhZO6
DSiDcEru4SRAep90w5RoW5NFYIBKm3fuvA/pH+XeLzHgtyPxmpj9BwcXZ2RmXq7WMIS1/mkv5F3z
uhEmLEy8lWE0uBk0wkLTqDpT1kQPC3zJk/hsaIcEkPLkAvufPbedaBrujB4WTNhymU2yii3y/6yG
0wlJCpMjIuhE3K7+orgQhQJEo0RDSSh1/5Zo5WYU2Yi0QhylYZvuZz/4ra+ELR7OAT33Z6T5Mj7q
rnAwe1R+L6dqa5BgxpIpTosG3zOAXxsZy1iTf2IofOoPFBJE7HOxsyuMVk93P5TmbrpnLO2e5vrJ
1D5VvjwtHphKQLS+OnZOLxo2nPxn7sD/474woCgHGPIH6bc3CZodZejA3qSaD8PyvvVdayOTq0SJ
1AtUSMiTMDlU76961pTx+gklMfxgSNiBjux/B3fg9ebuKnhctdnJtvLGDk2uu8fiOKE7R24MrZu/
iznlhJH/ITzCb53ui/Kbt3rdeDVWtF1zXlmgBJsAsHM2+bxo9HrU+xwsh9nglz/bnId7PIxH3WKL
+wxQN5SyCio9mvOyBcBgoalBQDXJQBx1SxBtgd9IM2AmuHY9MO44Wi+HQZY80k6EMd9H0jyZCWmT
ZLJFvpPvoVmZONDIEm2h1C4e2vrT5hqosqaFbwfQ7OAowWlwPNk80Q18TQGye8g2CRZMClmyYgdV
+sAEZZ2tIsTRRWhQEWOpIig9LEYTmWNRb8Axs+NK10jURHWyIraDDKN/ZoR3u7g/Uk+Vod/UzEsr
uV97GMxB33yEY0NdLvsi/SaGUnJ71IPqMbPtOufygIWCvekOH8m8WDQu6NKW0QJsQXgtpZRf2oTw
U3OAvbNTyPptgMCXTHehea8MqDjB9LNDM++b9jDItl0cUARi6JBtff/xVoFXA4/wz7GFeVFUC65J
/16sbckbgJs5/KpZ7SQlCLrR9jsBAHhd1ev0j4zAEZFQjEukF9lSlEhw7qGtrtj6eBRuJakJEGxn
bvUUO2uaI067SKjdw3GXui1RqemYs568nWei81tI0YP8HDgFSAtYydqGHlhCVNHl9Is+VLT6QrJV
cnsgbB983HCi7DyHT/FtYzYKIqez5HP8PpMxToQRFfuhIGBEB+3aPuXL4IV/Z2fGOkvB2180GTjS
r/qUd+ClJAO5ax7znVYN9OXo5WAxBeMCvjmAJPXEGywmAPD7KCrA4E7F+zWO1C+SSnvssIHHEq1S
kTf7zQabmz9RdilBo4URZk2GUt7wwjFafgryKUQ8ntwGNJsMOLjinjfLqvyuYhr0KwFl8rWwWzSj
2llPTGItr8pGCuKo3VjCGuK937Ob2Dd7Hbi/PA9X6MHsUYxMfUlS0wq3M3hSjUjS335hJqdnWq6K
7ND8UeDiACer1zwBnuUJR61uowJG82yvGZArT4oJo+E1A8/pPBUqfU/T+T3ivbPSud0fchk3/YwF
zIea0tKPwlJjakTnSV3MJUM5d4/ZQ3bJQ1xCuJSSzNoGxoariSJVt1k/nmw07bLRsqg82pOXqTU3
agrJUBjNgy0d66dPzzb70h/PmkLkgdQEM6gZwGBUATRM5WNujfS/JCPV2dcludVugjS3BqeLcRd1
YbCn50wyfAlqnrHNogOCEfzPgPYJjPQa058oJLX+bfm00+IMOcGVgWrsI4CmRGbcrZ3AejBPOLL4
T+OiUIiXLbf4XX0IkHBrYNZVqRHT7ItANwvqF7lvYtVB/1PWGXvVOrGY26tX8ASnMVfzyJeU0IYb
psK8ToKhGpy5oiIiFnbfKqz9pVpI+og42BNelnacYGeBXXRCfqbqWaKSTZpkYxJmWUcf4/FIhYBh
1JHNvtjFShwd7mwAH4gPqQvpTKrnyKfSYfxB/+q2UNRZjoZZbzMYr7k/9OIjPOWQbSqHSOp/RAim
MtsRj5reD7099l0cV24ZQiOrxWZItRFI3G9a8LtTvv7PZTqQLfhw1UT6DsXi2+VvoMQlkZX4lBRC
y+ZL6JdTQpXThjqhwSdsrw+V6E8vY4ctHOb/ZpOeXyNr0A3+A9ApjXARSNWsHEjfMUxnYOJh8Onp
wh8eJEZZYlneIH9oipEypn7kK0rkKWhwJDoev8jdUQZTK9/CWA7zGbMxRChzObkF1cfYcUPtm97u
MCw5GooYf/4lQcW2JC0EnjdflNmB4BPRJrxY6TlqnbTwInZBO6CmyFP7XoRP+zXaaH+dVs2vHGEj
SaeR8SAtLT25W11XFxME/RSRb8m68hb2w5OplR6QwCeWzqOM3uU5kL5NW70EqcjbaOfKvtIpt6aJ
3kdDtQwX3mDVWmi1RDnsppdzfzUDVH7woe5/SVaD2BiAewSWh8OhLKd4iS/JUu8MtaAJPu3fNfUe
3QYj/4oUZWXMB5ZYBy2KvvTe48nHlpFzErkrHEFS7kUWMAd47/krfMxQYgnFrvhxoiTsVdeafRUb
6njEH9jKPALq6gpK1YfsuK35cpR0Yo9cw6K6gTZISYNU/nbJNHxHrO2K3vQxW5CfA556Pbgv+93P
4w1EKjRjU9W8aHySRBZaU5kSf/gNmXK69gJQAij2Mi5EQvV6zwULurNOSNrl9H80sik9/jAlR43M
B+BHA0fysdVJe6RvS/T2YwM4hsetkxTclDTIIC/wDXk9eO7tSOJjs7hC6ZZ8cFbs3ahrafaIQPt1
Y9DPaMcLxHNa5Lq/F39vZmrXE7BSLsr/kUros+lQHasUQdOuDbV6+YYx53mjEwzsVZ6SR7cgERe3
R4A1w+iXEDHo8V7cmQiHLb8NWE8CJQwt5Y3RYuDims9YttTlzCmQ224Jh5MnpBDuB+ekc4e8oCmG
ZVu0MboBM2zZiRR/QMkXsXmaDdbREgztvXPD8RKR3AS4tgfnf593YDBM83WtVIS6eUgsOrWiVEJk
yWW+AyPkNcRMz1/jxp8DC7HonbPAFw+TMf0pkkZDEeyyLSA1VzxlJRd0knmWV94S8aZenuTbBNQU
Igd36PPWx22acn8L/2GpCZMuGxDt3pR2bsDp14gFPzdLpxg2csQ+N2b5RgjcftkC8SfYP2eIw1Eq
RAKzpaeZSrjwI40yCYve8xP47B1IvHNc6X6T+pSThGllNGgGSKbE+AobaezpSPn/ZwsBncVWmyn+
aaKkU4XCh2vbomGm13b2W3wH0EQCm2K9mUCkziTYb41uieYZpZeX7ylTmxSQxCqd5BCguBqG1mDC
Uw/f9PegVApEGE41U+MCicpxWpVZ399vN1n0ENDCQEkHpioKFRlTQzx5HmJMPzv/V2DIvg0vlLPp
aK0gxUeJDr9rqwGUAnmFkWmgWhQcj6pEIUJliyNTGn6iSdOdzugOeBiGv5ylNb69DsrvP1+Xop5v
bTlhNEdFc+uaQLxSZ4IQrx+soRAF66weZH5kgBT6VR9rLKvslWBGsow0Yy6Vb2AF47HhUwqPbJst
iAT+D4F6V7rZn+MfhDq63GbTq0EeJ0BvxIDwGq15f9ESVy+DVriL+QqnN9gg1LxJgW0H73+v8BBR
rzdgH6+ADORdDG0rOPookq5iPS8LYLZcWNJzD7JQpDbBRoGoLCzhTlbRlzpSXrWxExlujTJQP5eP
WPgA9xvx+QtVV2afXR7E/eKANOtoPkjB+x8KKLdHUaN+wCXMjHqxeY/9c3FYgtL91zsVwjXS93cH
/IigXV5B8ZJUcZ0JMmhboTQrdAeP/qswJrOXGxL8PiAMksA4bjkzo8MXQOREjypdVFfSP08OL3w2
7tJl1I6UCjKhUYITJQ1MrvbxIdt4lvehAdUUl465Tfv9XI6g/CVnBSZrjKX0YBfUbHoIu+t/933P
P398NxFujMZSR6TD9ZhRCbdno+WMpnqlLaixYcoRcLlBJjnN83NLxxFId15wGbjQydU9u+GQry7Z
snk2trOasnKLIacw2sa2UOYYSBdkyuUlS+iAG5ZJ+sF1GP+iyKoMEAjmg2+tFZt8UUw0Vpdi+iS8
Z5KymmK5rzDcREug/D4/Xuqktur7LiF/0NieMXBlXnaJTGgVAQanB/qf4+qUjdiyr6P1qeiGbQRl
WrNoV+/XtyVQySSQVxc5UpTs6QWlP7qmHuS5e7LHcSYWYjZ4HK7qj2aINJPL0q1ZUjjC+g5xaOuq
brUpf7AWrb7nWshup/5O5qCAIOFSrrBcwWDHT0IGHlkDf5UhWnyOJu/a7/kd/UXZ69r6UCe+TGqT
6M21VbJV0Q4afNS37739MKlV3wnLYKUzSmzu31Lkt3kPLglGpp/J31MpJOyq0IlTalirIv3v7RcU
7FltWuTnrDB0gXsK7bZDI0V+dYVRcrLV9CsE1pgLUXtGeg4ISbIfDtsORvAYCirb9ondZQx43D1F
OMo42UDQmyhfxbC4LmH8ut9tlRcpTaVZLt3Lidlim7aNACMeugt8ZrqI8iGqIt6b0mFD7Hd9xlNh
dWpSo6zH9NDa+lMIKKBIaiFbN3yjd75t7FsSpMFF+vleaSPMwX8RHlXZmNPjpJVvYY9QKZYEfLn+
2Y2EoLU1EGqiidPvfsJHHzRxn8PJKOWrViridKguffbU4s4y6/QwnCZb6KXHx1ltfoR+aNwPQB+v
agXlBndNRY4MOgPBSyzTzV5YoMjo6kkTvYmfZ3mwBQAolxGldp+Rtme6yyW8LSPDWPsKk4T09k0X
sE58Xp1rh19DJdKydPGkWurWp4p86w4hkfFx4nuccEjS+6z8f98UHVsUbQlqnzlmv0qv0TvkcHqn
GCGkw7HLlbTENvzqYkT+WyiTVAuKc/jxEnDjB+xaAWZCYXfEWD10op3t64CxWxe/ITyjQAA4UdF2
wkxeMMCKK3qJ3kIIPeMMhr4ZMZe3surjGhy4d7HmDdT4L2JsMx3mzoytnpQvjYs6BFoocJRFO5gb
O/v9YJiKmKFt8jnlxS/6oqGGoFbcS+9Oz284gj3Ex3er15OHx+qrhHvj6B6EznsyATbNtriA8RMB
N80xIU1KQo/6g2LOkoefv+VbE0fc0MQ4PoP2YzvvV+ygK4LDGwg8ovDa4C/5kI8XMegHVA9+pPa+
bJiR9o/l8oXbSh30Yx03iJCp1DlvJyLBEau57wEz4laoALVXjJGdA1jYrcfwGSdJyuuYJTqlh1g9
vtLSlFdlu7fQiAqsiiyS5PYyiu+A40ZIYz4V3zqUFicZKdB7yYKiTLWUGID9C6FYtaA9ZNMsvz1t
OOkVonptlo5rDXoNL9sZzmlj4aFyH1VkRRJnOz+8/A9GvKuT/0OoqAUz2UNLm2FkRh3hC78U+UMq
+gVlnX+UlGf+1N9Qn5jPMuu77EbLMKvF8yiNumdDDuR3mKI2MkAJkfIVcm7/6WJ/wdTDl6mle/QM
OpGaZX01b2Wx3pr9dcoueHAZMLb6++4ZaD0OLPU4HhAUk/e3pQz4xymZwWXQhuPbr+SCeZ6xzYLM
/CGqdPZKaVVW62uNbnVl1mNanTMOp4LrIkajDnS7J8AdCQcQCIPfBh4PTKmEzLDjfkbNiiILUX4L
PqhJtVJ/KFcVEer0FVVXzNNOCypr3ZGlhysjUc5H+odp4NxqIRixe/g6JNaXDnjhUMY2/Ch/bgQT
ZAz4le9wtBdNNxi+HSO/klK/z1YK6Yd4v1yfqWbFt04A4wsa3vFmVZU0EXsATd5hJh8LV4RX3p04
jmz8LDPd2B5cqwnh3Y4SCrNG+NKlJcoyVIE4ovk8w0g67PEnv241OK9OTxp4+mjyO7pogud/8EZ3
IR+Y9X+Gz/W6B1a+PwyWI7gr6ztjHL+ENCLTWRGu9VA4nI/28q7/0GaPYhOPXMbWS+Bxe2jzMbk8
K2nec29bsLi/aOqX4ow1OmtmPKDu3b1gjXnLvr3GBdn1bB4IgC70aCjx3zhDDRzJtlvzRoGGZsQO
l4BaPiZ0MuYkKNSN2Q8DX1cDD8MwfvM8h2FFXyF6euS63MIFyvYH35xfDBbpwiO3kjDhBqVz+ZQ1
yIsGHvoZKaD0tb3nv7I08DDTMne8KpYt8q2nksIT91JU9Z1DrghCa5id6jAqJgCHeDTnaRkAR6oF
YW+MuGTC/uAy8kukpasPPJsnhJG8ueYyv6i0my7LyPt/dItWU5rPvtaPPXXJP2KQRTXvKIHFh4oK
a/JqFsmZmZiFbtbDSbW3xhRh07iBcrK37UvaSjHvAXRzNLz2JuuFPhuveD7B23PbvEBPiuMF67GP
HnYKPRUukmTMhiHg1rDcMXk3XtGr2NwOmuIs/85PEGOtMY/dWghHL6Uu/5TSWVZ73MJXwp1nsK6V
uR1hZBe9ve8kVub5w/VnKpYWh/cxkAq37cvs8mf8PefXTGwDgVLN9BzaN/xofCIj2jmKywu8AZHS
A9NdGzB1gfZtAFWeoEnktIbnHGxOQ4eYyCp65k87/uRzsHa0yy7LpNbh+uhHBgGBZUfs0jaj5Qss
QR+K0021JjKefbNRm3Fa3etOL25J5TJSfWkqRRJTSgP/924igcHS0yWMP9qh/LAeF0YOL3Qvc1df
mtiVdKsX7KmsUhjXz79PiNIwUzbywyR1BEzE3MRF7hyVvu4aJRL8Z68Ut0G4K0VdJOB9bgG4M+IN
rZIsXqhZ5odwhkAqVH2Ai46zLsQNOzLJ3BMoOAu2xHXhsLPjlSBjNBjQObYlpamQyO7s/uwEwIqy
d0//X9WQcoT5JKZwaiBcvs/k46sQdApht3t//6IJRBS6LVq6Yo3CAPsfkTKw6R4w5tb64NsIolqf
GAytohmJnRNAaTl7u/2qHDer5rhRyJfIS8+rfulwKx5ObtSkL5ue/PXo4mqXR3CJGB3C3ZgBxRkk
Qp/PSTiEZfTRERsO5ot4ssfvwU4cvdxoazp/kC+NZ1mrE+SUaAjL4zVcznXsa3FP85ovzMXs7oW2
G2nF699Twm3EOTsIOqhIDFRNpdnHRS48u8X/AI7Um8NZp3WIHMOwlvJ79dtN2qFxHmXRmIiFiybG
OxxttCkxQ3k2j42sO7psyCiONW/DeDduXQqexq0fE/5/poX17o6k9Ic/5szREtmCcSYyCgnB15M1
aiAR4SIt1rMO4wut5puh8hALY1+d+XHJmzW++LDrATa0n7ivjiBll3JBLKKx67rF1lhf29Tk+Nmk
JdGOODUp6Ij/mbD0GYJM3YqO3w35SGL1gPJZPH2LyZsdOCwGnE2p6F3v9tQyBBtT1U/U7Ryg3ZDG
FH1YkkV8aXecn4HxbLOY6iwg4wQ34tPU8DSbmMVGcrgKVvUyTxIfUahLgzZP7T+ScPKL1o0PRaa7
zpSWikhMBRnzk5oV2TPNLj4q6Vp/FeMMRkMRbYHWI+oIMdqb+BRDYJ1SH5skZpLk7oYfZ5iFU9PY
iPF8k4DyYawg10metfQcZkF537ZekDtuBlE1pR05k5yDM0d4MY5Nqkjsw0F9X9VkVgnZCxoPRXiT
oTn2vh+pk3bEYQ9iQZV0vK3e6n6qJ/8uNs1TdiOXcEVfmtGhFOOQuxxzLhCaIh30BlXAgG86tSm/
xhcxW3vdR7kH8Xt3GK+j+vAU/6guBgsrOTd0x1I2jdPnReL8qfylhCkSON0vK6BeHtP9EzmO9Dym
XnmlszwSqFi999Tf2W6opcd/2zwoIGxFQaUtxg/5rFIXjBqeMkRQse2zv0NZnY+UFPx6zvw9qdB3
cDHVweoRRT3JedUJEYN7HvgRIuIFJn17qh2pUCm5eEnhZAaS5BeIi5Lj/7lAJ6xxxpfX2vqkOJNz
OWuRp9mcZZOH0A7gHemIP0gA9NdI6SIwEAZzbwDns2yzI4ljAIhGkhhwm00Cjfvh1+2ewKjayqFr
EBfaPT9jphfb+jyuGtlLyDDNB2XsfUMZ4XJzQ5GtDXmEitVnrcJkeA3Tu6fijNgRvYCpeYhb/U56
CLOeFNicpygOMCV5lvzBeL5hucFXUQ2Y30q8ISHTVeG++HfjHqW0jBnTaKsAoN9kSns5MpIhwt9i
Ud6vRucglvNpJHy471AkpPoTH8uZ/UexCnjMqmhUXOz7oNarnqR+dRQTYvnQTJZfwxqvoY4vo81F
6dVW+d4LsGiKKeJHDOIFWzwN3wFyr1asIqQ4F+dq8OAkT6OD6a6LYOEElrDHinU+bFl51rUtMrzP
Ya/WkhUzJprFCmidZtUtr4zsIizjBUhERPoDQnzZLnCODe6LNU2z3LoCJ0MtHzppHCTYD8op1rOV
CsXVsOnmNisLDw42aTL4ZGq5yOuMYWUxSsLOP/5c4ghWKrjOR7jI+lxPfHbnYEHCm8RZLhfzLtGP
49NceFUbCJ3kqa/G/Novjj45rocueYgkL1yuaOcRo33ToAlhptomsjWRYnJugRbKZ1qYuIIYxnck
Ve8qFJ5wu4UIsCYOgb0XjSWd7ZpiTW0VQYxIhdgF9qyvyjAl4DyMVw/jJsDe+P0YOGC5M31XGajh
JcF3NrQVgdlyHZrj7aStj99W1Vwi87RzO8sx5eJoG/QQJ6JVIs/uqsyuI0V4zBOw7GcW/0YK0Gfz
5HPHzlonS2EXMnRVc0UuMXViPfVyFIPGegQ92jdUzEAJRtKggIKAfDfmULj0TM8ZmLddb67e8sDJ
BJfZwEvXfKCEqAghUsER38F3KowW8in6u+4V3U2D9ftccsJLtgFYgSdqJtTkLQx26kn5eXFa/sBe
PXJub2lJ7CYnK7uBX33ZZnuo3m7CID/Vom+zwd5hOjas8SBhBGjoeKoCC0o+aWpd1+xwpoF+9ZAn
fllGalWK+bOPsVw5wrJkhQ7LPZcGvxZmx8LEs3oI1ek+Nks6o3kjmRD3+J50RPqyO3rtP3tmHXkW
xg+VKJyeFVkQ3I+ryUeRs2GeVhXoBJhH2A6rtEbQbEyoM1MVw31+rSaFwIZMHePZM3D0tV3YJu8k
9rw8tccO/jlMwSGlZEo8MNcxXvHFswZQAufLijkclEVfhkjNyBDDv1YpBu9x65+ii+I14J33lNv9
ZO1TJWXfnRubN7znxMj9GTr7/RpGGHlgz33V4WtgGX0YAyF6ocV7mDO48ZrquUHGakv630AR9Xpx
cHvgPLEIIK25M+XIYhhHbkJh9h2nZrEktL01oTSH8HQMd8rPe98xLLbhmAjsN2JVGPrIKQjiVgJ8
mYnKshSFDddmtAPCztpNqEIsFVwwZ6q3mVfDIA0DavjhvJTUB+ATqX1PRh2Hq7a27Q7/LyxoGp+K
HSTk+URmG+2XG75dJBzjLPBVYy8AdGxX6JaEYgChNK8FkHjXlWAwvtz88gZs8mWAbTZLx2NWGGXK
n8Bfv8/LaDQ5gu4VV3D+IxuQ5OfQlHFf9uqNMmaTASV9guUZHVBPwrqk5SfnlAUQKvF8IzdCqkhn
vYaSwznV3dWHMKN6OzGcdHqhfCHA0wRXMID33EY5aKi5kKooZVftPjk2L+h45moFiXGDgPVOemzR
KIuBGmOMeQONZ28y205oSKEBcy5J9UI5lqAT3KOtdSXUA3O2pTALddcRcOv/Lfkb2NQT3TDEY+lv
rQjrFrvgyspLTyBa0KKpXAJhm7OqZwsbX4cWf9DptsS7fpfvI+yheXbe+ua5/PxbN2ogNBSprKcS
1AGbte0nP9FVKS2bIrvb1EYfkdkZt26GPcq2e8F2MX5RiOyxZMqr39ibD5y2hrUQKUDwM2a8DBX+
mS3vy/jXD3RMULFUdooEvBe19M750M2mKKkFKLMglwMyWcaUX66V4YN5Tr0q9e52quXfitCe1XOm
69TqQUYIqzBIkfIzLvoWy7Nxu4a9B44LQEqcCxqnBM+JjY9EUhDNvP1u0IBiWmFv58h0kY7CqM6S
Ge0vCLwZB9jQlX+lOUY3f+Q8M87uY1+eHaQi3A3wXuIVVmyDmT+UsSy+v3NIxs2GalHYrPkIV/R1
KtWoPmFw/jEoTqCaghINQgvX0kxm+hOprlv3i/IT29yM9fVIZM6WRx7mvxzju736XbIJaye+K3rS
ucyZ3bAX8ry9t7uUfim5v1zFrYGqcGerSb8QgFgDvg3Y5IpNR+OeCjLA0j/y+5sOuN9TE0iqORJV
vIBBF3bEDnE5M7evOYf0Nj6vjCC3AE7uW8oKZh0GPLJq2dZqLoQYVahHSV7KYTpnmydX06Y3YqWT
e7PQTLbbGQH87exxzf3vFcTEfdGPZqgRFrUv0QvPHH07NhDfH3XAEi78KzJ7NUU4MS9eRAtYET+0
Vj7RYSWD0s0xnE8hRuBaCPM7YbgGZLewiuUrkOjkD0I1zMhjiMPgTpHIDPiC4OzMk6zFbPKYHeX9
pJqd7gpd2oDXmVPrx1x6I+igMkQ24w7nnxfpX1Yr4rD3rANzL4q7Unc2UZUOkwClEW5cckjXOJVL
tPgS5JrAVwHXmtzrxo1tqwoULc5/xtl+Vg7sGsMkEA7BvqEbZiP09k5LxjGS8c0uZxJxUhndh54q
dKsOxDd6+k2WrGLD6tet3c0D1o/35BlYP7l/EdeajK2xgaHS5UqC0eMYsP6o/7umQHQ4eA/CB08g
//TBZO4FvU2ML+KbramKvPbJYwsUud7pofn3Pzn1Sl+QTNKLsAdw2+moCZzLv0yKyr7AqZYN54LH
luVCHkroSsbb1IuzkaH/tYP22jiMDbrwpouOKZFtB6ez1MLKZTl39CG88O3w4lVAso/I1YnKRuBm
iDVG0KQAPn6rALIHRFaiFmX3+xCkUEG5JQINAI+CcW9y3sFFfVXB7j/v2VvxjY56GQ1tILVj6znH
PIPW709ss6PjRaLiKAsp76zBL1uHp0Q8ZxmFSlSAln9xLWZ8+CCdXNay/WZlkm/DZQjv0n1MgzT8
Pme5jfCgivxG9IQIxP8kzqgkvS5ldvy6Mt76zWcUQ6S5IEMASDosDWJ9Tdk6r41i8BSdwIcds5YZ
ItZqBv7HpD8N4JI0PoABAS33DgVbK1be/tLbyHh05WDCWuONb9QmiHJk/n20LaJEDEgTSh3USPE4
Vu/cfOUrzoodOmX9HBx4DzujHqC3k11y/IjijhOU5MjXev0CKzSMmSrhNf9oQvG9kxwkxrGQUpvH
1KgHSq6v6JkactjmHC6oX3IHPZu7ERn6IuCzE6ijamuwdzSXTFtM5gJmwxr5sURTOGXrLPWQBrJ+
yATI/8NN6QO9mZ2Bvq7xqa1lhr4tfS3yHTLALazvI54pZEmXJywqYJNN1RwT1+tldpSx2flq37PT
hHeIHt3lbtC0i7T4jROBQ+mRF9sUgc/qIxwSjGHLdAMOTfhDVRXtiHoKYEseqgyRBr7RuTAKYE7W
bCLQYVGtLACAAvZ6libGoGr0PK4QYKCgLWuqx/Ln+sZgz792XEygp0INSYYeSEfSMYJIiUjv3to1
fgLg8ShoazuPrL3vQHYWgmTOqGYh/JrnhO9kyd0DNJtvGM4xb1Vq4nromfgZqazVAJsl+M+0McCP
XfydvKTNrz11sVjEoDLfaXNpTYBuGaE+ghqA0r7Zbk4HZIatug1xxyatQzdcYaCc+YIISBGIaKz/
jUuDOnhQ8B5tTZR9EUog972/r6zt1y+4Dze+xvAw4pTKtzboQwWBpoX953WI0lbbg5K1vo+GPcOM
QnQROndFiQMW3mg+G0INy0eOywEqR6KAx2akmr6QPo9z+UxncJ/qSQZ9BQRJgxqBWPwxxkMH7Gja
U/nusj0ktOYoSRX2oHP37s6Vl9Q7PTqujqQqmpDIv6SwK0S9c1+1lbRGC3oJH1K22pgp/WcnW8J+
1I00aTp2uTlYt54ds1AmhrqKLwRpsMPvZc/MFq319Ma3ppikvNooqzh7es8wlX5k4RcBUshCj+uj
/OzC/ZAC9lLwzJy5q03ESxPtc6SR9A8Apm4gwR51lxIuXCMAZA3gKMC+JpIEOc4DYQ964j+JN9T9
3MNCkKXC7b8NEoqXtab2Y1cxdB6p8L/lEsL38Fsn3XqRbRF9eTIA7N7Q4xsjGX2VmskZRlNtSp5y
X7ztsctC5PEoWhC+E9rF9gApTeZXrXovwpJCa4FFcxbYd0WK78SZTCuL2jiSTQK6mA2NU9yMYslA
HzvhKUyZbdaKeAMeNTd669/wFvadxWdL/Zz5F6bYzXv+SVziNcN4+sAimn3ATN8D3gJHq4dgH8OC
OcuG9v66PC1eon4Zbmj7tSUPYXwVBRu0mH11/UFzB527HPjbAWFPSBnVMOkijuO2cdTsokh+ur5s
H59vttikpGqg7wYSz+QJP3DmeuuN4vvbTznQbNnHk+Vfqq+BhbChEZxno5JU/pyeA7OVspdQMms5
rWL3QoP2ShVmLKeN2LxvMIXS3pqIWkSPebYCUSMw0fVrAdW0+BaT+F5AISjxxRcgnsZ33GS0n4Bw
Kj4f4iTtlwFCSKyarrNsFL8v2nNCzg86s4B/15Mo993kPekEpkv6DeJLHRr/fKPU/t8FBw7DUIY2
pY6SsrmIk9+qWGe+PWOuSBFBC4+sEN5HcwXJf6CUBcGfQKDw8QnrYIAHbzb8UJFMdwZSQE+cF8dW
Qv/7e88UDIuBkUJXIfDU+GQRRPPY0+a1T6u44ImZHYiES6Z5AejUeuZDA+C2WC4tJ4ZQGJV2GE5e
X4CQk24NSxEJm5yLO6j+04PRzdj1gkqk/3hFC+eD1PLyNZIEcybX0Qpd9CXzJh0exCpyIID5fatH
5hKkEis3qMzjVQSSAywaVVj2qo/OHlyUegajNdqaGBPzbKOPWRcNp716ZnUWrcJqjyfh8irMLrB/
O2MMIsuOQeV+qLUAMWtL3rJLZD19bDy2irVmZmUUtWcdN7MRZP94G5x2/goHTKw9O3J2Tfi0I36l
jWzHoUEJTcPtoAKrbcBWY5JDJ6Uz3G5DPo9XfJDqEBurL0buWc5DNCzVjZI8sy2TJ1jEXBsj92+N
NIEN4wcmiRS8TJLSpobHhDZPkzP3L2aqh9wIK2j/P8w3RjqRMHI+bZtdlHH0E049Jf+FyGEabbsm
Z/a8YvkNnXqq4GxKap9k4clP/HNGf3Z5U9agw1dXVmiWSp0rE6dOnbcNmn+rCgbZ3ftl/HSxLE7c
2PzX+/oJoz+hUF7Xt8NclggYVNQTMX1qSvvbCv+44Ys85iswIrBjKGygET0w4G2v/IYR85WGM4qS
Q9sgt5CK59nGy21YpWPMzT8+uAKrfCYrqUyINRcq5KN63scmKIECzbic+lMn0/lscUOp3Np92gAv
HkSUqlpOMVqWLpednXl8OVQZ3S2AIVprqUy/Rg2CSyNA9va+e5I1Etf8xONwGPru5TlV67JOvthV
TzHg3CwAD+IIkeAXpAuf/ThyOhf69Hn8uFj9RhbF/Cev9PE96IqAaneqDM0c6XpCr4wjUlhIGklP
6i7qrVFlBJSuS66jfsbBrzxuW5vLSaRr1I3Z5S8/MskkKnSdHNRQjH/3VlUopTDyWzYbaknxoldi
+Pa/K/P3d7q4GEoR/dof/j9D+1qrUWMiE8/884sscNzXnb0cQtSbdyRKe4uVZ7ofks+2CuCLA/3c
KwFLaHjPk8y0Al/HUYqWo9kbQBorXwdP2drptBfsUqjiRvOJL8S3c6i/6mF0qDyiUVmIG+Y9wq/V
MdAIXGfiuGziXRaycmBAxbFYLBF+BoNU+ZEtlsu2IvGF85bJmMrXjIflRvrxJ7KFtgYKpRpEfN40
T4r3jvo86KOKVBCDG/lhFkiD8ExX56TRcktJKY3bt7fyJbbRihJqG1rVjR4a+9QHdgaocTmnvTGv
efXo1u+qmTHCzKwKIDf4UNIyISS9oSt91WdtSWLbSWtbbOkvJNiZ9sxjE6LrGjdcjznUpNvpgbnw
1TDElN/4QuAAN2vmJ2uBT75ncpiaw2FBdYPuP5WhPVD0KekmCRQ0zSXQvUPb56+yL8pj/9BbOtjw
fj5oCAo7XxWob6XUcQcWPCIW8Yb4DEku0s6QkGxQpulyR3o+wSAiBFgOJJcki2gHe3JUNuxmLoO3
udy6+Vbh2i6nyn+k2wrDnEjVmZ00PJII0fVmKu1SPdHCA1lh4S+l2n1MPD4uB5QnLZjV3X5cgK4Y
+m0PGyBQr0zH/Da1FmAX6OFA4CqShJi+MWvrTlNI/gCBI76a7eUWeSBUNBQghi1tmV5I/XL5QuqU
J33Y6PCfVfOd/Vv5qNk40/cLlPviCHEH4EMupl6CFMg7MwG9gYyxiUvpn7g3epKggK9lpeTfMih2
y3NxPPEHzNCsw3bI1gd0CtQN+J5ULoKGWjLdkdeo91EoLzniOP7CKGZOx7QspCcIZUvKqekZArPG
XnCNMpvGyRw0sAn29NuHp6nnqZY0yND52J0110NWdH2fTNwtYN/75wGlQltVKk6/xjlOVO/5C/mP
w4QnG/SyNNYDaOvymUAlRHoKD/9OMiWUp4bI/oG0M1AJEXpf5lSjcilwKqtIJNi54+mg/qgqiYlP
jUivHxrMq+JW0kY5hpOyurseM3t6LkhCpp1MbmOSo2Zlp9RwxvfjdY60NYC94WV1o23rDtYJcKO0
n9eM0HcSfTojUCSygui1LNvC7DrqzIAtxKOJUWZa7cqear2SMufu6P8rJeHJFzdZJFKAcobd0Vcw
ahUEC5LQQURIvz3bCroZ+4eb9uOVwpY3W65M9arsXDhFVSAde629Lcnh6ge5LnSu1NMH6pfnasuY
8uQPSPU3Hht82E+kIE6oHkLlH/O3eTyWg5VeavyuAgGyZ+/9Qp0ZhtfEdCDU0aRUiKoESDkQ711R
3upM8/Xx1gwEwFHc7qOjxm8/IwOnmixtR9227Z/ZTU0LWJul51+Yx2ViNCaGzTAAASPWNsf7ub3q
MHSSq7a0OpLD3UpDQs9Fe9ewfB7e9OQZ9vH+MZ7kMpTbbIAXb1l2ZvWTrYAVcboQraYZZZgd7mhb
eafa6hnC+pJ0txcjojvXwrocB+P0Cu0vcMfTEI1b7HTH/gAE9Xs2QZ/nPDfND8ZrGIbN6RSai2fM
hj6ZX0LWkuGvSDAogVUEFdkp0QJPNoaIwFCEgZtAbDR50ts7RPgjZkhkwJ16UHF1hbVLDESygIYn
Tdqj/4XFkgtFQLly8MJ4J7JQbtf4HfwzWlTPENvXR5eqENVXb4J/74U/a4cYYfin8mkIc/rhvhmO
zJeq0DEKGgJX2bFx8jwjorKkXlj41kvxqzCEh3Swhr4BCu1fjnaDUMIl1unhoOh3zdoOUFP13n8L
/Jm6ekoKY1Yf+UwUr10Rco2hFkZhgvi3CYMqvGTABXLMdpcSQJrksElNjyP0eShkDgpAl6iPku+j
MjAXzhoHMNMKHoV5myNh2ihqWMT+VITwOp/Jwv0JXw0SV5Z9PgH9lmp8FfUHUvQbm916/R4DjuFz
jxWn7gAyknQDTAGLGoauZSgxNdrfkRLfUx7HDZHLrH0iLScfge0g7IX6ar8yJ7tI4AYKSmqSQLAL
xoQ8KbUSbYixBSNBA0x/UAhzVKeqJDrEO9VUlrWHiToNiwXpUJ31YzyAGjiVLgLrIG+CV2vMPEBH
QFojGxD/qjRcNO2UdsIXjcqsPNF17jKvlHSZZtt2yZx55XeAINzXVFm0S0fxLCFswJeOvbZIlb7Y
XgXjQaEA/qUZvE0rIV/U0F38K+ovTIvpOl3/SLNFpoqIyzYQdL8/qQGwokBEl/Tqxge44KkLn3W6
aESOLITuoKH/kjjUllOtq/kRKMNSfspaSZmQXjeLriEOa2KSWND9/h20EBvaPr2pWQ+xvW3BXPOo
XTefNH6TWZpvWcuPMQO0lKtKsUynCOxbFekr2++qYjqrzD+86mW91sYwk7uNPQ5FOko1qE0ZePXU
XCCUCr3SGY1N5el8ywhCXGsgxElNYsWLNoTsMdXTsItZ9FzS1GY3nxVb2veD4RN4qAe+/IyINIxG
uU8BXidx9qQF/SR5GPSw84y3DO5cWlg4K+pNQXeSCpzCfbPcE0Wx9POGtbGZyUfo1gV4zc8R3Kf1
rczmBOs5sWrYNwwtYi1PVkuGjprPFyIE1s+7yZWyE+5wDHU0JPu9rBgd7B65/xAh4P+uARfZJ4S+
ow+OIqceNJmf/KHfrjWx5ipKrqo2kmxLHdpy57Igu9DPzGkrfk4RuOMZt7t/gHcsHwrqZSy7sa1A
CwtUiySPvCpJB3rqLfH9RpMTywxxIRBYsYphc0xuMlB3sdUnPQkjIiuKti53GHunOGKoOaZevc/2
qgiZPSJBGZnS09qedgfp72EmDg0K5Yr0RnXycHUOJBe7GmC9W33o+DZwBPx5PPWQkjaM39xSGFbM
xjLK37yA24dnVAJbloJA4FqDItA2peDGRJ5MJWOOATXg4ZpnUEdQg8yO3aIWxl2EI9vrN7V8/L+L
H/ZJtxBkRyJCdWT1OKAFYvXSEMANuBzM7SpVQY+gUgtAVIatTqNd1ChMLdYoabdNS4RsmubG440u
XNxdMiq370LM9aokxnGSRGbj4mBFaVx55IQLRxM30tfO63Z4IEQVqWGDbd9cyM9OAwupb1hvvR/N
oUw1nqpNrT9n7HsBTNZUd7dF2qK0eiS+Mx75pacRsRfTLj1O7DUObXeDVgvLDk6ZyyPTrQ0J1RvL
0OqWbBtFZccXEY36X+L4cJB4kaGCCZqXOIKU9IVlrzaLo1iA5Wbb55w7w7iZp00BtI9W/775bJXy
afr8Gp8NqwdQj5E0GETuhAzSb1p94T8DkZuZvpGCa1vOc7RAHzFWtx+oTWIxv3xTlcvaxIZKhpQl
bXGytKKxCsyTpdRANtJmpRajBmYvTyo8GJaCH0KoouNKnn6HHRLpLY+EjHiAQnj3BDPGIDDgIZ6Z
LRXrFgiDuJvpY7E08mfb/tlbYgDbnhcLVaM3THMXNarL21FggnvQxS0rhKlwfSHg+WDKuitTegxs
WmXiYGWQSBYfnTOZ8m0OdPQyPsvQnbOJjrfTY3ghkJUdn1bSbsddhDGb7tQ3cGStgnFS7PALupWQ
pfzvUJO8w3GzsQcdrYYyitM8CDxPYwV+oVxJVc/y01nOZbqyPH/x3V6W6nDn4NxgjEPWb1A+X0kX
IpG/ErIeuvKV7L2BlNpjboSG9jMnWMZ1GHRetXauC/OSpAsBrDTOeh36wABqDZXHpUqkRk9wA/wy
VMx56McOZhkhrYF+EzFAalnKKiZAHG8yqFNQXkjL2iDc16YIUAm9VoOyQ+/ryaw3dl2id1rjEB7J
hGGL4WTUrS9NzBBmmnyuU8W/uxDNqv6JEpBb09tLy5XtwHDfMPZ4rgoacjAm3eiFymJpbKf9aYyE
FWGigb+FA/xKUjCMDyw5Gf2+SvxHhmF3LRoe4DOR9uv0K8M8jYkhqEJhcvtdXwnlbmbUvNZQZCQA
54s8XXsMmp/l0ueV+t6p9aYs/yfHQy8M9bz1BtIcvsECs6Kra9K30IQtwtHQ4WcwusmsK/mxBbqF
j0eDDgn7W+GikWlaUz8d1nrvdY1o47aSpXG5Jbp5MBgjZiTmD+EUFISHFwv6uCCLovEYv0q70fmU
PiokpuShnV1fNV2yLKnxlz0gFnr19n5d+IpimVAMDtDvdt8F1DypADr+kUbRvgPhiPx3P3p6AFuz
9PdRToocY/VfDpeLwQ74KOJ7+2gpWxoBDPLoAxQAaDpw27IxyQCtKXL+H35RCL3Rr6A/4XhtVe8c
Bg2Tzxmn61sjZY0ms3w8ziYmCBdPfCxQyQKQgxJ52ujsQG2vIa7bB5F3c/w3YYvk1TeS5DO7u4NP
Y+GvYLqvBBdQ/v6CCQAEoUiNAPDUPrs3VBIUnpVDPucDKMAF0+HjU6aI4pCfoFR9HelkJuUKGW6u
fmhsBgsrKvoweNFFYk2CTP3tAhC4BsYPQhphASYBGYTPdngmvCWgHgXVE5KsEpjuyYCKjQDlkxa5
KyeZ0BE8G4OmWzX1S0zCd4hN2oNx5FnjbQtkwtuEJegp7peMp7DcSA0UYJM4iBIaj7Q/D/jdBTgb
S3M3lgAFTT5m7EwCTHXRedCV/4uO/6bxOzJHZUIGy8x2ZM17XIol4FvUBGRNXeVwuXP5EP+bU3mv
3kQQ2+4jOXrWxO3VRFWJK0RU0iYUsWEs4H6+3jQNj90qZ3Xkc5iHizL9y1CuPaVd5wTKXP7VC8PZ
VbehNGkk1q5a9wrD8eP2nSemqrKU8WFT7WXsSRddMB81mQcVb9RCsUCYgt2aZ66WhLlUSmoREC6h
9IjBKp+fDiWA/NC8BwlOLi4aHFmc9bPGdM2ZNgBgPPf5MsgsZP8RCZXDtEHEkynzrcErZyvptdZB
HYK9QzqDy46DlHlK8SP6u+8Q82CRYYZez8PSUAWqFoHYS4rQIxIXFEVuXnBRaFOXOyI8ABv98I+W
Kou1c+hCYukZLKXVdimW4MBEQwyI434XHi0JNQFBmQJepiqMQk6ZqTqN64i9K6ksTHscLQcVGovx
OEXyQtjIadoVYmEfmmP6n6cW6GLm5a0tEslvzIpQ8KECW9aq2T9/5pk4cr8pgo0aqS8xjAXc7oXv
tij1ZgeUEyqKu3ydZy2/LNpQ3MFTBQfZSJrCpsOwzrV7p1IsXrtBZPAxxdEJ2PvRYKb+Um+bdKbB
tpmzNr2TMrz5T7wreUhN+CkoH5H1FbxLi4pOtPJ3CgfD977yypbKkz0A3ThiGJcUCePAfZgo375R
fG8TWDdZI6hy/2CVyX3SSKwYRIjobT09Pbb8LD8bisc4c/aV9iMV2ndidGXwPvMPDgsqyHqdGihN
UHIJQRm9KN4VCpf1R1eDNb2Bi/CDXx7p8KmEKNo4JaKDzK9t9Xh9P8TWO0egoiTFmF1EOCZ1Z+T+
DZcXNyOnDYl7+H9vqRG20KFnHcCz950gxGGKHRWfMFRfaTf/Z1jGZXlfdPFQW+Nq5ohmXiPvPMhM
wPcKXq+2x35Og1z/IaIpctZ7fybnJq4qG53HurmqL8ujydFFUDLZ2BAM8hglEpeUmFEzRcBj9IwH
ADhyK1IgWMQRyuhSxFRaHaJSUL3Q9TFlCbT+SiKr3Q4uGjaCabOdjYV+aqn6ID5iDNvJYRVVbNuf
R6npu57sbkbMPqDFWbECsoVSgBOhe6Q1VZ3zbaVmo1R/vuee+67WaDhtAa2o9eBkN68ps5suDPZ4
h+m0Pfp1Ve9nCS5Sc4kfASzeIHhIkcZOrI8+7Xq+ipNXAgD2seB4ZD53VPamwmM82WnXWkLP5uGN
kUauxFyN5cIlb0c/AgbY1smB/1K5i2ODtXaagn+oriKzme7OmyP9j/ljwzft+bNO7cwQ8jRHWv5E
bztB1FEtbcSEAMK5akJITFLnC9XT4qy1yLoyKaWIX4S+4MocgxtX2L+F3GaCh/yjYZQP8Ko0gNzd
8moxDq+LUZi2h0TGsOy5s9PxGN+vRYOiXeya4ymWlNJYaL+9XxG+PZHmGmp9o1t+OTAUHhPSY40N
ruPUYgxTVsSFBAVa13a2qyqicNn1ngQn2LUD9BhvTCcO8yypg7hvJWsrFjrs+x1Asxn4fms5ylDS
W5QH/UYAzSRcbcjkbHGWKRcO6oN+cAi6heM+Dbp1yr71G7Bd591alMUZGsTws4FYiRwC1Iw8iGns
iSidbMEAvyEBlaiQ2p8xEBHzJ+Ez1ph//BpcLP/cuG/7Qsw4h1RKCSWawWnKFYSRUKql/dD8pqwn
MEbETax55pnaVR7jyObFoYH4FClTGkNbAfXJOAy5vaaNoGxSN+x09Yptx66gTdBMwbk9W3gKs44y
apT2miDvt/Hrh7W+ODXRAKVF8ZMXeRF6ojtwSp6VFleCCkGbnGMWX1t2Dlfj9umeiRuNW3A2Aiac
6Bae7clbpBSNfa9UjP/NLe8Vo0js7ykX9To/5QRE0z7zZuEc25eJJA3uf/1pt3dgsgBAy7luSYeZ
shJ/40I3QkO+q0rnjFiyjSLqTxv0X+XEfCVtfiknvljq97NLgpdg2D8RwnfLOPDHkHwbupOWcmuc
eAfBlWdgUGgpcv5ZF6iYVfNiQMP3oCGFnXzfJb7OIgLB2NBYCflzjiC/wfea0ww9HV0IzGd91R5g
YuWWtx8wL81kd946QMjJocdXA29ntzgwRlIoRSdrgfnPJK2nrsR0lC/4IJLioMvkITAY8tuwaaKf
aWxxZDFyliZ49uXlH6rT1G2RZR6iuP1B0RkeyJfJCKLMsdh9EpX2be9hVKP+VcLxLpggYk6DLFWQ
bzWAhQybSqGmM0Br01LdG5ndH8uuGGIdmWHNrstJ6d2UoVOO4lklGZCepuM+zD9XVBRzh5MCxQYg
Kr7myD/X+kLx2rrUunDc5ECFLKfXDBnZo3DfzO+U0wgAEI9FyWQ7joR091GgKpfxmRqPDq5M/aSM
N9P9qKv0/bZHGtAx6tfihdG1h8eUmJHiMpBlTlTZlwQ34hLtGVpJSaCdb97bNS/r3eTW3++rYbsR
sRowut5sr+OH8DqrXumXHgCQvzMMNLU8Gij83c2V16ghg0xG3SsS3jW7lCD4w1nyXcvPrKBTY7Te
PMLUekLFIbsL6MLGUUnxSqRl2bXi5C71tHiXkDIXdko2gy7nzAbqbl6anOtfxfDOq01jXjyEEjtK
tgLLzVdGD6y16cqNFTUZ/PQ2wpxhVovUdSdNMFlbOlM+hTLZHPC2Aj4wuAsZlkfLF0KDr5z1Hz6J
CQHfQyoha2IwZ8zGbl+EHLLtO2XQDGPRAvLsHjyTLFawWL2jyRDJNy1kHuH3kqIxBuRkP0avHCF4
PyrdNVcRzp3IVyMiFiOGTDyB0mqBKR/GTn9mRCtod7eZOSzjUFlaXnaGC3+Xi5fjYBHzs4/np0nM
azgjdjo5uhRuQc0HVYYK8R4G7KWbD55eWX9h+ZjspT1Af5cMYEVoy4lcbz4SzxHGvfVRnEQbMKsW
rTkz1RExabBKqJF/fOg1cp0yNmoem+uxLVGSNXVCrlRYO1jVAaezwJCF3TMOavVLz07KNPAqI8Ct
mucMCHxITMuLllPBFERrZQd6dYtkWGJyeeBvBr5x3zpjKlBNCo6C8c5xVWBnp4wiVZKiq7ux1Vij
vXbTZbzSNs5hCmfywJwd6TQpfcIvffCdj+r1kSzpDv2QVcgVhCvbFvwvH4gymrVEtGZDX4a18umI
MhCVj/xAtCEQHsaszZbcrOfDvWNKl7V/LnNIKEqOs00K7K5LCrhYvx1u2PbjOXZTcT/8Q60S71ze
5Qz8CRvyjUXwxhrD4Hb7YN9J9hWhUymifvPlah1CdlK24m02EML7S3lBgaegr1MiC4zgPTms/xAN
t9cJiGzSV20I06jKXrCrsoX/v7UhI4hHnVHCeS7I5/2AtzqRQBX75VUvc8oJ1ykU3WJst4vAh0NY
bc7U67FenHsit4/fD+793jbn073LOKA3cvg0/q0h9AEOZdeP49u/ZosUdep/4ZuBkmxmWutAjzM8
8SAeP06p6Y9ZqS/oRRKDrRuuDYW/ynzsn3Cs6fPlWbdyOUkPU12tDBGCUxgI20ZwpfIexhzDgol9
Ztk7a3tRX25Ulhrv9kdv3RRISCr1pIHU9wAKQ7wdR3Tm3PNRsj17c1pw6dVPDE3Wv3tPkG8la7Ao
ZfeoETndr3qkRTXooSuoTx2SgPjTW5g79FqYxdif/q8IhMvrDeKiTP1gq1uYuVA2iKNKbuXA1L6n
xnW/iWIAUzds19ODDkZy0y0CQaGk13d9SGo4+RUAY3MOgR9KrWc8ngadgYSOjnQaXsU6/alGBSDQ
9OjeIexB+xATbSfp8uiSl85SODYXS1V/qgzG+3//ZId9T/HEwbdtUrGPZCVuPNchjP9IC7midDDN
AvTLXk4Z7mAD6PEuUh8SYfMuHfe8S3ShQpp9sWcvHCppl2XTGmd1rp+TAnxAGMmblnvCrsO9OZaU
eoNgh1NUnaHeKBSb6vn682OSjGSSwcSW/4WgHf0xPueHYWq8sNhZR81wGMvJz0eRpVg9RrV9Xx9L
iVeXPBgq9yGKLSj3w6X+FOwl4cyfL69oSIdpWp6Zv1JX0pojk+bqijBeTBX29iv0KoF91Z8P93WO
QkQXBMcEW4ij5Iy3kiVs7+yubcQDphIW0duXaxx1WCjT5EVAQQrGBguZ7kaKdd3MC/BOacoyHtR3
1fba/H9I3TAZrIX1vnQDFGgrLAGxL2nX/b1pf76ne/sgM3p4PtHySotAIdeg7pbwP3mCOTIBExWQ
6bW2EFCbRCY5kyP0Tc+3RSS9MMUwHFsjxzGlYMfbEYm56WJMhds9+q7Zp794fk1mNz0tdUwEazYE
D7wWyDj1mLp1U8LhqfoAe5vBJf838mfX+mIOg+5vg44OTx4tBdQfcXosY5aTepAlPrGyxYBpiSI3
qucvnFuBBJlBCt/Au3zyeEBm1sp07Uc5sliFt6DddQHF1Z643yaySMpieRzAfYW2YkNycQadyqgv
HqdZiTIeb9KBDIUwCfQjBgVj9mhTkHy603rUmpb4NHB9HwSc4GgdJL1lCTS/ydZQg7Ah2btrcjOf
qTmGG6XOKGTu7siVQhixRNZC+1oTWcl9e1ozqyinUliVTFb5kcPSZpbFLA/c3C5STXQS1Ks2/7hQ
kNVWOjYX2q+V+W9+LpM/SGkCH+X9fFsOCCZcBq/X1pt/az9olLebMS9meoMWR4xqMjESamxOqEfW
lskb3s/WG5jG+t8DnWQejanWVhWLQXAYAOV01cRAA/7tDRchwWrCZ1sNZsoQtqqeNf4Cj7fYrFVG
RiO15uXfJQrSWIO/hnA/5EUhHj6Mle1D+4knM7sMf7+ZE6eeelFuBFrjxF5h3nUN2Wf5XKEOq/2C
QWIcCenyFKAi91nw8qPeSAU9WbewEy2qtN6Ic0/FGP3lLncqYrETo3g8s7YABcwnRlhcxtfwM1s4
elmheJHpYLiV/T2BG+oHF2/GIjrxDTkLeGpOrVaj+TlXtSt/qBViCkRYh8lGBmmtQGIojZXFVfZk
H/85RhIiBzSz2D89rXfmfhENgnzwSHYFskvcJRhQqtRKpsXP2Y5Zsx08KXMEmXEFKyIWGcDnsUWc
6jrkN1WcUArqYDTta4NGpwkWHZzfNwcrYUe1sRShAhKjvpLbo9uVus4k8czmuLpVZMd+FhrgN6HD
UlhVGrovlpVkMT9jB2cjrgzbTMIcT1EViI0KJ6yW3uSfuUY3Ry2fS1w88ndExDdDRS9gWk7i4FTP
tpuMWf+CaVo0PHM5IkJPvoT4xSZsdrjTcisyty3yMMjwRlJRYUwJwuDN8OTG4AGzgcPcv/8q2DWM
xK7Y3m93Qv5oHlTfYqjxqIoU4olk5LibNj9m5LnpsVIbsUgaN7ZS7LDlKsenZK+N4+Z0A6VWYSVU
H9YCU1iIJF509ujRXEdQYGrQskMcOB1AYNFmOmo7jaW+3I79qpYfV1edaSbVZ2ANWWWdn1QI9GOA
Hos5haRKsgRvV+zRTV4whwkFgoXVFpbxhZUbEWuMuB+I4m82AbML/0z6Pn5REFplPJTzGlJj4bYt
vm6tFES/0lwN+31wdL8+ZrxtMXAohM9kGwGSkQzrXDxDVPX4ia9lMva8eEpLMGlok6GLvfZireLD
kDjHyh6gNw75zLyUWsescD54BWwFSrumkZevQ3pE/bcMaNt2XAltUFGU5dF1fBt7D+ni7vUlKDhD
2v2qhX5b4OPHH04gT6sqUFNVxrFE/nw7EJGUojhWy3L6beldPnIzK4xyKYRAVp7XtDSc9AMvAhOv
TMxYMxTrEgMZQyHmkrDX9GK8AZUIe8rU6O8l4/WF3ecwUe8hxkZeZtZiFBQRExLWk6z2/PMByYpP
kB7g1rcqGysELUZ3Tdv9g8tG1Mz356apuSUj0XWYHjwdGeYn2kV/gdlFBzR960UO4Nj+584lfslG
pIDATe2tCVKkhF95XEoAoFGFzqB8kkDT64Zi7juXrGmXcaZ8rYPa78a0HBpqlMTngW6oXJxk5fYU
gr5or5VReDP54+cU1KDWW1baxmbQ4720qD1Jsc2f6vznquX3KXW8s0UJTUg68eYLa3VWWv6tKiXj
w4N98vtPWZ9l8itsUHsG3Sn4pvkIiv/BXsCwfY12A6ENO7wPaotPk+XELG0k39O7OkU7kycWlRcZ
VZJACjiGQy8OybdvuiMKRLEWq9rPmxV/UQSxxKkrDFQ2Hh1OrrgiVFRH2VCTmDGvmO0B49lHXETo
mPRY8U/KECNCWWV5huokE9VYEluEJHGkLgCPGj1Pu6Eh67ItRfF5BJSN16R8yzmsAawoaR52Rvwe
40KxJ7Bjcx2dzr+n8PTtZ17vBA753XOUiygGZq126RBPlPZ3YT5Z/2Hz7Ejx6ucr8RiKJQrbq2CO
vZdWu44uzyd2wwz/fz3HYm/X38fbCz2f2+skZZdNa7HYdHmcvylb66o02vL2v4sU7iAV7GTQKXd3
0/ouF6QTxnrjJanqkPtDKQwB2tjIH7Bn33WIWOXTqsx/l6I5l2a25ZHPWYYiuNelJ6sL+bVgJDvC
PWhuphYOPQwTS0lb322HmM9rcz8gvuJZOr+rsrAD7zi+S0fKg5IFpPqN488WK35Y/hArBkqvwtLY
rO0dd0ilevUEyhSPUwlR3miRw5nopVXayt70MSGDpK5Y+nlV1jZEvxe6yoMY+i9YGQuNOwblO0e3
E2HQlyFtlHoscmGdB80+ekMx9xlfwVyRyrwE6kcL0oKnkhy/v5f/n6w3gcMcWjwopJ8lH5J9HyMs
ZfuBShwZHO+kYq6wmBmwQ59qB5pzmhbLpTg1BCn7Nyga8heH1sud1bpZd6bwQN+eS5yn5PyxXnDm
CJWRtsYVfSrC94RHDPoIoH2eisPssX9AQKrbjSba4v57MRUGLsrqpJAqQaGktVQ+4UeaFTvxFn2Q
IMJ28TmSEq/bUCzygx8dt15UtHI4F/fH0y66Lh3IN6xw8gfpoE5VQu05TevFhdNW8p9eazkVNIEu
Rlc9RFioOQ4OfpKUCNh884q7lMVkIaGya5HRcbdcY5iB0e0D0PqYgF9ZFCtye8csU/KCcU6ykm0H
akMWOXwrwkUS8TM6zuRM5jsvbKbm8UL2CcruAe0CJtO6nKcuoXRq/f5WFgWLDQYrVrBYRd1c1+FL
5znPiQPb5gRnF8oRn8iCzOP0KisO4G3m+n1HoLDQ0ujted0xWxhhH5afcCrag59B5HWe7Mu4KKim
24wPnjv1hRh8zcMVyauEqbhNuQ10BGIaFupSRa+bMCGJmQ9sBfRo2t/tPPpQrfvxko/hiJC/dPpp
zYUactzoAF8RviQLMnTSu7BvZSG/7UiThnU/UwDqC94TdnbBHVlVPfihLy8gxKHUFoE6TknhwzBB
zApDk2JiCrmEJgzT7ozvq9Mcq+8RhnxcY0ZvQYik5Kf4Yet2t02hx5XvTP7DCNw1+f2wZYSr2gL4
hV5XCB3F20zU3pQFBx3kAaK+AC6hxXmwuIZjNFDaUdGYb3sMPtut3WPjm5yKe1syoJPTFmttVQaB
2xdl6x8rfkLbQzja4Vpbyyg97EC/Llw+zkeBy/dgE0YA47uJiRVWBfBol5gDiVlzBZmNrzlMxK7x
wn6F1hsUJS9hPPyaCQhBu7PY0vyN7pXnzgBoe9QIZ53xMh9bwrps9uJlYQu94hREhn9Ch84pNPZB
tCgX7deXm+sPdOzPP1wLs2Wl8qrUNvs+VBxmB+hTnOzNhQZ/Km0wzQhLVJZGoEW+mG1IyiNoEYHs
bp3/RqGu6maft3gEntbkNGTyi0/BFyqhIGFnemQwU6KhtvYSOWVRhXk+5Pm+f7sw8G7BrXIqgeAS
uK8Z1GP/DxYcK0XPAvgyaRt/OIRzebNt1u5dK+oZdlG/coqg+5j8SMCWZJdGd7BRSPYqDaHoVYf1
lI/vFpCV36WsrC6K+ckzQ+g6iAZnK4mgMzYjjof4k8r+A2siYx60vc+CciSZjusEH+XJjjd7Tomm
zyfPBThSjlO76AlyPqWnFxg/rcpxXGtxlFKmpR4I9FdldgPfRrPiEteaRPeDTohY9xVNBK7xWxNX
W+he9vzJWh1lst/1zAIXwxiVjNnlAfJHPPfrH3fiNXIf2JqAMZSo1lolqVzj5XATT6Wji47zvT4U
l/LIoKIPDe5T3n7MX/+lvSLUyDnEjXhBJ9uNRJ/iKxet/Ib2/4izmWYOGc8Sf3WHI/LIGhS2PSbz
v1XULVDZfT6s6vsdOOb/P6PEGALHjxS/Yjp8HaZW9X82mHMCdsSa9EGd8WMRvL7Yd9kzTmJ4SJP7
iKTBa86NbqgzeUBo15y7rghYyfF21DLI6GR2XH8G3ulY0JIy58kGMKPIZODpeRRL2RAa1k9mUmfK
SbCI9/8JvIZDaVqVPwtvmaSctuPy11X1U5AhH7vLUad8IzGUOoVwOCYyUEzcQKlIKUGKSGuld4kK
fKTeoH3gMQgAiQuGeGAirI7xX1lz+v9nzwsmYycG5PVMhx55U12yr7xqQBJyMUg9yM6LviEdD5SH
hCJm4+BECwhiFu7wsR6tp/j71Fj+OzlH6bXTUnq8KcHuNGsbyKqBe8JtsIHG9Vq4eeYSevYOd/3g
2hIOGOv4ndxhe3xbZ5fmnecE3rYoaCOhRu4cPUEbflvBaFIbSCb7IZ+WELIzmyIoVNj58HiG1W7V
azefnz/J94P/tNz2wx4ss8GugbCdyvZioMNl/hV7rV8MpQ8qH197Mcwda9WW63tIB+TcCoV6Qq84
54GYYOdzSd9xorjJnZ2R40h4ICU+x6xnp5gm48wBx4b32eJm2geC/KK+PNvYsAgVpu7dKQYtRD/2
nMQgGqVsHc0jXvLkdn67cD8Pta6LPhufMe6O07k2Q9HbNyZw59XIE88A/SBONFKKqMkZYPYi1xE9
tpFQEYDblRfMBX3e4Ew+ZCGk/Wh/xufof7i+yJc4GzgbLQhF1IUBK2v9zX+w/6YeJxLBYJ1sC1zI
NwO/2aF23fQfv0eWQRVFUVESbfk6VLhkvw5D04X5K9kM49MScvvOMM2sGL8m3/tBawOM0Di+guFV
kSt7a9KMuUreRJE0HLEyBzOzrHbpJq5UKbbnhbpgmv929MgA5XjVvnhAeurIMex/GbCdE4V1G5zS
AAaKaCAO8bAtxiKwS/no5GlleTrbdix3FLPw7rW3dmdE3Y7f1oUd+JIuiMtggjGnq3mvXNOX2HOg
mfLuOsQ4SLCLmQSkN9EpoigmVZy/ExqxrhhqLSmC3aZPETw0sbR/NaRL7xBFCx18phiTHnbJCSYY
wznnhZp+sNEMJWnW9lRlmG1V5Qd0tmzEvFKqkJLPMDBGjH6DtN5lWnxTqrZKZEnTHyTdwzciit+X
qkO58PEzyyFS8MRWWyiX8hOyl4649sDgdzM0DVjbllB47uOyPAwJhrN/zY64RqtG099m5vBV1Ipf
j5P1JdoOBGr/OvGJPcaYFotatqOvESqE0R/3U3uGGKDgEV8X2D1xgGHmSZkciKzJ0xgOk93c8QWg
GI0JHMZzEVrMsVT6KwrPGOLdhkH4NXsv3Su2y2Clq8vFY/34TbruGGKJg91QbZxBuy8nr8gyhCwH
qAZNyx2DmERBpFZgHE88vjC6Bv+gfjfJr7DQAd3Yu6CL15SdTpXbx/m0Bjj+BU3vkcguvh2hWUg9
xRNTzbx+5nI9DQg+qdo7tlAAmrhH7h0w4GTW2Q/aEgJRcCktuzWf2i7VHkSC/Hon1k4d0MZnT5sw
KKpGuR/hGEkM0OJrFCPPdWdcFNCrRiRfvGEiu141HT2m/lIsk7x6yE8A8Hj6JcCWy/OmdhSlUdc4
79ANyFAY6MwSuVTMSf4PlEQCAvW0026JQKbdw/O605DBmyxljsnbISVdqc9eRn1mu0Nv6C0nv12i
eOO5t7y6yml6B1QuyiGjUInVitDKffDpiOzqBgkJTN8bTLZzTc5A8xV+mEkHr/v7C74cpHmTX5cB
bj93H1kKcG0tS8boqETiHeW7fV46fb7ufNV+LZTA6p1X0wRsJVmbfZagwgIiPb3aHVX0Hil076Q3
PyPk7yZSva2qkdM4GjoS3ZIOjnKpnGFzpfw0NeYIUdF2uS/N6z2yb6M3u/ozy1e39FzF1/zN84+n
Zf9abt4feimh3VeEElgrB9UyGE9wouY1f9eKtD2LO7hyk6L9IiHw3ApaMBisrBkF8NNIxnLFt5mU
zmxlfphv2w8zeHoBZmzXAGA8OZn1ZeHWy4wzgWB6Vr3pu0ctOuKkxGbyADKWUYDaUxFh2nByGhCg
uZOt5U2orn/7U7nSx5nBvGuQuqAXZEEWsQvLy8Th90S3yiYj05R6yBNz9jR+Ejz/7OmxBOg2puKC
HrzdrvyxXVBS9ChN1qhpmnniCnPCXnNxL/SqwjKUtVCd8HNznub4jNUjAKP4bShAtiloCFkeBsIW
nWs43TV1ZK1UBCkuqJjLO7mbIS6CZj7BrXgeGePa5/pgvbr87H/r+DWvD8zH5NVvflHLBcWTphSM
O8OtyOxLCrSjD6MVTZUN4BK5sKPpMgC9seX1x8yNOPR91nJIAfsXn/J5NYR8/FMzq3SI65p9FVK5
N7ZA3UMf2HrxagRt/GuOZISHT6r+Jx7WI4v7S18Zt1xezcJkV2SfNOoNWFxMvo+m4GicsZ1K0kfX
bo1xVos/ReuTs+Hnvobyecd0Pxs4YuJKobebBXfY5TMSfar4IKa1lAA9tNgV78/zMq8VHWYOyd0k
HF5sB0+n0CRxe/O4J5isyEbDp6W/limtoXVnvmvSKlrkV2nEImAcHXvo+p5xZGN3U9QUBrdPXyWX
cibNaM9ZlNyg07p/uGXUsRB3Zi3sWaW2Ubr5nkfED52efuqqXmtg2/ZI76ISkeTMag51iJww9+DR
ob/5t2pAyLVj6uFSCzjieGjfxG2I9zMCWvypap0AWWB3a6BMLfCWUUZOBWi0u+mEX2aRbNA+twFR
cg2SVdvi/dYnQiRKUJDq8Uvo6i8A5xErLSO20gEeP5boHpV0Y81zFKfEGgbkTf8+9TPsDbl6b8ta
m/O97zRlCNHNAtrIMIa4PP6W/pNUq28S24qQXVzgOm4hXpBF8QRhHqIBzEeZod1IRCtAdGuT+c7T
4XSEsjlB78VhYOvHelBLADYL7he345OQYyT8SBsTjOFPOEeoZp/rjQVVwedHmP0y0vEwBC79+ZYK
NqkjjpoI/5/LsTVaCGwvcvbKNGuNSonFwVhZheK2KLsYD2NCy2gT+QoeZjUYNFO3odUTqjdbZmUE
WR+R5ejYjKh07sDeBGFVoa3VJk6q8CdBDND4v93mkL9NkWe1oZ9PblarxFr9j5x5hb04+dkQwPO4
xNkb7tT+nhcbIoLx0EMriqSl/iSpU3MOZ0mDjTRFHHMykAQWuVszJYOJ1kMyX3lb8WY3+i3HGCi7
r1KkSXuaRfQcRmSRmbc9xMjfngnk9kUWJg8Ti0ggXxyvZIWLyh0rQm8HW+XbukaXHOE/HHJ0YjlW
Ul5JAS4FamGU6SLysxGKcIRxMT4ACcp486FCy4ZOphBCmokxf2gi8NZdZp2z9Yb878PkhTNHgRLu
Mm5hZ8vXU/MJkRcloVzYoCZMxowxn9blB6WAu7LpXFg2XnIh7Kl2ziyPN28tCIpb0ufEPnBY91Ko
muJB+PLhCu7cQV6zvxRUT1wQU6SLtueTgumabuQLiFEHarhquYh4s5n+vst9SevhA2PDjehOG2fF
UD7Pa1QE6BRKKamsgr5VIn6Z/6yVfVpbQJEOfLCDST1Nae9APpDD2X5zFi6yLr8lGzYQtgKq6hD3
udDG2zCRprw6i9s51xT6lRrWZ2eMcmITJQPFzg//H5k2/Xp2aB4BbBLg7pqndC4ieVTfWyL4oDdX
2brhjOcA5m+oCyQYeQtzzRp1ucnoajg854isgfATQbFCVNRyb3u10RBNcAOdvZHwy72zFBFbccc3
dfY9UK5OaiFY9YqukKZkfnYaDCS71/nV64YnGX7A7v4YrUpVIpSEFy6Jl8dnFbHBuzr7asjDUAZz
RQK9n6bCaQDGdayvc78C9VfLG9avuIdMtwGHloTaHqNGxa+Y6jXumnEMzEKbmIGnhY/krXQ8UPPy
8thBI/XUcQpaev752Tjqp/01pBAhjhsgkvcoW4sRq96hfLbeA6Meg7tC7NPFtRiFH7omQEFatSGV
dzJozeaxdsRhRqawub9ysAT9xVbNMtlWSQIG9lSIWslO6jmbc7G5jx/tBip6O2AcRH7zgeaO5t64
qlovXFUW6D5NYT2lEZZPYMiMUBxR18jSUG5vnGlaSUXNA+aIaxAWXWiXOZxLfuS9JtlY0x+lsU55
dNbsoevQlXm7yl5q6r5CJIJH2/dkcenuuQ9mfwTC3tT9nSNtjqiV8VWr0wDYWXr/MyEgvqvo6L0y
cOjobzvvbWYAoHNyKXvCMtHqSs+BK3cyQ9Cn4L05/ANxWJCDzQl1qXdlwEmeMWZNFpSVYnm/0KVM
3kQHSAnKKDgK+mHiR1641OPvwcDtsp9wLFf/tHPOZG0IwQMmtiRRL9k1gQ78CNBq9X1YMP9hvyDh
7OtmIz5gcV+tKqTr2zGYxbYzofhldaQx9NOQ6qkkTA8HvRO7bIqybNUysTN5vKDTl1vtAY7Yyy9+
CKQVMXXUmFOQvP/VrYgVKBd3nEsbyr7zobjxq3SySiZJ81MSVHSs4YkK8E/jPSqXwae06ahNDo7c
t5SJZpSgLiGScEKu6NmGmUHm7VRSCByhrfHlrM3xWxn4b4Ibv9fUIlT5soZvsGabl7lwJdd6mu51
YTS/jRDkD99m+O9KSAG14Hmmwl73iHOS+iecvZjcGsL2+xsC94urc6l/70gt0+AEtvOLLHBl08K2
ILtJMM/OxmmEPz3Ktn8v+4dEbaZg94uMXZLfS6q576zUAuSNtn75glZxqO/8mH7l89ZH6WFMoE4J
t1EVe2ZwmaOkFzpdb0+8Qyx8eHPxIFmI5JS+nSy/lvS50UVUdryDu5StaMKyiSdE9oy0+3hYxGzD
ezOATVu47gyvgnsr3/dgM/8ppFtTUhQi0ek+WGlxyfDn/VnBmZwDLo7JbBfxjQlSMBn4+nQvrpu6
hdySWu5BnuBKdKizQJqCymlaT1UhZWrc7ZW9eWkSFTNB0eqX0ZYNc38x/iJ1lR6p2swJOUmfH05F
P/l43j8PBMARkdl/oRLFkz9j1hAGLH4mWGJb+iaURWok8pHh4v/PxcqDy88lXqwJkVw3Vl2fSCw9
jI8MDIojO2h7CfDiuJZmBhnYARS+3OIheXpRNAGtwQqzGpOBEtWxNuYJBeboRB9P5tJ+i59Y0how
XPvxzVPbFaD+bK0iMHK1J8dRmeDUVgnlBVzKFU6AAP4pExYqbdo1KpXyg8M5ySbJzyLqIrBMnJBf
Jy1l6Z/PNEFazVzKN6xzOrZpCrLPWjZi/UYyYFkQkQqB3d3ul82arYdHUt2J8VNm2t+/15Yd9JmG
3EzSziWG7MsjeJL4lyYA8beGpPamXgffxurLESGb8vg+boJ6D5cZcYQeP2JaEy1ZhE2vhv5b7huZ
ojSSB6dKHsnFGjs2wjennQmLbpTTSfkMJooOuZavoxWRUxOYa6Zp829/bPZbjXTLgDv97GUV5AoO
0q8NMIf8CLYT3SXbmULccwzXr7r/tiMbcW7NT5ovPwvFhIv8ac0a7XkBwqZb3Kv+U5oeMyGeT9bH
7Sz1pBlv8EQ6h/BiypeVcM4H/8z1KvTC5KAGiKgR+y441jrF2N78CuGkMMunqNgQd7cfc7Jqp2Gv
AsrF4+Qg2dzAP0oips+2aBu9LOCnonbEi3ZrekkvXlqZjt0/1izZLkRMfFFW8o8pX2WK/XTknbjl
wgdOUQfjoWgrxXJXMZzjcx7B4imcGtfgvJiMGf0GEZLuYPI2yH/sy8FoyABgKpxv6zidRWqnSJ+L
nFbVrh4ROA6eu00VLHi2WMPgOzjiGw0bXF9+e21xIfp6HYGL+xb452ryAineZ07EN8MqA67fJzhK
aIS0NjgPMvfACXUuRfCGQg6PXOVipO/+nqpgzo/k9Cp0FN0dDV4xtjx2ozUpBzo9Sf+RQsQljE3S
ltQv9WfnPo+H7fcG0M7Z78jgEOfkPKeCs7z3GdkS9H6JfHhGc2vjGymRPM0nG73QmajvfYoVbyP1
MIkOBD4YWS0IvISvms6Zztb9C13+lId40mTUFtixe3v+RVxhhpuAsdfJWs5m3zIVwiZmAS2P6r8P
Orff+jnRJ2lKbKWsODRKKShXqAWxI10YY0AcxJbwm8s3SCSuftjRU6ls797bJDEzOV8yN1nBa3na
Y4fGhdpi2vXmd7z/YUkgbtGgBlUujkLuZr8bc+UTsppHs7GDaVYS6fWnRhZemTcULuru9Y0tmb5m
gMy4AvJv9QiTCtpinjXWZrqAf88GPCOq9CjpCoDJAqHBS/MT9yqn8a5THgg6sTAvxnPb0WMwbUh1
PSe0A9dymMgOqyxNd+FP3z4PUk/55PXaUfkDdQQTJbDwO+Jay2Cbgu4CguTlK8KVi466Sat6ehk5
Kab7aHzuRlUGvw9S27n0EE61/wJJzRXX4KFt8ARf5uCSBvsmZGKXQHZD59jqeE6tUA9hoCiDUXeT
Lv9ZM+e+g2YXsAcx/+GsWNOy8ahuVd/1y/4iYx9TMuJlSnktB3A80wwQOzrY7Ym01hIFwXjPmoVK
sndDQIZby2ALn/kVGeVCHKIBZL0lIBo2Qpw2A4mz7glGfuVbshpnDi/wTDg9aY9W6XPXcIfDFQ2C
ubRRUwdj5/myNwapYVr6yuP/xdTfXXhRjspaSNzOlgqb5+3W0ekkKeJcAZXbLnDll97tdtOQT5oU
c547LsVDZCcGC1DA/Ke5NlqqKmsghFz44uNK2ejLp6g0vSv2Db+agj8K95rtygtiHy1msxqUWx+K
U8ozA7T4kEVCofayPjxIIlZgfJRabwfX5b19cMxmmzMOgFlh6pM8KSlyWKOp4h4/MtrEOmoSVv+X
FunbgnK3nwyTefYl3x7p0vz/dnoMxe2pMfLIvUwFBSgNJccT0B+yx/uvSyqoUcNUuwQS0zrVt6Q8
uKoVd1oF9hT6GJwpY/JfjcrfK3iGHabLATpsFQuZ93sejONPOzwR9+wbpxghv7lQa0tvIQqM7Hx3
rEKjg9VvlJbzaH4Mub+CUJEpVoXCozotW02v/Ue2orbsdPM91R/BRrBdYwn3vjS9AV1J0kRuAy5J
P38Qj8Oktg3w90ebePW37KKK4afiR8hZZJt4IJAdQw1i0kG7aRJg8bR5Hk/XHna0rI5qguKLiFR9
uEkGQWyEd6KpwYdgO7+gwjaflc4FdWFENAMxg1Z8JOEUYAaeknEC89imBNcMpTvBx3uxPU4xuiCP
+2eD24OvjvrkMnpMPvqkGQE2MAmYyIOcgbwwCY7wNh05rJociIQwZEZxoFa9DS2EDcn84hhuIUZk
H2OTLIPxXGuI/16N8cBfX7jZj8hAZtI1SZtWGw9R8jKPD97ipbJP3OAUx94w4hej562jnRrxa0j9
8YOmEN10TrjanmW23fHa21lV+GtSSewDr00wP37D0isQOxxzLht+/kGW1UWmZm08nVmov7HP69ZC
LA2qQghoBi93rMHaJkv+xF5IWE2VDasRXYq33g0PdBhIILEKKo+tlx6GDu6enMUfzF7EwNsVcv6u
R0WmbeYgnJW3elOfqjk360HONoYQm+mHEHAlRjY4nZWaeJiVAxBoq1HRmEON/tQzz9YaqYurXGFT
Yn/OIKAaUkUgN4QNW7kOwGcWTuN4nb3fq98b+sN/CZHZiqjkalfVP5H7fnxckyLIjmOwRVlIkNc1
ZYn3obR1uhE1pksAj/oMtDMNCyF85/CAjScJrpJZPy0wLr9gkQnKF1wWrvOFb3TVfewm/8KRkptq
d5d2D6n8VTur7SuvKhbVxrvl00NJ23396g7/U3qVMU2PRUma89wZDKKH9BcmbVi8ZwyhR+LZJsA+
0qwt44f1n/Gm764K9AKuSI4EMcGJKU9l846wQZvJj0l8YyxqHLUEpPH3VZpFlFkIUglpBhW2pGpv
GUdYMS/3LEPkvgHNvB/8ah2kMcdgUJBunIS5+hkJcL9WkHKxs1Yc8VtkkVTVlB9pVDoOsE0zeUdq
jnrehn6OsqVCo64o+mytuyyJ4ycfQHXXZfCqIlBXx8wFDdVDFPpiicK31sqbeRysLX91Fu37b13M
TuEk9uE1gWL1KY9FJ2dFC2fxSz4ovHJpTY4zXHkPb3gfQQXQyFKqva9S/nFX+WgB5heGpkWBFNBK
d4MLRwnVCgXKM5JTWMx6A43bZ8dzkJijFzKMY7Tos6u5tC51uKEsYZ+X1ssGYhqjNVOVgDtwzbYU
qwjgPM95faCMjtZTTST9E2aHtEZ9Wx8JCfGdgPyptLchE9/RQbhE8uT/AMj1r3nPNNIvyijQ0Pfv
1s/ne4WLjFpWUDtK3HfBEUtk7gAHSFiDgzg/K7iL3Fx66VpZwPQFOWi2sRvq2Gz07TCTi4mBW6xa
KV2GTIiC7YGMKvmRu0tZ2/hf/NW6ClPxuCfQV9Jpk4N20bNhuYXM+OGZNiomSEcnn4SK7Js71x7Q
gX4tb8Nsqm5mP5yBGJNq+iIuoLAMey2YPUImm32hRg5+qcKWp1j/9rC8Vj7whcPxFHcsvfjZItNV
3fRVocXUmPwoCVBXFHrHEnhzj9hqruUBksd240RJA0n32ouQiKk4oDOsatIQx2lyHFwsWllYGRlR
bgfIEGUqLToK3rw7BbUpnqmqy3RSmJM29PyyEebE1L5/bglrquXaK4pNAqekp5RVir1fhML14mzj
CyqFKUrvvjAG6JN5XFR1ZtlO2/RnpoIsCB1GMaP8F3yoEXCtLNuUstrIY1dDJg+S6x2C00Zy7jci
gG67ur4YNQVCDVcDW4XLTRhXSidO8Ywly0nwnn8pXzt8H5SPRlmfYR7lE+dfR+QH+QlQIuYFKDjA
Rimqhv84lreXtf1D6UKxBk92hIVGJIHjZ4qYBXMzkVXxj2FMFUpWwVbP+GMyvtxt5hUQp5FMfYv6
20DVoAJn6NL4l3iLpu0Zh/4ttfE84iLAGXJuzGVH9pnbWs/G+6Anbl6oHSms/ILLU+7ob7PrqM2M
CkPf0VimQoQqQQhp2/NmMiqPVy5DKySHBTlbJhqVA8Zgq/hMuhRFGTX9KWn9OD2qZZHqZCpCnOiq
iO4HcOGPHA7tjEsSjKPNrj0XQr2KLUWfvanFgvBoXYk4cIfNB4W10cEjV1IeByg8dDcW6XVpu1Nb
VSRQ+51BDtI4zU/mCmcZ9Tg8qxElcQ/RDDZGhsHDBMQOuWy7oQxVrFmTN8313MNhi9q0ayBUNVln
CUHP5b/qlCvUyKxwzr8LzxF3viQpWwFXizmLWYQ7X7jYDQmj5vc3jpy3sbp3Ymao/+4dKMPQpCwm
OAPiADuhlNVxqozsdLVIPLNzt7FbS7ZPX1gTTbAS03AbMtUKGTc2dMfjePNyi3XfvcFvh+Byi08m
juIMDy+qaGyPUSrhhgtfrniV6ButtCAYuKmNRwvuhIUTNpLjS7HE5rRetANmnZFxb3r2emKEnOFV
CO1q9DoePO0hFVY1vDN8ZF2i9Hi5E4gK3oeMIfXQ9hgXucrSC7G8oOAGWyCZ3AGgkn1NX94B0Hfv
RIeLCe8oS4WphM6Cpb3mIY96fDA9MyCVvXmEE3Oizser9MI5TfY/kM8zW+g16qKNG5Gv86ZH9UGH
W2GDwscff9RpBM8hRztVtP4RQW49nsQYsG0EwT/m5bXEdoPjPui8KBXwcDHS/OcFTc7u6VMGHsMy
5s0xKntbD3Bu82fcdadtIH3OIZNVtweoAk1FI46A5LC7MwcfTwyvprTcv5OceMVegD9iWumnoeom
o6FjQ8bv9/gV32QAyUHZwDbdLsvnUzs/7YYYPh3W16Ru74twQ5Pr/pucJngiHFIdkfb5D194WPIG
oCNe9np9ICGtoV5369xdrO2wrN03iI+mjhQjvgHcUXwVN/5sf1kqtcy4bJ/RjQ6NAbYJmFPY9/xq
1f7CL/3EDUYBATmqGG0PE1oKILaohYKBCB+AQgyOTPRM/J6KmDvWEK0qQeExEOppn5fAt9gJLBFb
BV/MtAzdKlbbbaU5haDfu3BYpHQfVWtugUaY02DMd/hyNN1pZEas4XHQ03hRR3GSiL/lC0Qetl/N
t2iaLqE3snvjxnw5B0o3gtWOKQY4mP3MXusO3aPS5Q6rKZnHlisGpfMXzh2lSqGBBa20eQuqH/b7
dd0tpOvcvO7DhkeEn5BlN/TXItmT2EEqzn+weY7XUEKW1lD5cH8SxLBPtsTYtX30YVYrcBT0Sn0+
1gBYCBDIFI9SXPx4mzc+6XQWolAi9C6L/nXPMkR1uNQ7GK4Yi9UB2M62R6kg4Y3SMOYE8p02Dmwp
oi9xn3DO++BIsS+41vhVRScITUWxYgQO9mpsfJxK93/jaTnRR4NeXcQZaP/35nkoEPAVewx/8LJN
RWtAcgnKkfd1ucw4YlzZIFSvaV6DdDCXHtYrgvm0ujffThTRI0FHSUkBq2j77qUP8qY6Td9+NASI
PU7Yqu7+3JbRGK+DLi7y81+m+j/BZVk+eAs7/jJVFX3SDfDCAZiQu8GD1pkmcsV0zxizoKcePxE3
V+u9XfNYaqnJDmGQuT4PpgHT7SsVOgB8E+Ai2iVMiupuxSU6U9Wopxu6qKwZqJrH3BVoHJThzhwP
sv42DfCUCBzieNtEpBvunSiSzLyPS2E2x+gMEGkAX5f1uZfkiyMEfbBpS0vo28MKN30yhZKQsGOY
pHWzlihuEjaMtPZBGl1GfeB8S8LkKk12inZxBZ6HZiwhS5hYMeOpTVwKOrwqpwrS9ADl3ScNFAcr
8CXSO7c/uF2mQ3MWKnSGXDmQcStggyEH9YsLg4bvPXKD6OaJzjR1yDOrjf/X70ZTMX5pe+3NCMh6
cDpOA2EIfU5Im328GzV+vOuW+/2h3MUhoGBm15bsLuL2XWc7BMuRdbWyfouvY4dW1kb1uuhoHm2N
e/aedfpfFoPZGj8Hqnlcci9gU9DUOA9fbefkDN+SXZDaH8hdc9cyqQ4z14xhnKuEro3RQUFYLBkV
2zLaSUiHK3zU9O/a7gg3Pz8CAnYv7sgTHlLtN8UdkyxN5B3hqyvbKPtDTeEJm6puz1+0eZNKyD0N
IDR5iNNMLKrExOlXQytyW/Wj88vXlVKe4jc7tZa5f/FtnBxlwlyIiaV8SatcKtjcSE19gBAhJ7wj
0o8pOUMlOD8Ejj+j5bcA2SbgiljuIJBBNgPBmginNlQCSRKDpf6sF/vjeMUNuB/5T+qCBnY5LZmS
h0KcPTcDCry4bcR2K1/uk5GPkKazFoPeSgmcvHnvWOk/I3qUUgHxD9nXHWDZqmmx+aWGDjZ4S0IS
vveeuiFuCzw5raOX3lWGftns5gD57HDpx7uSyCJh2gvnbKOqt61ZK0JkHFUEiu3bdWCYy0UGY1UM
Ls5vCuehBg0zbRpJ994krdhpt3CSk50adfL5+i4ZgEQPNR0gS7uS7vNgRIkKih1S26vBIvm+B6BL
S+3qS+pG04ixCiu87W0qBGZFBnxWJVPghUS7XfJr48JfcRgbEc1+A4xq9e4ZgOdoFukT34iYfv0U
Kxr7XXkany1V0aLuevmiy0mulQXQEJXhv7+ekpNQ/vVUdl+BVgD45VmRaSwL2GfRHeZ+wY1lB7wC
EUo7czXP/97iIhEAgIxh1GQnMUHn0Pa/N8l8ZdSrJszdpoM+dXc+KommjsDhF5dwkWQxGQCuWQ6j
zS580MaKFPoFXyRTutBu/67xCIARGFGPc3iLT/X8CZjI2X4ZE082ZG6OJ2mdmNDu2fBgnLwkXqLE
ix0n7ZoZSlKZEj3lTv/Af517Wilw/Af+CwaoJr+1VTJO5LntzYYOoqBsOQRyRD2syzxblUlDq8Q+
pGmp5znB9yACs9WHlClGJIx4N+BD1y0VwuGat7rTeMPgnu04vIPrLx9nxsinr2dSwj3cIJ58gDRU
2KAw+/2CfvFwbGlE9tgKwubX4MadBugcXIjJ99CdX+zCHGq8F88oindkfAvoyXGM9DH+2tdjnA9W
meHiw7Wpptpvb3x2QJ24/g7/ytOd6L7sncXIRs1rVrf8TCws3OmVxmLnpMZeW72XUSUGIY8i45Dp
g8lgq/LYFw1rl6sr5ZOl2v4QmYEZurafsLN/FaVUfUvzy9JHzfjic9ngLgcrZI/BKTBcgqvKQZh+
lIdA7O9+2uQGzF+GqyqH8g13tgx4L+8PNQa0Vl/8j6DUkNg6vnEeGoiZh+KL9u8Uvi8MaqPCbRpr
HdgQuPp5w+OK9YZ5rr4JNAwOK83A8+r9B8Yq7dliKBqnH+u96IQQthRbkTQ2cYkMNJBrP/0Z5H0u
k2YsDo8l+3AMcAjCT7lcK8KOALdmXRkC8fMikgKoyU9yJX5vvmpJ4Cy5iZDRcgZvISasx4RzV0Oh
DOjJhtcfx0pCttUxNoYuqu83MU4xOuZP/u5sh4HwM7+GxojZPXlYDmIdx0ZJYwUz8PntTZP3Lgua
U+/AD1DBJhGRHvsv59oPU4eLHPp1FBph5Ym71RJ2giBIu09a7W5rnt09fEBZL6yBkUH+0Nzha4Nh
Nlzb8lsZOApatF+iOqtsq2qwERkU42C47SaVvv43JHnGjpp2txDgoHm7SsH8+c4BblgCoL2QB75q
xN0lOSy08iN0RcOtZAodx1Jrn87XRU7ocO71cY88TjwXCN+iWF9c8d7ryStGJUGxrsbOmxRUrJAp
cDh9IVrUxTSagyHl0T1IKIgSapfPDbW4SRW99oSQL9OSG3NribyB6swz7u16DBpnj+k6ErocLudS
J29+Z2HlzhKCUqRDXCDqv+u1kB3xfWAkR5xtZpk/dkMkEbKPGo7qnXuFzIGR34jI4wyvL9+c3z/2
diiqag0+qXctO85S8MCdwD1j6wycOnZ6onCyF77WTeaSP0HfXig9FBk4uJtAryr4uHkMYYbnA/5n
/QU5h2/r3l5UuqpgxyZ9D8S8Prp8YFcdqRWQvYCSQUyCDAnUxdYCR1ZFt67KSPukTGpZUb98RtEr
mhnPa7j03FKVWLuu8VLmlrPrhBKy3qQ3phrc/qSDO1qax/4qGlO6P0Wv99vvCI+iigvBKi5HbFJU
qQA8qXiDrg8X/tRPttjcBs1L1n5NNgJT1ud2D0KmKBdY/fjRyU2lWO74KN0bfJHpG0fozbQPPXJ2
lWnRANtezHNh4UGAlgX9mWGT9hFp2m3ubLcrOjcHa7Ppgwh9mFomMu+VcLVkRzfjjkvbhRzmia2h
KFZC+wn/FtFNaCq2wqaB6RGcgTOCNPDVHhHl+5g6VBxmaYvrbLjhDY22cCB32rzoQJyuIzK6+H/G
+9k0n+XjBqlDvPPkAFHcOTYVSMIDdIC6pTb+7DfENUR4vfPiMGNdalJDKxaJIAVhsb6rks4EhWmj
e9/cF6gTDjQLkuLFrRvoRisi3kyxy2Wsy5vP9r3F9ott+v+EQcwKCdAVscBJn2zD771sKFYybgeb
mrtGMGuV4EGZ3vDFXgdtfkehGYYIzRz7CWwkm+Jl9o1iV++Q06E3SFW5PRti+7uUm4O1+PngLkug
TLeoBYyLTG6fdu53by+mCYYsDBYD5EcwQEDO9waMz75oIqIchbg3VCNhj8PzZDQl+UNwnPMd3aaX
qMChb7qwXQa52E6PsyH5jv6TXU7UpD+BmRR2j8vaEbJZa/9vMHaJFFXfyQ5RIrsE3REplZDkSfNu
8znk2c01FNsaW3yuommSQxAXkiiDbW4pxqo/rzQkHTtG7XnPbegut955RYBw2dWmf/bnxxbrCdVt
0OumMdvSSBpAoxpSKS7KM/DBJmdMqZvEkXCwLz7vNywjiltn0SdKRomDb4TchJYftFhi7WOFo65J
dzDrJlGnmbfuZTiojBoXbNPPGHvfZuybaTdHclrDueOSRPIDB7d84Jg+N1vnMQfK/hBKXTqh9y07
wwUZnhnfAbuf2hGVIcctNw7O9K8zKFaPowmVAF5Yuv38nFFShZoV4FppqHcdwtirJzKNXNtPfInT
YYa74lCYj+fztgn2cnaibO/dpK2FRifPCEsNeZHTqDCKkgFt7sUuc1wzKWrcqhGBmYac24HEXKPw
uPqbvi/QUIePuxSB7jnMEGmwlfp3I8PZpxUnDQarN8Kl0iNVs2MhzwuAkwdvEYC4r2AdTlArkycR
2NgMs3c6pGeiNNN9kyltTq72tmPZZ0DXRbTrmyRtAkDzOug1qyWyx7ozqoLJaMHupBi7JC3sa+hz
OL5icIdZi450gXKzuSASL4oaH7GrQLsC24CVruNl+3/DJ8+jLJhFMTSVA+RrVy808NvfQSIfRZu8
uV5TGHJndrgDtzm3ZM9IRy6btsLr/5LsiH56dcIMRoSQnHSTXokwOgppMjSWRr1D4YwfKsAv1OYp
qW01dhkcHti2GNB5W7B2mMO+n7keR+H+ftH4ZcIUoOIehMm86DKaIPSp4/cOgEfJIqhKnzdWKA/k
fDK1WvPbIVfOeWLEylrx3LW36priX7fyKtS4lI+HNs7OKu6jkCnnnXQX4yTmmWEeek/BIkdJnbOV
oe8jGAs7IjZIkIL+ua9J7IAl+rZMWinW1CsGJ+CaXxOiNUrpzfTy5r9AnSdOk+ZXqJ+f8/tSuF0x
wp/gVn7ZmMXOtSR7skTmwoSsQyDwqtolB2qMZ5gOAhtUHDGXtfXuj1eu1x/+wSq+iTAl5JesvKGb
wRCxaO43c9halaOrXWQebj9Gs9zpbgDKhXW9CLyp0wqtPg6M42LZlOt91ANH+WMAHTgRVuBrCjO2
2QS3Djki/P0OmjFR/1RRMKlBnWjOLYyFqE7Gkm3/EJHqsR3WepEzeK6hAROKOAUalbli+2xToYOk
MvYjCzsfiGDvtnXJSrGuEJ9O6TMyWiKX4Lm8M+FH8beUzTTp/W2DAi5YakiylQSXAutvq+KLsdql
TUYQivQBPS/lwApdby5fkHDRIRmynaPXep0F+E21ajNHIu7XTgE+eJj58VX0TUqRayMc1TteL3iw
B/PrPDTFRUigDWlqXToNvC6yDHoKZotRxM135tRMzSPUy2VgEziHhkRWsuGP2xO/OUTRVyKN7ziy
Sw2EQimznyv4YPDTnkSSupO1v3nuyK+dStq7QNEOMU5oO6MGb7ILbjpQdrifVJysyPayKoXdpZW2
Y2hkAUPB5m1QdImMk4MM/YrfpBrFxFntgHY2GO/WRtbFh8OSEk1IsK6yF9pdc8MxgXW9FNs4qhJO
vQOpSqNOr1BlHuI58aIPcLilq7r3ak0Qngo52k7ivSCUZqWw6jh83MYig7PPQ2CDF4RWKYww4tdX
pWu+CAWNlh+T0KCFoINe7r5va+ahxVrjEK3SmPxhrhOMC7E4V8OdCpwrhBTWe70Y1+nlvXmXNsyz
uYp8gOfV+XPJcZQrgoHznRQ31kIMVX3JcAu0wwR8tqss5NhvFVoFuq0BUcZSiqcU4W6PWnDL3tpf
kpPU6KhkwfoRoTPucGDiZOEnbhNdO407C32z9KNZPdvjLSkZ1lo8Aq5dpxakatdYsH5T9sTzbWXJ
OOfMeNjIZtpujVyCiHrrbMekITGTlqhw51/s8p3SIj8YnuebaKt2jyA5+yWX/UOmJCNhmUu7BfMp
o2UQNCVXfMEPl+mGmz60089yWUWYU/Q++tkhGA9wSO2GlJiQcvLt4xzzeYah7OtWiJpwak0B+nOL
pjgRWmZ8jRXBKZtcEz18BbfIoG5O5pEfy1ObSTibDeh3jOvRhs97sbtMkcFibyl4carPmi/ocySu
uAIs8wbrG1i62mwOU2223LP1ME7Buv3bpVZo08D6s7I2aDy1kfD7EnxXoUpvd0+McYS02xsM6i6O
NOthNtZevlJm8BhIJmBlg41bx8PM6n4eriR4D/DDVz64YUfXjYTyU/Q0A2jv8USaomvClXlXPvqF
MtlqTfabo8+gcEpPPFQDQqREFHERsT25RFI4XsQYVhpN2AWzf6yhPx7Tl8cx/BeTDF6l6BxLvJ1H
937GlNtSmN90++40zJWEK1XfpJTqCGpREhBGQx6vbBD8Bk/KHTr0GGc8onABmyE301B33epy1hPb
A8gvX8AGi/GQx5TUNfUN+H86vSyL9F9Qhdsfkv4qBlBuPExC2+FVBNSQG3mBxDJz9EMz63XIjscV
eWUhlMoI161PTPh8w8lzGL60MJ4IZtmOaYavHChL6s9Exuc+oOF+zMPi7h4gCmptSSFav/yv25jn
GQLOBnrG/x9V18Lf4tLSXgOb9PfY7Erk638O8RL9fMH+Ra2A/IaIZeT20rbk1P/KtyH3QAN2MNLm
eue7suYu4COpdi5Y7DpcvqJefplzjajQGdQC97YvPOMjT4cL4KimC4Pr8SbgWbKuLfohvbK9Ifqe
s7f9inuXSzp+sesk8gBJWEP5/6KAnKYHrCTVCt4L4nZ7vh8WAyffeBeUlXlRBY/GC4/2H99pHZCS
LjdEyQlrm21BMwECBBv3lGz9zhLSV7/Y1nltxz93C5ElsFtf5tu+kiQvGv8oGB+NN28iQ2I5qBFG
+gqkZ1jcAu4oHr36O+jr4TJod8e6paVIffaMmP25cuTHLPFmIojUJj6axVRG37Nw8md7GrctCk4I
h8htZrf/qsx8SH1P1xwYrZhsHsMYYI4/E2cyvqIPEMJs80fy06qiC7gIQAZqJ+NvA8Cz1CskYgUd
vcOeLbwaIhVYwBIFE3rniFHZ9/gGv3V1KWqDwFvMhqJyXgU2cheRB6T652SDG9lUC1NPvaUQkKf5
+t9/DN4BNQ79c41zHL406AnZmfosH8D+CEd4hHZpLp265lCmQFo0MhLdGLN0vlmFHg8HAmLSIEMx
sQINdirHYClW/n/kL1LRfCnihyV8Q6ZbvN6Umlf6ePYI4fbmE0MVw1bt89bLdNrtZg3J3rOGkMsp
7kUlKtcnb2gIn1OMsI+SoYGty83AmA7pTdqVwMF8tJjeFny6zBnpOzGoGfmjrOcZgamJhxhMa70g
M2WGHEq9hEkT+wMbEEs/7Vq/7xSzKch5fFj6yM+yIzHzsUN1pZ6fTpZE2DW/vEByaN+/VZe2FvYH
muVdCmXSmFzqblWRSfGcEbG/n30FRaprS3RVIomkoYfRsYVxch0R4l7EvR4gx+A7A1rItcoXlMPZ
UzWZiN15tkUp+hitJOZEWejVj+gZE1gma+9q2bAYe9ttmL0wGg8CHZy9zaNTvOFUorDUsqs/aHoL
rrLxfkr9NbPTpgJ2aCTRpPD2GgZ7oQIhFUZiW7ads1Ul80ftFFEL+kOewQEg1G1NWXQuUGeXawQt
rrFfCIfMBVwz8uqT6air/Q94sawxDKcEvl/gZlPjn9EKFtrf4PhomoX87Q+YeSXNweLdiFWcUp+W
YVIlpt027+DJK6T0CJ/wJe70oIdWfKglblpFltGoVUZ+fnYhWJglDVPCE3msgHbTVb/O8a7gmvZF
Wu9ilzpOtL4mwAOhvPKksz8AGU5eeDJuaWH+PdirPs51tbVmdjniwV4rJwJBIRN8b1vanDYzMuLv
7AvpIOu1S2vLeQhQM7U7ercW3/TRqd7X+VboRRPzKVEQiNbnxqucn+U90R8vYcmxuvGLrsDTBBSm
Y1IbU8ZHFbvQKpTcqFE6d6p89HeiB5usPqb6RUUq7fp4Bkv8l4GrMGOdyA2es4UyQ51C2eJrAITo
9oRTQuKtg/sQ0xKCd9uCU+UaJe4ze95OkbXLPlrwtIgZnocUYX1Sl/1+z3POjwosgYNT6OiIdqQi
q/BZzIRGBDtj13fBHTuBf3iTO9sbSi3cME1KtNDSw10pxMigcvPhGimJam9qaDNRE152qpxngDcn
Yu+Ggqf/SSfAOgec8MuJVNxS2Rps9b6rFn5gb0hb3lxS0wH4z4+VUGe3PLW2s1GsdQgAakbH5M2H
AxFlV1+h719w4aQQN+R9tsKwPOk7it4S5YlmZmd7ERCtXx0Zl79ZMrmGwp4hkgUTgDF3oUnLWtEv
75BFtBvIiyYIzsWYpJ4t1nhgLS3bDaJxfXwRxF9i8dxv5jwBOdvMdIJhPrl1UoWS/a6JJzkbBIDG
UU7EivdBpYTTX9nYrldkvt0LF90AoLF0WdBLaGMccxWsk6qld+9Sumy6wbLNs6vLiEW+L+kuUteZ
/gc1nN0WXUZx6wu+76vlIVPXhHmKI4Qx0XWMxsyVoeBoWEHs2YSw3QhE7TVmm289BMxsBDQm4I96
7Jncsop5XoF0llAt4P5Kb7cv2DSLxhUK3w5qZW5UoSmwk03i9AYmoRL2biAz1/bgN98KzOnZ8UoN
6xG9xvXq4aGmcgZVeSj8N9OX1XSDVVN//em4/Gd8h1oz1r7xUs29ou3JKuHi3GhmfYmYr6Um7rp/
5W/yYInntZ4+iEOaburJj22noQYhACttc9b7pWTfilT29pekEejp+Li50bDJo4Vv4/9g+5q3a50k
zEes43TZfQvxF9PRYobCuI4XA48eXMfRgzBadCQFbSSUjYoDYzEI1jgcTwd41IZxHIoPL7uXVQ4I
EU1/qIUPKHMgMDWcgp9C298mkP4CWoNvJS8Abs5dJF0xF8IU3HVaWi+UWtPubbiJG+P6H1nT7Lkr
CSkPoB/2wZ+xiuFkoZXyhiJtu6d/q7xfSfQuzfk9eYuVgpTtXUVoLdwdDe0gUumbom7HyWkdV3DR
XkL/1vXJtgcMWE54e+AcFf2elyLX0Fk5OVZAqhEJnu/NCKAsief8WSGMFnuWiNOXZPtrwyRRmtfp
Hi7A2TD4PSbNuYnuTPphI5G7reuGvOh/q1oGG8BQ98IM5HhTu0L4jj5FgHVhFlsFMFBogoa0RvoN
Pyv/xdNsuSH7oE2lQrkTSOLNy8m+xMwQ3d4npwroDcw+x7z7ZTnFsh8/9pYww9WT4FwyRd16eJzA
SXYGaqiZ5bNyFM6T4/2fb8SocuK16Rwk2b7OqV1GhWTsMjv1ZOq8Bdj8PzfGBvc7CG/Y9Wt7dII0
pIfn/XwDIINfCWBCdEZBZYQcQXgylwl8TOTMKTE+jnglR5MVkbbEpoSIHSmrLgOIUc9IMUcPUGlL
mzJM+D1O2uR+4R5YleCzOtl6OhRVKf3gm3gL48ULNYmUucly5CQ5qfpxn3eOTM9cuZVwnbmEWgyq
I1PHYD0Lg6iGIKVxN6Mtq589guWDD14IYIZsy8p9So/SimAQr4T0Py1poERzgej1AzV9Y7cFF6g/
9b5Tigi0Q+jnafBGxwCNjb1aSEFQ/+Ff1oakol5tgfk9wsMy2ZpOF/XpcDKWZgFGyOhu08TvzJLl
UorhZdTSq/98G27Q66PDmvsFPmCS4U6rPczDENavRRQ/hHPhGElXfFoPkLhTCmERgPinoDHzzh9y
K5x1ywCvn3h6bvyOs1oWe7jNm7BboG2Zn+hSvhDgL3Da6THmZmJSHT3l/PGvm4ZtBlBcn7qjE9ZC
dS+335hIJBr94Ptuvn+bs+VbmalvQnnEJz1bLvpqXJ3HAQBM/Sjjx5HlrO0tJ6PyS9r9p9HJSybo
q52teoisYJaOndT8jwr208NY0DKyOathEmlONICSu7KYKont+0Lnpd1w7GSX8KqF5W9gmOhwCZih
RTQ3In57mrbyzuz80iouOAjzhT/wMc06PeRFMA0Wp0omKl3epd20++/8kBP6CiziIt86j23eK28b
iPuF+cIwB/7Fzkm9ucAR1WN9CJgpkompjMAktk3GTqrDLvVLlckWorat1SucT4azk7zWmw1ZBo+M
Mf/jd+pa7zfXXJO4xxQ6QLVKBaUFj9CDrBmJRKTBmgWdY/17zFoTDNNB5ehUv9lIcYEo7w5xIwwF
MVSyCOhSReYXqx1Q/7m6n/gAgBOjv9DM1pnM8qZn++n68CZo+pp42WFDFZb68A31wxBNoAkmcQF6
xJ1K32yzLw3JbpjStgX+Q+RE8s01j9/XZN/gMEMYd0xMuXS4KbnaJEPTs6UDJ9yuEBsfx9fCl9Po
jIcKu3lmwhLOLPDLjthOf11LmC4+fMeNeaztD5DyAMwtz9X/uD2HaCV4F9sEVnStSz6fTYl/MTX1
6QcT07SKQM9MLeBFlr8kGOBpI35qp6yrnnYoVvlDW5J/gj5MIkiVFTQ0YAMpXcovMD64E1oZQdbw
OVDs5pEyLnE/6FWGoMyDhOSvEpaRg6OrlwSpchCvujofMz9L6bTlfgcdCxnBhX9tNl+LdQtIGxmH
rrGzS01xxibZs8kH7JktqMfSb2sidvFXRpxXJzCs0kXYDcCfqJ8hM0hDdlYcQEUaybaPDREQmquT
J4N1NYZtq3RWNZOa7i538XdsVzI9XHJiaCxMtJPwtHGxsdnZpCCb8iZi7qv57RUlw/W2yGG6rO+O
zhKqzyzEPn0/OiMCYlxjsiPm84QRt8juXcZa1P1lOxTLoM2oV9Xzx999eOxl1V4v92rp9prjNWhK
+SAziERabiMC4e5tN6mfc3dVOHHpmDVBQceNH0iClzFCtsxao2CosSmcvN13W8qavUhm1vIhwdKP
OguVGawTiw3gu7ye09Kjk1DJOahcrIKX/dO4H2tRBJbgg8UYvkkCI7zoWCX5oA56RBQ2YESHxEeN
Dz04198yC3G7yoXt5viUWMcLOrL9sXpyoo5wlbuxd0CgTq70EGLds+seCtuECld5UzKWkfHUrehr
7CaIJTxuYfXMdRq3ad8HKfxJuo4CvywT6cVb5nyMce4TxoxtmRut/NzP2GHQQ1F5tflTgi4nrQye
4biL7UvoJ9P5Z1ApphRTe70zvGedCu4oIkENY2bT44SWPPkDLcTMeRcZhNO6BE3zoWGj6ldCW6QY
X9o4TamBrdfmrAC+p4pwOZMHlr+lRhKg8A6ZCOgbmziflwn9NfK9mMPyB9+GTDPJXE0JXBpDGXQV
Y2jBQLImlTxXi7FANWtwoot9PgYmpJdqXQXJN4vkSMmpTie2kWf1w6g9tVMSYktthP9rfe0oJ8dq
KQOlfHEWUgSdWqt3Sbr4ydBC6R8k5oUZjIGTQKSh2yRMuqioMbGC1q/MMopTPET3NtzVQU7NCXcF
UAcScNSB6qkud7PuV8Cjr5W9GIzSU+AMYkbMrNyHdPNBYa5ITkAUw1PlTAPJmysJss15OTMjRzqV
hySKZXsyAe5QI0QysSIxazccJ6cLwX2QDDd4SPTB2+WoKeD3OjGSq5Qdlgk4CmJ/05ParZq5qWE8
PWhOkkA3crtKv0l8t+gkU6pPoGkJ/xfaLSt7yMFrDJ3vuFRQs9WWPrWfkwWobVBJUA/rAfQe/Ma/
rF8lc+HCp8QlloExLW8V9rXvLf8fpeILwPiOWkP4YMkVZTkb9kirjyxmSAzi5oD5NoVAiplW6keG
Mi21vgwyB0UpcWWIKmMl1t04DO/s97WCfKpC8mxCcbr0emv0Pz0P0y75Es0tQGNv2uJbrFSviyk4
kJECarY3oL1nv55N74pSnGwAbV1tjWwqcMF1iZRUTlx7zm4vVVXshKG3pubUYWEkdOtyIDYPtk/j
tFWvH5ZM13/gZpDu6vftg45nvmzWh9NFrUkAs/xKWnewtjDJiNOE2iF/7zhuujW3H7JBSNU+RXoy
hh1yUO+RWGVSrB6Crzw+9unvQBIx0LkcOSKI+HrcFR2NADgRpibNkVhEN3jqTuaiJTFXT5FFl9kC
dRDRZdefiKaQEStNzGm7OY3/K3kypbdeXcS+q2uOb8g9jje29/Nit25zgFiN8bg4MzV+t5a+UfzO
tIFBpm59BukJeopZ9eI/m+YSkoTmzaXzcxvHSuD2aOo8qR6OeOFU5yZWq0HZn/RzrlPCjH9IzfV2
yyiY0Ni2GZWCDB8SRMh2Ja4Ama5JzpLcRHIjUareZ+/Nu+7Cfw5/Z5dnbSVx5Mbz0e1gaVf9ySw3
PYwKU4NJudWOG1yYaLNreJgrj7WngIDXns2xvy5DL6gYgkYYy7pAbOW+gnjgxZ8u7YUINGQTsa+d
jrE/vU2/CByjeEBVCKLopys5cAUd1PKFWwK27JByQpBqZVqFSqyLFUUSuEjU+ehjANndGmcdv3/h
YSJLaN/gTyWhjnRoutbjrqQh5YUU/YUIWeTgPWM2VAXSF1/VJtnkbYxju29zVWtgcrH4oy0ij7C0
LY9kpICoNQXJZtKleChK/N0I5hqjU0BoyD+52kP1hj9c36Y5/uWWx5hCkfatLIHAXi2m4Rkg/dJ4
5v7ZXEhWZUpAwrhnAzrzb8g6wrAsygMgiqwFJu0dsvA38RrJT7+RqQL2lisW8H/zCo8tTTp6lguT
FjKtn2v0if4LVWh9Uz+1FgeAFEGdZvzMIEsVW4rhDxKCH+fYiCtkErzoXq3ABuCkOPq5dPGLaKpv
DJKP5ddpsFzm1NKHDgP8MveRHJyTBbL9RktEOjm+Vlu5STCSMiOfpk/AJn9hhbPdUaerDekDwE88
ggoN6NBzNNEL+cBjw0rKMgDuUkXo6v8PYHx0JgLOC11rPhFJJfzR52t3Qu0WfX3jaTdfJkmLj9dA
3eE5AhG8mmO//wwXvU7HAASPPr/uwIWRt6buOk6EBAFH5hjdKWZ1BkVKD3U435R7fHCqiWwqKfbI
39Lchx2h9Ptj41eNKi6lIbrOQ8S2gAoTdRJjVKgUpZvKuMzaHxh0uUBcE5ZpL6QCP3fTM3dJnom5
BJkECnRRUj0X57y5auJvQaNS7oQoza7/ykUDvdZKa2muHle7Dps0LyxGkU2iRK9y7odEBG7Noygl
LC1wyoUTknI6/HwtJxWRp43tjQIAXGnfmolcfzmtcubzoe7I675prFjmKHZoyGc0zg0dhhf+nLwZ
igNfFJamo/60L8dNB2KY7BNZ1yrvtPnD/rE7ER/n0jCCkzwDkxA1XnmK2YH1oMF3E8dtq2QIbbOX
Ufz3aHuB/5FrI3WDBpfKsMA2ysr1eT1WMyETkmYc1Scm8lBmc46BamEPegaoz5oXq8IbejBfnLWo
HUIlKp7msudNi26bRCv86vN1J+Ervqf4XsTWyfwb+4+AQfKwLP6qgZ2z6KrCb2vRNi+5jzbFicSM
f3N5yB05XWTCNVAmjqP3K1VqGbF6bT0hhi370VAMxYpd5izpfoTouRbAB44B8oSxFLY+EseqamZz
0Ist3v+mR23x/zkZ9GUJmFltKYmSNXTP1cR2+VFqlsP6RJ0ieyjdzdpEasWPJmKg5ae918Rhq1Sj
bhCPCSP+f7paGInZRxFPabIJ7KV/j0Y7yWTcBoK+r0ybSKiutYgb73Xj0SNQedqYPwJEjs/mtFn8
KAsucu0CqUQFo7O+Le1qldiwsjHmx2hr6qazpoHqdBwfD48o7hpSHFuCvNsfF/zCWy2MyXtrVv8I
XRgbV5UmBl+iG+nH6791TqcHEBwAT7suAwvFAsS7UVR8wkKiwCYY7He5a/FaSkc5eZklT6ZzH4NC
RRAqq5Zi1DsRyEgtHkf1C/7LS7dETYWyS459mauapZCbMxeyVSTS0Vg5a8Em/VsENEfrAT7IOm1C
bPAaTwE6Tq8d3Gzd0acTsSxw0L+T/e/NWvJgAJX8NSXdAtOBHhpAt65zLDP7Z2kCvBvzKfr3hQjF
S/auRiuHlOCyIGiZqJniQHa0QGPlHsDdrHlZUNGaoJcATf7uWO3x9qWoFLur9xyamIsmP8Oz8YrQ
0x+ASn7NRaKKDGVmR6SuMMHOTX+BVgIvkWBHiGnKC5EtAGfyrpHYiQ/qNiz/IgGSuWt6ibB5Dvfu
9ZDsjU7izKYyV66Cf6/gUx/0flhWFGO/SkxbV1yxpJzC36E5RNpfLfeo4V6ZF2Advoux1m4PfqQB
Sinh1JXHztACjSClGtECTvQ76CuVXvn77ScsXUHC7RLr9CfCjgFEBziNXNFMIg505ZwrJ8Do7L/y
irYO/3CsWb5O5qjLF3z32cxb2bsWa+ZbmOsUf7OQZVKdHaTe9rUw7Sukq2/792O5F+zRlmtMyANH
eujITmbWUqRap+BESPpebxqZSm4LYN1YH33Ejp2bB8JL/RbEJ4I9gKyUubkNu9hMv9boYBbj+7CX
MMDVE/yZAY8jYcVwgVPjVz729w5e97ZuTuab7CxpH6MP3CHMpzq0prcu9VK2pQ2AtvjZ1RAM59Ch
a8yFKLLWj7vN0dHuE/+0jHleMq2Fgc2xDwBW++5RUQQi0mcM5qefX8ZqOnxb/98sBDQD2Gw0NNjp
W1dOxe0DgKbREX8EfkDDqmZSUkTX/FbenSR/gWQ/guR5n6yQvAyvaKdP8AJh01VRlLwkwAPEyFBf
V9F+Pj91AHtktGdNZP30wv36PuklGBeHoD97F406MBawgTObg8L2lqB5hQ5jx5tFCvSKC7dbsiXP
wWp74Rd8yidCjTV8J+A3kE/T0rbdC1U9EUqgaRJwl9A+/0ZdqFuCgwaHlKCHmHzJVYDg0rADAJVg
Eu9AoOTmxgMfAw5LpF5NZJjhiquWJQ/EPKk2/kmHK/WTEqFidvhYN5YnXBYNedzkytyVjJtHfbA7
kudV87eVBi+ZinGPlex3AW11me5Y8272yiPo1VDQEjAdXKbDXYzIBVsw/Z5qPPxc4cK0KAFMiI08
jKzqRdKTseoOtG51kf+mwREsch3nlKP9K3jwlUmsjxmOlf89KR9MbjSjHHMLDOtnn6Fm05h3mlPu
yyR+RgQH7TSN4/zyjf2slybhV1FNuSWhw9n+2ihUcEr5IZC25zmP90alTbbA+QHH5ZiIYCaC7517
K7EFDdkJo8TXKK65ICuWkyitGBOm/E+TlS8B9UwqaKrRDQEDfls3CMHzOHw5vDy7zXVHoAoBPv20
vxCCt5jngrI+QilfIYUTJ4Fv/xZZNUKNiBlMMsPgnzNyGmUxFDZInwaDaighGxZGVisUioIL+1Yf
bd6zIyRhM9qBxF/3/EHnDNyJdF8bxgq6ua/TRCk+oVhKkq4bJkSDjZa7QMTQfkVmBGtA53LvfXZH
3YYtW9EQYm1RuP/LiLvuzzc8PGeHyCaxYVRsR5jkHJgHFeHGXkB4BmWjhgH73DQZ+7/Qr4bRa092
Rrc3/EcDmQgIIE9KDkizds2Rd27GcHBLLce7GZxFqp3rVOBnF6vkUs3918ZuoYjnmyneoOIoHLAp
k8EVR/bfU70xhERnH08aON47sB4PSA3/yGraL+UqhLanAAvk1D6veM+2mnUBd8gGgFyF+ZmGYrLQ
oPloJdOKke68XDxxRcWzYn5UF7AsmrTOMTEAMhRXF26Ap4F+ZZ34fwr3pjxA9eOFju4HOswlJwWE
lskTz5deqEpsDaONEktBib2Y6VI8XCdrd0tXzY2JW0S/xZWeRG4AJoTNlxq4GiwUtAG8+3kdPPbY
4vYqlLncuSrsKiIv1dSSvyGuSRKGtMDPGwfXqfmrQ2lwTWM/ooeU08scCPOHzlW4iir8bheB4jBN
UjMk/tntRTu0ZcQ71xlbo/vVj4a1Mg+lA7Rszr03+s9Xmx7KVD5VYj9WQSAo7PjP1Z0/uaJAyXcn
PG8Zzgwd5kk2dPXtOPHo89uFxFaY67A3l/HD1hFMnLavEPlaMezP0pT7X7g/Yaj5e8R3V62ARKpa
zoRJo0UJXd/onSuVR/rRrrCarschXl3wZStVTQ8ch+qSkvpN+HpOpdLF2Q13IbskH+Ag1VSPbP44
79AN3dMKyjGn0xQTwxquylSDQo/exmyGEBB8trwDOGoApTXWI6716amp2BzcVA60FbEsJyEHjXlU
r0z0BY7yqSNhmJesrHAkAULjlzv6sd6pjt5hAMiQp+s+rajomIGCjGkCcNGibL/Om9SWw7NcynTV
z4iMBbjhpJJKY8zQoqKM8uLlDUu78rH1naul6YGZhLatbfY+widPudO2aQy+pFBI3lMvcQxokRl0
k/GhaMV2JRrGx3sBfbktSuKxAv/V/klDg591JgXtaGMDRdzwj+X9tOh8SctKXMsJktSNo+lLfbeN
ML1tiu356c4E6IgGaKio9+sTQ3ua9ITpj+GxZdQDZTqii16P5AIPBabbvxprBKpEuAxSMpyE2qpS
O8EJkreww4fpyddmTOCqQcf32BIgGzcPXXBGBS9JaxkypwN2LthWqZ2cKYGX6uY73+grW7Cdi6uL
xOUlhiFiYj4vVa4jXXx6dvhs6G6jxZGS3fHcriD7Ho3mmiHBtuH/VY8m56bD2j/kFTzkHkvPZ/1Y
amoljfOtV0JajTcvvKqRpDbt96OZfcIP+8wYYwiL0LaUypSF5vtz3ZRL7dwP6HJOuP6QCPbWI+AA
rynvW1Ztjt9e6V/ca1JMfC5PVANZlSP/2lK3E6PIvGDVBkcTAGgnIb0N5z+F4QlmBHCvTBAFNuL1
TD9/Quw5d1xzuF9YWK67eF8vkVJTkS1xmkNjSXO065FSzBwwkY7DvW0VLEUIOY7o9yShny41iQjn
VT+pA8e2zHfrTNUWd6UQxqMI1zSNiV2vGyk1Qfa9JauQLrHayR2KmS/YHNgWpAQltd2g/Ld81dkH
+ImgIlVr8FkVB9b6zgHGPPsPqblxQR9AA93+ZMf0E0LIdeW0Hk+833u4N6yhC0gzIyxJscht7NaO
y8cHm1SS39exaVxxV7K3RaYmOMSTzxdh8WROuGTF5KwhrteM5n4smw2FU3kRFXrBODz8AsLw3jrK
t292glpvqQjZG+uNxnjZm7U31GP+G1RrgPMYSj6YdRsLCUBBqDt4ssXiEZhhcOXaxMrUz5ScPRgJ
QY02JWGX00eNbevosNtCRUfgaav25uYdOUJPMqJIU0xsuHZtEkSCiiZWQfier2OhYsY+GNWyq3i8
soS+syYOZDowhp9Kld1IarCgU8YLW+tFBTyWEZfeymS2ijU4QFE7w8BxO0+ijOkGJBZC3OE08p4q
KbKX+5uk2GtvRwdaFMTni7sWf7wvNTrDykszMNQULGPF7v3eIZCXjDMEqqG+ReD/XAvMcADJY6sY
3/fu2mmf4Abk4B0BiN/uErlM6eIokC6SkQH+cN+YabCq8ml6X1ePoOFsbhL646k9eTS+407auwQe
yiR5EPWKUBZ61VHfe5r7ChtTD1vYPhOZDn+H9shd39gHbFBE2pphK9Cudc81l5Ljt655qXj15umy
X2jwPTcMwZ9Ha2FvCsxF/KatKsZH1lZn4bFRTEiUat5nt4UCa0usvly2T/ov5iLzdkiRSLPwOVdy
J6deibUukj16E5PqF/U6cMqXCRdcxrs747YHWqit31KJLDGrviGi0qZg8byCmbZAOvr0HPeZMs2F
2KfPUQJk+chYu0WIGizgidbhKKWnycLh9YuxhGxANdBSXRdL4a8sqaqcOzbqTGA4PtwbpGXVGcLU
mrhmg+96cvfzCXcRw9inKfQeFS00nBIyyHrQtjkkcfBhvklD2K+LkUcxX/1myXEguB3bmvGcX7C7
5Ouo3mY/CVIQZFjpwBhGouehSfNxz6y83pOJDYSvBBLk11EiP/DJoUXnP/FfCpiJPAiNbTKFwLeQ
AniaitQC5Nt6NwHnxb3WGQNOa0uBsVZyS4BKQfzZidnDzrJAnFy2czR9Trah16rNFqpe0WW/5C0X
U1W50oHT1Qf9tyeHTLfJKYXZI0fZnG5W0Iii8gsEsa1x4PLo+x1SPABsKLHDDqyc6R3ZylF3T0zB
ZGtd7U1uqSxWsISz+OG2jUCP1GxS9Q2Q+sfBYZTlViNNtIOh9dhX9QyfkwjO427lalaiEyp41MBB
Jwfec7eiX0PeMXtXVXWlMSU9sNLftG6+AIH9fEqLeBKqNGep51u0DFd3Emr6UhU3Ac6innhlb8QQ
wmZ/SXUpn1MaAZZ6uxtI659TrBiM7auZWXcFD10Nt30esUMzBe/y51NV+TkhiVhA/a8aFbrMITPL
Rg7zhM7vCzxZawHPjnXxBhbx2LhoxlRHyrHoOG0a0FES2/QwGHm49ZT6ddxojuTeJB8UgWsnOICM
sr3YST0sfKuvi56m9nYlqygP+j6wCt1AuXMdjwaB36nXb1AzOT0KBdSIPeACqUg8fC/BeXm4OR23
WjFPG/g/1ol5XpM0bqyIMDjIUYsDj8Y1JYUKPfZMBWh2QIiNiTwGjSBUkF6LmcHydDf96BHMkmMS
EqTomCRVhAMJQy3wNHTXQ6g4ipH97c4zMgGI0nSzgm01iAAdPkBvWp2mc+Qs3ukpa5WVsxxXIsi2
9H2tiVX05CxfElYU7SR2FQdR1D/4ayZThcLbxHl8kAEygFbY4cfATRi3nDi46fsG6Q/2sfWNR2a+
DxEiTJrph34YalzMqdELSCKgHm7fwoxSaLulDWqEnmvQPCt+wYrg69by4SDPKMEMxDV3mc0G5KxQ
k/1FRKCVFiZO6DxJX3tpgyFUNc0QQkFo9gm9HlBeugwH/pCYbO47Wyr3YWZ8w3hWWU/DlYeW/dCH
pVodhfFESALn8wepxsF/m+ptjiGJD0TwpgT67Y8GMgy8LRDumz9ffQaa8vrO8rNlfZVW6WaP2llF
PAgGHi8ptvmjqSCtNXCk5OzGl9b61b517Om1UGS1emhW2sgmLshD+1dzrZ84bfUsmlbPSr6X58+t
MPBM13qhsiFfH7llkVDaL4Qj1agquTxWvjq+aCbvTpqJofXGV5kN/UIl4QFHo3ouxJnhgA9WcOc7
XQ9qiC94n9bPFiFlBfPvi1OdSheD7yUvha8oH4LwSkR40s2/mTRA8n0nReI7ryR0/aiR8vsgDPui
auZQ3Aaymrvu3oChZdCwGpHf/Sx9fQOXcD1oe0sGjfHxtJlrjZC79bZu1wii3IVSZBT4K9F7x9AH
tQhXDOLerobmz83WbK+Ta2VVlndLJNwR3WhNtGS8e2oLPRXgehTRGDQ3GQgvbXsx2FR0KRFffb6j
Vm2xIMmZTF8+xvjbkTy9/czMuDsUBwG5kmX/L6pSUl7Nt7hBKFMKrHCqZ2MqCce7kdKyvbesdcDP
rYtMMz1dMkY0OCAIoB+ZiRdXns+wxppM1bAiMDt7fRhNv8sy8XXqPlSzszibomqYTQUe2k++qQhs
0bxhKT06Nw6beLnYjhBLMzqy0Fa9kvllRI0unKbJpx84rOV42LwAuVpgwwqYZZN5PuoC10jk9BrY
nVPQV60SXm1QjSNMbXrDXh3Weg7x2sNki4Z37VPTROHRcs+9ceVUtYqtu0vAporTFl/60Kwb7uXH
ZGbXlQbp27uPOrMkc7vvEtNLemQ6PfKz+k4y59qNKwOeOPrWk3l6B1mpwsE9SzIQErPhqsszJork
UfbT2T39noPMVXPHnJSieqg9qOillGKfLJ1E9gVhNMtkLY0HrHjhvc/tmbyJP75a/IJgn8Nb0Dth
qb/BUc96DXYT4HXz5gQPQTV1W3v2hv05ymL8vEeofLxmK7m2xDBdZt3ojLymhjFKHaxCX0quaVl0
0ckKcrjaivLtNW1AnlehswMzzaAu5lN+YG6ZVU/wkJP4HklM7N7RGtSayAYQXb3gTaMzg7mmedwR
rav5Muk5XFdMTHHc3hv8paRd2a3Omol7akY0LYSKCuEiZhKRGJSxQ5bEbTq8tRhmN+f9IwYDKI7j
sAmHBHQGMO/fClLP/tpHGwmUsI0o55zk4shmiFhb1D0nA1QGbXVVHShadn8DsgzC5Y/xLzk53u8x
y3oMl66zX52efC+qRkWjXaleqkcAg7BnQqPe/00ezyRjnqI8DkM/7JekvGJqvoUGRMQ5aME6tIF0
JZPfxX0Ridyj8/fZWSIVc+X4xshcAHQ086M7OXZnC0oxg375tCGjYxHNPlNhB8IWhKlOu0nNjSD7
i3Xn57S/EcprMU8Czg+b83PqgLlTVUXEWCau3EdBE2h72xw4DJ7KxAxbv/DiL9zJdX/H+Vpmmvqj
4JZ/QRkwTIClC4mJr4NdV1RwdEo+pNJy7fRen0oyzjkM/Uda5xSF96xPYRCySXwqW//NyQuDOed+
5iGA8P0RRKawyFKD2yhmBdfaKc7sF2BollA8YQ3FMWUKJebcuor0OFZf/w69cY8LPTtdt+8SZGLv
HAR+v919S31fiU/e/8ZRDcut2A3gTMXjNeGAd0VTlCEwIV2Jd3NsiA7vro4vxt/e7BBPwFHaSrIR
JlyGhwarwZXhIZUPmgjYuXM6rfTx7ZDzKeQoA44S05qwJ3YAa+M9WMP2XF3it2vx89j+t38BFVpC
0+zyCPpQjUEqyD8Ppp/czNIjasXtS0o6cmSYUTzXE1h++ZeYaWYUj7i2L4lySLFAJgGYAsXa/YZ4
sQHIEtKu2Sv2PD5D7P+P/ZZS0xUOHwWWZQDeyYhj6xqHiJw4HKPmoj09N65W62X3hdjyojogcdvL
KlepHKbEI6f0uMozJB12E9XAKgRrOEL2aMuRTKgF7q9kc0XR5gaBzLydJhD1L0j9b61GeEGxNoKC
Ju4Dc7kW/FtUR9qp3dJoQw8r77rQvE2LRFEthqu4NlWwE4lBQCnSLODpdKtCI+vmDIt/Es27MEu5
76IvHTYGceBMc7fkI6ai5YVbKQvKCL3VfzL5pKUtDCKNpDzPvUm0varycq5A/7hJHUG9vUEY/Dxk
15ajquB9XmXICZEYnYP3ULLQLabxYJn1cEqym6aQFbmicpCSvmCUIlnp6AxmXP1XQRUYN8ZUCH+U
4eBC44smGm2ksVFHVcFpNrIOpcqhs28/Alao1kfuoH14WVNr4e5urVHEyWPxaGkJTXUqiq3jCc/X
+VsF3NS/ewt9VvCjGsHWS/Rsm5bkU/o2cZpbh+lpVax0vFBouJ8VQyag48OOXySjaacoIbPRK88l
WLhZLCF86UqtHMNCFwzElutd4gA8QRcGRb17u/RrhBm+70x6gqcbEzbQbe+oN79jyKUqmIyhL1Rj
OWXlD4ye45wXwYWSiTNikA7nWF6rOU26/jh587Q6o/ntbcbgfLFE0XRpJPdZtdVVB6c+QHTV7iCQ
l/41M1JVtRYawEnnFP+WR7hC3mhGX2mt5mnHjEld3AXFzSzcVZwGfjGvhHbyh9ZHw4T+aoX8iiqG
wbTAj4DNG7uIvNuE6JOORLyro8Olf5l/blz9TVXJ9LvNt775Twqx0j//i4UtoJXUgt4s8Pcd5bST
lQBdYNJBXVmzMbyOD0jMZBUzrkpowV+vrvld/M0YLyf9WvBWnc9qvG1ByWxf5KhHlg3LuyjFNI5o
NsZWDf/Za3aeuLTN2z2VVADYO0TzFqWjbEVDmSxNPC496Rzn4bc4kNboE4sjqQLMkld9GXYVVLrT
HTQ7SGRANPHibG1P+2LlD+ocX5xwGPEfMAcV4LX0slwwyEENLpzZ3jvp9WcCOIs+G3fsxZNrY3Vq
ctGfT1klZImmwB+vykHP8aADqd2Nm/I3UFWBjlKvu7AD1134sxHBTpQDSOzpmXoRuWWP7junCNDw
jsx14C2HWX+qsioCNPhuQqMPuKVEy8nZj0tkL0rh60Bbez1mrwZ9UFe3sCCeQ5I9q7nzWQoAdgAV
hRqFJuHwsn+FPRvZF2tbMAEvYOj2Iz04AoVGAkAYnRS+LvcQnZRDRR1aG0dhdTB/8R1U3MuN1E0v
cylco6KetOTWJf1sZpDmDpJLjtYDRikJzzKTayN4gBGtzUktPKqncPTPPxLdrzVkNN4P1ZHoWRAn
SzlR7Njc1DtiHVQV9WF3ZwVRjeEHdq8VDs24UJqLVYHKEjJ2aRYLrZcK6U/NP8y+s0XpkUPLaSFD
OiE9uf/2eZWgd3oUjGuDU2Ysynw+yxoRGEEzTCLxqW5ccpiXPZO46x/AX3302ShqWhDPPg4sZpgG
fPWqMtoO11/Tw6HU4lmSXKijSoWLYW/EEnp5zjsdXfcMfyxN85AEn1CmQLry1UH16N2esklmxeCq
Hhycr41IT4YBXi4vfiSGCzyYLrL6Nf/wpLxsOa2vUdFz4HXsepAxSIQMq8gXUDF8BH1XOEBbAY0D
K0RFFYUgdGpsJvviOAtxV3Xkhv92lNAECGj8qTXXINhdRRcYJq0c+2S97tKZhXrfc1rHe5lNl3q5
qo5riXibdu9y1IP2QgZteWALHLnTHgWRlYKfcBYwL/H5gsRGTlNMslQd5hhn2i0BQVcj+blpwIs8
hG3dJWvmBf80hv/HHvbu047ME31KKcwXkygLRdMTa4m86RNBn4hPS+poSGx2Gd3EYDjVV8NUgklB
H8y3mV+5JVVrJx82h8kZn3r1whxz9RryF0E2PhqKWWCHorY9CJCruoGoQPzyP+b0ZZM4wRjV2bfD
UcLGypXI5mQHJhIAgdIZ3GstOzzW/Ks7oA7i89lZBf8HqLHDA0Ugse8reHnNo8RwgtCL/ukf5NVw
iO+ryOnuxZ4Ly/2XVlcbq0qrKeXZl7/URlqI05JaA4y48VCXGQ72SLR3G0F9ZsEzibjwNi+ru6fR
DbwaoY1+6WOIK91XCZRTti+lewCZvA87pIUTc59+I6lvrelR/1wNawn3EPy8GDJa08WIhV9DvNK9
7qz3frY5rCF9cO9fIHUxFNmP/O0kDO8SSZDYX5Mi69+GbalDkKo3obLu6LhG6E1fJIyGJ4/baLph
y92wAsaaY/q+bKhYGJyOgzZBc/JR/cDTwKKecTK8jBzE/AqPMGdR6HRfWRegAop5ty5PmkwlzyKV
dNG7n+CvFL5l8s+s73eEShQYq3jGNinMic/nCH1oH+Q/wBiQjI7Hd7+bE3AOwvtNJl7W5y1eN8bB
RvFAIMA1n+xN/uTk0zGlt/mzqVHrTHSrP4n3ysJjW0gJCYTpl2CJIoXh9XnK7gYbj0sq2tnVRUGS
AcYlj/w4ST4UqgH2J3eJeVu3Xo5eg3V9bZ6imZAzDqXqjJVC6j98g46Z0P8piOkXkWLXEZwY08mG
33o5HVqyGyE+s9gQpGEhOmrZ28Z7l+o9FpJBMlWIYBgdzsgYAnbjQVDkBm7w/kXD9mM1VqwITh7+
5QBtp0S98eqxCeqZyO10cIVnRpbFgS7TXGWaiwvlxOZmGlJC3bXyYu7d2sSHwtvIT/6on00c4CnX
l4jFfetCeDIaKX8jUzp+nZ+Se05O/c8IBucjX19pDE793OUj4CGOtTvzJTB57r6hwpcJPsLNadk9
WcmDOoXFZMphryRsqH+mx2aTtrbRCNmSN1pEYI8Rdesh1pLD/eQXC5ID0CJYzT2mDEgeYvd+fazT
N+NJfJKiUEoeMFokHCdCK5/UO1hSM08F0vDXeUaZJ1f8T9G7c7Cg5atdK2djA07XDl4poAPYnHg1
pXeY1ZzxfA2eBJDFPzIJx7WCNJIydba8N4n0un3pFF8Q0+oyPkWOneCqDAkJpLBUiIx9XuZq5vvL
6vL9fvCDbUxzfnP1drxpG/TlDTffRwLiC8AG1I1VitRa4xRR/3um1CeBonPr4k/UO2d3Frd4x0dl
FtFlYG9vpjX6LD/7NIGrqnk4nXClOOblXwXA+wmdZtKQkIMTA017HdH7i5tjOmYMbRBaOFqlIzAz
QCdFKd6mw3ggsRaKjkl1JQV6H1eXCcTBGDbO2WSNl35HHigCwPK0KDmVGdh2JccfSwmPzJBR2S6Q
ApQQ1LBNqZ6OBXCM8JK3Q9IawHbP8YRn//WDbN5jai5brjTOOwGJ9EnHb0O/9AlBl2F2Z3A/OyIl
pOGqh76Sd89+Ku1JAHlOywkgGGwdPJr+QKT3mDLnKlRohvNsKSF88cZYLOXwK2qzlGrX5/azhNFm
Xtt2qdqVhAAN3WVhk+SVLLd7cFbf4BayM8/7zz34A/l4U/262I6K5SWMVijp3Zp2xPH1SnqaxcJ2
GKq0RtUfWI3j5W10eT8B8TY6eYW4Vp5LR+RITbQ11LHxtvsGFMz/+WBCwbX1+1eRN+bKYxDn+6so
YIPWGFAV5YfdQc74OKBfWPNy/l62nry8ZMjyzaPjbt7+ieBl538hjbjxYq1OIQaeeFr65ASqDfz6
A7d+jZoNGd+PYEP5kGcSRl1DmOjfibb71KFBM5qkDuLnu6tVC1CDQHMw11ZHf+g5ViPCjWkBL4sK
7qi8wRaa61xCOsYH5sIZbtBg4y3zAhXZrlgwHkZ+ZD3WbP+QdyUZHsWbrc+oiwIGCI9sHObuUZS+
J6Bz0IJl6+KKBxoz1SiRQGGqiyhbe5wif7D/YYkzcwVA6pc7KLvOsrsVnY+8sUac/Wl5OGktqdr0
v9aZYXQDBn5FcsPUJnsgMMNoBZ2D8rohV8JfxIyS0stTlBwre84Whtm/yYlgR0NaCwmEh/8JVS68
QY6vGlnvgJi4ceMAML3NI1iB2r4mrL2mR69FyxSMZvWFQX+hkBCM+I6E30c//rDqYpbmPwMY99HO
4D6BJ3jND8HHC0icM7m46JmRGbG6+VS4hpWPA4ZZdc3wxX3kSKL7/1F3gRlQlCfRE6Xw3Tzrrja1
21Ai6FaAovM8RPMnuZSJmS2rBSIZzZcDqTlkONKP3mR9W1trr6n4+dceZBeaCEf/RFpRyiI/t6lY
1mLHwl6jokA7mi652E4K15kU3+Z1MyVnDEQYv87/oZYRPBWMJCxkE0y/gEyalJNdzGx5cWds234C
A97seksxpW5Y/oL+35YVCVZNW7I98EjloUXOlCgukKU8wwYYxTaJ9wHb0Ffu+ZmRPZhSVria2ZGJ
hH7BNkf0jqwNqcJJm5V6groUWNrU6aNiBNXY4xa9L/l3/z7pfH41RZ9uX83r0juReEWJ9XTHV6oW
H1nt6iFoa3NoRdvmV3bmK8e/X2uv+4egGg9EoQc/FmAi0lH5f0+KkWi5UU19CEdF/GvmE9hUI7Qk
/Z5gXbwW1Aw4QL751IGZaeWXx/JaTNqyANJcVKrtUJkcoT/fSsVAy8kZronqqpMV/DfLu6CqEH8R
HgpIrkXyR6eaiFRFjVhzj8webZawbHIEf//NlpIdsOoRwf30pJDfOsTpxZrFDtOwMSmzrhhqFjzQ
lKLIBt5b2iCfxJsAOf2h6CED2hVZIMgPjFGrIUR8pGZiSRVcBmMG0QXl3JTCbeh3T0rdx55cFjOE
NoGq+mkUm1HBp8ZWWV7YEl2aIjCH88kZ483QB6bbWffZnMs6Dxctp/ZTTYCc0WO6yMV8KWitPOz0
mKSINZL+onjKPrgtiNk7pYXXgGfy+iU9bJilhn2XrX8C7zKP5j9a+hEEHhf2hAQF3+oxKjgcmLvN
0GWMAzjdmMIZI+LTB3kTC85sGF8liUOLdnd+DhT8Pv9E2c+KSFxsFb5epiKUGiZu6Xk+xS1XR1Mk
nfLyFk50vizTm0ZrNPFAxePToLaAw6Mm8Kvkcf411QJL5RgNTkvJ7YfQinoM43SXHbn90a8We3G6
YnO7nseOE8YFgldlGwrg/YqpExZytxGGtvlIoSZx2dDim5DqBNv/Z3aCQKqcchLD6WfMnivjRQPT
cTdrCjM2JqBWibJEnkzipCXty7OcxmSfgywEFZcEwhHZFdMAXCydkSZ2lxk0KtS/U0uvvlUE9mpr
ZuvgwCllY+GCBl9LxnEijGfVvq9B7TNfxdYWHVBhUNWsxQaws1TZyBIc/y1Ut0bUhGc/00HDkHNP
+u+klMx4tzfuhLzTQp+cJibRE/75rnfmMZEprzDojQ7lMexBItgBKqkX+BQVRGVo0aqgev+3QLTd
h4HVtoTHbFjXojlsLY0YndEWrZcgu9bXL42QA327uB/UjCC2aJecK+P4ke9WxLp5S5Zui+HUrgEj
noeSsjoTjA8urHnzxoFM4JRuevfTK0YVAf9cd+VS4S7xMMcKXE2xrZphbeN6E4JsGFAlnKkrr8c0
36QGiomn7aAnoPWfz7pFEqVu11oH7Y99xsDMZRnWxJfNyC+U8vqZg2fg8lfmzpz2JgW0jQxXVApo
9IlKVA9L9Rxsob+cafPZXhPx55VICS7XJckA5rPUvrz/vlyYHzCEnYWceOEGWPg3uQJrVFB8N1K2
ymGkCZRjkE75PzbzmZLMpjzMXy4qeAp9Z91d5wv01qtjYEyWsAWxEbjnkjPTOiskmkVAk9JKHZd/
qurYWSIGBYv0QiEpFNk2mw3lK/NIUkUxoM41BtMccQ6flZ38eMfodJjaY3V3rUEY338xyABjjp9h
ZdXz1fbgStxJXQgzTI07AB7j8HCUvmZuMLg6ST2Wg6HNor1Fk7dpPCj9EgwcCZZsawy2NZ5JJZEA
oJZNgKICcMpa8aEs6Ph6lWmAQsbWKQ4TgiSEv4zd1FmaIHZ2o3LMyNlenXi8lYDEMolyD3Z5LYn+
mTUjZdn8ZAZgrh6UiUMnqiESZydJgyLqh25b+/jPN76CTUyDN7FC//kOYR4j9YqW75vsaM3bxztk
8K5zboJirYKKB4WLp0Aj3fhqa9cD9QUSRCn/sT4IW0NX3Mj5CRi6KFiQ6PIat+sjkdwm0AUznlOD
BjYBBxX1NNNYQjl18KoYh/FKnNUnU68h7HuV0YuePonAXxs6APxotMf+cbY8EEdFpeA07a0ZD0NN
Fa2LK9SzUD82dzvgMhKmxovgHwZB6E41BHtlG1kjUl3ZnPXUdNi0/i7Bpqqos0O/WjhZn0snHTlV
Hv7NiYluZ3goFLPtiWYxb+RcIAeHnB+80jq9S6VKYlpSdTkP97Y+fVjmKezMA/pOiRjI767x0sJt
Ru4Sq484KL5/IjLJcTrv3TqkZaGkogKoqghK7UwshX+bZv0rUfds9pic4Slof1ztnyunzPIK4GEm
d06m6+kOBe0izJJUjwPNktyghQkxSUwxXddeEHh45j/6DIy6tmEKiToR2loQs773ZeDem7RWSfFH
Pt3S6NWS09uDM3+s33/55JfIsaD31YLR/J7Iq0bJKJ35cV0T4kztGiErXlrV8JaYSfrlNAzzLPI2
2IiTOMIuMauci8L+rTx7YQ9VSvEKuURblpd6NJLRRaENhH0HU/E45HDUKvVluCw23XPu+Kt592/S
YImWXQ9zhVnHAnpcDVXutwhu3W8NN46HfJ//iMvvtd/Fh0ITml456WLT7jlaz0C6V74HdTabQPIO
aMwkdyYlb5rDrDD3heIg+7/RWI2kTEWFc8fBnVWdjV32vZjE5iykhNDvWPqtYpYpco0bXtK5/vcX
x3EWKWwdnZzPtkZLjIWApn2Iu0I3qfpQ+noBx1bzxEbfxWP7iU3w92ATcKqsMcoaCsFZnoqWsm4q
M6rZbJ1qg7jIjModPu76Wh6A4HTtAONKR1NYpDOQTyAuBb3D38Fk0zmBcd+IJ81z3hEHmexqKCle
myIE1TFKIQSoZ64qOXn5QnXkwn79B8dmZqKhVdoP3CsCE2MOj9uRW9edeHyZnTXRumiY4RAPvGXF
cV0tWwMCSCKbcmYG1DGlyFlHozNnT5/uPUyqY8CCcV21ycfMdqfBAcSxhPgS+zA0c8jhWLHAoUZ9
B9R0Kv70BVXMywdWVzHFVQ2inK+qMDTVaTa95QRK4pKupEa+UasQw+mNYbKLkS3UyUm30GTzIMvP
f8jv39M9J8ygTtTb/6ewMN+w/vDY0vEeOFEOTt4QSZAb5HPE1QzQouZ5PJyGauJhf8IcO3u1GBZ+
f/2x3R6ilV1ZWpPmG2Cl0eVgZrTPT1wtbFB8bfLn0rkUfFlvKAKW6w0VcUHrRruDuFKdJ9yoKJWA
v3nlwearxzh/AWqIlK8q45ZV+qxGuFPKbKFw6MtsHBj1Y7ISVjh1wPpQPxlLA5kz8B6MuYnwFIpi
eOgY142RTxz54ScxLB9k6JxR7M4iIJte2byU0bF12GM4jYwk+o/8sjIvBdASAykG9JdFEovKZGA+
sg1HLCzqvzwRJyqde8OI6tm/VazWEyRHSikDTSjD7DS+CJuq6alpHxRr1ayCcTPyEybCTqd6inrt
imLruuCQLindC7km0LkX5zTASCF6j5nsNA8+PxehuoaA0lD3fSUOGtjVvXsA+wcB8+jNEJnD6a64
ASIPMQriCqJ8XQYedpWLcoQnBDqSZHmZ9leH+Mja+zMOTm6qVHi6IpodLFgub0cLXkOsEPojs6Pl
6FnCHz5MDkiSoMXfRp0/n0m3hOi9WqCmui2/IZmjsg/mbu+FMtZA4txMXilktqW+fa0NjBWpxtcv
7bFPGqX8Rkg3I4TYWCbiTOb76pqMTJf1MfNdudo3n57xNXiaVPTAN3hnc4VFMAV4nGwF21InXwr7
hg0x5go9hVQI1FrGlEVdWF2EQDiZvzN+dy68LAhsLdfupLPWfQElRPEbirOOrPZgpSIooD6GLofL
cyJanDf0yk4lO40ol6I11pYg1VvoJdQAU8PIDL6DNQkFryC3o/1K2BHftEbr7f6eerXq66LDyoDF
KqY2V3yN1n3bULROQJdo24P+HnSWkRLapIKkCYwvObXNTV79HfV3GVKZ7twAapiQDbZjJP/rTE+q
msg66eAwkEc3HVr9nqX0pe2Cb07+673AQxNCRxbqxMcpeJkaJrTBbrD0DVtynY3JEGj6970plpqr
/5eXppU6cA/Rw7cxHeJNhYNSh7gze908UkcswA/j6oxwBVWyBoA51M+fB80Ssdo3z9Cjf4x9KCIc
hnOgqiwuj9d9FVHfF2aVyjXjD6ksEmiavH9mvVLXFPuo/txu26TqEsJ7zjJRgIFnCehNBrqfL7z0
GC6Iusq8ZkwJB3yDmFvlxIBsKRQDsxV/BWuqwKIyOKwHHavunJ5V/TeapMXbvzmJM1DX7QyaEBEO
OACwJHZ0lERdQPk8sn/0btmegXPspIu/D0+ub9SP9GBEO4QZM5rLbLVldWU6nXyT+nJVyNAEnOfq
oui9CEOr2ViTCLoU31Mo1zaSksSbTBI3rqoepOTl/Iz3aSeBbiU3J/H12j8KtbEzEOezzYvcfJio
HHd/UEnlae1uW4Bh4KWME6bdzpU0R1GJPUzWouMIxyexk3UijVcbVQEtyJi3LxJy39TFTl9hc37f
fwYw6Eqlzs/6xhu37Li1idblwapE6PDCBCOJU61775jNm6TjJ0Mkb7Z0MvYxyt9rxpB4lhfUTrdG
Xa9caEttAbGkPtTslTy6ctZViDEZlHt8PcuLjlAZQ/f8Oftb4VanU4gsZUZnblddxYIkzP1CU3Er
T3zUbSQDG05bmrTWLVGRfEwhtW2j5E1aWoUBfI9zJ5dxVRay3qsdIcFD3c6u95LUFhQxKsUmbr/K
nZiLdSoUoFRk6DiBZoVboDu9D48cZn85qOdSPf5bg3ntSyF6rTpSobH+RFgZBtBJOXMYlwdoE4Sh
JNulodr3tCFr7Fi9lrGJILdDf6JlMyGHsIjh5851UdncH+1kMjao4uJM6dj2D78+aencMEZdJ3Ge
Wfu/6T/ecB+8VNuZ3NE1MkByA0aqBSpDfhgPaJ+alwFc6z1paUNA+kiSXAQjkPQbVbStnRbh/uAe
YOt5sIQiE9F7PfROniFBAST1pFO3mcafvGfEFXt+42LrSmbfaV/70lYnwu7eC/YsFQ/Yj8ZHEwtG
HQMyXnO+LdF/vsGTQpZzjCobOFEMqmCX0Ms804J0OdLcsOrnf2h+v5djisMZ9MIfsrMw2V75BPAx
2Lmnte8x/Sae6ztZsCM4GrTPU5WqhU3OlFIWu0xQn7QvMVMC2Kkd/v1kn7ys2mwRtnbd5wIQ0Z/F
MNeauZJg0N+NZWsWW6og4JjpATqjQOCT0XBQWR2wEflawfUr82gGb/bxPLXZfjCppy+SjQHW+sfJ
Szy08LGLVPSRMPEkdQksBdaT7b0aygo8EPnhzFbkKRseHUFy64i3if4Tybs5n7qLQd0Jf03VHU62
KQ+/YFBbxjGb8PtWPGuwONpC2h9PMKeAVVGwtnhRA6yDJoPgu4dglxRG3n8x47gF+zp3bb/ukTG1
hoJ0wDaWjQpWzQRowsbrxsDDcGNCQe36Eq55fVxftXXAhjn35FBhf66fYIjdIQSmX5LXYvuWMfWh
KsHi1NSrAwDrKufyfoS0B7YiCELcM5+/lxnXvUZULQEs0/UvYggH+QQxKH36EGziJs6I+mr21mgf
cI0cmAhO8RB1EQyXNxqqGmF7OZtRyRuaFH6mbnE5BfAjW2qIdlkF5d5+6XEhR+9e1aKUtGiEjo04
BeWJrkDglVvgEi2aYTfCsWpyDqJGRDLOtB3D7jQ9hZ7QHHzXWt3tJjZgGXPs2p6hObgutM+bxjrQ
ekoYeuR1Rne+AwaKUApG8x2X17H4sTgsVr1PVJrzRvrxgUpqtf7xh6ZKck5UJXCycN+OmAPtiWJu
CmJvH2rVcEtr3msGnjMM1TYo3SvDZZRFzuXdIvVfKYijUtkGWVhEl59ZxIQy+jwzA6rgDdI5yyq/
ryNk0MwKjYsHPIyVwHSKoGYIm9HGjpUaP6YW76YUzqygEi9JQYuNRdZKKSp9hFroH6VF8pKUFuX5
vW7bDCYY141G5OVWNvG9ZmxfoPreNKke51eiCpL+MFwZSbA7ycgQY67yE0wI6IcUgXOSS4q+8Jhd
6eDtFuXpKMOWvDqMXWgLvJhxFqXhIrBfbbu39q4ogRzyNN4EsqXqzpXY7jslL+2b37+e2x7G49LE
BmNMKOuobKl8VW1rUHdvKd2MLwcJD5//5/FRJclTnjEuD6h4f304ll2ZyJknYjSocaBW3qPNXZlQ
oDjBjJ+TftqpyBYf8Tzn1ZNRxjkpNQgDIBQwoTKSZ93BU6byZhPdR2/ypap17v5z35R4UnuVtHre
TtShIBe2SDwfL3IuW0n1bKKnzgJ8VAaUmYGYDiXLloy0M8nKF9mY3EwvobBy9wuWLSoPEyV13raA
JNRB2mBGAFWie0fCCyv5jqIeiVr3lvm0IN9VPXFOjfXcN8AIkTWEzKh5R9gFFwnBe4WmsvPAptSq
4Yj2CJctr3VPvOfgql8pLcneh4U8no9KzVdrEFyCT1f5CSr81jjqjsUQ8e/bfpYgl6XfKF5vksSF
nWIWK4zL3yupLRiuRT+NSVhRKKaOWxOUYoyoL9lPglSd3E3smfaU5NXIKgMzuk7FmutcAfk1lcdh
7Mv0zZnqyxZTvL3nzyE5Ifho9wSRYJR6ca3FNVQFBRlVvjvrl8P7JB+bi16I/Ai3TD86DbWo7VwY
dEDjjcdnYv5W5ElcVhC8AXtkTpVBUNABMzN8MvqjqOanZgVh4oy7aDiKPXWhbcTunVuwo5dk0Dab
n82blaZvYPnXMKiVKE+jbsMgiqVnOhqf9vXf1QvrIu/XBNtCYVyz3+KMEw74zxfBasm9N3bjOM4w
S0nXCnzkKlfl5pLQ145kZ7HH1b/bA+pTDuTrsezjdd3wNgjP1yk/HrQiUcabMBihtQvm4LgMDLLN
qiRsYKE8j3+JG4Ap8EhDg3aY5Ux8oUUF4Ca0GlVkpfw+XiSbOQ+wrCKgoggcfLuhmMoNlkomVpgy
WSrcCdhe4txY5e5JA19TOyxbUt+cVarOUf9gY4GqRVvlgKEndn4I9kNT12jwaN4JIsvQglrAhR/3
+K/wiI7dNLCpBAz7hRmyfYkRDz4sMNSOjmE5Ynt6RLp02cUtYObGHOzpDwmykZfxTrnoA6cqFvU9
6t0d4g5sT5Qm23UFhxO62V7YEZsecpNsK0ASHj5VBjZ9KMeu39cxPqT1YrtETw1vZw6vBFUlSX/m
kpbeZ5BDcY0Sh9ICczj9cKoV4trr0xIHFftn665MPR7914b+x/0wQayZ9xB8twFoL2VOHRN9FWpv
oEk7m/UKYJCQ//nXDQ9PLygXP8WqsGNGPntjs42W5XWukqqX7ux/9UPFIs4NAFScgawZ9WusOxqR
OBP0shoqoiWAFAuTAKJ+nWDnRQAhB+X3rRUOvmP5N/bBldLYpFHe7A8XPYdE+3R9Xp4+tS0mHGBj
iQJQkeT3Az0jPzvsQ4D0MbZksnGZk1CfL3PuM1cXuPencrKNNfWPff3rSzyXhVAoFB5bN0ANMca/
EbMGrv1B044bLjm4KklcCapHBDOZGEOLJ4jQg/hyjMDkDB/aky3D+5QMLwavoDQ5lNkbDEb4PfZ7
HN+iixIHiVa/GcDQb4T8e3qu0bv9VCn7p2ASFvlNa/UKDHjSTM9B9T8CXiP9d696VLCZiMyxADFY
iov9dIXbENbYWD7bzK1b0tAVeEEKB6uxDbK1XZSNr71XFIipixEQs9EBW/Uh25O9S2Ceucnwj3vl
yBxMKYhBmICjo70RIHltDcLhjo7hFRbVIJ7uFaCVaFsfbEFjEPtIbkD5WpnIW2OzvC2OSF7nBehZ
lDtmS42gqsZvNIdB+Sgbg2ddyI0f8YObzxCTns2Ge3mdgi+qci0leto7nvpUC4NTYKLGvQjM5sAs
pQc06tea/zY+Vrk54dWbbaZ3OMPZZ1rMlMUcImM/v790jYAOOmFlMmGKl66Ub0LbYT8Bi2arXbEZ
q80dGHhuREDkHf6RwYw0HDtObvAuAPAHePHZHVOkVCMd+HlpKnX1RxPj1OT/zS054J1DAhhJzFG/
vqoGJ+Zr802SKnvTQUtOU9jFWEyqfrdGJvb4S8BF+mMSsJ51BBJARurEPXHbXXIO/ibEjpOHyawf
Bf9V+5RrQIFL5VsANbSxaOlcdVNG6xppkJAnMXwXikSOVVCb2GWz2hzKezsy230dVmaqke/zUkzF
EIDZSotDAnEib2v8Moq3ElQpADQYSZWmV73KMGx06vlg0vHnjLdN01TkJDzAc/ImTbThVpV8mlW4
fBleEMjHLtqQaZA2lX+KdUyPSEWE9RfhDp05s2FPXfk7k77LGGl9kvtWYd6xySI/y4w0P5OIhRNl
0C2EA48CgLQWDzLU1iG+V9iDGd4LCGvwe/bksZLIxrwUByakcaXjnvZk70cCnSTsMqgG9WVY0h5K
bw/Yoeq1vOULOLdQNOuc9/cx7flMoroolLUVHW9wKfmd91R0fZUUx1sX36atyAz0E5qmRI4CFxy7
GcTLb+z3Rtqgkaan+JNXxvq8a9VoVkCtHlFw4CnY4miTjmQ5/MDPIkKYK7CKW5PBM0HUWCOKfjIw
gBCzFO6otND8vUrXuDk1B8blPq9HBf4iu4pdSv9HGRY8aO0d8Bb9xJVed8tOG7ROSWoQxdKTqqyn
jivozFQ0vFxzLyqFKeJwo2oHFgUXcgouESOwS0zYJWtXHpAEo8CGfjweNllfoxL+Wji+o72IUVnW
HovDKQs7Ms0tjIfcwkrQlh0TjGeWHsCV12oXZl1veIa/6mwFYKKOK07nYfyHgpFAvd8+UsuMysAL
aKDzyAjJwrpLJbHzvhivnDpHtyEyat8+0B6KshPx/UleCIjRriXpz7wIbYg+Jkajwvr6IrAA5k09
i3dc0U8kD4CxT4Gz4PtbFsZLMslW5Pv4+PiZWvBOCpvivaFIJcZTn7fbSEHxxPJMGhBCiTSDqcOO
ZW16JmQPMicKycR+7Cz6sMhDSdDmWUx0KCHOov0rUMWq6dWCpQiX967LZDx1YaKMMi7ADVG3lQw6
bMfloOK6Y1+oed2qDI4GLLLNFyhGOwaC8+zt/gd+vdROTjqKa9FICZLrwXfQmQDYC4I8SNpic52O
oOOmQXyAJe5RBngtVb90Nx4a/PzVCfYNUJQGUoF4mg32g1TOj5lrA2at/Ud2MTDKgqIe//NGBC3g
FLjAAimwMKfsNd8OwpH40hWg3dCqvz6T1NZwxdEwYO+swd4JjNnBbeWea4HJix64ciCBXbhumoXC
HbrvgN0/sZW5/DLEl3/M3b96JJLqQJ6+pxF4SvOGev+z4YB1pZWALj4ioVezrgnYJI490GJ5PCwK
XGE8oqQysYWjLyhzCvFGrwyK0Ejb8u+0LbXzcg4XBb9PlT2UClTfA7uf2WCl0K0H2YH996bZwXby
RN8VEiivhOWlsdFUbw547roTNyUUa6qBJYmfKhwmiMQ2Jk7kFMQ0HOgKwLXqy6/eeqL7A5pwKKwD
GWWiNcrN0RT74V6BSFH6U3++othc5xTQXw/9dq1RsZKoXclAdDfcokpNs0JUHDRTmT0L0vAmqzWG
dLbLYC+5LozDQ7krG3xDscSRjKJqRvc3H/OY66qSLkVizAklyKbtXZj7JVYMJfJmXsX8bkSH45YY
FqV310jaA8yj4dMZVDAnhUCquULKH5hXxxiCrcrnEoMVEKQxGGwEIzKKKrXqFMYZkN8bpSXGz+Qa
5p/4cL1LAJ37/lo2ofueUhSQP7oqOuwLLNE8sLZeMwac74JN91hMaLB7Iv9ZT+XcXRu0oNecoW6y
2wxmLfXN2xGk6wZpqWfGsY8kmwN+sd06Z9Y99Z1XADsLW6tbSiopxc0mifMF4Llga+qX8JtYOAUO
4YVjrjTu/nyZYN9Og5yE8O9CR+wHi5TQTizW5vaNNCZemVEbII5II9LJoYR6/yQvpaOs+W+uKWy0
tIY2u6+KG5LwQEBMSYrBk5EB17NZ/wcGcB/1r+fW/34os+Uh2tFlXLYl0enq3MqPGDNEumgIntNH
gFFncK0Al6Q3qygpXU1mL2XopJs3WU7VsnEgD2oGNwyKjWqQg+rxdGsjCL5pTQ6bHkdh+BJI7gPm
Ue65OjRdUBG5m/NJP2twRyMeyfNZ6rbIRLPV8FfuHoVRs/cJ6Ms4E0tMzdsWajLa2oXhRXgeCxt/
wEviVSfGEpFxpLsChp9YHAB4IF4tmTcvLVU2xPq7ANuDgIAl/vc/CEntP78ydJJWAqfOKn7lLpiH
2+PZ5BkCuy0Wn3NsjinpycD5TCFB7JP/6WjoTTwITsmeX+o1ZX+EQ5MorGhqkvQ4oX1DLMdyRPT5
mUtA1LyymYSd3tNQDD5fCQXPu02ODwK6pM3UwanV/6yhH4EOQhjuaaGHmA28iGmUFfpOMvE7QYeW
+KLQKzQIJ+tUKHXuapU1DRbckiM1sX6pcqqfoTSgAJ190uVVyZL2pwq+oTCdvOtHZKXrxIr+z0cX
foo7Ww5nwAtwAmg6yeOr0oi0cmZ100UC0dcSC03S+LfTr0HVmSUbkF1A1jlzcqnlRuNZG/4wflfI
mfJkiFI9Zsnu4P504NzSnQtr++9TpBJ7wdl5ahHAxORU+vtDKpNXczc8cNO2UbLttPpowBo7DYgf
xkf1lvER+A7NPKnK4N9CSV7BwxEZsecGoqgQiEApMZxiALScT4C3co4YhFA072hreozVVoV0sPJy
txAgL/Re4S3O/kraWzEem5WR0uiQjRV8BzmqW98kId+/1yEszCFkw1KxU+/ZgFxu1wNlWXIH6DHP
rXIlIwMHKubqdCCfSsf/1VrQuMD5mxlsySrxUlRizi+92TtSbhv94yowo2QlWiOmWEt9TIhvQwV8
zpDFDfY0GLWrZ9U5rCVMtrQChmlitYq8798ZwFDDmZnRfDIa9ZUd24Of404R1cJbosVo1agsHbSM
o6u1o2UsYGZqAdVV/pTmOgpXjTxEBJKuD+SMflYYoX4fNAJAAgkdrmfyvPNuYqFOc0GD7eBpw/HK
GLMPqf+CVgzmdplDVmIU3BlOm9rixAbhrbkOaRICIKOzhcLr7aw6gl8QwYKvpBm0jVUEOCMMAqob
PmtzkSnYVZu6TCPPukxjSYFO3E36rt525ddaqBkH9ocziLHsmRYVumRlP3kb0DhBm4EW8kCOZUfQ
a+nZ26MysIMc1wHrUwU3cf3/Q2AX+SFa+X/OrEbGeO9QP0mJHk6T/ZkN5TQtwGmAP3eqtFoy5ZxL
aeFVu7Z87WiHPP6UWtaGdbOU+PU8PRxhxtfJ5HOZNi9Gd6m8E9k609NoeKzvUVXWJxy3hGxQC2FU
RtJvSFPS7k5eISI45W+xLJ0X/O5yK72KjL4axlVvqqUs2E1kJwxyckxgl7M+NC85ZVWWPFoyBeCT
vwMIlv8NdPWBkfaHHFDj2SNzpYFElqHVyeANEBpe6s/sGd5+uYqBOVb9WG1aXQ3/FqGynbsLjDFT
+8a2so79FHqzgjctHucNiEiVZKR+u5OcvMtPnI1sRltIw8QgeJlt30fjfTpa+5AdOQKU4k9PYSk9
frGZJk2T/2dnBZi+ZnFs2lWw7uggNzc9x8AMNeuRN+HTmCm/WY86Yo8N0SNnwp2Xd3bVtWukZ464
hFBsZFhJpm2QJnmD3zPAHhzUSpiRl7VTgLTHYthB+udsO6oxWzUOFRQimqbECBXz2tRwZT6HdQPq
SVT++q2swjpFv3oW9YYda8ACieMYLtffFzAZVdA4J/Nd+rnfcPA5pTcuLiJi40cr+N4yd8SjrkYx
zGBgiJQBc+KKgDcy/L6ONwI23w1f4SpfiK0dWNPa8+5t/mhkU99kCFIFyCwYf7ksr2OEGuCb9JcH
H4h4QTT1ciTtljDbqQ7s0m/Xv3fpVysc8/IOfQPwd7KZGWt1ifbUUmv4FVWidiUYxjqZMCuzz0A1
jEyDSAa90JSmYOUQ9yGkWUbvR6/MV+89YU36lrgfSxfoOCvehdFEzKRkosuqBnGao/0d/GcfidC0
c74WD+srM4ZJBOSQ2S27GXOzxAZ3fdcHXLtnZoyaD/RxhIhzd8sQ8xgLeuyx++++iJil6bZGFeUo
/TvJvr8GlMS/XhgzTETuKlgvHb7P0Xq8SKu5wlf5lk/XUS09rD1Qu/KNJ6uRsDojz2oeffgwjR7N
paMQU21LjAYrxdPTAXqKi+9gxWergBOWpIbLz4CROTqGQwyRdwLznKqyNrQg/7Cxf0XfqFEE8YOI
SpRV9so18YzMjKthlj8oX4xzmEV6eghu0g9nj82VAgf13fXzcpXmPQ2pJKPuwOq2Gxiuw8cObGhd
PIsIfy2sncG69QBLfgoveSG8NX88jcpzqlhNoFpR5GYJl15irvzDrh1FGQ0aKlmsjYGg8/2W0+CP
LgZ1XWv1xl8iYIuT4IgNlqsDGfYFrHVmjbYvUFgtCjJWwWWrIbjyldgbIFV7XvH9gvjs1/XeDvS4
0m0BoTJTF5iYI6ciqeoYqNw55PSuEcTOLBhGPGSz9Mag6nVcRsKaDhqwssfULRdEQGlYY1UgP7T0
yphnY2VPivWCOzZPgZA6BRHtEhuiSefgaVfS0/Lxk0kBOs8HGcR7shzMwvNsGNYDMuDu7n/Gnusr
b7r1MDUdQqo1RfHcX3iC+o8qYDhVbPdinfR+e4iGqc+fvhQg02YqiOYL9XOKoZT2IDz6X2Vh48Qd
9kVD76j48EO6bM3UOtq/DneV9d/rrMT8Ajq90FTrDwhfJK4Hq9hvkDzkUAf55JUmSvh0w1e1WFuG
rPs/+2zGd+gIycjFpFxRTBYqfuWtesyZO9JbgTOvDko4NXrdwvxChegKptyo7viPLxCv7qncR2y2
MUKyr4irbvYBOL0uf1TnvBA9/z0YBHZvw6OG3QhTaVTARTHw7kB18/J9z0K4BrrKtNiR7kdrs+Em
1RbpvZvjk0LVOS33MRBHGkdYSNdKZ1354cUaqKWy4gN6+LEEzb9aQrAtKS3psIAzEim9n04H+Kdp
RouIHwvsIEU4eqoW2YkjGMs9pQL4J9E1ACL9ncoEmox/tYEvagqtRAOJg3/mnQoewJ/fjsh6L04L
lkHyY3TXGOSy7I7Hpei1FK5z90YNxmjN/fLbaMfIDCGA9lROUrLHZmqP726ISv4Qg/n0xlp9Aykl
/oDwb+QwM/y1R3T3PlWE0THBMVuosayg+V9ZD+qELj+oH6tHW8BaTw8TzuCCHMKqGMm+hAtiyJxp
CPHexZ940UMa/X9ppv4x+t0tWCwQ73zXYMWIB43M2WPa9IfUwRVuy7YGHGMaFXaNXXhSwWrUzKcN
g1B4WihYvReBP8HAguQT0FBRgSdcBTtqfQ2ZXXbF8JyFt6vCnnXxvxjJViIHqGWbNiM3HfccQWI6
ktIB8DRnwffNHecr/OPHXXzeIuzz+jgXs7S0XWcATumr3AjS0HcrJfhj+73ZjM+BtEdZfAOnIpAO
u99d7aMPvybHX6d1Mj54T1bOifz7maezfITHnHK6mtP/7fsOqKXgeeOSPzhsBsYO5lt9GC8WMNag
6eezJlwf9CrJgQ3j2L4GxTyEeSPw3Jh6R89bnoPYbiQkT3FvVjd4GQdBNelb+W3E7pEB88H+mEVg
JqiBA+UOasCC44dgFkz9plFOh/0oIxv324a2rTs005EcCd+MUCs5GBkPEJZJNBnvkAycTil7/YLc
NfF0EjerJl92lUvbB/IvSJ4NDfOY/RMOuV4bdjnCPKK1/qI4Dm02nhnfjKKffaOxWl18NQAvRkkQ
dfaS2RcYM2GtscgjpEJTeGPDioXHfh+FSXqwav2qoUb00ieJipUIBm/S++HKqithG+sE0GgzCII/
4bhXu7rPuFcN/PiQldehEtAj6DppXOXPCicR4X53Mduh5S5H6VeNfRjl1iMZTzutacfKN8FzcWEW
kKTFdwoX4aBIT/818rOS8Nno94hrMhipJX79x5pCv0fYgh8Xt1uzfPP/mylrbgPzKxi9u0eC42O5
gXAkloMPCm/B1CurbHN8Mo2oSyqpHjWAdsJIV3TvZIxRMtQ1RbmlR1nFOXg/PpuYc5SImvSwiT82
PJPtVvPi6y6OeoyKwwHld9zxvdqg3vj2fd/J7WfBrvBfoRAzd1vZ56v7/r7xSzNuTVaACHORZBT1
N3X6ZGemZOtCGFoWLlnkoqp/j7TU/jwPKajQtSHU/FNpjE/JCKn4vVKdFjd3CKXGuzRbW1zoS4oC
+CT+7gQPEELw1EX+hBDn1A46WsGSB5x49NnoLGP/45FluDEf31ifUKJ3RDC/v4IsO7KlVDID2Y9I
TFnvgFOpzqEzjLuoZPamLMwuLHNTIeZTIfNaE69Eg1fAijZW92ZXXxqOdHdhy4zVFvqSgJuzjOU0
g1qH7VoyIcB0TFlH12XYOBbP1NQ30TjDwinyyH11l3rTMuQh4GgCVj188s+jH7+I0gTfJnneAR5u
0Dj6dkjJkDiunLwe+71igsagemvWkCrZW44NPYT61RjE54wqwNTFbLCawYHnsfV5e/dEllwjjwT6
q4QDfxOC8e7JTQd3ie/pt5iHEyI/5UozGnXzaUq/yeY9wQ1zuBH2JSeyttmqtMMgMdLePJu9y6Yq
bHR+MKBLu+d2QHCNdQKlVfV/caHNBfsoyn+2krqD4w7HUYSmlEmf8/BUM3Hv4eeaGrJ/nr4lsq4D
wem/ugKnTqmMYlPUZfzVioFOS+X+ROZU0FcTwmWrxBep3OVFKf/K8C57nElR1AzhMdf4f0kOkp9/
nZTxA9eJ60nGNkWDsrgZhpwP1d9BZhCNz7EsrVB7w+pJggiCu9gH79L0X1K+wIlufXZDdSrGpFsS
TwQUiaZU1GKwJKT84kPVH18L+jK3JZqPLX8nHG9M5w9m37QFrx/d2OtokV29fSk7UbasEbKBvdtZ
tDsol5VO+Yuo2flxNbvqe8eyQ4zpM6My+jp3ePBVaVWEmUzkb24M/JphBDp3f5DeFhE4TtiNQ6w5
JKBoMlO/KOjahy19vyPuQY/QlU4VnvUChIXRM1SZaMUCKUCzt/7lZwXNBgV2EYqE2Cnxe12eO1v1
oOwzJ6HkbH5cufwg0fO4qS7qxlj0kAzrv7DGMsoKn3CAhrTjS2nQDZ7jsQc9AzeqivgrNcSB0VW1
zlAijVq+EACsgzDFw6TKtPuMOQtPu/I7/mKuBOcPhfrOj29evQNmPn0RCqjrmpJa9afTLnsJt54r
RsvyoDL0b2N8p1hcMqhYJYSCSySQ6yxgpo3n13ilE5ZU0NmVoi1a3aOoPkDv/h5tAxLOiusyGbfW
TKLzg3VNRj3P3XHnFNCFdR963/nCUkBzFTecTp9OLnC/aTgsagaO3To6ZOpHXz9hPtQpqIOp6E5n
mQjshWLKWc5U4hghM3G3ZsCWF3y2MKdbo+T8a2lqBknNDQ6vlaR2fQx9nqVkzORIaBQ/++k/lvDT
6as2gi7ky1W0xzLlrO0fE9Y1YTs0HQvYGxfStvLdbJ6TUWBA2qGR4ECliwrbd/tTErm/XZhpkfH8
khO50yBCetJxK4maSA8WQ9T3Kn1jhFyM1TbxhGQOCqfIEWBp+pJYAxAuX0xqEi6chl4miMBYnxAF
V4MiyKk0sR687i7Is6M+Bef1zqNGvm46RhGB4el4scAmEGHHUc7kWWLV3u+digfWqJOi6GiNE7WO
1+O9slmABAy1plAG03nb5BF/UStaEHBBNSjMnk1N/pk4UevizUOkZ5qgNMSRWmYsD5/NsNpKxEjf
x7mSb2rM2acb1fxh12aXCKv6OJ11C7f2uHHIuJpGCAvyDlkvh9Sj0JV7eHmCQ7fOm4V8p6FJv4k2
FMLt7Q0m3SPvE5IsV6lMHomZKlBDrICgJN5b2dYN2JoR7+nO/TtlswZ+9/go4DXuZCI/J/6nDFyd
8MqqQ/FDtHPSwEehvTbOO6pE9LznLIKeLBTYYk83E6swtHRc1WZ7i9mIfs0PMnY9itK1v6ILBjPp
W7TpcQimCwMKl3qk/pHod0tp9jWixq7Qs7LNCd+Xrk2pNuaWRz1UuLfaUyTzfHmr+ScCRFZEM8+K
txzNGW7VidhDv8E4YVrSBNkn2FNRx2jzGG3roIau2UfFfnPCXxgS0ZhBiiR/HdLkQi5O08eHlZCX
fY0aZmdQbZoivy4kr/i4d1LHPv3ong5/WawDOisofz4LxY5s795/lBEUsLhB4cXMuwV20PR+XDEG
hpyQ/V50y8n6peYDsqX1v4afABUbNvINOwNl5ZNVT3kAvWS3f3f6rBB0SH850ulwGSYP8Qp3gTz+
cEYDPqwLZPoqZr3ReqP6QsWUuUrDJxtDGYP7+Q+lbnC3rC/RtfieV/dqTYYp+nHMwOeHWLzXHIRR
W9BcuwNz1EqeIdFLvmloMWFqT88wqT/jKkJYcEtpP2r3jOC4uG3QTXXVCTPw4QGH83CGIBCPW6R9
gznxTVDk4xYMpVClNXxBi+fnlQYufMh3qktYj2H+lQR6dBchpxxyis2CXDUKpyJlRD187lH2kbm7
sh6jUgbQaVIQZcAabOBFS6y8/nIRbyy95JyStZx2gakB942AlvVm0BujnK4XW1rw3B+2ySF1slMI
8Ukz+UUboVgJtjBukBNUK42wjDAc1Aokm7NyK2GjeO562p8j1QEY4Eg32aylBpsch2MvGdnoieMq
neqG9e0VYdTaSeAhgFobUxdw/tzLGnPFbYJDCiNlrpIZ5b+zQ9aWgsYfqODueWtj+aJvchl5tycm
BrNvWBpWSL3SNq8lBsx1QN+wnKra97PA/J9sOR02kqHXdsqf/+591/CuhnJ3wg/pj4Q3lb8QEg25
ZBr6Pc3IUvUNrfHe6dzXAivlazKaBb7nLT8yJRArX1Q7LuJcWMlqKFYcChAcVmhXYCAgCBWFE7qk
xYjThVR2b9rRUNbT+zbMwZSqZ4TiRLoFY3Slp8+I9Im66wBnj5/Qid+WuIeDHZ2jtcG71sDOOxHA
eOFkMAEtw3IRsQQXLlHu7HBkQ4RH+oalbGmEuUhY1RzM1Jz1aVO3Y5jbTVHuuzlNZiZumZMEoy6u
SdlBRHCfK27+6R9Cm2w4fa9wXxOhWzHUdpLFZ8Casy81wZxi/aT4u0SlR5MgFZySxk9q+LbStNlI
VQPzHmvBbiN0pFYxa/HcN2zQsqFykMVpMpe21MOeErHcEyIkAT+psa4ec2dX7hy9VEY2yZ5Xyr/O
IPRYXGl/rGtvNl0GsGa2AvomPgxLwL3Tp8thQCOuc3oPwY+8SUaF45jXMj1LaaderW2KlAakNRQH
11uEyFKo7EKx09sxJ4okQnVYnfMZiGiIlwslRQBzklzSAMtG3q8RoDKVGBnWRTTFEyiGD+ugUVWz
0PSyWjJxwsOQXkMtbkWs4OsBRELNCF2Y6+6HzVzPkF8vEr1i1vjIgC2pPXzf8MeupzkSDIb7+p9i
11fcY85ryr6kt6WaMQsHvJp7u7T1SLrxQ/x6zXRbNQRGbCYDWMJyil1F+FEcZHPiHjy2EqOxJnOB
/RmSnP1JACXDSfl3svusHEE3cLDoAqdMYiYk/OdN5BG5XNh8e2lDP7LwmMiNZ9EDnWKs/jmr93HY
HHWJFOpy8tO4jYAaLlq85U+XnstDLf4TAXlGVMYkWmbh+qDA2BKbu/U2A3eJw0AwQrnpFb6u+IRN
3Bl9hBw8SAp+EInxxNv2nRYYzuYd2Pi4vLSiKo8NbYZ0trVAy7zGSPw/OCEZj1ujkZPFD33dkYlu
eWZ5n2QxOyFgbU5KwL+v+XXOTTvqvGPWJwm07RN6qPH9aRlFMN5O4WUk9LXLm0Q8O6HHtWWuWfpy
zoN88lKkXsVK0k7/AP5gmRjT/mNcHoPtOiNyBKFCGjKhbDnBzvWIM6w8ckJe/LtHe7nqyHagbOj1
xSK8Ik4UimcfRSAvtoG++5FisKJ0u2Ux7SkezsuHMFX+05sxQntFiK7xA7byqAVGzN7t5EzRxloq
jDwyD66m0A0RGYjRGNtXSr0OwbK/u3izgvQVlGofjJSuEBkFbb1+GtOIMAi8GIA5THfdyLeHokkk
wIQsm8pu6b1WxFXDK/UTwywut/giisziSuuaXbVugKz64zEs4Q3EhprMvzlF2mvDhMgbY6Zk+Xjb
OZf47+3PsVGtARcqxADbKpqKm6zuTv6ITZmJS0Vt1d7YBf0FD0OSGJ8+kOP8XPOBKBzGEhUZtPyY
HNKudPa0H62mJ4JyJ3AViMBOIR0SdAkyhad3OO5c93E1qXt5XczxZpPi3owJGq22dYNZ3xDVFpbW
0gv6Wy7VBRgGE941DgGX1ZCIscRpy3qdiS8Q9TaUviEVhgndmtYM96VfmF9DcZ+5ZjOAJrK9niwV
x+iGdlvn9tWyEYHmLL5ImCudKK2q8COk/F0z8WF2TkTyhOWg3uWAQK0w8lIJeLvlsNOV6lUoQGv3
9W6BiXplo4lLQ+Tm99cOevtamsLx4TgxTBt13oQozypPED5vUuwzo1EFX4Xpk19H+eNwh8zEJCf4
8rLg9mzhT/7911OM9o5OV3LRUPfw3K0tGQBqwfZIgEqIwPb7rfAgx1HrYPenQvaeIzBR74Zx+i2F
q0bBVHwrg9QVqZ+KA91ORoSF4EFN3mM5D6+ej6bujq9wqVemqrbN9LOj+1jIDqmLq0XwVo5b3IWy
XYwUSQUmFw/yPsgp2Z/YNnCioWWT+22ZNSXK+1cW1X9DRi7Bofmk/DW/KCfcdaNoP2GgqmOt3WO6
IKF/akJ1NxiuZjXbGymMrIsb6mXoty3ZCP1sIPsapu/hNAtRdCokY3ShzUPuT3YqssnD5nEqykO7
QNHlILryw0+vp9CPFaGs2EQ+ZYW+d53zSbNiyAMfDeqJycgX5jyUqI7+JW+rS9j+PcK7YxaJwoy3
HArIDsgzb0kv4EoAadKp1BNo3It5gJpOPd9GIbSIhNCiFX0mJ7zVjMOu3PoGceDoRS2QbfMxb8QC
rNvHt+OGr77A9mrDMIzm5gIANkF6hYe6KccbUN9IIH+UNHK1ZSOFBMJqvfyhTKLM/YN3jcBj7Fya
0NYP7Xv+akEiA6I7buVotEdPJ1IlTuk+ypdMmC5lkpb/3sp4y61IO3vCUycOkoIKLVLa+Wsqi1zW
j7qsJmV2MLVyWmigLiSpa1bGRFSQZelTXox90g4+d8FstEL+Y5Q02b42kloT0+Y7anOzoXijj3ci
ZlQTCGPq+VmigU+C+2KN07eoj2mU5MUXhl+JDV97NriqJ4I6E9YnuLdBLYRWuaWOKyyyDi+1NuXz
Dqgnm2QMvkcADWaLtOJAz7k/TfQpdkj7gFGYzZ3ry71eicdFCqQ3GKFQpcstW2GGHk17QaFt686J
QI7y+xRHDmVneQIb0bFDoYJawjEGYmwYbEln4/DW/O6H14PMkHeerwkGQoC2AtGweSDlmCpryrRB
Y2ZGN3/+c90Hs56GrbBDcwoIIU8043D2OF4SbJmkFP5kQkhKfuH8ijNSuvKg1Qeo3A+nIMfR00wf
H+HgsAn0ExYGSa33TZXvi8Mdae7oYdpg0zNSukg7U9zyvMMHj5XYTD4qKxY0oRMGdHs1jMyeLElR
/P342HTyhpa3fITYXI/EnWWsZCCQ3XdZfHeB+7p67EatbnhgCLeZFtpfgyZZNvJrr1JDuRGF8rOI
DuIK32pI9iMH8wsdFSsDgJFXjFvkW5uST2+mwbu5oQDOpxIn0EVX5NmxDXY6TcY52jGMDRSixSTg
MQcXvvTpq9x+wTWVPC5+ujz5nPLgExRZVEI0z9GesnJMm57NRcSvyBzZcH+5DIOS1r3j1rBfWRJs
CmSmc/IlHmt4Z1nP960D+HUnX0Rao+HtVeg13JkTZTEFi3kMS8CU+d+OqvyvTkOJ6pJyik61j0MU
4zYN0rEvO5IyJOLv4SweRHtmVrBYgKutoL1x2gX5kElK3WL9tQamNKx6u06ZocARoSJRDffAMncj
L/FCc7Q0vGrGXYryohDapR780ORMLrnr3XmZ6hnCY9kbiqMLzdcDdYOVx1pxTIU8+4wtNcs0RnD7
Yp8LbjNOUURUVzTJz+71xFLfEIEzV8neIBRzsl8ezvVRj/6PGwewlsBFFHq+F41venZx9OI8n3xu
sFFRduqYacYa3tshF/ZLDmcxzAMVHKhod7XkOjo1BGOu2Cq0gP7L3vhQcBIRV7H88wdUvl7NJRv8
aXx8ryloAPAuf0rsPP/7UVcYnmdCT4aSE8jHJN11Qyztalo7kkW4cRHEEBgciegSD5zn9pn8iyQ4
uS5dDOXVCny2vWKIMS7U0i6Z7iU1t0lwt8aa78dk2KRXInlo2SEapx/atcTSEbzAu0pQNr/wIMDP
gxZaBh0XeYsXQWoVi10sxcoKD1f6PvhqRaSPpYoFIRnDNPGsOwjLm/XBpvJ9rp9LrHjaY46qildD
+9CVBpwtw7VbCLrFoGal5owmRgd5VejOI9kKwFiZiBQ9oNz7nvSsscHhauT4bP4DN2i5iyLJ9Anv
5G74MMTM9pXdnaT/1oGoyNY+jJGg94D+S2yApIZYIRVZ9xQmSaLARxMsp7pG6Eok1e1b1Ye73Vjy
04dgt4jSlvjrn35/1R1/GaWlKBVm5UQ1tMUarkps/tWqk8DO8Id9zxjYVwxeaB+matIUHhqvq/nm
qqMWjDBUHcSBM1xmQOK0vgm1vciffmmLiSIEN414UtvD59FBqWz+3rAtHCBd6a82stj7Sb49ohZz
NxMu0JNkqOv5Sa+CLgoYI+/i/F6BEBeNMEJlALhgVnstHAecrUKYuBdF8yJ7hgPvY++3KKz6Vz+v
CX7sOhOaJai1Bx77/FcfiVX5uVg/HT2ixqwVGCX6l6OcXKuFkJEC0gQfV4Ngt+Q7d/X/G/wUPNo8
mkJXRuCXrYnQGdv4J/HHAWIPOamMuoBOYm5DSHh76rg80Zg/FkIs1h2eoGy7+bFUKv5dSWVvJSWL
NPO3xKKd8Lcq0v43mliv8gQsLaXErOoP13qZIX4hRem4wKmmLTbf3wwBrhRujIPq43UWr8w0e4bu
UszI3CgURzoN365YT2m2lma6DFy1c7Aw6yScGonaVpe1gxDLVty3yhxS6yF1vPYDa6rrRI4Lnsb/
azdOLcx4CB9Yc69j+28CnWiroyAFBVt7tiKlxsk/saJ2Wr97C3ZhqlSSLiGdRzXCzoyjAWzvQGb2
fLuNQVMfaPoulNBWWlbeKIWFKgl53f6a6gV+3flgohwDEjGTfpSydc0/43JeHxgNU5HgewXg21Hg
3h5ogw74Hgl1heufX4NoAiXOoXZVq3kACDyGmaadIfj55msmlwyO9LdZSUKHZyxmLCWsydYZqSCv
dx57lggyNSzeu7ZSOU97kZL6KT/q2YGr0KD/wztycpZef4GvW9YI15tAuclJL+R5jqPlDfb5ztLE
inOguxMeV3e+A5KKkFymJUz0MGKeGtEFKGNk7/IcmQwVUedhLjbhO3dXTKvBH2GgxJpmJduCQXN2
Oqb5qYvNUPYuqZj4dqfckukQZp2jPb5wDswcZYMEb+BvOgfBSeOSn2DKN7BS1D+m0izHAHKLA/8q
r8RfNUg4L+bN3wLWhaYpVVZeLVpoZv4dk820Ct6pjFo+3ep6E7dr1ZkTVBw2HBqXIYBhAQdqGDT2
LwHil7r9tySj04f28875KyBcTzFSeVC/iQuNdA6+uqqtlm1Oarc1cFNlL7+DTjsND4oJx7rHBUqm
kWTohzpRZMbSCPRnC5NSsJ4iaCMnOuZa2ZJCs4SdC5batqPILbn/Y2dllIU+M66o5Ikab8o3MSgR
1xYSAkEkL4JniZtJlC/GZT1r+nllWRePt4CqQqINZz4QiZRSXzX5qLlivM7Ms5V5F5oUll3peboZ
1xKBHFJewf+OP++hAqWydxoK/DaKCMfMjByPSP1gBCfxTQKq0VabVdioEgBnUfOyNiMHOmXOgJIT
JTfMFVy971ReY2oVb04PKPzbe6AT9mPntaj73PUpiL8+GOJA6vGZynEMJrCKG77vRFi47XWFwRyI
zJk3KmmlbbyvSZ452s8Ylbr0QjUgHqiRP8MSIfLyfuBEuPsWlK5CBgwgHlycKDKzGjeQEN2eS6nm
F3ruVBC6q73FcHA/7+rqxrmMKnazDiDL87U0X62tSg0DstCJd5QsbG4dmWaJcQ2Bt4rQ8P6J+vuv
Yrs0oJVPan7+nwMVtxBqvaDVt17PZzlEej73BVifxbNACG0Hc2EnYyt9meO6Yfmn+Fyc1rMQGHDI
Pc7EI9TV4nJFzWLhQj3RmLqqB0ePVZQxkuZ1D/mHkfNzws3PD3zbsz7ofMwOPLwmhv3+IMrPG7nd
ScF0r1bIrxq4u5IZ5YHnZ+1paBstU74sVNZoPfImS7h+U72oCx3RhVW9R1GTz9ndTNcVoG8COFw4
fNxy4uFpSSaPujDYuNE2rZFGyuY4VWFcncz2COL/j9L97N5WgvTsp2xD3FCG+mrazzt/v3wRFWlx
xzh3hxVJBkPUI/VbqRHnqf+DsmN8+WhMb3JIHaQ6zdSbH6b4pfrzEgu6+lWRdg6t3DMtj7mt+Lme
YHOGcHw8dY5bmJyqIWLqkXHEy/BzaFBlGx05f9ngD4Q1lzNQVSMauWb91SYwiq+vS8YGsDf+8+Ai
IGmDaM1BEof81AvrrJi5/uIDpPdaihzLVyyNq5z6bq3XGK+faEAoai0uQuIRq4Ti/WW4oNMhbkEc
t0n9SP3Ur7tFS99IErebAfgi/gqsikEy2/i6fCOBo7kNogVcYyKN70JwnlUMu0Lofk1NVV4SKd6P
muBY6p3cOscTNRI11Xwgw7w3cJfNwdjQDeP/4FkSFz87lrCNxtbBh2OmNwqkrIbx63xymLRtxwuv
nroa7a0ZMqDDSGnWU0OUk43rb4URZ5RHONMtjQINpuLJnKP3kKnYPCEiXf8rzD//KWO4XOaSveWY
su4Ai5RUewCwXO3H+lQ0sFpgSR1Jc7Zaknmqora7ZX6LbLgbFJP2BWM8i0BiDkmE+xAAoU/UFG+9
Odm06sIK3AM1oug6os4b3UbQM9wIODlogpX5sj6ltYgCt4B2qdp9XgFIl2yMXqZqOXGdRcYqd2Jy
9wJBJ2hrOqT/rMYcGd8i57PtH5juslbyObALTJ8wHWjMykBP0y5v1SZdCVm1NkQgWXO7TPsY277b
FY0QrwUjznlb7qciMD/Q2juAcjIs3RXftUcAQfBj0tHyTG9NBxU7qtv7ttb5MmNU18/fjgcBCyBj
FQdo3m2TAG1O7b2QcBcIAZQuQu+vRAF/7BpCrGkBg2kyoyl8Itx1BKD7lrjl15yt+B4n1Kp7mh5G
f3cp6n26xB+DWAInE3zBbagjxfZKPoO9OyIJ27vIFVdwGw7DK+2fqXyD+l3cS0M3sE3Byz1L8G1Q
HrY/W1rdYLq7kGtmmsqTWITg/oz5JnOH/zOmjpQuyWHedyIRChYceb0VCasP9RonCqIteoZaWpWo
HQXBuYB7isLxBlXjJ+aJXBOCaQPeoodfwREv1yV73/fnBzuDp+9x6mb9zt5yiiihW5MJUsHWv8qx
fEKCrIqUCT+2/vj+/2U9aYNFu35B8E5FmXSADLU5LgkghUJ91pk57opRRkGnrPc2EVgur3jgwJ6X
C4FflRq6D71wBxkMAFdRCnSqDhQd3o5EBCRCsF+PYo9URcT2dQ6f3ibQg+FccJrr9gJ5VnZmCNRo
KSSqR5Ep1IaK5WCCMt7Hzvr72EmeJbNkA5/KXeBO+efDo9Gl73LBFcBjl+X+tqFTQXXSfsc2t2bq
0CV0N+9qpa4YAUxCmTmgqClXZ0piMyy2ALLGjHYtylfduSKBpCstQ0ckgOnYRnBJcl6eXtmTDNWg
gJTHFMIsu87bmbItGLnnLZ5sseHVJfaMtLaDFtFVAPHavzf8CfP6MK5bNLjQvq4utmA4q1tYzVpE
orzSHjVgVO72r8hxnCKfyJq7Ii/a6VUNWTF9irzKghoxGpgmxllfOC2Q+74q6Ui6tO6CLE9SDg0F
azmTPjC6zlz9RlTXH2eKJqxHpZlCRLfam5RXUvdPPRg7rxn2fnABXHEt41NxoXPdL+Ino+WBUs/4
fIk7JCSneUgmOnk3TGPPAmyiKTTDiXKpiMlHHVRtoebAm8i/AeuyTbBVgayhwBP/1aN6vmkJVLOT
EX51i8iJYcNggBSFnQwz8MBOn/VbffCF6A7VrGJbxYbNbLdOwMpWIajjPoN/pvHE32Px8VOtT1l1
H865D284ZrdJa9hmsVGaW+brSwOypPsCqAo8Z2NQ6s256cEtnCPyhId1YP21XS2TxxwNBgiHZ6eM
lm7ST5lKasZdLSw/mTHdUHCFrcxJQmHyfhJv5HIak9Z+F7w2WINReLCjrNts2U/vC82YmFt//0yP
mErGp7MqdvTTzZClhMFlyOSvYKB4VUSXJzm/3QW+HIOWLy1Kah0Ut3Jt0F6KQZ9auReq2mEG1u2Z
QYXY04cTTC0KwZm2BNTV+okv64KBadKGIka0u2lFr69oJkF1fn+MsNT67CFFZ9Ujw6xQBuE3gG8P
yuBeR63mvFxyCsVvWYaqKZwYkByduwWHAS8O8esAzEXeoqr9CNWghOwPiPWk+3qKXMpa28tP3sQx
qQMJDhGvifHU08s762cmIVmCB4rEdfORekRzOCfNvtsCpTQSCQjSVcyMJyrI6Wj0+B1D/sGrkz4L
G2kX22YXTQgFDtssfEu2zYVkZ3QepGqSxmvGyDE1dB+/3feEDV/oBvAGkazlS31qs6KnT8O4C7ei
7qwbGVGTQyTSph63dcYZObBD+NPepKtJBwyj/l6+QnbhKxLGHBKXqGSnkB6dAM96MDY81vtSvUDU
5WiYwDrocLL9Mo1Y2pP9VJrFPteU1Hlv0flZo0le/DfL+VR1n2bl0NceXBH3mXif85+NlVw/1w+N
/1u/0OW0MZiR80FzvRsZd6J6z4BU1doC+dxwx7NGmQCcMeC94fOW8efOMEmkAUK2fEBvZF9qgtJX
FE73Q7gFi0a5gLTG83v6CiGzSATMhNgYEWnoiZjRfc9UUkU/FmHzmxIL+tLS3ID0z58ZMbvhs0s2
w7p7MGLrHcT79PsrUyC+c4HFol5Xj2lsTc0hjwmajAjvfR7MhVgxwlYh1fEDBR3/+96gYEWs3oSV
H+bffIgqbPfvLgWXSXFxKRxANqV7/eH0ySIoAOyl668pCmv99hbJl+dRqnxTPa1ev9uCQbqNZgis
GpVm0DTqW5Fc2K+Zh77DcS17iEA10b+RbZBTIEI3QC5Jl+fY54WQvpC8m4JbjmpRuG8LMMc3727U
0WTDQJ0lRf+nGV3d7MiH5z1bxyKCOfTmRVjOz5p9q+r5Lfu7fxnJFnh0kyQVBfwLzLz3wL5dCdYY
6ed84ovDDcSAoJZv0diUXQiJZGxVUh2Ngr793tuuTOzl80OMPOmgdyDXgqQUT9l5CQAnBDVd4RrC
xDBPJKbTgUI8aD/69rtG3thM2uwxSItrjdfXGu8gXwrPw81jjNwMmLzph/I9xkw2tYNxbuwj/J2t
jX5rt4eGnSTo4CFgq8Eu+00mTTCCxKrlznvmwcEhUUf3I4FOLFCpBj7lSzDZtKfuO5kMZ07iLrt7
/21h0ol6SJX5kJKtGtWAAWLmL2oQXp7HCuQtUVHzOa9jwfE5y4eu1dHVJOJHJmAyy5gY0pdoDu3B
ChMzPp02MlJ2h//Wpu7xbReEXzMikJq+/NN7MQu+4Y9IvVw4Kipc9nKN9UVKzI59iuAJnMWt0uU5
XdL0R8U8FUC39wXXiFrZuB7W1FeJ6tGR3IBXLzrhb463gGjlgTyjruu+5kztP9U+uQ0ngb7ryWKq
xGsv25cj8lZXW/ReussO0oCAZBClZUgeePOo66jim5JOb/zfos/az9Fve5msOikVicccJCLwazVi
MNIfzq14bZ045UdHyF4bDzExPH99ABspJ48OGqiZYBtEIIKcWI61D4URcXOIV8Xf2FWYvAXcyhwI
X5lKj54B2FqfhzL9muYHjnpXdQtInWF8CuWuGKPX7HHNwZDhfO7f+aq0yWeMQ5j4hm5/6ttXXiBj
QdIlvne5ECzhbx9vYnZ9ps9Tk7e+bnKYfMbaQdkPpkUk64gU+5TNXc0LzLe1P2KIv3qbNn5867pY
HIs3aXJiHkVaW++Lesgygyhtgiu6HR9NfkJ1dBtYaIRiUKCOhd/gqQvxdnF2xrXbGKxuUHDtRMsB
T7wFkKKzHgu1u01CpxVrQdP7s/ySdOStmgi78fz7qQUf3+S5YDovMv21p7vlaKHgTlo671z7SY1C
2oUOCWICleT6LloIxqRYdxGx7Tb4QWBAiwTmwkvN0Up+qjWn5BSYa14bIgPNgGqZo56T91J/eZaA
WAY+C3UzDTevqsRdzNXwEq5767T/iUZ3Z2inhHNXQD4qZJWtSqvlzip+UufyrtPTKV2+MyJWua4d
jenNyFbVCSkw2pVsdQtX41cG9OytEdp+HyAugENPiPItKCofrJ7OlcgwrxQV+L0DJ6MemJYwDKXR
8lmOe3mzWMTvGDjXB7pfEojre14vLogFeLGyignSfIMoapE87kxsRsABRsvJM9epW3ivnqX2YIq/
dIdg1zaIfbm3ofGo4LeOmpvXJoJ9ofOaWF9jnkVrgjSYh6a7wgejk5I6zmMQPB2Y3mcu88LsSKDS
q1Kcxgau3mZDrJJeyXgba+ouDX9B4+nuIUyNJApAfXlNOhsGSvMsIHzRINvcZz7o1huEwEr4l2x5
nr3VLN6bPIrikMtpGPWl1ZTVlRnDX2iD3cKcZYkAoplCgNwXzpo9VxTXVZjtFx2UqR7GKZ/nm9FI
942na3dvgoQY3BExXxRPcJNBXYom1PrTei5GI0v3apdtiUGF40g2EmlutYG1W5GQlOZsR274voaB
MR6zAULBNwTlU/pCK1MDAk8Aq7iORt6TNqLvDQ3jnJHLXMH6cg+/jFblT4I+w865SlsBorGxPBn7
+yQ1puEN844p6aFPEfWXayJpTiixgUKtT+OToCAtp4FGKO3bVA/CfvbceRSLteKLRQ2inFaXKVGE
q1LbbwnMEDBpOXrHR5diMOdD3y9g4EwZlyc8TO8McY/KlafLhwLRwkUnjkMAwm7qsl2cOsbB8iUE
lF8lSudQjerD4j9bnjwhZRKy15P/fgYVLi3gRf0Ev8Me6Zj20mQyIrfUyTMtyEnDB18U+SnLjrsE
RbDzg4umoebqZAN8XUHb+2Lr+QCIOuGFqag8xs/lhsGMoxSzI4xjiZiWq/Tr6V41RMk698XZrfBK
CVyGgiHPlndLWKCNeJ6sDMAOhl+y0yaaA6CU+T37m9sPRtkfBQgGG8n1qPu/6GaKy0VxAjLN0Yrk
QTyjoj6UsYYlA5Hue3uju0lzjIHTvoBTlFcMrqXnMeWZqdhXa0rSY4ASVKhWsccKTHo6+dbykCB+
6M7QLfGzucxPqVJoPsQj5uSCnJMRRfdLwQnSC4bCKroG/ubxAxuLiAH/vCMT14dBtGofk4NrPd84
IjGhdVCS13w/FSTducKCZvNh7vwBRXPJJv63WwCm6gJsKFz4d86Py61PYDOrqOSSJhjOEN/aIq2l
KHn5BjngWhvHt2yi8yJkhoOuc2r3L5/AfE/QBSh5J2QHWjSAlWJ7N4JtJFq0eDGHpasyOhxSv1zc
3ubLNuoeR9XmKxyh9YQKLTp6sWDDdw4z645gJFQoemOGJQdipOpSrZZWj14zR0VB6XTYPKxRGuWw
nv+9eV7/qpzQgXOReMGtnVgKI9siK3LFSjjEX0UEtJRtwU0LHT54eHw7qWccKrxuhS4KlkQfOSxd
AYfWa4979TMBNHNEnBwZ9D9MXCuld1MyP+cKNcHBLvzye40kabeplgOIyFlgD72O0veOkQrIIOH6
qbfS3UtcXfS9XwP/Td8uhud7l+CgsyVIhkdJJQHJZOcLmi1+xDHBlJkae4JaRKo54yxjW7Z4hhm6
q/PWzlbiDiIncd9GeHTvar+VW3PhlBj4Ny5sHrtdeuUOkBzXQZwPtvi4YZuFFLvkV8lARd5Kjxq+
AkfaGnEQqLn2rfd+IhZLVNp/mBZvzg73CrjowcBZqI0GGzod2k0m6yTgibVEHUh6UZVJ+D3xe6Ik
ZyV1dLFF+F9zNWzgYxbekeYEGJIFEyDOvOINqjVO8WmMtu9MpNeqwpKzoNkr1MexZtTBGMdhaseL
vxX7JRH2GcAnUN5yhGnuRRmjob9OZTZV023AgI4HlRsopvwlQTrlzMPCaf0j2yzH+zC5ArNTgtLm
cuoyoxgYuB/7qtucKPGWihh4I+mTl+jjczeLShNpKKjKBOv+67YVaOloIPG8VVH2e5xYbvQVVbbU
cNrwtDwcnUJW0fPaKg8fNjsYrKSKpt/lDlmYDzAZkbRDuybEYiuU56mKiBDtlPFcQcYgopuhRwu/
bOQjr/+bFFfzg3aH1BK+GTLAS66hdh0ewYKqiODJzm/vZRUR32yiLrhWtv9W0LYt7EK4P0pdvm2F
7Af8QMktXJjsNI0SpP9c1+5tqFRU7qVsjUPThVo8eSF89xn/qKUk8FbIugs17VrrTHx3Ej6Uj7jZ
zH7DWdoxLAYctJCajAzgbilI5eZ8hOSyspfChoDVdLTDIxg0GZgIS24WLptGTndUKXEHycEh+Vz+
Um8SZzFofe0Zm9CGNUPMW/EnWH+Q3V+gEbZv3BxxQW5qTbJEBrkAfdt3Y42Ch88nRck3AMW8XDMq
JLWtUDJq/WkSA1fJtjalFDEnkkARSHL5S6p9VKNhihxDv5G458KzbcgEd8FAPWc7JGfeHxtF/BIZ
t6slTw5HNNZCSevgiuiE2VczWJ1TBV9gJS8R62Z0h5ilvUkyS8Cpn5+bgdczCNFsU0iek40wLG+c
6H8vua7b0ITB39IJeL+2++oApiqSLXdyxq9gs/ut0vviuCqce7OmX8IuCVJ00uGzAPUWoZSIB9/G
sFdxZpA4ZqdV4qRl7DMbgC4jJqkOK1fVYxRZ3Ga3d16EC0CN+vU3UnNTANq3RB81nZ+uuPQXa5SM
3geBGXG4qeRT0GIvSiFqmOYtAl4lfsyfStMmt8Iz6gKqfGmK2ZQ5nsmpj3kqbDf4aTqOxSSgV2Rf
xiCN2hbZfbUglhGaXSx+RVUjHxsD+jTsrxG7TjaHF7/3bMFpwHK+Mg6Mo1jgjrtWdyKRO9dQR1Iz
tRzLHjrxGgp1GTMyOUTP04/uDmN3mIJ97kaAZ6BcGXDELfJ0sNnE3BOytEQc8H+SjQQclPKqXH5+
CvNYTTQt4JetcznwpuZ0JjJUTnKO0ChXdlAhExzTGDUNBVDHt+ojwC9c32eFrwW4gs5cvjAh9kBp
7tU0P+QmdjXtvVNUOJWLRwaZPm+NwHabDswYT+0yjymeJ3vqrTFIClfdwbszL0Kbvo6kFQ80lEJo
4bjZfYnBtID/+rixg38HgZKLCu5PC8KMsO6ewQe7T5LXaYRcXAMWwawIlcwVzWgfBeCqYXPniICA
D3OlLSukOTL3ra8ulW7F+QSI7M74vTgnEVXwJ/wijBFULH4Lpkmh2X70QB+Jzbb0UxYiorwtiWxF
ks5g+hDxASCWuru7EvpiQnRBexrhT/S4TXGrTx0wtailipuTUqY8VAAaD0eZS+mJz/1KktDKfw97
2eTHo2fSYerfpNUzGzObnVAKLwb+f+ByufBzJSH4399jvQMqxG19xncwSUCCdCUoFlLWZA1wZI4g
pcy6SCQPsKZkkhE8u/GsxrDrGYwJURX09Qvw3XMAqLEZ+dQav35EavRjM/cuaESpftwB2P1ZWiV6
r6oCfdpO6TlWr6nOxvB+ebomFkgzpqBjqt8/XNs9BOo4D4n6EBsBYKa89v4O9/alDvALxPUAkiwp
vx5aBwqynz0nJKTkCLXh63ZLlki6OQDDKTNHPsLf/AhARNAw8/E/GR6v5xZ3STtWAJIXBNhrG70y
tKGCBUSrWHI72EeBHrtedvrZJhY6qrL9BafAQABpaApjLe5dg/TwvGufGizjzeb2EJKNLjJwqjEn
RHsmgujyO5GY2c7z+5G88cjFSZY/OYWF2ydcZ+0Fv6k/oPhv/kmO0ZMG0QTLG8+l9i6yPoVogsjd
FNp37qxP5WpCAXvopFknyj25k+9OstSi8z8klx19p3eOH4+CsV0lL3Iswj/WJA1+00F+ZMB54/Iw
seAPHyjKCRbWYkyhPG1M/v4hBq23LiKxYNK4x+luEq/3Se92rUcKtRDSL34j4tppVTidRONk57Ek
Q4BvJQS+BwNOKYkl7ciUiSGjNZuSDAi3zIpr8INFofjcwoAHDZDpRU+zOYe1SJ5ViMCMTeCT2fwu
+PqVdR8WeBJoJCKuwUlo06JpRdvdznFHKJx5P2IeUec5Iyd3ryrAaD5nKV0DosX07BZwsrydVXPx
gzR/VvgawbPVIxXhFDWKFIpW4wE/J1aHo/geSzwU7FcmROTOaUsUERTybcNdKBOuJ5WtdvIv9v1C
5slG+Bi19mcJQm9IkQOYlUrIcV8PvrEzHa0CY61686rF/nxtkEP+QbPMUM7xsFPh43tR4PHLIJTM
y2E22Bu2eOmYYbYRcc952zeouYmA6s6gpJ9lGFfr1X/156eu2eVbG8rMTDogaYfBQzk29oLaoD3z
EdGjz0buRoE6QuRICkuJozw00c8IEs400vJSADM85ovKFwbVVjwF+FGuiqfavdshLt4xPbuY8O1n
YEqrvSlDfgyxB2fDemTARsK+eavBo54K3oTUv9tZKXO1SjkvCrQNc+ebsNTGQOT25ErNTtKhLu++
7k26AMBGQc7CMB5yzJf8nj3YcJJ9juNbWP142K6h0KSoGJiJarC1pcQQZ2YZio0rXnqyiVqUEeDi
wP6E7ORUH61S+1xWKQArDchnfPp7uuHTOnoU4dKrbu84fuW4YCNwNwZT6c0fZ8zAtig2dNdMGIBu
FYQudjN3crmAsn7z8+P0uJ7KDO9s+UeOMckSn+Xaalg6GOc/jFXy6YTXtqR38OeqQmJbD8bORmmG
1VNbQCi7gVcGAl0OXx9s8hmex8aa1HZq4pUqhUuOizjT+FQPdwXWwLrb6qKEmgHa/6ocWxVSB0Fm
AIYVDW5z/YLOkkyHb5TdBA/aI59vN5c6OqZ//LHr4HZJWo4jmaVuzfz3ly3n5KhkbsF8LhkA1Isd
rkXsLSVNQNDR6NrCghhWZWYukj3m8MTVWbpgByarbA1ecYsApwOUZ+CsB+QuKzAStwZiGmIs7GbQ
Gs9I5dtaiuMuvY+gNT1pREgW5uI9/amWty6S+W4XU0TLu+jLZ2/hDlWpE6Efwggj0+pfLtY2Rg9W
A6FogmafnikLUSEOuiO7vZYhCp8kB0XbfB+Uj7NhjxLkNYak+BCo8M9mKjLy7dbwBUgQKz1eNky5
vVBoi+ai8bCHC5EzCunBf68bMDRWOZ7mE67Cb3Eiju/B2eisYKcU38vNpV8i9pOKVPbp2joKqgMx
n+aV4Hi4M5tHeREB5RTQRSbLJ9qbwgzlAvlFXtLRLi+qr+TPppqG69GAI0RD9WhIERpvBmt0ptrv
e4OirIjksIa/4R2GGPJjPvG0YoGyaVlQycUFJpvIz48slbeLMG9BF3lxMHmr9hr26F6uik87eAkb
y8RAqyYZOiNotBN+W8xdZonx96d0LvxUmOnCQ4zg0XsSNKkeCpgWiDBintjmk935OxMh4pA37pJJ
4oQ7OuLyvDieA79VdFvQLUxo13WfJdYcnz1GjKADA5MnpJnTrmEvI9nefKq45NX9TqgWIBjo61r7
eShrdK54l9MbMcsvtu/6O3GQ4m4ntdm2xuuyO95EcEmgxauKuBEGTvncPoxsPdVZ4itoLE9Jn2MW
kSydnlw5pa/lwZIeQOPmdqyiYe9b78hTdcrGeLUQ90oXfJhMqP4LBA5mNjOe07MyqLs1BHSx55kO
TH4iyFFtgon/SGSrHWPrLiOZy/B6SuKezAkswiaDoRzzHlgXa8x/sYcHY09sLaU15db5EbbsNIAj
Yw3YftWXhraCxWho0u8Vd6mdsvNuDbfCEcwL8S3FZQ+VkpGKKcnfIM1mN+rdrhRV2oa/7rZikAvo
1IZyShe7VGMCDrL8zhQ8EI/55bHTdOmVNEgaHJzj36h2noqVYdEyCd7gr0lcUgJ181rnQJngzwiv
9f3wVwjBvaNELU7CPKmRUgTvNkf1DyquZE2Ch7noD0zHtFDhXPJnBSNniBCPl/VPBVTKPHCx0dwW
IDvpkuYA9nHFL+Ylj/89Zs9Z8WhhNZ920JyNlkLPuUwXHLNi89feq0vP7x3hfpjQL90cQGKXt2QU
Po9FF4SRfdkfg4KW9/6uVl8Tze6rHRHEHsoqPA609gBehAGbtKlituiuCkGZKHmnKR4iTNNI75WM
qNCMjZ/uenjG5NtpoH2Xb/MW5Pwm1zCsIJrsrM1zZpw0eI9TT/g1zgjYDcC8q331afoo0ORaGSt0
MXsDTsDAe6j9tmAXkwNG7z1bOi9Rjr0UAJlQqSq/LJQtLq/iyYcu6u5SF6mxRPvyN+caP4jZdsI9
zbkAsNU0/2PfNrxjeAH0pmZXAdzWqD9CbWUS+iuOZOUrzyEs1xxuoowxa6yZQELWEm7UqVjOdNaj
EtOasskJNhy8877eFcEW4E2ecu5y8IkZtaCjna/tZTkrJl4DiXERMkSDFgHZIucr0dW/Jx5TlenQ
YVI8BhFjzKkFyDPEoIJVUJz4WmDBW2EHwe9WzUSrrenhq/hsAsGJ8Tz/E8bFYh5VCz0PNtKRadGV
VOsSnEQcDIGmFZR1vmpkoula0Dc4JeHOfssloMMnf1M82BrmXVO3qwBFVpfmFgsvhZNA6tRopdse
EQDk7ExIZU0HAaH1IiXBFmqcfnk6zOoZLzq8o0SVo+nA2FiXn6jr6aIUE0vA1MYQVIzxlL38/zeS
pkyJ5xPzYlDu+olZ970ck36kwRoILrg49z1EHoj8uWc4wJo3fiNlP0iG9Umxql1tAHtzRiT3KdWA
eSSEEyXIsy6+e4yu1Yoz75QjX7E/pMlpYcho1TLQi3RGkQaIxkY2RVFBBnxzefgRi5Ww5IZ0ZL7w
yQqiMI+vodRmiugmWDtbb34xlB8xcprPGq6ryT5bjziG355Qx6gIEziQyen575ihi6MiR5gDTWBW
ZypSohfHmIiJzaTUz6Xkbaxq370ZtAsZ6wU5A/rR6vL4l80Zq4ZB59r02PrH4HouQ3+M6xoTNl7y
fv4OKLF1Bne2VwMtpIINcmWuWAu0ZRMf+jUVHzoY93sAAqgp9d6jFYpA+FfiduUK7rOryIaQtt5g
bi3JMrXIc5OXhi2kmBucbVhv3taaxBQO08w3CvVbKFsauTOMlIal8IL5DyTXODdv2YXrejwFp1JB
wNHoLC0dj6gDnC23ppQicSPnXaoOfRw4wQLB0pNEn0d8hoMbSyouU1xgfYDFKaDQSMdn3bI+fZij
69AVXr0RI5Y835ypYjeZoPVL86HCAjOp6xSi8xjgJ6v5BpSMZEotQAqyOEV2oRHI0/Bnr/bsJ3dz
0UCCAvFIeUNS60fQn0CzyvJLtBGvBqAqkZo06MyryxUfB80IRprWr+s7fzUys9CswCpF2bdH3KYw
d7AsJ99RAEl+HqMEpwqk+hB6EPwfBIYzKAVhzHTkUxmEY97/dhO7dD4xQHWqLnw5OdlRNQ92yWS9
aSP9r7pxuh+vU2wWyCb/2LTLGJvHR8/bx/NcLDaGON6Gb3tJdSQH8LYbOgANeFS6vmYGPY9NSsdb
KkPOOfZSKCcydUMXA7LDakYPPKytBc1DzW/Jw4ITnr5KcHKfpBvF6N/DZ4qrUvnhQVb+IWQhp66k
lTEiBFQcFUMEJ+JWpdtWQ4/YpfBsiwPAGY6aUXMEgTuwckSpI+dbUcFxrNt9MQB3GWafDr/9cu9y
KKoRlVu07HpRCWxdxVwXm0UNn0pOdswhAxsnszsrH956fwivOqcI8QihSU5agZzvWnoIeIcl9Adb
BhCpXrZDl5WC3oPTabf8uOMnKbB5+BDZ4nPWMrJgL60lCRPtqqleC0Xfwi89NIjbZz8BFdThUT4/
9+Vh/tCvX0PStB4lR1yWBUl4ohzR+8WfpEg1/hJMpRo8kcmWLf5SwnYsf6o/hb1BTEI8wJBAf/dN
9ltRyAPpE7LRNjbgPlsFjoNs7emBTeVVRsNbjuuttWd12q1Y6sx/kQ48W9AjS77a7FSZZc5lCKLQ
XNcxJU9IcJtC/Vzm4h6BQUypMUzGvfOgPUreSj0DfYRc+CBrz/V1iV7RIPgvj6zj7hs/yQIm64vJ
8qvkKlPLs+Qh8JXAjn+44LI9fpaJPefS5nMcI+9WDY9BHsMJK/FnnLNmGbRFuZ2TYh+y+j+9ZCeK
ifj/6xBZzQAUJ4Nar+nea3J04l9IFLD5aSJNR0TX81a4xC1eR8aA+sz5hLy1DHGPfg0PH+DecDhY
HOt0aojnkf6cRFHnQ40Tl0nROGk6+YwLihc4AgKNFFSeQOP4JRL2AqDhj4SeVSkggejRZSoyT/gP
STrw8KKPqqqoRs8lP6CV4gG3WUecDxmVZi8sL6HCaAgCe6MGeu+hP11QLRElGQzudgMkOxdOzHds
UONt6WBfKd6UX3wMfq5F72pSvsJKSRrPEa9ofwRR3aap6IP36wtMHm7cAnQKwkg058+Iua1yu7rt
53datdhniTf+uKfGwcnoGz6C0K8ejv39GYyr+xBQNyWPfmjVVkWqwod5jKfesuToiN4/uFGu32sS
DqL/cbpWzilWtRzA4MLitLxIZZiRMXriduJQEK/H+wlQGNTCnv9UC32q0BwC8ySga2ijDWt8iZkX
7yFcpxpRkrQ63uEfm9MIDG69mN6xLnTvC4Yfp71wja6M0XUEMspPoLjAfyXM2BQBCLN8GQkPB4Fo
9tZwdplg7R3a/VWZZEDHnlNp0k6gDvhSXwSmZcj4GOAdTMLDoP5DiIBDZbYD6dWK3zFJE2MBY6Kw
IskoIcW6jojnMZv4Pe3RyD/17I0+vmnKI+5DsxghbRMLRTMJRNPnuOa619svAsOxutniNyg0P+Hk
NxOVgyAXendQHpbgLXNMj+yLe/NwKnSFoOEFmzIY2z0o6VrZw7hTnKDagemXyPfLkzobJz2CSuXC
+dYdoT+SWq2KjZutEXFGirm3s9kO9ZwvzSrIuqzr87KbNfO6zSo35kTt9Nx8XqtmQfIuhtOFysRC
S0SoP8QngBlxnQD1wbIlohHalpC6vwO/IA73tvpMhSt4oYcSJ4GCbXliDkSBIPpim4dD5OTRkkYB
P3krTqB6u/Bq40JNJUEeDf40g4VStcNXdMqJBT6Fi7C2Xp/6eh9uNwyC+YT4jsqN/liigF6Ktmne
7S2UV6C92vbcFXW3XHNL8wVc6rXUvj2cf4LS/KlANYsrPaNnomoB55g4r6isB2xncpBusw3rxq+2
C6f7G1YPWcIX+PeYDxNWaI93Iff0iC5qZnCQsBxyozKjQLCP49L3fkbeQpNA2TH/zLyTiEc0SUrY
BatW8gbN9I5Xqq6JFf/+AhdVgPlJHMDO0uunGw/pRNC35hvDHxzflTl2UlaPgGkhMFO1lcgldfGT
G63L+ftUqKWnfW0vh3W7Kw/xtwMVH15goQSsA7HrSvkZaod3nj1HjS6pYYAuyMKlKPVzSBmkU3jt
lxv+vVdrRFT7GjiW298o3BL4do64Fs9Xc0aLAI0MQ5489Nbwsv9XrCdo9Os6QcVEFSRGUS0vxY0x
gbijfk7N3az2quQPxi0DoOQDizeEnKQXawa7UTkGGMpQ1t8q3ffGE2qb4KA6nnFWaO7msdoSUeSd
6gmoZpwsclJMcJGMl2UkYKs8+H0Vy/NT7ffFrVE3MlYBueXAXDFZQTjBJJUUtQR0dEZAEqTnwWdm
6wdTXBeOZYGY/qES3cFWAcQZxSJNHQakmaTG9R9TFtw/fZ95BNwLY1uimLPyQMjXzw/XbqRg5EsV
/BvCSRSqWo/wowyz1WXrmX+QFLU45N41yWZl0qaABVjv8mGHjZVbu1bY0ZpUnFxFzN+FjzhpnYzN
69urse8oc2ftoCCfkNGc01R0lv0nLTRPF7dFWxOSM04WuPPO8+0sp0h6ZrehtgUm+5CwoMwcfP7E
QKnFCbWus/WNFB6j+OAu1f2F71omrahBiL7aSsXv5h+znb3Jp3De50PZeJuUTd9jHcJH72OjLW26
Kxjwqz/TxlNw93gAsFTr1SZSr6zhtcIUVct0W4g0ZWNUHc/SdflFc38fiolj2wf2OBJjyreV09ef
tl4/ozhXTa6ivxPMAx6ERexYjNKCX/LZfW9bvaXMJliR9djodJWXgSTQEZ5ndbc08bWC3I+E9C/n
zvc6XcWLwufnW365nQXJl083R3XjIuFtepn7E0NaQ/SjhKH/ayhWliI9Gi0Yts6xickMkCk3mCZF
Uh6uOROo8NI3eunNnbL4uWeFAnl9Ib+wa7izNgqQ+1bd+/WTS6PtTtMkx9UKqehORsLaPHK8Uqte
u2nI9mW4wpmhzZ0tBcEblD5PAKyIRz0wQRxCql9mta3Z7wDgnQZNXZ8VgxZ0SuwveUkE5FkNPmkK
xNGcwiDNUMaB/UzKcVgzI1kSxVOUgULX1BrlN4Jx+0cGpqkfvBocZm/SAgSUy37uNPPgDarCrdkQ
8jYTKXP/8J27VCMxfyvHCKPAKchf3nS46aB/kIejzyfTj/F3nWtxnbxsb6ucmpeQJ7OmxEPfBSNg
fPk3dtgzCVk7DAF8MawN727PZUIQm2D3dKG3u4zlb+6eKyFRL1MjyLEhIBcvmcH/9URMATIH7NQ4
2m9PV3LauhEEDAF1mvrV+7d0WLld3cFuFxJZ4t7ae/iI4/7wRaMuCJ82TsYqXJI331EaiupINCjU
Cpwl4LM0oIzsemw2k7iTntDPdJgLZ0vRYAdXOZ4C13jwN0KFJmzyUJCi+Ydoz5NWyCt4ze8L02y0
wsqRLHhucrII/y1OrEIBNhFMrFBj3OrtzWuArHvSth0j10xEOXGOOZAr0nbS9zZc2+MFZ4ZlJNRf
dEREjXAmcJmbGcDIn8iiYyLmy1Jar1hd9HFqe877yZ6Uox8sD08Ze1T312Vo2+2Rsm/q1Yfv+tp6
gdbxvdvdpX1d6nr8MKXV6pbTSAicEVedg3hSAc3wq8X4itW+lKWfnQ8GQYC2hdCI1lGVDToTI7v9
x1zyBWinVqD1s5ZumMgycHHdodbKeosNwpn38Q5NVL3pwbOUxlZl6fRTHUnAuorURqi+zmb1eHjk
u5tIX+E8nr9mPzfoanqiuPluqDgeVp2YF1hWtYMN3S2v+RI8UQiBlXVtSmxMSDeFTxQYEOrTIyaa
/zTrnEXlgoSMYT/1CIVVczuRS0BuCyTIcV2QVwV2t3UMTzAhxojx4YZ1t7GWY0CQjR8OdPK0Uw+T
uICOFDQ/DFowd+oPds49gCfz0pR5kDDyAYZYE/iGvDlM9KhVI8zQcMua/L8gILud/MG4Br4qcTpQ
6RWVjSiFGXu0XK3FTcQmo52bZ4jali1hZJdn55b8606wwIpp1Wh1NRRZSCCjA+oF7CwwjNQkfJU2
shLMbpz6Es93NkWqvaSd8WJhfPyB0r2JGdhO4Dtf4Dwy+h4/3JBKMm7dIUvdFsuf8k/PbQ0vpAQo
jWNud7iP+kUEfqgTg1F6aEcC8N9QzKE8JWtw/wybPzkuleucZPzSPBvxczvIC4C5Dj51Cehhl7yL
Zmw19Jn7l7StX12Q5UurWCdMcJoZKre7b7r5jw8MJkGZ/G0MnA0aeNVtS8aGBNj4xBDZx4RN5/hN
Pb88jevIHkb6vc6hALa0S543Up7td13OAw7e0G1ndw+JQ4Pm0nE3x0GaYLM2G78F9L/HUjl1vIU5
zBFx2SaYG122zNmdfoJyrsUbfshyDtDvIHpwjJIsjVViQn9LaWvEhStkZoEppmT8ffrSQDOOrKGD
MaZX0vhk2RIoMnc6jyweInzBKxxFBOMBMxLWyRSicXLdrAPmnXvThng80i9by2YQY/oZW0xiLW0h
wob/05shjg8jO+NTmx23kFjOGxhJ6mxCa+eUaDxaqtLO8BFwjVk/TeXZpd7RIxVvec7VuB4E0U3O
dqEkY78TDnHKzAdbEA3pQQBFQ8oghXDm07OUiCxw73na8jDf0Kpgqx6ig4u8UCx64FbCi0uMN637
OkyubqB0b1fsvpgKoNAXbxKSrpDD76Ut60dAjYkaXsoOfcDugVYyp+vSUuRKTlC/O3LaeFOD5/s5
a3Hntl3D6+HX50aJE3YXy29fKD+S53v5hq93uNZnbeoy0N2ZFxnsL8cB+zItrRzwDndBltZgHQc4
+7FQvUMQcSLoZVcTw7cAEJI3FB9JLxYhjhVNYqUrkKtwk75kobWW+vRapOx0mRVNSnWvr/QICyl/
6SsDFRF6Vn/aBC74KR3KwpmVwp6x+55IouThJbL4ILlpIkw4DK/2AKuuPbIcGLjoQMn3dTAMoAQO
U/lJ+52XiwrhpLp0JK0Il8Hgols20X5X9fujxB9bPl7+YEJARN8Nf+VQ77OOJiaBTQajrUgGl7Re
n66C/oMBIHkYqNC4NoXWuBd0cTkZCqD4/28nLKV0hRrQzFGzLSSU0s++TsrG4r2P7DNPqfVJhmtX
/JUrq1JFSUicOnHrT188udeYghVz1bd4dYBaosnR+Vu6Fq9ot6ZsFRSy8v/UGFLdWKEi/PSUQNa2
y2uS43HBpJNnDnTpihw5eKTzANdBS3xjrUTQnPnSepaQSEjDfw5u5WBrGI/FDWHcGH7dicpfdh9Y
PyVruFGVhHYfdZ+am3USTYFk3Upvrlto+A+u39QEr7OzqG73WqG5YOI7DAkaoXa7y7WKY+mkr+8Y
NE0sQHY2y6ZAJoMFNDoOE7LxkG/9m1iorxUwpmTrvm7GBDWhnWA8SoSHDfIjGJP9zJuRhlmG/1V1
Sb9ac/C3XNhAEKg3smhWS0miwV7xPqhuBUSRZ8v28tdhOitooE2JASDi5kLHKAGpGsyTLfgR8hQN
9r12rBcsbt2Gw+nWx50yJihJajpInNGtrqQQB0TV7FJfQk8MXNf6B5LU4Q0z/mubIHALV1HWDE1k
xQe03fHcQC3Jq9xfao0+Ht6cdKSwzY3WUUuTllpASU5UHksZe9m28aC4UUYZBy2NHweqnk9/H2Gz
AZBjs/Y9qGM1eRVVFPpKmAgxV9Cu4cc9G3Q9cV3SbAHhcp1aCwoB85R6Yx4fGrRjRvD/5ZtyUKAA
wP1fMZ0pZ3m8mSfogLCBQddGDCIXy6CeN4Acas3EpBMMf2mEWWyvyd40VIt9asdTFn1i1/U+zx8v
sSPVgWuQIN+QpBGrMD9KgvLFhTHD6vxtjqOz29rjIlWu3wgkVlw/7EQffgO7eN72AycMgx/y60QJ
0o8HJPMvdBZyIk06q92QHwXjBTOJp4u77sfqiAMXl0iWUB3XWH/752CdZUsDS+9bdiRI9l3uVi2s
ZXbbGV0mVKtn8b+V6a7KKHAijEZtTBXIxQx74CKqm5KUi16xux7v+MBAIqbyK1wP8U9amhv5ImRj
UM6KITkq2neahe+G4QfBRTLIut5cmVbZyPuxZdX3L9g+dEaJu4pTlCKU5IJ8n0y2eAdMFR/ZMFH6
qcOWQ/4kQ2naIVR5hzqM74w/vzYDtzC7cEWFV/m9w30i3c5P1sx36CieItLezNgS2l6Mi6irZ/9O
6jZqSj8yBFaBYbQbJzR5hvPXO7/+fwLmOZbRzGBJpBaiUC+ta0tA8av+5zUevEpOoFGNyixPAoGB
r7ddxowviQ2G4BqO2tXhOOn5aooQtFuwGXst6fI7MHucj+eGvSQUoNlx+x8W+xRdOV3OOlN16rML
BSNJs5dND4lLaUXLVPRJKq6Vvw/ef1b+90ZZ7vsBr9wkRTemWb+e9XlFTpwtNmV7getv9qV73rNS
FZnfWNo241ksiGa3+UBiBmvlHS+ZKP3lg3+LbJ7h0WUVtVvCHBQeQAyH/85If3MaWblh23KgwqQA
6fVBv3EGChTInNqllGA/u4hgV5Fmeuu1ERBrQhsQf5wAEr65m3sz/AC/QjyWxz4Ggpwrer6OzpD+
3xCCUSCzWzrVlTTekqOLvDD7nan3MvgFRpa8osMGnGR0/0l7WXS4d1BN/APsVFcbIe6trw7tIN88
7cwv2AQ5mKxFxBS7VEoDaQUYCrM8LNqMFtHv6erkJltRBTeqda1qnPmpidKDzKOKI/bne6QpJNO0
PWZqxMURDv8k0HC9t463K2wRKD63soaTmj9TGC4hSFyEvtni1J64k0agFPHUGyZiRaBg/PZRxLxU
x/uH/46Th4IxrlMrY88U5rFC4t59rSdOsz4ia7L46VsOFx4nAs6FN1b5YsK2S1tByUD0djye5vZk
8q6BLYIF+Jc57vyEwc7ccPmGodoKprsuwPZe3vutvwUQLRO61yKhPMnL/KMANTKYhHNmBzp2b3BR
W6zop0FtGo/NCJ3BdBZKJOSZsv5PLcZz9YM2aSRIBtTa/LAvzsCouPU8BkGvBrF/t1YpMW7euzfE
TOg7qNWwewaRbVD/yeyKFueyTqzVc39iwA2sao339akmYY++HVD1p/CewY/F94RPWVNj2id0ZXQr
4XQ6R0XxaKJJuHQPOmPnVrUngN4fgTxpn/kHO45nIDTFXrPxOhK3mXneB5xggt6JeqYgdOC9oWz6
39DA2I3IWS5WupJ0vqMFgSXSwgDp22LJUEP4QOVLpmXGgTLuADObnSJEtZ5m0NJ95jRAxYxgVvfx
qyKrtfUXqiLpEP0BHXqaTsDEY4nBOik9s+iC+gd1VGcHutMsXlL+bP3I6qCP5W6ujlX8KGJPNciP
zDZ49vM2r4is6G5zBhUxRsmUjP4C5tjAb9qm+FNDtXUEJDClJ6nzfUYecJ5bt3lK+C9yz94YxhTo
8kmK9DmYDI9+pphLsvLy4KbUiol3TjbY+N0Uj0LpCaqGUNYMexm3tTaEs3JgO/y7jGt2YjZ17TDE
QW2JASVc6/Az/6M0oVQMpyg+aWjumE80vycUpWYKgv2m3swGuTx/GF7qge4ejb6Qoa0/syA49scx
24IfPJwgXJQZHgiXs0sVSlt/uURjEfSGRRgElfNoUTiN+y74wUXIzL/kmcI/QPDktm1IIGJ19VaK
MZ3VFyJoBxZk/YyyNF+hmS4I2dab9wDH+JFkpVZdBEI+iiZOaPBVKokn+KiEgZP6BstVKMmw+65U
n1e8KzwJn2kT92YTdyg3GOwxBbk52KntsWgex1SYFTkqo+dVnPcsZM5DAOwyfHwf85n4CX6yvrcO
JoUPAINrhsp/pEwKvu0dt6JH05kQxEjfE0HYjhJX3caC1RgyzofVonldchlUCsUHeGFrUqSRpzZx
vpHfaoviC5xiw55dPImMpoo9B+TbwiRgxgw5+iSB8cQtpjk6KXwVtPIMN4xyynbQ9IP6twm790k6
EUMJcba0d8GKlI1MdWAdCFipcOrUQo7shOSBgyT+MA9vlufDsPw7w1OvDxnVrTiMPut+LRtBxem7
Z6VZrS8QYJIq6Zq0ThddfRR/yVjz4+mDEGV8lGE+s+g+ISnBm6+e3fLQx/0UAjKhfGes+mv7FedY
FXFf3MABPB2Wru2RYSzlGJjKit+YvbuEGiiDmeIGe5bEFPQZudL1LGVCaF46aCgTQ0XLlZJC438p
fZ7q4KpKojn7p8dLli1S9d3eq283JJs7B3eLYHJOKReWTIAq9GM2yIUy9Kq3XGTkmjaMI7NXSPWM
rI0vzw+At0y/4EzV+WsTEyHuNLTPOr9EjFXA1UJajUY2q+iFkg6oHOjJS05ElNQQdTdZlKHqmBaS
SbEsrsKiLWZ3I9axh8zs1NS6nkaThksUMKzz0BYug8GVgJvSb+NljZszeIxqGOBe1l4OR+RIlW13
+ykaUYv8nB6gKRmsfIsd/lEMyf7xov31FBfymu9CR/v2rU5qEi5YbHaueElE9VEumFmL0QdstQJh
t5bvXNfdFAp/Xi4SbUBHH3xmjIe/PGUySlr0CaqVLWBvrkaPRL5vOh/a4UV49vtG0V/31WRSI0kY
nfTGVBGgJqO1/hL89ndpVRlHXito1mMSb3LMkP1ohsyXW5kLKc/nh0VeZymHiLlD2odYqDNq8b6K
4r2kU3RZ5ylQJ6xvf3Ac7HsukeosQmn1ur3UAF/3BPVIXOHLVpiETQyADRe/YJ6zzwhQu4ONzNC3
/vwZuy4mKssw07VR6O1/04UrCf5ci/luoZb+DPP5o0k8DdynBuVAXiSdEUfJe2QxrVlufndBa0Sz
XQZTmYWj07tT10lUb7q+m1otg/keq/Kn1g89fBXpM8kqRJzrLyg3DaCRhyWXynP6mWXNyl9/siXX
u4BbGQkDW4zeDPwydRsk+fM3UYlRFm1Bi230ckxcPBm0kbnWpwFWF90l1HBuOogyIU+WN1Y/DObc
edn0qN0N4IlRnM4Izak2Vru9pKfqyZsrIgMub1Z+/X12Wi57arvBgLnspgF5SxUJMZik6/O2gxp5
uxn0l66PaNUjtXXzB5l4olp907DNYOqj0QriDFp1W/FQPXQjWEtQ0yd4YHGbpgh7jRzmMGm+sH71
7hEbUvbRYDbsjMGsCr9Y5pBf4b6NG+WxOmIYc7/MU4UpcbH8Q3lxYEPZaVTk10qYLmDudCZqOZID
o/TfWY7t7doJBds9PsWTCW/bqOjhITeuwt4YQCO3tg/saNZkUZ2hRsIV5B0QMz7jcTqT70ZhA3ua
j+IhBoJzxWEkK8//TCLFZTvCG7IgykZiCs1gH8AkXjLDcp84gM8QRVDD3wW5AhBMauRpFnOKIdqn
b2rS7QqVg0GRntrpH4aVFtLvQVHEcS5tbnM4bidz0n3zVjjrvKYngI26baD3+aqZ7tAk9lq4nWi3
Z9qz7noedp1wyTOhgspiULbYnDDT7ngYr38pAt1InYK/FiCyEyuFlBeCOYE+x152aPDSXfL5yxgH
uq4UBuZmqafevKIt5iJf3C0GZxSDGI2GaAxzOsoP1JoFV0ngfYbMT5acjaES67tbqALeG3k+MQoD
KpMP4bKSXe9NQrmWJhamCmo231MMLG48tOQijoX1cP0FLRdB2lLMS8vrvWE2yv6xQPqNKhyyIBUy
qHH7jXfsY85xoOB9zQ4fpw3hVBrtQfMkLCBJRIxteJsSSX185dYwqPImYTRlRNDsFpEExAwA26+K
Ur94ODAAtACyP+kJ3ea05V1O3TOcJnb/rKaDBwFVe/RPnfd4DD4bQXMUB5BPT7YvjteAU0qGGkle
FMYdhgnGbzgf72LVjPdYklYMoUQkkdgGCejNAlkhBexyTZRDyxl9L/G9BNdbchKNWk/uEBXKNwF2
znjqeApao/OjyE8WOY8fg+DKyXZOt0fLGLEu6qi7mSJ2j1KVAYt6AtpEfUgYbmNdiiJy1by530rs
R/N5eGySqczX93xR4ct1cR/c8hGChI/Iq9Z5EErItFJknLTmFghTHYVOiTvYs47ZH6/lnhvQTUI9
X/C40sMbsTDDJ1h/eq7FfE8q/toh1YywOiuxI3ZkoW8k7Zvk82vaOwcJDOC9/dnZHQnOSZzMqW4s
3o4rwBWm0XMiiIX7NUupVreANMi0WcUtAnU07iFr0wKyLctD5waeQsekS18ZXgJuUIQqi4ge/97C
BGeLEyKM6bpBuKTclkgUaksR1JPUaye/uKsloktY1UdO7pNpxJqiwk2905QzsMUgrfoXOC7B8JTN
sIaaR4cMUYUsMj5mMzd8cCEHjzGAEpb7srdEgxdtih+6BiUjl5EC89r2r1p/5Nv2Er6mJCKoOPTU
vktJ14kS4QQ6MEIXBif3vSnXzURfK3u/zymY5nQCax4LgTW4sbpNOiuzAI25kZe6ytGN0IQgzXpd
Z48TpOQ+o3Z98mE8x1aV36fA+2lkhPWDGabLMV0so/KukIASk7qmrUzM4AwodM+j1AD3D1DYEwRk
pV/zIQoZ8rRYthBO/wPc4X2Gd/zR5xd9200n7hB2h+6PaZhc1lBRuQA1F4NkeMNRG/GXNyx5/a5M
NaKDyHYpfB7hWR55TNvtdEOSF19mZfVeCp+IPMs/yXapaHmjj3NXiZj9nZ98Ahzon49dfjG8jyrM
BLdZxV2uyP112ooIzctrzafEGp7QMVz5bfyZ+LoEpohkbsq9e33yF2GIrBLU7jKpMj7PvEV9Isru
hnvWigF+WASo1WbjLpbxvyXOd/w8M212bKzPSEBI1FuUWpzNb3zzHsHlHsG0z6uHvfLpqce5BnaN
DzASkSo7MJP80Cv6osIXRJChgxh2lZoUufVuyyxFVrovnChmxhhB6Hj1iCjy0DRRUBLuDqMgUpFq
G1o2PmrbhJkJQfrta0etOmF68XKgWH/9C2iqFszglb6E3fg1zKTuNE8w8WazlPZ5faXSzzuZonwj
uVwsYVovViUysQ2yKdVstZc6SN89kfvKS00N7FVWJP3xzTReIee09vwMhEaUwPX5Ot7kywWY2eoL
BeLDQyaS75wQBxsZVVb3JEmfosWEthM26r6jA04xIbYs+vTkr5lhd0sGFf1w3hQoZ3koKLZnKTrD
43CvGfH7FvoBYorp3VVjUUDSD5NBerQKW9OirRfABXhzUv/5ie2WWqYOG5WU2+7ZjY7SskN00S0w
LgjhHlQNQEgmbUry1lQ/ArPs7NHuyyFKZIPKYRh3iC60zfqkNtrEplTgB/N37kbBJwiGd6sxoWW6
YXveATMZBknBmgdF6HbdBt4CzxpMPdxH03Lfhp/SaPw2GPl/GjUtYpA2ivzLigMnl8ww9G/TMqoE
l3VnmWD3p15EhxLi3pU8K+y15c5SbI4CMnpfgAYbtLTHluYtlO2r4QXdZmShWA/Req8kMn32UcJ3
kYoe9hra0x0wDrCb7X+/kpLMKKCm7WftRCHUVS70TEU6/hjUEjef1VVWSKm6vQgxZ1/QT29oCBhl
lMwb8vfKpj0QqVseLQviW7YKPXyP68DI3dXzHLeQ2/3JMyF4X7wYXuQqg/WFlesLzxfHAmObOvH4
gHR9/ngSw44TOr+sI85P8NpFnyldkBLudKGT2eiRGkgTILhHhicFNi2u5YHq9rj+QTo7SSffGVVl
X7ykIWHlpVtAo1Mz9G17MHg0TuJ+jY6qXIAuq5qznDQmxswCHo+8GtIC6p9LN2l+sY6TkoyzkU7i
J2YdkJroyUG4coQUkhdo4V+7smC2Obuj+G7T6ewo2iNzR7Rv7gaFyL0Vn0dXTmTZAxYA2s0JWYTT
H/YCdbZ0JlhocFoKsUHHlwXn01MKtXjsL//ox1BhtvJazk2T7zA8+sTigpIeCF5Vg4Z5jq1IHDY9
OhCVkv3sJaQQ3z/KE821pDOpEdYTnL661FzyKbVvL+J//R2uf6n4TlavOK73LujO/j9/ZDoTvfy9
jMYbnc55hMPOkNuuAVUmMJsApiU31alI0SHq4lll+ZXsbxSlqym4aN1cBmomMgk4MGWX8zG39irO
vczttulGhZcPwCYPevdBzvkAYvloMGgdDmEqIt2a4SpReXDNOdTx6A0dzZ/0Lc7i2oKCq12srMif
KDLO9wMxHWX4NtJZFhAQla1Dd4UOPzAussn1yiFO4Zp1xbv/pL5tH9RqH4+/FiXXDjy5l3RUijSa
m4/F2EEx+3xEYjqAz4JXJ1b5bYE+6tTFgH3+281PrsR4mp+WWfWk8aMkwMWp+sG5mAoACptjSnxD
05xExL4u9iDXhYxi2Lm3yTG6B9lmlE+Wkq9nCr+84EJVyqvZEkc+rDpdhfaFh+2fleXP03B2Ah0d
X4ZYi33+RQuigS97zAxQAKMbiTklc9z1AFFP4mFxQSFoEfmHq28n4PW1ORLKwG6FW54GvWYpr/2u
DKlUP9X/Ga9x8ZhlPAI889k+RJxtG5tpsVa/NyIoLWLdYPj72VRALhUqoyQCvo2Hn4LeonLaEx8l
P27/WGvoGlhmz8M1QExO5l94PNA4nOkJLAMO76LLC2UdymD0p0YQvr85lfZfxBMZE0GQIVPCI7hb
DYTQoDPc+qpANoylTO8gTNjOYUTP4a8Xx9BWf80d0WgD4BK7XEERVLr2NG+emJT8AlP8mvlOI46o
WyF8KlWCg62NmqYo8TPQRmjnXihc9rkE35+WaC4EKZTI4POFCCRMOJJIyGSG6Bq8MUEEHXk1D4Hw
ImXA18UdgCYnX8gTAKiY23zgAD3dtjZrhKRklT6IOcpBIPBcp2g8o8xOFki2tQXD66HFdBOoq78u
du9ySJE1P6d+pOjijpQxy+KgjfCdLmXwz4DpRKYlhz5AiL5nQTxoAFztfuVmPzpyAVAs/0agzoju
Dp38Gpn1H8yAS5EZSllWlVGPVLnZ7ChT5eR7FHM7ngX6zmApzGad0SxOiYeMQSSGc+TWcd1wZ0n7
XcZOkal6vkcU6EVY64c2DxtvKmiQSW3vnbqX0gNMXCXTJcjAM5T+yaLk/bTEIchrifPqOtJsoU7e
bu0qdbW10SB/i0lsTGei3JX/BaT/fMIUb8x3U9Ovw7zEWS9cT1OtPeMHNwpScThn0Jj3APpDYqDj
eudewhZ/GNEbHuc6YnxQFb1eBk8k58r0nnwUdtFLAzf3Qn94kc1D5nfWpdED8uTXE2M0hsyT7Vu/
cv2Uf0frLEkB/GvHaTB4yJAok/BfHWHaB39T6GaaYMdsVJXi1RW+8FQcKx/zQ95YWxWv8KMb4eVE
QxXQ/XUr6XBjo0jAq+oTJcI+iHj00MR4ogw/US6lDUTd/7E1uTB0q3hxiLGwDpg/R0Pj+CKGWS3m
frG5omqg71h202lM0R8N2RUptE/Bj+8DcxnS26QUe/oplB4LMc/pcRBQkTfT9AUsFTUGa66K+/ce
SGnHWB1uTDDit41q9V/OYwyHCScx7tizvLh5V05KttJoFwxtT/G71f61XiLpJ3BDQZnteJSzQxX9
Lew0psKWaKC4ukppPXTZOGVq5C+yV7aMrL5oW1V1Agq/M9WcmiHrOhHUqtD62pwWLIUWw6q9SpNy
L/KXZmvGn2IpDg3gvYgfDxo7WrX6mzYs3BAXKYU2DAnUnzCQLR2y3yMCDdwyXbk2MSYAGGW0fmuf
oQm5GbsROYcLadSUF8PteUwKbxfkqb1FNBusbBMChqjqUevypukW+EiwkAkE1qDyyxRH1txK4WgY
R+MCwAUJQKB0xYhILdr1hWCn3XK8BF18iKA2UerpmCd3woli+SQ48jTY1RZm3qK84wUkEusFCRRh
jpvFaIy5UWCy60jfhoNQ451qwlhJ1O9kyW8Sfm0E/nXoJePdEv9bfsDYhtC5t1L1Mt8oPUuWarwp
rxl/BvUkbQVBYujMTwmvMmlXsOQlh/u3jOybmR9r+Rl8pN407SMXRGpn8612Yr9kGllyOCyp4bH+
Yu9JTcOVARdmpRnlZEp7fh1SVNfYomOU8KACdKfEvr9Au8DYOlMTwp3bRTSY+ICvRzdIImiWS3rO
Qg/cQ+TBFQ/2rpgPCsEJecdTVub/hFsM5FlK4Qc0JoGCPs3kBz5ByJxmcAaDZf6vwnQXY1uYshBz
bTagNzdNb/tQpU34AaRQMgRNYTGzbKpsJOuktb0+0L3nit1/KLhk2zUvFK42jlGmVuTH0tzoFLd9
COJm7qy3QN81TI8LDlopvAxFPS17QEVX0g57Gwce9EbgdMW0I8MYubkPw2gfH31RaM67mqS6yw6I
JxUwd19oxxYjHBb7/ZZ0DyUpm9zJQR65Y9mtpvJtObtHBJHRJq3KkJTvxrLp5VdKMsN9+qS9pbRT
XkgWEdXWngwRAxbtR5cMHI+5CXXiv/ajYyV/9rjNKtVHhj4RTpATsZyUJG4KQNq82ERRvKRhBgaT
DUdCOv1lO8hFl/4zDkuxgORZR4huJY+ctQsA3MJqhMC/xl7tiYRzcsGHPQazbiCOgs4nbu0yru5y
nzudy6Rm1XDU/gu3o8ffeaTj8TiGF4TFebQkwt4re93Y+1xpdw4s4SexoqD7vYYjIEcy1QAY9mM/
s+JTpA6C5gisE/KIugLyvW3/An+kB60sRmegH1Lyhe/1lK9zfhR/fy6Mm2Pi4+/TjZvwjV0/LwAR
IODi+qqIGehbsyNUgahlmSz+HRdpXXCD4Kb7nVxzIv6F6laufXFmnlySPOigXvKfRWFWB3/nzP3d
7i3vncmg3MuHoUOT044BcfnNzOjMUYOrEXAJaUeuD4BAX6H6jxfgAxSKxNGfBS8KXAq6S5qJwIxy
bWS7Vw0t/5+aclyxrW6ulKIuqHHs8+tM9WHaLGAAXvEied4zwY4F1dKGHOdwpz5VoaJzQcnCWVO5
x0memZAumwMsqQoM6t0oslRgLOnbxjlpz6EI+B+OHGh/nFFs965A50jnibc8LlVG5pOnMs/A3cI0
DCasINHZMkL6gHS5QPIHPMe2o0duJ4v35LzUFqh3xf6pNMrTWVI5d9fu4qVrPYCekGIH/bWATjLo
LCksfVd0DNxrnhz3GEBGyiHmZTfKst0jTeFafOO7JgVOAZdu/yIZ9sXnZGbjN/aaibFfpKQDJAWE
UaGLA3daj+yJV/wL4WVhB+cS9OKEYTpaX+ywV4ce/Yel7Br25NUPFPUkSHFJQH/yx/8mX0zMvOY6
0PdPQe69VF6p8BNCMDkLSJiHXGMvVbQSAb7jeBXyDN90XgjB8IWy9gszXdk8o7nDwL7NMf4a9qTi
inwE5pho3q6pCkfBxC9k+Z7SryXFYE6NvUXWslTsjohgx6RDuvADx0xBd8It6hQVfNJLqMzhRQkG
KktKHOKlTuikTsPU0HMBBQBp+zIJXTvng3oyEmd6OrZ1tMe7SPoknpQb7Oy6LlnvlkF6OftRD/9C
0tuIuIE5l+mBJH99+4itJBWAX/uahPeDBRcuHlT5ppZTNfBW7tyasWCMWyCfd1FoxfFGTYtFBDeO
cXBLEO4BacZETM3b6kLGOBa5lot7qwD9mM867tGhC62iyoHxzlRBZrwKLVsHNWWy8jM37JC5POPT
ptbhrFzmBp5T3X9S+W3nlmBWfTMg12G88PzNeMIIrQVl1dHknJRJV58GLAT6M8KkrVl7cWiD3Mxr
nEIafG0NeRhKmr8nlhdQWHKu6ONlblUxQ8M5Og/3c7k56NVgAMdTCjQJsdfOofYhh75FWlM57b8M
9J92rB415Do7za3tvqw+nxad6Qg5csVcWAtJzaHzhgydX3FuznrTjUY+muC0i5UpRRCp5OoIoXR2
NoXgZf8hm099w3V00YcOMtkqMFMyzf8ZLH/fwSrDL8drW+/i/OwUBS7RhUBRPuyR+Wx00qE36SJ9
Jv6TQp0n/lPaLDm7sj59Lg56GqN72eJfwldBlEDxp/1xoevzgb0gne8NGGU2xwixiUrdczbXSB0b
+cEdbyGdNW48fie1yU9WDkk9M/b8W51ZpdaYLyCyfPh1RGW7WYvdebVT0A3i6E9NpBmHWAsmrtOU
kid4UU5AN4sJ0IcUfG1onz9gth3OaPrFJMz7SBhMMeC2ZDmyysjF1O81FNfPEQTjbJBCa+iT+5kO
qbogAZAP1grRi7kYkPav0gZ6DjJZxkK4rsfL+O9QrJXmsFQWdl6FMpKBGaVREF6nfwn/xITVCG7M
KsQCX1nZXs2+OiqDuWYyhH63c3XnJkr2uZ8E23C/Ec5yQnF4zo3tstCsC1Bf9uFjy2bu5YXnc5Jm
eJEPpZGFHUtX9Cj0QA1PR5yDeHtSGmxMPF2dyKftpU1lZFUZNEB8mWlzffF8fqjxfVJqlQAu6/D6
X8/IXhaEV3qBPBwcKpo45pwNK0K3pVoF0eqL9+HuZInzyr0zCFK6y3btTwkhFCW5UfXPDJwAmBIE
nuXKmKRkli/MSWKY2d2ybxPLIh8lz8qsJRyn3SW3dDqOv8x/P9EGNXA+js8IwGiSmr5pX6cfgu7r
bUat5pxmKN9wl5oh+HKihCfogkrD/WwqTD56la9unTRVmNfXIwMwjzS742l8VoL2QMrnn6r/hN/V
FWd/WOoj4zXjGSUPaYieWg19/u80U7RSP1P8nLF+LzJGQsMrScBPTR0M9PG3ZbRVGVslGVsQdpM0
gJXnqOS+aE3lFBhg60ZwKxu22ntMJzi/X465ftdBKAtIu1gIzP1NDa5EgAoyQ72NH6E9+xTND/W5
ivEylkObzLD2wyOQ7WCBdXDvdRL/eHY5qQaNRqf82U9cqBu49MLtK5Y0tLHxK5iG9cSn3E774oY/
mayHz8Up6gv4DwdE6dd6szb31sw5F5RFwlW2HMgtN4wtafLLryat6O0+353FC6tFpltqmA7hkHrg
6TnKIRhz129Mm4AwlG8+uM3xA7ez06eP/FxjTf8NMA0qxhIrxRNY2h4OuopgzVRTyuSn/PI+Uuwg
dLQPwzQLwgqn+pGZ0lp3nrECZ64U5OLEIwzKTAuQ8JXKpl0PTrMOMaaSZaikDOJl76K1v6D/688D
1U3GC5yvGAwCKX+umLU8Y/5TXgtwkhLpaRJ5FxGL4pP2jWNK87bkJ5fn4o+H/UKKLGqXvrrDYRbY
+bcwaPoq1VN9BgBMkxVQV7PPUa3vnK65zMY5Tj23Rj8Mjn03qaH5H4x5PaAPls24CXEwpLVlOnj/
fiuft7NULx6zJyzWpy8qMR8I9F/gdIrl6er4p/ZooCUnrZd1xdA6lRxiOR4VxsO4HwHbhRW3G50B
gkK7YyhHrVPyQMC2K6TghYJF0okj/+VjJ8w34c8CQrznqy0bPq2406OV0gzhJgK1VmjH3Yx/75zG
4tVHdIRfpTtIRpDoC6UgBl3kStUphKDF6+GkDEPqc91C/ulKVE4vZwAp6RgETO9zBzC48THF3MkX
BJzoNi+1gH0oa2vGcSuzseysRBmBpENBAGjwycW0WowzFISa/wNfxmBTL/wpnbbpRnU4fcL+k7J0
VmDR+bQm0r5ugYnpFgwX6L77UFdiCHtv35sbPwAUstw2qdf0RbAfwx3fsqv6zB/Ic+OtOZiF496t
SYoZ6UsvAl7PzqBVfbhQpKv7Wbk2Hhr7uFqcrF+HRb1qvIXoUUwXyqxAwOdPvcluCaYdrXTnmr16
udpiHC1KFVU7WvqQxtXy2YtUubdSNrhxFLLyQo+ttAEg1c3LgR/ocA2yM9blKFROczL9fJ/CFcG6
GltuWQ6y8MsBuljfVb76vvmqwtH8ouLoHubagl0c2EeAISaCDvohSk9fqhOggGSMXG67RFMjIMUl
PH3AV2/XwfTTi9mOexdOsLZfBpRYQzBTvNgEMHM1PoHV43tS6C8VH+zWY7jqrXAaH6G1M+XD3+A9
jXWF2j80rAIbbVE5s5/CmniAC7l9ZjspCFTxGlLJ49mby44czbXbgWU5SAoJK4X3X3R5kEV+egzz
AQZ2Oh+5X3hGxJ05OmZ+FxYjo0po7xEF8Au2TXhei7F5HMNqj/qVlyveaiQQdg1BhYsgrES7tA8m
tN+2/CMp/Ba0CvWObUJ6WU0uGUFlDs9xflUhLWl98ZtyFtf9YTr2mAsKT9NoSfXdj8dLkCVlbXv7
MXszSFREFTXa2pbItnC6rlZ5p3DFO6/PObAYbnnIoh9J2ELpwG9LMRcsWZhEU+jbvLu46Tf9z/Ty
UnGDhGT+MlwiPrsPCRFZ0zDSF1KRIdqenB9bGnjecqZ+0WkJfz53fWmA6S0Co6FpR/zLMX5UmHCN
c/5XwXPaEapeVOv8c0WXM9qPNbo/M3xOqSN9G4Pv38keu3t3mcSk7GkkhxUabyeYE7zSSU7mSBrs
wOU+dKGmbAEIqHOos2oSJRhFw0ls8O2TPqq3BE3FPVu/WzSFwFIUq1cPPIPkLLIviNnc9FtDjx7U
gVRPZ12GpCZN4BqjxXMnOVgwMrsAzoNCFJ96gmgBekLGrDhxhQu9ke5GZb8wpRhS06r5xREcIMQ9
YOjV/rH8eQD9BuNG/ZhFV6UYrz9F9wiudnyrkI//f6HqginUL+waLeZL3DALCAY3+44Hwvh/ihi2
EuY+bnVu9M8kGseAfgSvtEMiO6nuTK9xZa/GRiXQmEX5DBrJO5VPn6lvR2R/pFKkbQke6qGhssPu
xdwuwuo8s9xi5IAU+BmZwbWmTT/+3W8q2BR/7V90+U6RgzrsDWKu3ul5RbJ2vyvgyttRfQV888/b
lLSlnQBbHuFam5KrXd8u9FqrghwRxXhveVTAbArKzZTXqOUtme2ImPiAwE1UMeemy88jqBEiGdmo
b4T6hWdOzrnOipGYdIYevt69Qxaung+uSI4IeP7V2HWTqpzFUX1VUORON6d8CEILbssuJm+vmtCz
9gFtfvucyfIjQSRniW7o9zMBDtUpwJShpp9uzAykSD+bWjtBl6YEcLuUhl3qrpOdI/46dICqDGNz
er3V1T7C/r6xL1SaLBVWgieDaFAE3OKqssxVMuI6RnpZKcMbQmtixnfdrs3tzoemHFP34vNc9Y8L
2N5GpgXbfUuuZ1/Eh6vH5QdgvAb7c/1QOj6CPvprTyBnvsotuMPZqhVlEYz8+FVPiK4gamaJZd6o
QpSECDETMv6mkq0DBB/5I0D6GSoCz906wxSQmOAj/l1lUQDQZPV8Ne5Tga8E7V4eKtubjTJfhDB1
YV1v3Js5MN26TJ0Lqgli2V2q5CmQW4ZmTIxXl6iU1VWH0lFkaB4pW2KusAFvyz68HcZ6e+i0U/zo
usdF4Z+QwXbIOSDSUDPr5O9S+JqwWGrqm4w7LlYjNfQmZEpl55MiIwAQNXA1lNidbCbvHkSx0bwF
Yr3M3olfu35cowVEyrDTjUDZBmkobFHhq7HHIgoLW3i3PZdhRNOLIFuMQzHFTmDTd+H4vgZFrDUj
IQFMikeWZJBrvGGatdqqX9Nrso4utMD6xPqP4/1UPEToSL13TlF9mS5MsWpbNWVk6/qDfv2HG0UJ
waX+FFgPAEyvXVw/FOMbh0al1rY1KhVissmDytH4MHPItMKTz348Cvd7JDfBZfkTnX39x0j9At3v
H1qZ0nxA4bmyqKliu6jR00de3+gEdfyLD+Kmj1GZ7dx5elTIX4/OICUla56on9CDEjqZKNb4fzCU
C4eJRz++y+h/Afjt9z22j83zaSEP0bT8ycG495T48E1RAv9ox4gRMEr6ykDm9BKxr+yc5DSYcTwX
j7pesQNjpPnITB3qk25zOT/blQ8e165WAECDigtmEzHxTdKlsqz3V3m6Q/3ehEyBkAYXQkSEoMSs
RnQjpn+E7vZK3n5H4MMFuaXxGDGb9z0vogZWhPcM+cbikhy3+4+dbcIxHVwM35ZvQmxkbrftWyBG
wpvE+RrwyiL5CLcKh1NKLXJwuBbsyAUx3i2noYzDc+3mV/mAS+mcU8XK4FyzUif2wGMjZFfjn97m
21PvO6lpApdCZmdzRbAV26D7lKlfmVsM59U87v9DMS8BshhSL3MLSoLa3XFO+PQRT5IC3v0AnMkJ
U3ibaGa4SNcLj4j8eX5vRtsGzznwtdGa7L/cp76ZgvCc4N3va9rSubYyJJzuMgq55caOlJ/sjoTz
9JCUBVJ3o/Pt1VDGQZXUR6X/2Q+6zHejYKXRVC21ik8DVSU23IgEx3Bu/LhEDdlSS65ST0rMMcTq
Non5NrJBbYm7P1lcz/d1qnM0cy96/Xv8e1LA2bDuzzHLf25s5uZI8pqkzccdFoRRm/BJQAYCAFXK
3oTPHaz+pKY3Cbymz3IGnJoW1n5ElNMHOxgRy9n6KAdvTHdNk12YCPsUYpZhdWhNt4RJD0isMoO3
+uSNXfAGBTBRyOmm8i9rVFgGsYe1rWHd8SORwppUE5aYcdqN8BzHDEBhh08+O90AtC7nhdIh1rh4
YOYJFSVwST/JwPzHitQYHzepanM3EWb++9vu5douWqHgZZQofsPnejAQ/k0MHDHA/LBcTRc+1slx
DCbMP/kjMdR0q7GhySucVFsCQF+Y+8f1gzrCEj5kZaq8WOdo5pPuLWYfjbVXu3TlleuEjJX+73bz
7Mkx6yc6SypUCz+Y+U5Znph7Jg5ybPzXw2qIOQRHSQ+NTOrZq9iigelQwHmEtUm6d0ojK1upyyL1
Bx+kCjnO3M96EVRfryWE8kwkJCwo/1axc+LI7MNLoEuP7/3RzhhymtdLV5t6R6qNDagZt6FjWEtz
p6ksfih2Zk0ytOhKrzkFqq94MEtH0QkHFQL5QfCGK+sjqvB1FhgcZ/z6He8LaqvJ5ceSsaSywjUV
xLzxuo0VAf4NnUSLYhcWLJq1MZX0XgNdcNoNtjVc5kTrADJ2dZRYld0QNHXlE8Io+re1PeesCv/J
N4H7djjJAu80yyXjfA14iYCSfisRQDjYT2i0WXf7T2juo8leXso1tr1mB5WW7L5N0oSW81b5C4LC
Ey+HECRGGQ0V+UFwFV2W+RIA7OC2nEp5t1nfS/n2FLS7kxEOl3JXyoP1REAW4OUca8+6QFlR+KnL
50Kz0ksD28uFItPE/gptfN0hqz7PUen5YPGAT5fYcFk8JmEr/Ejjh2j6ctmIA1XPHS9qJYnjMEw9
bGHzKNPj72z3dGuCMJhlljtvQw5s6pCKyFH+q3QkKg7sMYZjHdHSVmmRXc9K0qYb3eXpfACkzIif
tHe3iJ1WjPFvYltpr1d7FLvQTH9Gn86BGaTf+F1KW4AGRM6FN6wVCoCiXIl+ToxGMotfOpYC+GTn
1uo10mbbE2TIZ+EXQVNBp/XnQTOHYqNbYV2Mfz3LDK0pDjx80qiD792OHWnFxfTUHBgpwRAfD8Tb
wWv9ohwcsWzJ2vJYIR+hrEVUTW8qmqA5swI8lUtPhLH3i5nXmjiYhu/WQEcu9m9kQOVxU0mArTrt
aa7PWAJZSbA6zWxjFFuWmjdUsEO/qVYyHjIY6Qpl50CYvUMrB97BbZ4Ee6F6xIT24bzwPBr6JR1p
TI59k62+H2PEG+iBL9RYT60gUXVPGlmRjbnwI2VpmH4gKnmRjL/++qu33K8lJzGKg3eUlhlbeJ3n
Mdu+6Rb8gkH9m4m4MRAly74q+wRuaRMeqLUQnOxe5Atx4eYn6NZYLyl3aqEUvSvr8HQjmPnGt8XW
EC7kICp6JVtAbmZHitEOQLzaegL2hlEIhpmKX/Uk/aLrxpCj3p75KhDz4ayg3wPKpV/9PIa1i7df
moKDWLmMuQeo/e9qyPCvNGdlXFAA2pM00vnmNK4fFVxKnmjiaSwNK4Fvv851/9fd3ko8xJB61Bof
/0jI+P8ZJGtVHEQ5wrrw43LonDsAWHvxQFCAY9zTeF3suK1jUIAuq/EFNvS9qoG0lZJVyGYrK3CB
1GUCVx6zm7NVA37eePnctmSW2uNqjrHwAEPdtPx5ztBGhV3iRfiR2yjEvOTZby3dfYmjDkj+f1PX
zzUguiziN2PEKwwMK51VPEpwoAxVUNO8Faicw1fUd8Hzk01IU0mKQ4SMqJS+whFgNAmvV7811pWZ
WUzUMHkgCmwGzFazWAtlyg4JN3tVUFwWVv/d4V+3rYbp1Ovp4fioG9EhKSPJZpS+JbCVW4zFtXCY
XnRTZEhDg3+ISpIq5IdTVmmz/w4P2Ah4U+4PG4anCJ28eFgwQT7nyijwN0ZC3g4c5rNsQvQlV9Ma
DcAF0vKM6wsRKZV9EfsfM4OsjOzyNpp107wgS2GLshXuxNrWDvOhg4P4RdF1PTuxN3t7N1gk8H47
R9dODTGNdTIDnEy5EAWef20S4X+TByiJixtXVoUVi/q2qWgm8znATUXT0jZUxgf5LztnesDKxfJr
6bvsRh89l1d2M2yjWbCGm/ijT3l47/V88rzuARuPz5rX0LcRk8KlZAe6PsVFUyi1PpNZ2NgvHkQR
VDKViXNUj3rV2ax/uvxqwIWMFrNS5sKd3uiT8DJB8dWS84HN2tC8ciS5JxP+4qydKRnLY9urEMnz
QOa1F+6TCiRjp4OaC9mJJujMggERJtWkq/fQoCe9svey3mo6u3KWFqRSTRrYx2H0cMZB7uywUU24
DM0hScnlVqRFErLvjyRWuOGH+2FVDexZuZ+JorTtOifv2a/3YF74O3NXq5y2IOXk4+jWtJlWZO7g
sFU0sc4yUUJL+gLN9ylci2fMpMU/DUbO5mQOpQJw11Z9QH66A6wkweiHQyPZzVPolUs9rtjksHBL
1CZk33tmwmqI7NHcqUP0LYGQ1m5P39e/EP1qBjyhRStwq6b/6/4RY8UnnXOUSpvjI4L3xDXHA/FD
u20OSm5cUV3avb2bbqffP3t4sUc+YJR+wxKFbuHRmGBEWyAsYNdBXveCfoTTBpGaq5l4feGgiQ2T
HvAgbROPtKJpAaBJoBHJIi+CP8YY0grOfX0OWmI8dQZCbE5/XCqekpBnDrHXbOJ3wZp+kjBPay6x
VLFbhsDDzBG/Ubv8JsuUWBBDUtcTaBqJZ68VeyhUL2c0awom4AulEx8rmMIB5wXplfJuLJtxMRPM
26ChyjVbAMA6My9EiPD3MPzNNMOF1+9CaNpgPh8LOHt9oPDr5dffBuMbEwqeYwX745akGgwARFbg
KJLDJ4VHbF1/Y2rr4G19+D3AtCXgOgDwlvbLJQqBZsnS5B6ILxA+XzmnsiOdkdCErB7/qVcWHCz7
XJuy/BrHIstiIfU0qIaleESsJZ1vTaZ6j6KyeW6EoX5fQDdRx6tD95M3GtZcCcDvj7TbpHdR+Gnl
sM8zAh4DyV1qH13qEzXT4AeKAISZptonum1644vpIfatErq8vO9T3N0hg9sqSXhvb9tcRAubAqIw
zEJ3cV/wUPrLPr7++LSL1QXGe11uCf+PeG+uH675x3hqTsl6qLAr9pPV4fKZzpj8qpAcOw3AFlDV
hI4hddLo5I3a3D+JvRast5HMDIJka5u34iOu+2n+9cyXN5m/KUMl91ahCAE4gvkZjw+tunT3zEBy
wXsFGvfCQAUIH98cL0YZaZMQCHccmDIrEsdhtEuR6Nuj7Zu+L79xeKy7OCU1cxVE0M/dt/CqCInd
KgZQihOxEEq334XXkEKSn+ctd24UjtPCskT2D+eqJqgDFGLnoeboW8Mui3tbsUjlw1unD6zki9F+
vE0XVrMELaUBptau8JKUcQgEAFvaQMXAWJEgv5aA5Q6V48BWAqqwjI90bwEPqwEfanO2s8TkAdAQ
VJ4or/MR3U0h4mKA91DvDvC0fZ3TU33iddx2cuip9hxu2S0Ser9ztPaJEHkglg5OtuxzyW1mFaCj
UlAIJjoE92ZnasPA8Pqy6srFaDZjRl+uA+nclxAi8y9ERZabVaHqjE1/iPoGLEifPujhXgYJ9+Oz
CXSKqNhaneqdPoF2oamKKaVQbhBVJAZRS6SPbxdatkCu8GyVRiy/CE4iwgk2ipmSTg4IZMoIMdgK
8FwuEYK+/qjOwbMTOR9PLzyTpSDevn9qNjbORyAG8MkDQRw3+bbxN5yfqpxpD3KUaKzT6zzaWimw
z+duNRXsz6NC/2OO3iGg9UpXSQqEO0ltH9FZPCSqthLrnK3Ea7lbcCl8mStQcRf/EHh8V0I+VRNb
DIioZMyH5nX46WFIf7qJoPISyskYQSQQ1bi6Gs9lpLbvxYaDpxzSnUUf4lZmA7ywyqIPc7G7HFfC
Vv5yWTPQ1cmBjyXcFBEI3DglPgMm8qlP7eHDxYRZgEINto9avNVpPnxR34fJgs9Ohpw8msBc4uHn
//ei3HtVLysrZ2Gziu+t3YwY4XomzKo0C2tALcejEYajaBBxYham9pJWpBetQt2wX78a9EBOceEK
ZqBnlCsx20s1yikGultQGkZr9SrmKHXmth4hwJC77KFynkoBCBAtae6dZMdnm0l2ee8WNtEA057p
RSb7gBrEn5tFERSEMTdPuSXm1wDu9bHpVmqHLnM5Z4pJYx2J4/n7jM7nA1cGzvq/QBarUe9rzt5o
I6sw75DUOc0mto/+tLGarRISFA4QnP0Nx1/ENghUsvWuqWrWvzfPVSIY0NSb8Wu38qLLnSfHAH73
TGqJ082nLpz/t3P676d/0nOWKqcPA8EZ7q5Q2ViciZtG14ESHY5W0x4IzUWc6L6T89rxYHDaAMqe
+vW8x9o7O4X4RE2+LLqcSZL2Jc67A2r4b1btGSNMk1/l+zwvCfdzpI0aXSjT109ViLKnPuY3FPou
xufSQYKNkrQILBMk6K8m8Ts14llOWX/eI6U3iMiBGVKfnquTep94JdZRSn9ZtMz48XzT7EHtwPVc
HAw9sMYRnsGRCrFJxRD0SliHPoE/xM3a0MYM1YDpzSp2TUVi744neIj/KKIxARouh6+RwFVzDV0o
/HYemdEKToVsgaaj16jpS+ffFmzDQb96K8t9i4/EhiqcacG436iPTGpx7jl8qszT+BJK9movjYjd
3kcZyCl6N27EmdD5J6/GCILt4idjcSH8xZlHfSUttvL2H97lnULZdIkc9403kNnnnzR15TTwv5hg
uHzZ6BJeG3A5DSCsyjQC0oI4yKGrA1RcKMMixNku/3gFqcF2ixWj5QrbgWOXjuFhsBn4KQ2g13hV
SBzaDoADlkerr6jU07Pm61cONacvXvZbrlSVsiHUU/IwG4e+ysy/iK6LI0jQs+RUJM96/LXeSIdv
GAzPvQiiN12SrmNaeULC167k1P6y7674PTSuqsKvM5Sx5LVwRHzoG+MWmEb2cXF4HW/l5kNNP2kD
B/tLg0YjYkAdodqKgn/E+d+946BGgLJC8GBhS/l9Nhl6bI0b97gZeO6u+tJXtQqSrnSs+unR3ZKO
UqGtIoDSk17quJ4iiImg+n9qVMoMI+2LPUo1Nrhfwuu2pjFp1w07qydJpA+eK8yeYTcugGKQtJUa
Wvvz8FBITQf4AaHxWuaC2W8t7e3MZJgtT62gDqqjoNqZD3dpMfRt4Q51wpAxFSCyRpYW9twqUkzi
6MPax8VbpMdhkanupQv6uDU69pEGFc9GbYP5/Sn57uYwxsdIJH4k5zHnfmptUC1r8CdAzUn7aC/1
6YuyOHqrrOmqzwY9vvEBSywO82vMbpBsJC4MPlPJBp9bp3fQpzTppy+9yuXLaOMOC3989uMM+IKq
Q5st3Joy+DvsIw+75T3ckezwM0AVO8e4rzufkqKGPgMy40S2j7u6BTYpG9AJJP/euQNTyr4qVCJ6
kM8AZrRDawgxIOsUrXVs8sPuGoC5AcE0x1LF9dZCOq59NrB5Xob5hPI3z5Ri81kshTzInNiggE66
T6xFx6956sQAIHnW/yYKF+qADHS+K7N2OWUxAI+rwuAENouBrwyM8ireFH06vGxWvgt3nCHf43h1
VI3KU88Mxy+7xGxjTh+T+IG73qkqCC14o/4RRtTpYKFsel/C1qnGMril1FF44YEPAJorKgMZzX3x
O2JHxnoaTmx/Cek0HG0FW5m/6BWkNn3h2Fks0PYj2ZhOXLtjZOvrFJGXNK9h7N69y0HRF5aWxutb
DK1wTSoKQp/Zs6y+TI2iSXZ+xxAyNZO33dJ7k4ogrQGU4kGC+4Ta6Qr4gdMkZ7GN6HOJm0Xazapp
yTXSs7Cy+jrJ+Sh6CtPmwM2YMkEFSLuEsA5WLAd3uvhvx79wk0mUVP/8bC1wI7s9LnRhlvYZ4mqR
Jy+jD82xYluzSeApRJwgBEK/04c6c8Bpa5tPP0n/PI4XFFuPITIzcjFk3c7HsDFNHaZTxgBtUYYK
Z81wkgLW06ad0IXHdOYkichK4xSLkRYdzg5upjHHxdK1hNTtGnPE+mg7K9quZeeJf0RDApLIZDKa
tInytbV1B090AkOh3vTPoLpAcSlnQA7WvsjFwZ2A59qKF0Eh2r9igHAs7mJxwrUq5i30k+d1MGLa
ajWyoXf1OYwxOMUUaoO0yy/lNCjQkJAkJoTb9wCXyLedCaZkUAazKOlCeIOSC488QCKDwkOpMl0d
ABoLol/uMJj9Nb2DTzZahEmXgUHFN3OtPnFrttz06szFodCHeg+4poIIvZvW6a4Gib/WKb6RGsFP
sqrh6GY8qxbx97eoaFnAci1LtClM4Lbl+LoVzAhhg7OsLvESTxs+ROxEGMiLamiUbE3kiWw/70Ne
fUnHoAeICGNS5pO9tnE4NYTo87k6+Ytcl29tWicHzTEVKNSWX3WfxylxEtJa/kHxqEr5ZOiTJdUP
PDbFZcJZa0X4LIo7+0yQf/OPyik7N1WSgLisYpXmGoed9C7hImh0RbcH+I7GGLYhzVqF4vDgjxH8
iI/B3K5+vewlqW0ptu5qq9fawoc7xLv3IcE3i3AWBwVt2RJcjmeFmBHgtkHzY3N5KSyuc6hqxoCj
Njn1OLcYyNjPaKfrYrpsNMVfsmZe5pf/hSkhZWysDZfrRv4nDRS2AmSASH/WDZyghOysuiZ/tkin
BcIyuOwj9eUgcAfqzJJkzTemPl/cE3ZHzF2LtjdLZUsV+nCRNJUFWFXm8r+lrnG+eEId7vOmbMy9
fPi0rnUeK3+Un0w1aPYyB18SbvjzoI5i7pfKWHB2fkiDil7Hx38dYCt5Ws8woPIBMOod+uhVhdbI
ZKE5w6I6fGl5heJC+6DfhnZW00ECl3KO3R5uDqRyp8LU1gH1Dp67+8/sK2uxd+AUQDEYOqNpzOis
dPTaImabw1k/f89e4NGz6MS3l+Ardb8MTGi/MJie1um1imFjNYMZ0999Vy7yjOvkAS1d23NiYSca
7TIWxgZ2zZXXBQKQws2NhpYKvnrJmjvRlbooTDnMlpbTsG1ID9e1wwjJzYDeWsV+UQu7iYbvaYdE
fywgYAunmxFZqeFmNuhgLKrKAEIeZnf2yyMpPjJJrNiQ+Dsz4EiO8j3kWtPkbB31gjQPVjmOQWzy
seBWCasWN5HusTv+oTgkungzRltOsDy5CTzyt0QyrF6FmIOrj8cHKk1asJJlPay0SncXzc663ByV
KOOLe3BH1uiFArE7H+/DqsrlguRTqQ7txBsUIuUisZhNPXqqO3nNxrvj9KD30IQuQC/BaLwqyXbn
j2swh8pBhu9lQ7X99CYlmpeWs/ez4/j1x7zL+ZsNT3B3JKnfMt/6gI6go5DxDV2OoQbzmaxRIcGt
jSJsLzvNHQLyj1evuGyoWrIT/CZJe3COB+1Afuhi2RDpmT+OetRemB42rFyMFN/0guZm9OSDejej
jCX4dSjWBZZ6AkjDyG0TsZml0IRdUyWy3JV1f5kxxj0ZS0O+ZZHRuctcDmlOo3iruf4VgEKQodgn
pQeKTGnpKYcBxpZl+4mWIpN3u1xq1fyTaH5k/YU0zwc+m242WQcuBL0KGmzwLGdOkD+HkP2QRq9v
gpE4KxB6cek41WZ7EHFfzFv1fhQoV61EWPl4jGKyU0Ci2PbyVly2j5tmKJcKDl5tnOHWrRgj86zr
A/r0TDlxJDSckk1FBZuV92v4dh9g/lm5tIi6VrSBXR30sNFfyHyEj47so9Qlo+xt6JwsIxCyf6hs
hwYfyGoukLbFyB2Y6aDjeJlGJ2or0nukJfseGCEF2IBI7Xkl0jkgyYazOWDDLmUbKAtjwDqB8hDk
+T9bskeJh2tqFKeLWs409/CnjyFsRWLYfdaAHKs+oSljpYPe9RCAmNVwc/csv0qwNWfthi7nASGr
7zo81VBBYnabJxVAeB6Xq/Fou3vSleviLQS4mCgGQZDwbL09qtGEkQbuvxZaNz90KX3c9naFwmJd
1gFQn6IZ4kjSK7RJDqTyeopT1XXQzrkCFrKFEuHcLwbiaFLMG5910TtxiWSSJhBLqPrZJAgqYwUq
ZzxqtLLNyqDNBegPRrbwm9FMkfWkfK1hdrc7duU7QTKfQVae8MnceOvNEj1G4EWwA+plLeTeGoNq
RRYsg5OAvehR1prgtA6QZOC4JsHtFpKoG3g6Y7ahXR4Elk4KBl/iRYZ0evJfLnS19/Y4JEdfCrYW
ZW7XHX/8p1yS84+Zq1z3HXg2cZTKrnAve7qYDf/dqb5yV3jL9OO7PAuMzznLHRx7sWRZm5Prx2ta
s2T9V07FJkZeqdVkPF6/Lk5AaYtN+iZK+Gpmgmjswx9MpzQ21/m3KV31+OdYYs/v04JtLskcznp4
OpPLPp0mpEUhGaDvvptzYI2xzJso34KnqUNo1tL2P6NufHuNCCndhYhROxeHxpk9GUrP3y6mRrvs
PggladsgUgUN5jUDGYtjYrRX4lhov7enNcEWBKXeT1XgeQ90hGoPSgtKqP2rB5CSPl/h250NeFMG
dKoCLTckxR0W4Vilf1Y4Icbf3NlHkHIhb8CHw/twEIMlhVgIQISUciMgayVLGcpFYWZ6zO5N+Xd9
9S/D2MibtXNg0FPbb2paJMbTbSvGfVHyh83PoQmEAYKPwaN9z1C2N87VK/42hpJOSDmhg0CgF9wa
5hkX9rqQ0O7EUTR+Ap2XSFVu7btDyeK1xmSOKry1gbGmZZ6WE6onl+HaxJB8q5h44pspzKTDb9at
M/7xFsfGdJ+YQXVnryrJS1nJ8JLicd9vKA5Gn+e/RJ2JpLKtHFx63GszLNYiuv85wi0YTGALUDY8
4rmTwJXfCFAHuw9AAa7WE422ulS/GHRBu4ATDr+WBDQfci+Zw+XT9J5TOxZJMQQio5fq39n51ViG
0T90MH3Usw3JienEfKT/Eq2stuxBY9BUBrbwbIfsxhHIQ2pId6PonhFiyLsT6aDIelMxwpoMpNmK
W0aRsYaNXgHy5catAQigQ6O+seXYmuRm2naJ7CsYk41CEFiYJRluyj6TO9gzlf1j7dQk55+PIlZa
ENLyNwHVQGI1oH9LT9MUsL43SBiu26G+Myfy1RmXa5hQJp+LPWvhizwuHcAd9H28bUW7qYFUmWq7
eUNmOmc7BYAWt6PkyjnoveYueyR/sLsatN+LqaCFt3pVMlfuZWCH2TtYBeKaSo8riHbAbfSG0EFs
v7D6vkjw55ps9ceok6WXF9FWzJft9Vf5fdnMypsW9qt0KGiSsSasGEr3brnZB17h00y7r/7C3EoB
eULgzsIEWeeBWWH8x9XTYLzNbAJhs7JAq4AjUstu1/vlQblR+q1akTGHgBca2E8mJox3QdHnIBOv
/ArgvtGf2nLc+KRn9JpsTIGU3b4IzsT3zoMpDmgGvrxxwFC0P8fmnFG4EyAaypNUs8CwzBV4ztvk
a0s3HJy/yXYCfaTIfhvoUnTxvHk70+sWygRr8Ep+9L8yxnypaBn+7kCTVy6W/I3hJK6L9jkgp8LQ
vNvtbJOrM2tcXftNI7FwT33KLF3IxpMsqfhZgAtaYy9D4EO5xF9xfOp5cHpFKIi3XCCrjkhAQ/bK
E8BL27+tSEAvxyLh6+t1xJjnn7BLSJuaPHi4TrZi63fLD511xImohN8gdinUR/aDu3KDDohTE14A
8Jm1rMpVn0kf9UpGLyJaC6vW18G7PXmAKp9f+kdB4Dg0CyPvYyfkc0SbbcrG94t/4ftUzjXDPvUy
yHNtnfpMAhS0FnbYRDsxtUldE/2oPi/8cOYEUnBVCpqE+JhGobWeoPlk+7SRuY4yWmLAM8X/r58S
0N5i8ISsVRhGg5vKY91rqkrQ0xXTqHItbErkHYACPIBlrgHL8VzWtphd8ov+FFQKVRzQacfWgBbw
F7T9A27BpLsOK0mLKXuC2fT4pqR+xIb8SUK9geaOFB+uVd4vo98i4SPDmxY9dTgdtO/YUIZqfI6J
zO9EZrZ7Nq5Kr85PXI8vpsGWM7JPaP/viLoP7mzb0g/4/SK6PfYdS8OfD3DhcQuwVZqElWlH9NMx
phTRRB4dkj7tXS+V2ef+TbtJ+JFscIp05scIR2S+36r6/0nRV7mHpQY0hVUmbMiUSIQs2r7hgmUm
wQ24AcPxb7xnsIn8NafF0LfRv+YJlKwlRN5mvfeTSAONr5X3Iwk32MCV54xmPavuK/1nxrnXupce
fi04ocO6rX8AQePtKy8Xni1Xe6JqM6mLLaa8OOWZ3MyHwpzyEqvj99kXUH3ua4BXmULM28l5Xn6w
3NQzCoDG6WRZS4jR5xD9oAiZM3ncFwpSJ7fcpHhABg4FQyXKzt9H15TTliXwa3UO3YBemnIIDtlT
HnAJbMHrId4Gl9zy0gnkUPdhmZaGwk9HY67CWr6sCJTl61fMM/Xd2JpojXbzsXR7gdfGpdjdr/di
VysuaPxvh/Oa6yeEytsPbouz+26bnOYY48FdkGYEejPrRcLhJlE6NU2cnv8Jf/3vH554nVZYv+Lu
l0iOzC1oIpRpc+YndMhC9VZSe27k9kSAvrOzh4S1ojEqJ1LgFhya3/mnDzdVgynuK3OGH4+pa/tz
3GgYEC7kj4Ksgv/3DvgMeDGpmdsnhAXAgU5jAw8xo44Ykk+GvD3WonKMTVkxuZPQmLsACvPzLHFQ
5cGC7Ft7FVeSHEWG/H89I1WTOsumuvR30uN7984YkF099TRt3Cws5aXZ7vW2z7sFEpQBvVdUYk4R
TgiDFzYt4z7x5Om/a2lhcYG/XpYY79bVaKWMx0kZvbDLUw1ruuZb94K/miM8Ececfj8X1gouecXb
WLASHT5HbSFjKPF/H3lW75CX8P3POtGb8WAlmvb7jdGqutaJpcMI4MRa+iRd42Q49hqKBHrbn5/8
FhifSpaQ1XZg7D5PNf7c2W2/EPYR7NEYgWZpCiGgJd+9bCj4AEhwexutc07v0Q+39nOANzlHFWFI
Yiec9MYJ8T1I7u8t0NJtVui5eJVZFFVXNJIU5fy86ltBww4yGVrop9nPCy0QAXbyMkhMjoxL4KTp
l5n/FGgKFficBWf8J5ljYTICO/QiLNQ+sA9TPyBcGXCMZOPYefRAajbU/eK5eojVtMJNBx0+RR66
u4fj5939eMl6SMP6FJ3aLG1U49LsxyYrwiBgX4fwoFh7mFj3TKTDD0dNtzIZDB/mZO7CHRMZY5VC
6R8p1SuHmX2PkP2/Hg8adzW7mi1jIy8Q/nsLuddDA176XqXN8a/WrTw7Z7foxnNY4RD8tJPF8Khf
pk1FVvyMFz1hA4ijlEsVcyl8ByXgyj85chtObecxTBkrf8hxGYiOgZrzYrXu3foy2NFcB+nSvTCX
P7YaSsspL5ch1W4/xGdhBAmO0dK6NxiiBMZfNwLj+kuEo9vbWdBzNJH5OsRCi3n3yVkPPqg7EIq/
lIwUuGUO3ApzByhqu++3VgMFYSqTiVu8LdDWi7CIgAl8vtc8DWYUkSwqhqs4/SAGJuXoVtbI6O92
gajn4PYFclpEvAwd/wWOqrcCG3S9pg8DHNo/GbRdj40UwZ7O19h6onMCChn8WXAp3rRnSVTBPIeC
t34m4MssUSqeqT4Vrl+hzXmjAlJugGuJfRNApM/pj9MpvGaHFt07Xw2FRKi7b99q+DF8L9TOrN+e
LnCBt4UoSvvtLtOiKerS/OeO2IYEohR0NrIpDAr+qCwVdMFKafvVprdfyNnkLu0RDeUvVYYlaycq
vRp43737cvLqhY1g0Iru1+oZ5eH3bMyhs59taGSJJw0GNjIkBdCb+KbynQkIzF5J1kStFr2jjn78
2xmaJYvywQ3ep9sW4m/eS1aFdNyzUrAcc7URpGh0B9+RdSHcKvBIGP33jTlxWenA7lV+Ub9uoS9F
PHAhvsgu8UjhBcyx8rUAZKwl6MZFPY7Riu4d0C58ck10wIbRxWSTWR0P3REs8N4Drmp3xm8ZN6oF
EZE6jaQEIxQ2ckZjko9S7SgO4kM22OG6AYuw/4ExFGsQAixLXPCMq1JfeU0iYlOpd+GjU96G3KMD
CpACIU7h2xyRtdLqNkC9eDsqep34lw/a2TeT+832PJRUqdzMDRYGFtJVLCynMObfoQpiTPFeaVtw
Zy1hKYZyZVST5IIx0kPVoG1jbC5uW4mA3qBE+LQQ9LB9GjCBGh6vsySUHiuijGEF0y90vajNZV5B
TT6Cqil2Zj3WZVB2HCTxP7qyaoGBvj6S6ku3T4bBb6goQb9Rc5ugmLwqDvZUuBrB6iuWDdPYqO/a
cKlZ8w59UC9lQsh4EyU1Aw9sw1E0ZRTv577xdiwKsYcDn0b4JNINC1UbOlUPSUOewI/0s8twSx/i
2DzkhwaFC4lS/AzlNmqgnpc0XPLWW7X6bNnPbJgjimjcOTaPmqh8EajJhwN5tQRcMzz0GG81otk7
Sddl07NQqWD3pRbVZ3w6zzlB3eLnUNRbXTywRoytShFEaYPHigAExiWhGqZKMlTAWKP6sgR4y6cE
9SO/TMhjm8Fo1OqgmSwuEZr5Z8/eI58XHxJxdZxYzWBdqbox6WwJBokGBkN71g8IyS6bHiRQeLOT
i3FT4c4BVymTzjBFTfB9/KVesvgpmRYdd3LojAOJxjGCEWCbJ+AzuiJ7Wn4HbrRn+jqgYocSYy6B
bq7K4ETS3p1+VZwEbGG8mAKLwKEfBd806Pujn/pmgHtGjNXMKle6KmFQXdGT5zDs9Rnmc/3qhucW
Zs4f0eP3n7qI9pV/qAoijI83XWbEf1vChTIdQb+Sdw52y37I1vHaW90hBJiLzIu+O49nUFw53X+h
XaXjMzSrWuGt2XFsBGZ9ibVJFdxUxDp0A+m/kuwLwmBqlJzbfirPZNZljpgPWEWF0qhEOrHtPdKn
hknHyjvy5yHZ3sO09iP5S9TJUnWtx2zuSpwE+nh2tkUVm5gKnp7/UqfKivES+zI97j9/j/MCLQq8
QGOWqEsQ6TSCkKzrq4x2Mcu4Vy1dSnt0dQS6AJ2DbM5qlAXAKl/kBKiRke1yP/lcS2MCEu6EIo1F
NlLWbVycnDHnkijavQm/ckUDWRfMHnLnvEZe2Bp4bSgvhZnPVewFZF2X0IbCcHMGDwL5ObVefXMM
VHvzjt/v5VDxwTXLhwdkhrSNtmxoN5PxlV749eCadADGdjouESFSy/LRwCKl5FpSmeAfX6/PWQpS
abrMsjgTfCga0VmCRbK4WBtHvy4vjOHt6tm/gCjyd9yYJkDX4JN+atfGAu2J4MBAFdy4txKF5Uow
Xm6ydNM2+CY38K2h0ZO9Pz8pru1t+RiTjYLldpRT7SiWie90+uVd10CfIZ2ow5cEOVUg07WUHwtw
K81/F8bh8bu1ZsyxT2tNwn6r5TizhLCxpHfLo58gXFaUeRb7oKF3h0z8WU/obYJXi/zqLCKxZn/b
azJArHHwT8sOsF/LdMLCd1+CUswssu51XE6uAo65Tb7SndOOX/wfDt+hoG5/iaatHnLLj8yS/q9V
yfliHH3JHlvv9ta2ZpztjRNwK/dKZQraL3CZr76uHxFAUgKTCb8tRdi0Klj2ON0ms9Fi0+ZmTN3G
IEqUDodJZTVL3P2KXYUm4MTznF4Ee65J7vX2aqDDGuhDh2Ql2MHUTOD2nc4uNLZPP8J5JVIIBo8H
w46IsvLVfQb6W8ZN0tHgQcpKqzcLbE8U9STLEEiCFcTPolzebTp9TEIXojjCE37SLykdpbX0KSor
cagqYPq0i9Iso70daS7/TR78s70LbA1BE5ClMNKHWLg3dMUJjSs/xfK77btI4Ijv9uS+Sj3ry3o3
h1jWO9RJacMKlYcrQXQAOuHeLwl3eE7wlN1oP2LqFqHoWTJjattM5A3xLBTSh4YsT2ARXQTg+O3E
HsXgZ3NCabxN/AJkT1rCGFtken+6kLAjg75uVOSNE0mg+daugNW1iLOiCUiVL2IXcv9o4XDBjEyQ
qAgJ09d0FGl3OVx+hhA9THu1lXtEub4mTIdcpkEJXqNrLBwD6/z2UxoTzYOnDMadELd8uRqlQs2F
gnQkvg6AIQsYKJhaSznKHGobU9vEkyXfJtzkkB88IzPwUQF3AxZ4lwxCLajkEv2rXyZXzUc5B4TD
gbRpTtq2mEUz/vLh+/e6wQDyFIR+NJF0vyL351asAQcnjUE2youbsH2JQJYu/RVETavIOWrcmY5Q
qrBX4Vxwc89BWlyUGNAuUn9K1yEv9x3bwQzkK/OEBDTXCyNDyxVEXKgmy90qKMeT9jsQUY6pgBdk
n7R/uEJz/Ngs3f2FkfEWzLLDV5MjfDTsGrrRMdRtJROD8iFi0ybt4HESrHpmX74LR70DWtqmMo0x
PiHhgVhQOLoVz31JcOgKBq9DSbN51yB5s+V4oci/HqLVYSCMAJ2f2+I6IG3HYru7OM8yUjQfOwLs
geb+06IwwPkLe2/Npb3N7HNFivkiYLok8Pr2A9+Y/5k071F/YvigjcLBJZ6hO8j0Jn1IVIk9AI7E
hyrsIaeAbFDUncuhT4DYsXvh8izhauFhXeE74AoiF/6mcWp6Z/2Y9t13185qP/9SgCrAyLJiWIXE
LIe1Ybp+oQu9QvDPlSp25M15pWaKMPZO3ftBPgnjWcswwHtSVoruiG0QL0Tmp/qBymdz18PR1IbP
oWYdEjCsrW4IXyjfxWJvHcTgJvbA4KPn+bu/ECRUFxXtamIfDuUiR0u916R2FpGeTcXaiXcQhpWn
9Wvv1FUvaAFuX6Cj8LgLMHE86foh010+t5DkJ1lrqGqsgc/oflLBRhIDenc6gWFLF+7btxveZ1Tp
zCqGQUu4S1BHTwMbTn3Zte0aQsAVBBzXL+vRSly2TVnbtSd9pNhIckb5nmG3CzYg6MVrwwe/HCxY
+Y52T6mASyr4XzxK7blRhFqLSt0GnNMWCOK8vB0dclECx1GM/gBx7XfZyJEb7823ClNrbFYsVNhk
It1oe/aIwIBG8+d/X7y88zpw2NRVEqaMflLuwHrwd/jitnP8bXD8eglWlIkIFuJaFyhDqolKPg80
B0QZEVLAg/BuQHidmUvnBhRx2zD14gbK6XW0L/0QELSbOpNlyWFQRwvKJrWH6ysr1kUMgvti10Aw
DF2CeUZSYnjwVY6qpIaovjFoQ1favCqYyrQwf/wCJsAU/rYa5FijNi7ssIO+w3tazuwMjrruVvKe
x7JrIwDW/n7lM3j4ZPwMs7kr/zeqYVevjQ8zuqe7tDi+odr+A8R28LEABwfpdq7K7JRXHf+tpMc1
Ftm5I80ZJJDGGzih0kv1+qD5NDAKGm2lI80f5k7FD/icffKOMhQVTH72Gy0zMFfKY26+CCYQcNk7
4+IcPwU+p3iBzgL62jOIo6anixp0/v/6RUf7UB7eVDqFZ5BMc01ghs6ERhBn1UpD3KLvOaB8krrb
UtAQVpttsGRfwNNlQ88irVWKImD/XvgTW1qubpAPqEnazzUbajk2W9x11j7xbmChd7q2/hGhXQxd
BMP+7bbJpc/nb3dpH4hArW2AwAXC7H13xpGKFTNVvd8jwe8dT6KpJRJ9Er1mOTvG1HQavsuuH9x4
6jKmPALgBN9iT27h/y/RUOwcS0IwmCy4Eqtb/yv5ax9DyIwO5rjqACNhFjQyOW91HiFIQukWbSXP
yI/xBw8gRemqsTJXxPOYmYZ7TmrmnU5nvHH1r62KY7wfVklNi5+4QRZlplFe70zxfOmPmTfYJ4nl
0lcuXVq2OqBB8kI6kKGt4Iou0VJrL3QAgtXf7HzJW2AexX5Z+Z37IZvvEOkQHyGRcuV7BkUvgGhT
PKQmuz+8Gryn7bWFM2B9zlazvfniooBUWmw68gJgj7izcqrtKA66CkEqpQmEBI9KRBN7gBG2Nmz8
Iw1go32XYhUTKI0ql1YBW8TyLy+6xeVmsOqCMef6pFZPsIpD6DYiQDETjDnUSdoozUrNNnDZTdF/
Y4qFJ4fWkPYIxot2Ea1/rR87ra/7kraqeMQrcMvQgilpNZUa0jrxc10a4PqXiSFtpMGPLvnwwe5p
pVg4R6Dhf2MA/vJQHFCZF4lx2LNSClcopaG/qdXypjFS0q0hHkJuLJZqFRxLNsjuN+sU+UpePjzI
9jRSSmg0mv+sh17zTiJh8g/NsuDO+O5YcsnliBuJSAEGkgLGfYdnACYkvYkqJ15rGbrnYNX6o/8K
U7e1THZLDj1bwUSPWDdyLEjgBfv2gtWRZgEbx8kp4EfVXMoD5Us6OoWJ7mdKLpEDXAN6hKM1f2wB
Z7Z4ldwQ6M7H71n1XtgE4k8x6jz+bCNNP3SzbSz+02E+T3fkIWCPI58ybKQg07mPY/hxgBMzlT3/
J+ivnYhe3mXPwj0JCx15kRd8G774aY134mSBxV0UA21bjauEDqdKnWRwqufA2ejPRMfOZInlLEZw
pfoBM5fk0bnz77KEnTFtGHLXaiIXUac7PDYBIbikCyOgPWWvXzomoxZl88g655PnG+eKAV6HGMKu
wdQnpX3FkNTlZbV6D6pFISAVMZ5J+tA1BzHt2QqvweTbRVRp+nBr+ypGiqASF6PdByH4Vt6JNle5
c0VsOSNQaODZ1fx3DRPiJAI4l4cY//YIlV49h9rQyOOY44glE6kIDKFg8HCvp9l03wU+fNWFxizn
K+ubEQUTmaK3QBXGiHk2QbppCTLo8jkysZpmEykWqbKmmf4pHht5BkNhT5+qHoYJv5Oxc/w7Ap5R
JUNSsqG8Dw6lWY0f3/DkmR1tn+8yQ8OrC9jGeRSXqXDFTmLWNr++W6zCfsyqL40oQ4DdE/V2mIPE
/OvlDlCVR09PtvwdadnKsBsVSFhDhjfoiLDeNCIAMlh258bkOoj0oyZuqBKYme4y5GO31ZXt60A4
zRqPEVemFLpniJTaOX5I7CQj29qU5XYyzDSnmqiCeTsIyfF5wDJlSbZUH2/cOjQiCqV4ANlMGjLS
bKusTUiN5z0jzO7IxkC6Y7y2HZZIBudWiLUqgyBr+47SzMERrtkRsPAr3SMJbeZdZ3thetGjNeDX
YObT1EWOl1T+qwVclm4JesCyU9dsB1VjubMfXSCANBFUKgOHXmgv7/qiyZJ2gy96t8Wfv7bq9Wak
3CurGk6dHOILzSO178sYSMKemcOU02PYyqKodhV1zONKiROSmxNXVs90mQQpdSfTjqMfzzYv7gN7
jG4eanv2l/7+bQBLVTimOW83h5Oy5yanN7Zz+5aw6ouqb6PwmHD+sA938S5bzJSAVx+xKQaID4SI
dmDkujep9oEHP6McHrq4lSbwnfWBnHKC+XzEd+rh9KJznzX8NZ/fk9qtFYpYrYT/vOvJjJNpMjvk
9ElvfTfR+K2Ex7NCnYMm5H+t1sGFgnEiZAQQlTcfgYp7Fr4U8mthHCVdG/SCfXX8rjr8S6usJEfM
JuOR1F8h3tzt4aWaBZUE5pFXsJbRSUoZNtBiorkTWDkPiwA45oq3xabgKAO6cy4L8MxIbuadSJag
Asj/nvGRHK1grqmtBR/yifoo2aicRSmVtGNbfLvVY+sV5d6a9PAiSNRZfP/O/Z9eaVAtCxTjgquC
tQZvr7y54epA9SQ/8Wsxd69sDIW2U55a8N343nFwbaHopkA7tTfoZxMUyrBGSKIezkyN7Yjmx5vf
FnJ6jDUPhOYTwd1orCME7HsFkzxdTEgtUi8v0VxCSXM1UngcaS6yq9r/rczv2RO3DMdaUaInC0tD
iV4J8Ux2kMAxaJVhJQQ+X3aZg1cjKJcpwuzP/iCG/mwAwaWf3gBD2agjl6c7CqzQaN865kl5Srb7
WnrSB1PVfJNW6XHIS06j6JtJlKEJ985PQ/5//wiw9jOC+2hysviPskK5V3QmfBigdBaTywvI2GTv
RUP65SJxHZtFRZ10r/3MBIDDgPIKJjYeoPdrGqUc8kI1wD43pciNgkGru3dPYn+t8ZC/AELlau26
Y0+IX5K9e44uUdoDPih4LeBgQXpjNLznyTPwgeVGrnpQ2y4wjrdsMN+aBn7Pg4i+MYXjyCpLON+o
duhEePIAkkBc4i9lPR4BIh7uWVQh+Phv9PlyE+0nG7eWhHHEL8xVPfuHw4lIcAIFNxUcNBatj7xj
mWmAEfdm50/bXin/65kaNvBTy8AAWlylW8pOTxSkmr7U5Z0Gct1lJTvODFaFOnZ/oXtRqX4mXETV
ix6T+HDBrBNAnXVwOcAsMsQlzTCPTZLyV8iBU/fEPQO+IafX9MGdrh5Wfy5P6JKFCQxZAHYqnroK
PUdIxazbG4OJiD6vk1Kvk1lhyuZtUoszCq11oshUwMKiYb2z3TBvg7ZE9J0iVAUCeO5eVsAV0xy/
dVLhhZ6csHGeOBG5UaEcxVqe/ej6NQRQFEHDsNa5+geCnBalXJXr+1FkJTlrDENcowsslVq3TE/W
I/3M34ldjHOyVbmFY94hHTR7+KqxwJcDR037zPJwFE8AjiyD6lNcLjqsN+S0Xas+8DYaYFig0I/7
3UfUxWwXNLRbc/xVgqyvxHhrpiXSJpFBq4nDQLLp2E3WpOad2eWr3A+ip5xgjZ/4pLPjMQfvQw+d
RCZd4OxkQHjtatMKBxOA/N0bVhTgjndzUJfFN0r4oKvXXfwLuEqJZj8wc1c4TYqeGHgMv3WFXyRk
d4k8Pne1dgXcsA5Dm9uRwEH8DCj5OwmycmcI/vXKYT0ejSkdBuLts5zHgk+amSegad1LWHlfTCFa
9I2JKaeimWnuXhR0GX0ucaflfjeHMk03A7GhQUl9Uwbkxv7Q6C4fpVqwU6FHZdfRHiuVi1xHUYfR
0N3VtuGF270BX8JkUcBKkkaGDVpPCZ6q55BkSFu+geU9MJaE2+pw34SCufG37Z5Ym+ezVlSgb18O
mvYY65nZ92W1G9oABJ66LwmVHfEQ8Ma44gvEY3WO5N/maxQxWvCWHLt5t94/Ycof1ixC70ydRkhu
Ho5i4iWOHutz3IUc6uEM/AiLqknnDuidbbqDe0kR3wqHxmzE+MOHY+38b4Gxy1NfF3vnM9Tts0v/
/62Vn44CTWzXtB7Yy79eF+hOXegWzxxUFkL6nZEiNylyKayrqFC8c0kgyZ0ZUEth78kG0cP1Jd1w
Uo1pbfMz7eJztZhNvFYuJn+KKmVwa58/1JYPpJKAzvDRF+jmwJWn0KNBEOQoZmnwC2w1zxbtPBYW
rQXcQZXwpfI7/Lmtb7L8wjhzm2NULPBrfcH2KEqXrwQESmIYDPftyXdPa+ANIB0M0Xh7bTt2jzoS
xXWt8pBKWWW+fQYNpUJdz+wzkzIqCbpKRQWFbTVXJfMRhBhw4aztTxV0fQCaUwIItdqQoMGA3iwg
XbQ7+amjlVC5pW07PflcJiSQyvRn7EDIx6ewTP5cQCo0jZTi2cfAfA78Y7EvkyyfaZ8jlQP7px3w
3CEpQTk56wEUbsgm6hqahzH7k75E5b7bkYXUWDbs3USRzFhmaaRPqH4/psaAUxN8QB7/Pedgnh4C
p/S5i8p/PGU0ppQiqffcT5N/9N3vlYV4Ae5Eij/mis4d9NklCL8MUEOCeiMb6SvuxvRlqRGSEKyu
OcjFERkQBM0boKaVhqXhsnaasZCvmIqYKGqeR0vzeeEIUfByTQhDWaUVTuWKhPNj84PaAbQHn0uc
wHAciy6KFZ7nhMHoUJ6ZLkEW7F/pxPDWTyEKgQQTMCjVQmAM+gM7uj8WOUxAKxS7oQLTqP5rswjJ
RknBklVX96xZezSIHPzfLErUZKbgmKy/Y8HWRU1Hfmi22lV4fXqpBGNqaznvQxtOWO/YasTVvAjX
k5rAw3jii2azDm4wUZ0Aan+qQ3qMkUdb4FirgkF74aamJXu7IO8nnOEG6ilT41ePQ9cFkQB/qz0i
QFT8rQi8x2MUvl6B4qv3c1suALEG574N3o/bddx+v5EkiBp6Wvt/5l43HIHx9iz78XwX7M2aP9l8
+1XJld6dd0A1the44tYtT1/yTUZyo8h/RcD5s/qIyvdK4zNtIVvY/KA+cDHevXWT+ZJhzcOuOEM0
Si9KMNXs255W9z96X6O7TcasmTWZqgZYj/6jBlzTB/2sMDi8HiF5ZUB1Dvp7UMc2tFesS4HJNq+E
xGPYrC20TvuAKLSxqDTTuBV6NNeGz20blFcNq3zBmQoNuM/zfPG0ilWp8h5oC5osSQtSvoy1yvQl
OSoUcyRAr+Apb74789nWOdk+GJYToPtCJ48WOjMtGwqpDJUiV847zV4p0seHw0Bi16ptQBIWwUjd
0b6fCkZgnmn3E/QULvvEOfQHlTWJJ7pt77cBjNL4/gZlBYBwUJ9tykhthoBv4h+luBWqeobBrdMZ
yoct+FPXwU38Fm55bFexFM4+Yvb5HLBXantJs8mK0nIK3b8ANIhwKi8HondNBTL24stIv+le846x
KLVKYIDS7FZ2Fkhifr17zKG+z5zgAu7nWnW95Zv0odFg6MVnQi4gWlyYHonSX9MboXPYOKyUMCCc
5v7Oj+vdGmYoxF4vaFV434rNiTgHqeYeGwN7DWOHF+jofbWWzgPSMTzXQrWCw3Rx+HDqisL0fKpw
UbL5az8aXAPXzTNxC64TurzEP79aGC/l+qRWvO3YbH4aoSg1AEijDIccS56ebT5Kk2K6Ysc2V9+s
ISf1/iSaHslMu6pTUvn7Bv2a7rWNvkJ74YgEPxLeV5Eixtr8t9FTD9G7g/xs20fMN2yeOo69wxR9
B0b08Xy7UFzOuv6eN43j9bJzVQBNSkw6tfanWopMXX1Td7E/8WRSUsPnz06CO7/KOt+PPVwLq6FJ
tirENMZag8ZAlFu3iBJykt12hayJroXL+Ylc8ufTcHumeCSD56ZwS+lynKCZP5ld+7IOmdDNG92T
hdVe8dWEB19GhZwmEK7ANu1U8CTPG0Pohbkfmkvy8nXOUQ5meTAeb2c+1DCOfeuPz9g7+QQKcg4v
JiedGBfi3gfUIRidE8hRXhkm5l1DkBkWVUpuNA0p/Lgy2q3dXB5euBBeQKN8hYESSHQSLAM9/W1V
3aPPx8L3ClGesp4SCM5U2mu2y42jFZ1Jwpl4WAfXig+zNMIyJoQGKlQyE/GK5X5cMP4Fv9Y3jZ+K
u4pRovd6IniNbPD+ahXhC/5pjm+u3T/dn8lMOUKtrgEAkyUegYEOfLIrsG4JKjSyrHNfQAh3+yzf
fmVxtgt4lbUZG9gE4AOirAbbms5990Ns1JAEwwk17XtZkMsTmPS9+PbWA/vwsST5pcuOVjgtGg7l
Rlb9u8ugUFOFwGDqzTNuqxDSiQTovUDW2b18xJcDlGGK813acalayD10wu+cfOH7hLe5UXHZfPoX
UA/eWXsPIgUfzJE8mR9AHhPinQdIQv0MEszLFAPSkMIyxsNxuYfV4d2Q9n9TY+45qfFRZS6X0VR7
4nDCNz3ElUsSYk26LlafyKFM9TDtPTXQXta4sSwK9jmGIwnaZMf1AkV6+Lc/7mbKPvNCnNbZcdpN
AchmiM4GxHSs6whSGhkzY9B0cFUMqKW+OJ7uot/rMrpwKiGmuulMUd28YCDratagFW85iThgi+Rj
VLn8YvADidHOxUmg+OkheaekQS7ILhknq87QbK10PKCCInHGauASzp8BJNkr1tNnOeGuIhiy5Wgm
BrvDQFXEZlcg3n3fCRq4oaNCPE8gk4GQWZg8qdNblVeLkLGMdi6fORjMgxjC9Dan35lpWoUPBnFv
wsrX9TD/umfljEuJwMMSpxLhWA2iPGpDuGj/GFNGz5bRtK53MMAlKytEcadXHhyD9hpboyKFgW4G
pnGL89IogmsheBEvC1XuwD1oEVJWTMR62ykiJI2cx4wblGus76yLwkYtzWScNNapBunEV+JA+ecT
B0s1w5dW21qo0C1ebPYbyQ4anWWcvPe1JkQ9w7WP5SJ90HMbk+OwudHiTU+eyVk4T0GiC9lVAxHy
zfRwT2GepcL/rRnHb1pSjSpa5ELEPQZMM5qZ/FhBfQGpojGS1v+sECkHTHfsrdssT9pqtuwo1+48
T00taPlJkBqrr6xx/onKRY7rjjVKEZ4d+lfgfBmRVaw/KxzBWNcIalS/nOOjc8OMxBb5bPODqeIz
iHWVnmH3zhgX4DG4zftoc+0XkI1mKSoXha5yz0X+qv5xMB1y5oG74pINxUbP7HFxXLDnEvaXVeC/
sbBKZkdxNyDmbjJKkaK/03b5UNTMpPn7sxkHwtIJqmqo0Zs7RTx3evzwhWkwUyGH7LNgppBfAOie
Sy0ZWVSt068nmE7Mk+0XVahmpsybf1BJwYxN0wUs6FfUfAdkglNSnGJ4FK/WPKy5syfSN+BgM9ZC
Npx/bESKtbjx+4K3Q5Ypoh3YcAqQO1RS9W1SUTUb/v4kx/MGB64XoOFmHWcm4mWAPDivF6iDr+oh
BToCf/qwhVEfdDkhew0kic7t79JnPVGT6wS14eKgUWk+6fyiX9EE1f4DdzpvCyY2st9aRKcNIJJI
yhWu7Bq4kjoWNbPMLDfgsWdPdl3RG6LsFHhGHo3umGck8prz3po4++69txYaZn0SfQLluHUdeBId
SoxZvz5uGwy9XNteeof72iGlH6Y3Szb0oLGaIRXWinYdX0boD9NeRzrCUoeKrzuYpsKPIeNS0TwY
EIhKXU1kOCVQ7QUnfwYqdllboP1HBAlcF6c2WlXACLLJ1LJ5UJIGd0Q9MAs8CO+SsKZlIW7F4wTj
oII96PE2lZsYojvekdF1rYxyXu0Z4bzkQXjqxPVPUV8knTbSSvPvxQFBiuCMXFjmV7awX4BBZ65W
8+wgd0b7kmTJheQIHF3s06Ruz2gJsm9dDlXzIUIEf0rXU7AVzI33TFtyN52+0cUG4qQ/UZ9oodDx
H8q61W885N6pQMz8cboolIWYg0v0bqvhD02OKTJFIAyzO3rp7herznX/2F6aobsDhYz/aaplQ5R3
hdgJ1iemG+2Ks9b5jK2qA1ZqB1kqK3eNHWC+CPyCYtCAiTN+BB4neTFw1a+wPbIo6NYowEISqJ7L
JlQycH9uf2N40TcMFtoFjq/HU7KchrPpFv0Qd0qza8D5MeiZDO9HgjwA0M3rqOS5X3I03s2Hys6D
5/j3eQNVLq7OdfzJNhB4/zCDOi63HBw0SRhZIjbSgyLqW6Bzcn49kaZb7YLI0FLra/WOMNCMgVQi
30V4v+BDkxzVPw1tV1Sa/952qS2F3Kkud0j7WSWL1d6fTrFkGhzwzYxGpJF+LnyMmojnN1vTOTts
WusUEqakcR2EZgjpvyj96vyWu0zlyXmepEVz0WfcxF2RuufYUtuXVicK4WMVOUtFLtbwYU928U2O
e1hymPr3R+L/pJSome38LaunMXCUW0vP+exQ503R7CzNdwXFfY6nYQdKUqjAg7kyoJwM4KIkL1N7
N8jDMPAgHTZ9NREVF0RYEng4z3+pLY50eQVJC0RvKvbWWc01zB/cvHUMI5sJhd/0d2Zfm4W6xUMV
gUMeVtWBPnc9YDFkXsvu4HYgXwqSuYgt7OE1ALxPOBD0R2LMut7IsK0V/Y7c6W9I04/8u4LkdKiN
0c1YbinE4Hat4dXg21Z7Czlv+0OghKLkIPcYPwsdvOb4d3S8W6u0FKLzVuh3+gRbOM8ROA9HkZAH
Js98b8pbNjFpzVpinfQIAjwhknEJQGs6mccJcnXyTFhWw/dYhaD5nSzh1xWI3BAENqd3Sf53iBhD
zvQFV05VSAxLI4Xn3EbcnEyh/vXYZlhWpR20RHxK87uvEmY7CwzbgTFHVepmOkavs0qlayVa6kaq
sZOF5pUCCdLEJmlTr9b5gobo+IodIsaGLOt8i9wyGzcuHuPmxG1TftOy9o5/8vZvrTUR+4ke9nPr
tVSL3ExmKZxiTp3O7tup5bbapV+3qX9IbDI2AEFGGOUB+z+giP08LV7o2cnbapL0kKzMkvFvrcTp
AS52dl20mqazP61oe58yCJP2c5sDZi/KQ6uZIKOovl93EeLOr1tilG1ff87t87iIFOqlPleJMSep
UwqMjRD4fTqEcxdy55VHXMqJFXleoR/qFlMAEvaNZBwilc6zZPVamVuw/r76Up+Jxrwl+hTk48LJ
EVRlxlMwUbGFVuRDIZSN2/7aFbRPnQucp8b1F0S5UbMEbsKEW1RaZ/HzXblRnS9cahCtvTKi7t2T
iD63y5ekbTmxGpPn1WnQvzWop1zT6uFretIGc/fQLsr15nsLLR2mDpqZzUVxsifXK7U6HKEXAprQ
BMjyvLZ+4bhN8ik9LnQU2VGCqf9PG1/9/CpZA+9T0MYrYmqv9z7PRsyCh9q14vLhjKjLYwlG37p8
v9mxZfgQeuMmtxC1QjavZKHoKcXaLjUeBYXR/Q1Ur09OjjMFwPD8JFocSmIV0P6/0igPO7RhTEax
obeSH7pwQWizB+fsxYbhDDz4T1W32oIndEOSQVbhPg98oJ3//1iHFaCaGKcbVpdALzuKxx10ixyA
t87UBby8h071V4bbHWfJhQNsAL3EjCicKarnFZaYuK6PDd/bDBxArRzCBUoylUjKhpFu8Da2K/Fj
fkrZTk08gvpmqyJe2titUhrHgAP1mRFI8290Fcntlzp/9rNIG9HCGbsmwxDseLYK+C9ab9UmceuT
LEI57cBvVuWuI1krO0sFcYWC0hXR/M3/fuCsU4mO2I9kvnQFRwKih+PwlHqeKYs9qim6N+X7oTe5
BYvbwF2wghKmDX7YdVTgVN73yxuZjnXWpJDG4PXCK6yTulF0jo1D1rIs6Y8bOz63OPUHTrR9f1DU
xt4lxK+oG7Aj9O8tL1KomE9nEo3+JU1OfZRcaj5BZ21ADHAlGyhSv2/n43TAUI2NIHbVDOjc45L+
BaM0FdxODejw0oMYqH2n2f4Fi6p83OkIliwpu7TXeFoCJTHaq2+Bas1tfcX9tLUOZW9/pDPKPBjI
4XMGcazctnS/sr51zad/hv3P1yRCP8sQcTBGU3e3QttI3GAELU5OmqYX4iOySyL9//A7g2Auudk4
z2ZCUeJVD1oU2iATpUwdlha/NtlV4hfekrfiysBceZ+gg4N5bUSfkBYlI/DjM708KlhE2sDeV5Gn
LVJJG/sd7Ntv7nR4YqXdRE81TyqPMYY98NpjDXtLS+W3oMLW2rRQm/MCorUyOF4mbsMVmSy5Gell
mXSFWT5PbbI8X4FowazMtpAe+pyh9/ANI1tdfdI3a4GCyxD185PZT1crfntjYsZ2fHNgLcPCIxfN
VYPIOkVFdsMqMRb9ktkWMQtR+nFeo/+ChPAO9CNg3sDawGOlA0vXnP9BzAfscH/XHzbXmMOHGzX/
bYbdGa30gIWr8rkqLehMTCk2IyBtKU/VT5UqmSzNCMHUxBGPK/qFoC/vOb2YEMUQFrGxoef6ZEHU
3agdpFpaGkWv7/GixA5h682FokElYrDwdHMTJfmt455tAQ1qBvLIDWFQ8QjFhddBonqk6rnSnrEh
vqgN0WpZDwbAq93IagHVscQCTiK6ymJAOtS/LJIS6dIbzVXHiHDRnjPoYLkmzoXde14HczSTRUbc
RIZq2Jf0Z/0YU1ZPtWleuuksSAfn2WT6TQrKva2fmjsGnpLExUmQRy62vxUMutlj992Evdv7kNW0
JpSsIwbwFSZZTU5ctzXB1UfkWbwi8pvI5r1CxqkEq/mNZzkdB/DzOVauSxbJW3CXc0YHToa/ePTL
USGbXcQ74oaROk71lwGwTw59ft7kCxJSvufBNgqsbN+OwUDSYrWPmLqiyqPfPzShfCrJFo39Dgwl
/KbOPHkt7fhqIRzBv0fRshqTvGI6hjWuU9PdWvHEGDsfl0v39TZTCkbQP4xN6Uazv5GFMOufLGFu
W+2O7OVKwRXZLTbhNp7zidc6i6S46NyzQudypcf32E3ZolSS0yVok2hk4zBdEjrxtjAST0rHwoQ0
OKH5z8HlmqsCe72KRhXis5y8adn+bVm91ItUD1NhQ3NFLrMxYl7ENugGsZMmzrz/SWXqdl+KGzJZ
E3WZYlkBzHO84vSqsYXoFJKbIKRhBu5vBCbxH9rkwencaYJwz/KaZCw6WltN4qaeDhWT7lafKs7Q
jTSXaE+S7j0rmws8/cvMZ3xViosVcd8j2TVDU0ku5GZhoXV4lcg1oe7kcYh7mp2UV9k9V4CAvPLo
roeifrrUg/C3LhJlflb94t4VHwSHLOwIYA8ZGrNErkqF0T9msHl3o/Hp+oI8/GtowFXo3JjCsdUJ
YPBXQwzlYBVW3Yh/EZtqRvkOiiH7tPfl/lAL2aM30cpnmb0V5eqOAQZYV2etQQZc56ViKVjJBo86
7ZtEDvDoYR2thLQRO/DP0TUaoNAjLAbDJPq9L00Gkygqo9l7dk4W+X5hO4O2NX7mw0eBZFH/mqpY
rBhkD49mGcAoXU++IlKdBdLcNn0CkEuncTMcFSXvI+J1fFXltkC3nvPxMF+Xsgq/ZUs5bWkQdfn9
M8eXtCc895cPiftaBmGy2wJakWzIDDC/szpIrkAvY6D/c+TmBi9XRFfkACmj0UB636jIwGo64hO8
+YxHoqZwcx5M6yMBIPyuMvkGzgJKeFhSOWrjnVMStCKtNzAsrGOlDMvAGByGfbUxR2cLNz2kUdFg
kgucomcrDpIZ5OJAZUiDivlFfHqkTpjsEEVi5U1/YECbU/P4cdDSV2Hd/++RLUYg1eICa5AS9sXz
/UOZMSgQmb0qBcuau1xQar+5szC4YYLSxx2KDXgsmGfHvfF05upk5gKKquU0MFFPMo1I/tEjgQCU
0TFUKav+QzWoZI2odGrDTQLG+QZ3UHKP22qqqefPn9xm4mLU0McBnGBc4s13o7VVwrVCJto12sFT
jZbm4CLN9ddAWznwW8f4uZLcqDxzXpeo4szUuS79hh3FnYkCi7iSo6jm9LvBsTLuHjmS2hvPEcrk
MasyUwSmVmD1VaKf4/+CkqEXfw+aYApaSgwgBlh1oM/jKndYO3sEoWd7VkVFRkbul20PjVLBzjr6
CK5qH6zMrNIPka2aNVCcvaaC4sYbI1o3ewqQnBGRB7LvqVK3gfUHJD43iyoxWP1enShiLwYSk6Xl
Z0WWcPnKSZrSslXdV9WzcyiH9VRzDCjPrfjDFugtBEsKBC8se+VnsB3B4VhAb9aicRgk4wU19mXE
GpH64XDh7h8Ji8l81K482vNMFhiY9D7s/biw0U6VCgHttGvn7CshuwAnxCUO1KUN27bBMT2Mnb/9
VEATQcijPvB2iGB1VhSOCBnKtmz1qPi6aUFS3ks+QYscxz6OJ2i3dMIvqfODegxZyW4WJ8uqlefU
ex7sajQdZgM2k0bIeDrG7fFpCygY9eM4E+sCDol4f4DD9BWaL1JzGfCl62R3LseysMuweYAhibxh
6kPHObAByvNePRvl2vIMsFm8BjxriN1nxIQWU3ktO1kwsFKErxBoNnnazLRO/QBx6UUiRmn4kgNC
Ylw0OdRH5gBJAShorjpr2Xj/mzOf+6ETjQm/HNfhYC6waX5XvvpqFIzMM04zfF7RSzh3CmFXyFgy
+jd5lbwQsdV8NvyOk7FwgsJFKRQmpFcDcPi2NfqXLE7TMqXKQLXArEsEcdYsE21rpj381hXG4vo2
m465jJPjbRjt1zRCsEpagUIBsuAdpSdI7Zwd/dt11Rz6H4TYWTcLy+EQa61XUO0NS5Gmvi4gGBHX
PAcR9/DKzZfpwem47Kj/xZ28RFWBbVVXJfvHXAseGJtpw1KTZ9iE1rJQwGqFzdGqhT3uv+zhOIcq
kKW8K3hOt6DSeKfedcSI1U7awxbrNlSgk0W+vV4j0Fr/+Z+7bV2W05cnNAyyqg8eaDT1uQzaz9e+
gQItK1tivbFM40AragZD8yAHpSlum8asGks30ktCaYxahF5/DFcIRMBxv+VbSIi0XhEDMq/KCOnt
DL5YqMRl0Ttybk+njOUmUh5g7/+qHNK5GDj1dzk+Tkw+Wl0KhIkOwBOTVhgaZhn6QAoDxD+1zJE9
MBV8X80QGka9FrBRqaPLaijqDvMYx4hh5hTZLcSR+knF2cTehCx3pD/1xAOcoIF91t5IlEIBe105
Gl+H0CkIzMa/DJQlge4klj4P9tQrPE6PPU88LB1dmbErhlvSabP3l/iCM/wnoyJqPsRhwUKDKmBp
2HgSEc8IZpFu1mmUy/16XJfL2d2EqGXqTx4dZ9rp+3NaKZdY5SgQYVsA/dP8UMEysz8hIOWt1u12
bZ5eg6S1hfp0McufmeNSeRCP9D7XQwtEcpo+WW1F1Qs3hT0c7g8tDjpYPRdcwunoYjkNQ9YsCFiH
RpLO2TlxyOfS0rLzukGgkxPN/1WmBs1NmmNMOQahM6dTUNTpvVOx5DkIv2E8dOR9y0HRLUiVPrUU
f0Z+1NCXTin1LouTaT+MI8zVJ+RDztCmIyarUlrAvuXGkEaxFlwehGIX9jT9KKxjIVZ1NALzO4F/
Z9unvVaJfwEgXIoh1dK50x+iPaPalCeGN44SnIVRQqPwJyOO9CQC3kTw6uJFgWruBLzrUJG+QOjq
/63YFfc8mmUXj8e9kPr4QjiC+Fpt0InGxRTAbZNgTGYH0APhG+CLb9B1tx0fbev3ilKH9yI9h7Vr
FQgfLGPCinIuavBiqu32okDIAWn2CBbQ1h3vDxa1R7ZauYPTZbG5VjWPaux1XlbmgNm6IxMFZ4Jc
SZSfIQq22VzGWYcnwjgbAMyosZTnYWjyyn+d/KPMN3t08BaCjYCGGOymRXZcSf3INE1hE5lh03nq
vgPVRqHvY+Yx5gMIp3JEkWx2LtJGobOXeXLpq/xATrBgQ9zFJvTbXVKGfkHxcwzTPAKatf5L4Wxg
R1pgdOPEgdCsHbUhdtVe6qm7nD/0SGltM7Jw5VJ0bSLqJ7e0BKeIdUxyXLsYtrNV1kaUEIcNsYZD
koIVLsjMNG/+Xacs49JNEBZyymvOKhC9Asho32OdodV+ZpqBtVNqHRN2Dd6bK20XPe1QHs4Xni28
52iZ5BA8+KZu8nRfZnPzfft29QTN9jTjMHvyaKB9rhcgeTErQuNVYL89sVAFENwqZgG+//kGZ7rM
JVkTrqkzOC/ObcAPQD7JEU8rAkoMiLpMK0Ed7RoZ4KZip7yYOPyhu0fDXVzQxlo9iGBvXNyyXKY9
SGy7+o9L6NbOzpzRg5sJIuzWJq49g7oWEHbAcRW99HryNUbCnzwFeM0B9wM/YnCKG/Xe0e+HYy+i
6tKhqf6K4G15g/Um0z2on0m+72kdNohqsPLLf4qWHlk6JKCWv4FL33LKtHlC4wwZA+R+baXKcdwN
wi3McYcZ2t87E/YZEMrDUdLJG1dscZ1VyCbQwrTJv9540pd8cSKOAoEctnfrHgJVD7RuVz7wmujP
U3/ZXgovjL8BfS6UlGVMZbo77V5BvxFcnmiCwRToqYmOt9A671FxxImPr8FN0RpIBIVbYwLtSe+/
Fd6rMiVT6pNM1Vkoo5abCW7XMicGDqX0gCJqUhvklWnmmOKWA3rDWQXjueVlEoOVejkZvL7OTAiH
nrlGsnIvwQAt3g8f9a/1WXnrWMy7eKNpcv4iv4oH+7rj6WQ1eqGB2xxlxGurOtoAdBcrhqLlXlM6
0ULv6aMyUVOxFX1ijDHpKIqaZVl6VC6WhinDlydUWoEgIHr1G4lL7OVldbkpaVTef34udxRVOBUI
wsgikF0xT+BamGi0qodNXF8IiaBWDd1bxxzE7ftNOEfWniWjMV8f0C2Ro+ld4A+9zpT2Nf8h6HvG
DhArch7ckUOK8Wp4e4ixu3Q1kYrsAuihZGVxBrmYlzEWyhLACAGwi/XwsMCpFLGCpagmi7lHakiR
9jPw2vW3Vy9sfZWQEQL6THFXMo5cNGh3H9y49gSmPo5rpOk5EZaih7CdTm1BMXdHEwZslPMVoem0
xdZDT00GqsW5nFmve1k2WZc9SIqVekcVoiuCYlyuedZB6h1qojBO6/WyMz5HECNtyrBXal9ZnmMz
VG6H4YPDBOO/usQvVtzxV77+NO2CpYoMEp/Kcb7qBqLC1+lS6zVaXuKoK8HLy5jLsaMHsBCdOUz8
8smB0cnDXX8v+kDqi1uPgkX+JDT/8pJslCJTb6gE4xVYcYMTKHlG/cgdTWNHQpZjDaK5FTtqUG+5
ZEYM7Tf8VVw1IO2fyLyl6DL9WeBCOpwLEhD6ME2qNs3je6bA99TI4DAxUrvUrm68yfJuMTFJYRfT
hwK1wzvwUIrexPkaZOGR0wseWrDn+HO3lUNBGopIqaZOZex6G5w2Yxei+eNzWIjXs0uocRcB0C7a
EbqPRUjphcEk0kXYM/tx6ecYqOfE7iZWKT52UiiGKiogiCTg+mxtjtxprw413y18lYcFdNIkF1Z2
IlD2PFhJNGhZpk2BWkd2MQ0eNYTQqxPQ5R6+WEaX7V5Rlq+VoimbhVe/RCTPZIsdYpQBhb4+IYqM
U1pzEx0Y3sAqhJgIE2eGSguPePrGjygmdzxYp63K0jGbJVmUizJCtLYJHCKbQBSeFS1MSEGDCp32
I7VLWU810sNekuqd2qdxNoG+yXv61GTx7ot437wX96O248xxlgnwsLP3EdTv8LvAEmDdAhZ03cWW
hcygsGnb/3AyqnSUD7CpPZ3N9cAUB3Boqa4yp7uVqMtfu5Y1QEmZvBYoIVcT2OJldAxur7/kKx/9
cNYZKP6YPC6rC9ohckClAgoS/Dbdv0RL0Oe1lwOPHcWKOy/XlI/fXGr9NgInoCIw3U+727Bhfhs0
q7BXmcvFdR6FqXcoTXf1I65l8Ki1bVTUvIi8EDjZhR1I/ZDgsdbBohkv/lXirhuoGqecPG6ibCTY
E4NVqv880h0Su4QjUozhPoCn/RXxAyn71HYo98itJcPATEmmRHyqXV6KpAmu/QTxePcsWABK97d7
p8FROlGyOAXkK6d4nrpbiKRunmY7BgOOj1wT0GmZW0OpkO9pm0aYZ9bmYww00ipc+a5vpbsBcy8I
0ZkMYZ9sq8ikRYuWkHsfz72Fn3yA6rmMVCFR0E4aXE/4bE6oQIhU2p/00groaICi2rIeeuFekrNE
xqB0GCORnTFWUCBLhBaJVpNC5jt+ErnUGXS94G5OGU/mLHjDX5jWjrEcZG4Mz8u/yyE8ktppjXB2
chAofrXYE1FkXm1XJAECWUSw4uYHBUSc9lZr7FajEV7V4V7Bz9Dy8f/7+oBoGdLVBABaeRXRInqN
SBjSDYlETZThm0jYkP7Ca7m5Cl8PgTdC1HVIMpUVQLXP0v1+WQsUckZFy15GrwxUwTLo/wZUhsXx
/lQRciFoAPml5JXOEhqr+ISf64m4EgOU0CxpqY6Q8liHonNvV+tY/xwtXRBavcva6A3tT5Qc4xme
PV6P+FyjZ9xlPipo8bs5BbsmCxtkBnDs2qJTdiPekT2TYCMhfXEVL/hFWxBlEjK5havCdnEqJAED
7lhRJw3w78SKfanWNcdhfcggRWHekcP/ruQBk8FqHBPgM3JnNblm6OEB36z/SQb53eEPIXEuQXJQ
S5T3d0ebjjwwiKYUuoS8V3FYDR+ou+GVoMl28HttP9MybF+1N+dnnkFCQfaQ9HkvKWZVNzERiX34
TioKv9bU0lPYfhMu+Z4JD4BnlHEyIdnNY9zxK27Z8rWYO9kQQDjr4r1smKESTAORdj3dBfBhS8YI
7QVtioahvGxsmYaWh9TsMlaD5ZA5cF2ZutnBR9Etk2+lXYlcWfKv6dFDMSiLvFN/eJZjH268xk+1
vXnNy9mTzCkAdQLg2XxgJWqY/al/yZ9saRQlxexlotAMTJGBBH4XQ8qzci+mcKbYEePyGVajamnB
Hxb6FnUKXZImiIF8UKky5BTYtlVoawxhn2yfrmu15PDdzhtJAOsp0vCIbvZzq4uLYALKv3NvqNj4
FrCDqFtsZ3zltniSGztTWvLbtk2uo8BKdDt6Eu4SugaNPHwZlm4aX1M2e7UOhUatkBmUed7dviyr
p7SO3bEa3y1q3cbMFviTT7jJgR6uW0BtAtmhaw0PLjG593yr9cIlaWoNmLp1fQSMAcGnxnHz2vhm
ZIezyBAn5rDWnPmEwy/5JOLa/+9L8IZyOq+UUMlACTSXo/gNgQS1wQp3j2Zzo163/KV2VGvaGW8d
YS9W8Sq9ckL/TfMwZvBs4zYeGBylUqDLnB7mXAL5SibAgUG+PxFS2ah5ZD0fMP4r8jxJDcHsWnPI
IxI8liXnHEyGS9H+biy9FdTQ52gh/cRWGB5qTAfnOl9z1HTSjv93Ie0OXe3LuiDjjN7HnW/PvXk5
diQ33ocPMOsQVYGiJeLcij6gtRTPDg6aAzZ31qRa+XxVUWsaUwjoeFxHecrGVYvPdKapIym9UdKY
h/Aoura4j9mh+t8BzFVM9GpLbDEvEJzwMztLxOrSUWNxJXSPNbPonVIj5Z+Zy07ux/e4nEfVhNWK
c8tQhQkxVggxl+/a4/L2pILseCTae5DnpN92q4fdnFuyJz2a2/eVHSBAsgrvKuGuFx9USM9BmTvD
BIoeU/R4VcKFFqI3mLORUIzhvPd2r2OpeaQh8hllShMQoAJ6rvNmRRsKyROlmYrfvubZrUhAaww7
mtpYAnaAs57YGmCJSkbu9nGrf08u9G8rewMUPR91n40+wbHuabkhIRWS4kXETS6Zg9w5Fz1TCZTH
KSZktCOLyyqRE5CNfNJjcdy1yIFVpeBFTOO734eTg1Rzas+dnHuGcItkZE4T+AnkNe7sMgqZZfF9
h6SW/hdz8/Qi8s/9NdHHsqCXSs70wRIg7QUNdSk9YgCKqBHFYpMfhdOs1xvplmHl+AaiRzCJxcMK
3g3+ZETll+liCIyMT94iV9iHv2JKpq0mMj7GlIoPePFb1C9wHue7C45kmg0zIru/vxx+zlzMJZUA
weV7PWG3VNy3zZhcArVS3FCsnzjLr+5uedFWolR5b4ci2G1GgfKb3pgCBP6AeMPZfBRN4hvK23v1
tMtg64w19wyCYBmN3wWXr2OhYYX0TlDZZe14LSl4L2ej2c+9iLPn6+paPBY8Nr6PPlqlM7mNNcb2
hAuwYSU29+WOMFqM4RQBlZiDLA3pt5R3IyeO/URiZ9Tv8wNO5xNGz474+OhvkbSSJNA7NgwE80Do
HxPT/q0MJPXFWUb+gq0kP09hD3X90eM+cvq3eEKk6zKv6jX++Nc4KCep/ZO56+h1HryPvOPQmZAN
GARXc+RAl2obyRCqwSXhmXf8a9R5kR00a09ekeajLlYDsY+ZW48oCM7iEwGZvtYiCxZfOQMzZQd0
420vetszkcZ+7jm5LTqBsPpUrRQ7MCF5W0QKxUgAknzOQ03SjBogBnpoC7JnTpx7cPiBouITSKYf
41+cwIWecP9655CKRshcOpOAWaEabbcEpIOcELiHCk/z913ZzIqthBPKwTO3X8/yg1Ln0Rd43PiT
aU9lhIEAVsldFmKPQYMjqodNzRxRU7QTdiVZUixuZ2QDBdDhpWBmN/9dW6b7Fctq2Yx+5pZaZovV
/7F6Yngfy4HXWNsEwUarOaF9YTqTyYHNGqBm2hhSF9zFZ3htfLMtiw0W1G6aVJCXRH1/Flb9eU+n
OF2OeslSQGuaJtwC3m88EXEl/zQW3GCJogUNkXN+K/jLa5D37qdFiyL6/AgraN18KCMH1FizCi2W
lIU9xpDjomO6BJBAPw0JDaxDDyHbAcwr2rOaRZyEREadpek5MNGojmKR+a63NG3Wax6fsoKVvB35
cd6cC3HZl1W4Y2nzaPtxOMymQ2QUSVjgRNkR+IzxxbXPtnidBc5wNCVqFIEi97doqWo3YrBoYVQY
ZjJrFnLeuj3QIBG2BOXKl6/uqGcEKKimwZLZtjcSW6z9hptTbr7WttkdiM+RFPCuwJl68FV8WLx2
V33Epwd1zC8MBF3JKtiTeB125fqM4RAZXkSkw8SnQEo7oDWLuZhADpTZlkuuCZ0Xy/Iya60KxEyL
29ktpi33p5rlwpcq5VQzXZzPRI2yhvU7yipK5+cSfYuNL8MRTP/z8Ga+T1PI43yXLRZMR+dGeUX8
XZcrv8RdvMrZgL98vGIR40MsglNZ37SXrKcBMoqyQHWLQn7I2COFeoqvMF4AksNWZu/WqkRxLtOO
/JwtWyprWXlpWkEoZO0Kbn0KFRapvR5Q/U5+7IQCkh6115U3mjAb/yfsCeXeMoPANQ5q6jbS1OHh
xuaFL5MX7CeIy999UGtUrA/41tI5j9jrM4gEvbgsK7U+Y0zxJONwA/8I+ECNtPQrt25dylxAH657
WefydOW8URQVm2MVaV42zeYxOD8By+JOt0HL6Q4Uy4+GhSMIRRSIlJd22c4BPbJaruqZPiCOyeN9
SBevOPsQy3U/KmJmas9mkFXOP/qSbvFO3RVlxw+BXjRqD2kBZVcXz/Fqe88+SePUy1aLDzo6y9JO
+2MLTS2WWm0U9HsuHMCDF14n69mdmMj3dqSYUXW2qIFaON5PknIfAXqfQnOD7accJHzMOvKxJ83p
H7V24qyVX71vri+bS1icjltF0ST0hBEv0JISu3MlvNXeUG6lvO8C1AKLOynzIVnNmZmsPLhZ0gKf
r0Bw36x0paH32HOfZ/OKpAOXXbbQnNmwhF7iduFu1SA/dfR0CvceZyg/I69jeyoemTkSayZk3eMU
CQa+J7terfY4R9UQ0wOGXDTrTkc/pusAZgO0DrR6L9b/iPacn1orOdu7O1Wc2R7jMG59Udi4U/it
UhyyD3FwHg9JV1DE6g/aPObFsnUFLkA97G8Dr8EbcCTt5rugnaM5xFNUIxv+3rLSrPyTQPKL8cTU
J76q05Tru1x4WKp4bwzpQYLMsUx3J+YdwKrVxIsJ+4o3o+D4rtF18BUhtBeg/soPRC4RhaeCcs/7
sikloDS9KCPHhd0tArgwcj3REhUhxlTE1NDMlSaITyaLpLPgN1EiUogGZstQlBssTRPk0iL/GRPN
oNgOh8TVdIZrb66UscgLQDaFn5UVs4MPDvmvAkbrO/naWrBViQv/UA5M8BLpzBrWb6UYUk6yJ2b4
wu+McQ5vr/0ySxajhSLDGu2XK2+RC9zGhWHIOPSI1fqGx6KYgjRJ5Cx98vPFKW8xoUjn31Z5S+0l
JouYphcwh4hsLQu8Pnz1s5rTnPov822rqYKb+ANdITxelICrWwjodsMivDntRH64TcRxZFJg5H5K
YVlpqh/yrU9iiF5qafGzDO4nG14ywNnyV4gSZ7FdGx21bv1hb57jpS+2AME5eprzuf7j6FenAq69
DHTVBwe16KM1dmZibraxtsX9OWbLkBt9YrjBAFYzb9t1PjQTX7K1Fg1psZ6Mfe3VrIkuV/PCMWql
lz4bFq8Gg5fw2gNdGyox6qD3es+IduySsAu8nIXNkiRWuKxb9FkERheExPhBfPsREpyr1tM2jdzm
2Ani+0xu+ZFbxdqtPrIxcHj6HhPEhIf/7ejSOMraFxZihV5JNWcLO5FClJO/HZJFGEVLbUK4XaWn
w6lwBrhmzFlTpi6wb2okWj/QVMW7MW/rNCgopkdBibzkzBYGdybVVQj0P3N2O7Hcvrz3Lgr1P1SD
yBj3o8KH5k+EleRSP9I9idsY2+jB36mWqyFPkYTtd6IFYlwlWMWrjiiLY5CQj8YD/esOFexSpQmD
4nFYDHg565FwK4fzRiJAGW7d8POJR90Lr/PDz83VXuqO2c1dXDhXOGmhTYsh4P5XS6o7Lk3u1/pL
S/yOjdtJOYaQhbGidSQrqLQjPlVQPyE9KTyM55z+I1XcMJEKH4UEGr2cBiwCzMIpx+SbiA5vgTgi
8aopwTZqyluqZ6dSvqe9al3PeoW7k6pcvRCcq2adN/pcZbI3r9zqtJWjfvBfPyF0B1eANtPA8iN+
mndIHzX7QAWuQRrl22GXZIByYbpxDLz8qdS7RVCLJcmk90KAoilV9nRtMI7/aJiIKen9J6EzBeLE
9O9P8A4E+eNVuR7DB/7SNviEqpzjrAaYkHe+sq/0BW8xUIEWOMIn91zGjtT+xTVzuswneUIoV7si
x9GlbXJhmqNHOPmlYWlQoARGXTwOTwkArXkSb/VjxR8WRFIXozm0FgCegvj/RrsQPAFxuUuLomEV
PjaWqkMAOV7M98io2hkKK+3UG4N6xWeXGwzD1Q44yazGdx/oeHsxYL0d5BQT4Dr7nI79ASmjeOJC
yJrWiFiYfIRGGGhn4t1ZkxYY8GZhMABs8pLW4Xmi4EMN9GG9MFkVzaVxyYgfuXoyAbKGSYDRFbGi
u25V2gqw3PQmwWpRmqkLxaytD+XD7+DRu7uBRgn2tJOk3YE/gS+jKNnkKzlpyDXMbTsin0gu4CQE
EZmZlkUH+Ou638CJWlUGyO0N1nfXpm+OIxXgOs66wAtZdtV823kyXzQ3RTKOdOB2CCS8gr8vYQ0Y
WYXvGyzn8sOUfonV9NEwo5w1rUtJ48LHBp8OLjE9usaea/pgzhnq6/m/mSIfoqev69Cv5N7kWXpq
zowwHIt+EVa8hkwjqe7kA6Qhn1FfqPahPxNf3tpsDvsuScIB7Jqn57FAKPMGceCG3O6w+bBH71rt
73V/5u+d8EcHtbNtb8KBn0yHbC8adbxtiREWa8ELP6XuDoRpeqrIucK6yZxmV8+AIIO4dUoBmAF6
Ufyft77DM+iIpzelkySCcVUcJ7j7r2lg9C6wPMpk4Lf3ES/mqfbV7qsGafwvousPE3oWyEvzk00Q
8cy+RMUxPzYiU3hW5WuITQz2nhD+VRAxzQuVpTK5sp5L2oNBlkwuS0ReP/9LDGRk0a/AQsd3Bo4E
nX6s7PLK6OmEVag9ntLqnjjroMWSa4uj/x2u90RTVBU6xMzi/t1kjrh7BRIMVXiHgMFjZ5Mu8wN1
MpL3Az4mmW5SPAQ7576pbeSnG6CTIjL41Rd8OJ2VDbbq/xCP4PBtKWGjDepP76l2vZ5XW1BY7Bb0
FU6gVriDKiVYxzrvUbX5jE62er4hgF9o0IGbBZDHM37KJbK+5ZOLWTMYI9Ye69oR9HGHnJK17x/I
awKNBwD1IXtW8a0uklBEQdct+gmnFxvwcMMJuociKAnjq9uWioFkt7j7BrYDtqCYWpil3B4DyU0+
veBkC5Fq/5OgPbtt65XPTxuKlYTn652akwBLyKJymjshUI/chmQAWQALENUFwoLuOk2cCjiTU+wR
OXVedAvCFq7k8OnrFNC0s7n9+i3YYbM2BYLWblehhP+et4AvR0cSQ401rCIZf5Dg2vnuv0TvwC1L
XApjF5gAMro5W96wghwdNwiRupyyEmEiX6SKZrZXNOHmbD5yVZkihNzpBA5lJMkz4MwOhUCEFLs6
jkU8ROD2IKwXhXSk8F43DrPtUzycnDleP0vhv3coGTJkBdF1HYiOsQ8TsKa9x8LTlboH8R1WFRjK
wmoQVt2dLdAHxx7ZKM5zN1wRl/cv1XsbSCIKV+rw0sczGYRG2zXhvdUS3etP99tpQPux3G/X8CpR
nJoFE+WeebB9MOIMJFdDD0Qrzd5NkVcbsHNqS6I4im8TmlEhlWn5UZyGP86Th7y/dafkrSsp+31e
bU3JPsTWNtP7+G4v0nRv4bc/jSsz1DXQZevRNSkuHoSVW6ypFSvrz44e3XJQcEUa18htpRUIGUMR
TuvLGAbWK5XbRgZjbtmPWl0S9z2SWRBOHiKewKQwTy9rJDfKH4KPpSAT9juUzFFBPC7zGRX9jHfF
UUnrxKzkUfr1vN8t/CT1pVpqdBsrEIzZqNZuxvoWvIifRfyFW7psfn5Vo5pfV2wfkV9qhT9zLo7u
FnyeS9gjsByZUa4psMNhen6pVVTvwcO2E4Xihl4qbnRMn3LGu6FlX7Ei0qM/YwV78kH9HU20mDsA
hD3UKvJY9ScxcW8cJJMoWfCjUlE9LD2qpYcAjag/KJCriXU8yNJ+MU8XxMtmA8r6YCyx66U9ypAF
SuXaEqFKighGDIA4pYCKPyeA4lrux11UpbjgEapNZmgrVcrauKEPH460w/215k2ZT2mpwLbLIYyt
UAsUsaYYhvcrvNmKpVNhekARSHAy0cWF+vHGWHKpT1YyQOTgkL7/8XF3wDJelfb7m8Ka0Vit9DOX
lfTbG9jWUxtRyOXnL7+80cylvlXQuJcc4KeR4i65NvFhKAAtHVem4ke3fcBMUcUkV4tFXJWR+yep
qeZJfY3c9r0ewGzQRYPYDOdTbrfyEhZSPOWNc8jo6/TZGc4JiC+PCGolMJGtIVYARYbgjPjG0dHc
djDLjGwz5MSqkC6h4oQNhSxiOX+1lFj/eGyIahGAgLzkAkxWa4v7MwoSbKLc0E3zXa1qSkaUE0MM
v+eh2SIEAopOkJjPYdb/qHHXXbusHurkV6CjOyFPWjz6WkRCU1tdw5QUsZ2INPB/iFGnbBrvSBqY
okU8JG7JQxB9owjAakMpHZlXxucFZEpxolgERqr7MTNoiE5tIrjpKy0fjmhrR2jL7Hgw9TP/oB40
sFlFNA7DxSKzDkYX81tmZ+0Qy2oTbopBPClouxOPe8Ajh883uYlEKKuRHMeVYEvC1OZYVMyz/gZZ
16Sinsm5ZiDyhnbY9OssEONtS7P99iat8VPZqvv1Fe0115CoFJFWAQ9/FVAIx9YpdQ6kfum7lEQk
bRvwfkwre2a+a6gxTYkT/hk+azohS+C8QmnLHBzxbzNm1PtHtjXq1oyD5XpGV0FTe6Gd/AH4jr+x
smFrSINegTVflj+ktormR82VMYOR66aPscpoeLSi7jO2xJ4vvR1EGa9HOM/h20OiQU+IapYClMqK
+y9DwqWopfmKmHfJrHogaUFtSzNnwgxN0XIcQHg1+7xXAPrJ2DM9OCfeKNFyHJVeyf1pyrR4pFFw
n2Mn/WCmAGVZI7Sgx0jPZX93dGhosVAouFmrb2HdmR7DdS7lU4LX4CkErcm9btt9rpDt8YF8o7CP
yBgBI/cqDF3AdTP5OWeXuYs13plgpadHf2Dp+gLNuJrHVSNknMMEAklA24XjvkjnSg/V51Dfk2jk
ukCTi52TAeJho78qoEvDvytDGluXiG7uGHQyUKJMe1Tkqo9OcWbjWY03SjQ4FbdJ82NlVqJs9AaB
+XOlDknoiw30Cxp6/Q44Ih1+LCgYntLYBGDQlzITYzyplh6/GUSEWR1JBvKQv13jxsVD+/RpaMsw
s49Hkx2ColY+37m/iRWjiAoeI7oHzraenaOwRbtY+11dh+/+OYPVwBkFk3NmnLK5/keeGDtlIrSi
CJ5QCC5est09/ako50z8btsGi6ZItvYVDHepD1ZCTjDxF8Sl/upPg8/kAhFsZA3sXRtx4gmGsGd8
7EBV3zLr/aMGG1WfQEfe+Yhi0MblO+GQXTnUvd1RN+G0fz6XkkYuvix/pYPQk+blpSELvYQ0Jyzg
obsG89LhNI1g1MdieNPRIzinIItlx1PobZgDfPHyFtlO058AGCWU3W3MGwVAP636fV/fosR5qcHA
zaCtfBG1Ysdk5w6Ql+O1zmVtc6vOvBmcxgPsHM9bvZyqEVet1J6h+pRDguV2m27iZlqcucubetyY
UL8ahK6XroZnn+dX58PC14TQeQ2rbhdoPbc6tstbLD9kbihJq9lVkYLFph3a7Gr9SzHWVfoBrIqR
RXLijLjBeRHnS48yzG+6yHU/MeW2xJfnfTNrmm3Pd+fE8qeoI+PCwjvV43xnEEkebRisIdL8O6/n
RVPb9/7ILgh588taSXnqf1TPhb51tB0d8UrKYq9hcPKU8mtpoptRtNmnJQtVy13MsfTfG+YQA+RO
cd9T3zZdMS5ca/VBJmOhzr0f5U3gUN4aFzYTcIXoA4Hhe4JyinsCrrHNtvj7sm04Z0bG/3y+hMZY
V3ZZjxdAytqeia8oby5DknIgZmnBL/OmF/6Hu5ERipDzgscVKGjeC3EsFwa42gmMJNIp0/rEE0vc
vG3NlAi9TtoLT0/RSDWMtXVfPfrGbvNfcAOsAPq3ebBr/HBUSoxTIpireva+2KKLxSzAzD30Medu
g0xE9NSkTOP+YaIJL0d0Hpv6XYaCmnVPoscracl6qosrG6lRWuKfqAa/eqya0ss+42ytaSaBsLr0
aVFfiw7F8qcB4jgXI00+mWuzlXtAx8qAD1X9mO1ac1qOyD4inwzHpiOcEvCp1/rZAH3/DDk5tv4q
mRuiAfaXEGVKcubSzdPwRb1OjG5fyX5dxv7QKKGQCM7CDYr0atOo9MnUqx8W2nk4LguccZ932lhp
HgXSbSBSn4zNm0saYkrtamfT5NYUYFdl4sFMjg1kQMIoVpUnRYI2XbV1W8OEPZ9LaEkUsmQEgKog
UUGPFf4XVXUxlPaQvwV3KF4rPUx5vZQgk7t203/RYu/cw32ng27IE2shvyAoO8Cwusd5dd7bD+Pv
nlCuqIXJemYIZdrCkp4hg+Afi88KEYgNVIZfEOrkCNwZo2PDXllsriLo2GavdmayjVjwuSMUWSpi
9SBK3Yo18Ixf0mBj3NEVV+8ZYg3XFVGrEUvDUJSsKhHqyAvzFX+Za+tX3VwoBcwtbTw9ov8fsDlR
f+hynhZUGuaQJn+c4SHIPlqJhThSG1IdGtEqgGoMAR23Y+f/x3avZjoPRpX2N11q0jMO2Szw3VAk
Z/FconboP922t8nEDMGdeehGWi1VwMavg7ExypPdsmcIcC992XcDaAjp7HQmOzT6YP+bBjFr/VKF
F3vlNYyWlgPUwLwwo4Lyh92fQsk0YvSKb5KkUAbyZaarc4S4+lpVVrgzlURkIDkVLSw8JxnGNEux
i1t04rucGI3YuPc5zPYJDqE//DKfHKYtPyThzkQi/X+HhS2BOtwAb5WZHd++xLt/lshB5RqQzSPN
6tyZSOfYNtzN2Xmni0w05pgNpnbOOw65bEk/o4sSuzpCcsk8IYTvwYrO6DK6MmmlfToHEHW42a0O
Kghzlk1qnVHzJlLWDOZ0sc6JcXxDE42IXARoPH/Grq2MW2qpgdYeeY3WXIzf0DIQbocQvPUFFYmZ
JSyvTntV9HQOe/CctyKWUG8X5304b6J6SIn1WY6n4hPS/T4Rpx6NGBOhr6uReuoDIn9iEmUA/weS
WKMTRHP1rD6GwK52U00T7A3G4r72AenvyGank9Y6zfvLZUeYBZGtNM1ZXmsYxKPwsMkg1Pxyo39Y
RaT6dDSSrmHdc4DO8H05d2UPK+qSAad/aH1upKgWWr/aCUcVZufZrAR2ur1zOpnJW0W3zdPtwI0h
j4w1Ip0shutF2QLOay+dOi4SZMWl8MdmJ0bHZD6Gjl7uU+re0ICqN6mLA8qbkrh4Qb7gs4Yhohe7
a/3dFKfzuB5EXQMG1R7MPCXWOMIxykXb5ALObZvn2EvkCSpcmHgIucUarPAMi/aUos0dXzEySy5j
pQlFEfVU5nNiKMZFHMoEYfdASfEK3TxmNSIaeLis8qYDAUF8hPW3s7PBKFSnfNzsRgdgl4t5iKpl
kh23ddGaRbouW32UmkSOVmIAzjVSYTOWBbTqaReK4mALpKIYQvENpAAn/XJEyaHXMj+ysJik4wn6
4IIYtFvGioCEcBA/pesLhvlXNlQYgXbsNmGk44f80cNBwP+pboejSRtscdekhS5QikLiMRAg4Wk0
1TmSjRhfu6Ib+YEKgKxaaE4AIwLaY6CV62qEV53wL2SZyixKEPWUPHdGCmi5A+AqGz4f2tvzyzym
CYceNfYrt7x6jpCz1/vj7K4aBoAMxak+d+PFNlRkQLZb2e44OFFWH6NkGaPYs54l+LlwJEdPgGeh
dZ6o3WV62+hZGv9I1f++b+DzP9F374e1lvzqXaYEnhgbJXw57HlVlacuXiKdOG7cpkuQ2587zFES
5Q+x467ngFLCmouXluHa7TYrOVvQXnTjCEFDBzpW9mZYGFop4E9tBEPsAvsgFJQpkX1JCdUrFL13
Anmg/obaMREJYM51mqw5uq0jB+CWNrnUEBwMvICFKgogASs3xrP+3smPr+pUCfT+Df0aJNAz35Ep
/am9CNxVszXv8Z2F02t+o2YPIJwQv5Pn7yhs7Khh0HhMg0/fp5IDP/Dx2rKHxPg00DAVtaVPrMkU
UQj5CWXYa9OLppwZoq980wrwU0/rfLkwc3R7nkrxiloYSCXjXRQh0hjR5UwdJXXnMbYkZz5s3E+B
dinVq04GtZl7pQwt2SgVmq/3ZgsooaTYkrHi88pA4Jdc0MI0ndSg6FuDHpwhOkFtaQz+hPfFZclI
Wbvn8rfrW+8WByrNIpMxKxioH4/ZgzzAzGN1DuVzhighQQ24VjNsp5wIS9SqGV7bwMLQScazv3uV
xbqIawPOolaKEIpzxZw+puYZmrDVwJNMcsPIy6afJ3x6GkMU/aqC73yPb9dhg7E1tWYdcjDJkjbp
Wa/ecpf6p94fZ1yiV7HcKSoo5C9QP3+rzckSZIeJ1DI5xAky96yDXv8b5Xmy/0SBqIpDgLFIdhBH
3JDuqNo2ou42svc2P3Dl71e+qppAbvabLxJVvTIlFKcfb8XOuD7pLvkY5wuHWD9Lalp/ftj5YIXa
afYiMN7wpiXapHSK5DrRASePuDtew1+JA4Rvli76NdCM8jNLEzNDpDuTjoYOp3MtiRY1qhbDzhB5
Kqaw+mqlf4ShdreXwc24k7V1EwIxTFWfWNkqxtKXBvLn7KJ1xwZfqoMynODFoOZwTIOo7Bm6I/ec
CVjSPxNeo1pnVcv4T5e8jQzVn2l0sED3lcaspcVxmTs9Rn3jE+VxUuOQFu6v5Fft/uKt3IKHli+p
NdLdxAc361uJQhV+ccOSXWzwKXywmbaxH/dewSgFuMyHXOtcYbeg3YjG/OVFFwHq/stDQS0EjVoK
Xld7e8f7FZy6AVkHd2ODWarF2ngn5x8CPrmnckZuNS09B17w1RM34rFxFmfIhldbO6duO4a54Jl8
JiM5oLkpH8FGRQ8FQNvEcXJLROuLhCD1b8Lub9C5kNrdqXbtBFRodOwh73odgMzFnlvR40nbsFC/
7PX3/q1fkzqmch//LlHg/NqXCXzjBEzNh/1T8OHsOY2IOpzuAHAOpxzCqz73tVCE7ZvL3cljPoUS
qbG5ZWIUvWi+GTTFeYshtRO7IB1WzPwJU5+JOfmz1ledLYHt2+M0qk0F5MWSvICVlnZSRR05SaD1
B9RhgaW3sBYt5SETzIvpe6M8IKf7RXy9V5QHX3rZJLO+rA8+7OEerLtcSHN4PxEsocESGSq36EgF
R1S8MaBiFUlBcdiXr0mZ3lclE2/Tr4UFwkaHjIaKqq9IL2BLJiSuibiXyruol03drZ8iwf6GTZcC
Yhz8b+oejh37QkPKsFcbuHG/hZpAp1VXSlSdribuUQ0pRqOKuYYlIMoUGqooFecTv4NnL4XhyVIj
2ixgYV1sS7FcIlzjDEAEXCNP0VfJnrNb73p9j1CYc5Lj3uRIYNHrWImaNU/Hvm/BCM/cUYZ2YDic
C3xGPZOO/aCXgbGxXym/7Znuu0wNz9jcE825qO0ebEcr7F4Ytf1CC9xiJo91RgNjtkzrzLrBSqBv
Xzb/bWS48S0/kYrMbmTH2ECWG65n+BxMh86QgBtOPYqXsytldsugUf2S5a/iuBlNfivctqVP/0sh
ixLEf2NDSQuyDNyhG81i0IDk5mwgoiexvS9FZAAa2bBdtMDbw92VdgTp2aT8RLIhhnroQgX8KVgf
3NYCb2dy/4qTcpOXgYR61Y3TO7fQ1VPrajBAorYy1805W3O6lx9lLCJYQN23UatrnT8EeiZ5qlPQ
rDdjzbaTC/i+gPJpSYParIgZA63SkWOOaZrAy7kWMIDMLPv37r+iSLXRDBCM5/URSdqaOW/c2FsG
PHma4XaS2GMIJERfINczZXYqkvkEaDHOpYc1IMgvDBUEqvF9r6D746ZXSylqeH0qFzJZRLFsNjAy
uU5DSsEVk+lpBRA7P80gZRRq/c8sK6sCnzqv7Mp+TchTM1kSwQQnprI7DouYZFLJMc/hcxQEzLq3
S881/YTahwpp3mxqqMJ02UdZCL02T3FY0KS1KVg0wJqOUwLkOxDjANpkD8KHqdNiKxzlV5n+fBNi
S5Yhs/xcRUSBRjTZz7kUGdxJPsBTBZx6x3FXeA8bXsp+626qn61wEQQJILntopX9W5oQvNf5cOAq
bXNHJBhuVQ6aS+g4DpWz6d6s7RoUdT8VP87IwOrgYtDemhjFfFob3N8dNgDtnyiSxynJQS4upV/x
2cbV/Qbq3rixxfU/bN7p0YjS5fIsjpJTmi/PDoO54rSRNdxG+zGkFjnAqzDSKE1iZW8ZnAyCfSt2
4a6wvdFHEkhddke51CqWmDpS3iKfPzgymCRXcm6RBh0J4B3TgnGU+sv+6eaRvvhwhz3wumPoiJ2N
7hLXWAkxrup5rYExLZZ5ahU1QFQgtoZhJo9ZnFZ04mc4rD5NA3HAclvKYT86rY9vEzd+fyP/6oKN
vdZoeF74Osg9VPOH08TKR98uaHYH2NXUzM5Xiqu24Q/q7x8ae2UDBxbCA3lL+HQ0fh04k4AW9Rc2
+TN6WnDgyQ8PTgCvpoTnQsN6P4eXECqCnceB9w3NyxccpTLLxOvhYcBAYM4/zUTJtX6A426F5kJm
Ub44ptPVnraIieW40LtkeO7YbATh1HXTLr/oKy9ywdTJyNvGVkqAN5/wMP7ZewTyrBkVRimGThLm
rXmj8fmqjiwR+Z0fbV+aWWgXO6StoQ+pJcZNgxaObI6z3MIzcWRvMlGmmjcs1C6oeyQpD/ZLy9i1
dKDQfVhtFwRdOvJIviG23CljI+joCMjYRVxryNtGRClHT29e6W772GAOXcVSThmmGxAaZd0KOZ03
VIc4a45Fvw/czZ8Vq/YBQ1AIKKtRD6K8DUt05tOwLMyERSebSY+GiKF9T0UmYsZiqEzCMtPOScPz
FsVzKqf2MDPZ/7n6+a181jhBJpULMTk/zSXXU+3oGQcQ84Teo2mkKYu8xQN5xVwZunjbknJX0QdP
0ozQagARn9ZiQFsuCNzGhAavUwHG5mAFjkXd3QcNkTFIRBnJkXTw22BWCfaOoeR8KaFQDTvGrpLQ
6Ncyk/vIe8Wbki6YVV5tnHrR2sk9xoewwfCq4OJSR9Xr00hJ1g8bt89azJXgZTeFQGh8Uag2da+B
wH8qRc7tLCJxBiWPMV1rMDRmnUPejfN9UhURR71aZ1vXrx+uNOQ/x4o4HrSgv5SQyp9tVdMe781y
GiemGQX++MUemuNia6Fmh0M+v9Tgbf/zr0TsE+H0Jp1XJg6RGNOy6pUVHnYQpK9wamJ5NBZ4opT4
k6TpgNegvAEcROAjXu6iIh4hlOxXikQ+czGCCRT6ieBqpLgIPMttJc16kYeBTqVSRCzKxCbnDzT2
AqNootFer1VIqwbww/jsNdm4KQh6BgPJorJwTXirK5lJF7m1ySUAdmjOm7xzIC07v0lVvnshHcOW
vwkBpA903XGy0p0exZU8bCa4qxu5+9317O0Q1B5UXJUzCMPpoOWpScKPF8AkcUMgnmH622Mx0GEP
oF5xOEQFTSwLW9TKndMfdvjl55AjwQ00ngSPyBAGp/8UP6HAXrXKnKIjnRAaTeViiefJ7YrhxXU3
JzTiSy59T+p6k09TJHSq1uy63tl2TzevRIFU4nmUzG5ZdxuNi11G/CAWgqMbo5vo9E8cXaoy+BgD
iXulIPp8BIvJRTZQpnyTCwwI/1R95J0PqIkCqZtbYc5Ljo5NiBVMORLhKii0se2h0k1pJYstSqIg
9VW4S3b5GuImv5/Xyj7WwajVTsf7AOBvrcZpmQunpjxLVQAeSHGdr6Nc6Aec5bZO5G6nQHnwNc6A
fX3f7va0CbgSj0rKfcl8N7yk+3Wb8EyH7l6DUcvdGA5AY8l712Vz/+Jc5jmuUT2kqdjwhYFecmXl
8EqtaY61+2XbvYD69n3imwCuf9I4XepUV2vLcl0H79fQtvfP/5RV8su81nP1wq3Bg6fPO8dybGMh
WZ7G2+qUTkgMOXh0ZKweTAZbR3Lx2pyUB2VFjLuNUsE33QfM32wq3r+qHW4atZLW2sp9l0YEPxis
1cvkF0BeLuu1IuOs9dMmyww/L0B+FVaZvZKt5lhVym+G8T0T3DV+tG8c94qoFrtj1vnK65mRqYJh
uQKnLtNUFmd24G5O3eoGlwes0vwZxAHgNnuw3K2fBhlGIF/uqk8l1Qyuqa9HWarL8HYoDaE87gd4
292nwUq01xsxWdSbN3Jnd90VMwXF7lx2weJen3sgwUw0hC/jmcQae+1o6Cc+LQPNJyhuAqzaE3Ul
KoziKMCw5Ayu10ig9AQ6smpJu0Doo8fz7rx0lumImsyMOf8hTxPc3u6+TqG7NGUyaxITnmRiFr7R
Y/Ng56DpzCZBp9kv8W591p7gcL/eo3+k1iUzOY+fvPw9K/v7l2w9PZuWfEmjkmMLymn38l6JkOi+
/y4Rar2yuxyOswSR/GA8ao7AwI1/oFwettX22tqziIGX9wXH56jKoNkCo0glYUISwEVoVKN6Er8j
DRRVuPdbkR2+qoY4ZR9EZyfV2Hzy48/Aoeb4ou8hq+EylFc0cQwYuKkf1V2Y8P4pPO8yRuyWb8Ga
lr6KKbTa0B3F25sk7V+Eaqru9F0iSnSZVYMi4acBMY81auS4iHRsiadQ48AVNmscmJszrwVFIi8v
4TyDOE1MbceKgdmjQ1YCJCLVUyMtGalVHOEINSmtQ+wUNE9zyMDBxMKAZgUG2o1peAyVxGAFBIky
WOB2gj6gOiYVL5VR4L/E5LmYbsMq4akCxSfg2SlbxrAsAsl4zwlLLblDbUxKnAHTV3oD7wU1CZns
eqsoma+fW/aMpL7UYdP6iegxRymRx2W9t9b3eHj65qnLhb1lT/Ck4EChlkXxFT6E2L0c7pgaihX8
/Wj3/bzGIoxM9cXyLkf5/uSbpVse2w2A3T3vBd1/f7oOLbeVhhDU6kDlnd574I9U/Wuk6TAgejpI
eWQXG6vmpIPu0W9c61wRUnat180yxEhEsNUsfo4IKG22sHWksMT6waO/yFfolQ7Y4Cp48yc2WKPY
7LMR1x04VBMwUvHU1nmXWAnoBqjZZp9LIqUv2tC+E881H5SFgXr7idAduHpQcgai0YouxWpyzOIo
kJSoyf+C7GuH1/zOr7aMFGQPLKs8a/yPKF9etIKrCIDiPObSuT7yBAlxCk13Ldw6t4YghYivGwvQ
WeZRJLB1HE3u8Pu/5azaOCQA61GCmIQZbWVjr1f29EHJg+eTprEK08OlXWmEOp+5NDH1EemKzeF+
MJ6R/+tOuDYuv6LIlp70vDj22vnOt2LBU8CMnMLbdcs+eNA8bo0HdgYq6EGQHbXNUjVt/MN2ZipO
M0MjB6COAXGwD9Dsh73P2nXYRr0cHouGRpsl6QN1ZLK7nhqIM4hrGfeIzdTaCwcNTuZD2U7m9qpG
c77dG0Log4DJgkqswds9hXdrpClrvkQBPK7Spc1ZjLP4vVqcZtSEDWeYR+02r79nWJyl9vFOIc7K
QZAbMLpV90KJdr5QOGyibH+iH+7jI6H9A1s9Jk4YJPA+nE4ehJgdMlalxKGI5N3MGBYWvbt+aPD8
1yYjKojtu/rRC4D7z4rRCl43th0lBE5/ecDgDn2whxr+QvlXPEf3Mqxw8Xly7D8Aey+p3+pJlfU1
2mf9FChI6sA0XYCWQ+plfHFu4Z9MYkK75alBEiXy/ApVaFZw7KEVenvfWomKyWKjKVpZjrrrwj+R
7hdEjEPCmvbDAsqIc9AAk5B2UaWoMmtIztQp1cvR48Xo4wJbBZ4NSfQFAS2CClYiIpAR0VfBf9G/
e/+7BKT0KfP4Y4HQwpd8GzsRGePwxehXcDZgwpMMLSUek94Pnr/oIhtrRS7W3ij/akqYeb6bMdZy
nTNZijL4Q+xkrzTFXOv1jF804CYhYk08OahqbHFaLtDuiL5xk2vHtBGgD9SQZpu0a9ikLPk2MFmk
m8m5MNOFlAwbujTv2dmCKpAlpNon5a2R5v/OK0fFnGV5mlfJFy/o4o7Et9Aq437stVxbHrxJvl3l
dnxoLNzH7oXjmn0VC3YOEHcFrcW0IiSKwlAx+NkbPFxiF45lmiZhsTauu25UP9olsjv2gVDVxTEM
A0cGrfbFs2olonZ0AW0miMboPE0ZUXE+rQBG1T+/gPfl4FBWrj/u6PLXUgGgcbKFzB5HJ3n+8SGy
duo0Sq7nIlkRBS0Zi/xAVyozWvM6suw+WYTAgI1NH6B2He3B2FMdRgONrdvnQfw+FC/s+h7DuzI5
axVBmN/+1oipPQl4gsgDkGHAV9yPlwnuxaiLLftncJRq46upR6fMLzmVc/ODgMI1XSVtD7Yvi8g0
CMOheLb0xsKFPZzgjD7P8/HxUuziueS1BlgTbYlJo3xhoRfcNmwBmVBdlLMXHVbRsWp1PYzrfVol
rZ0r+qolnDIvvLGpu8Y5yKgkRNBBjAFTkreklunyHYgfkZp2pkuuooE1IZ5F1J8FccAexBObeR+z
GMzgCgPS+ugBWu6H4Ycpdq2eC9u1Hh2Xn2IALIa0+WWzpneQUJAfRLpUon83ZybIPmKDIxfpm6ox
EaaeHprmvz/vGNuyjpqeG7zzkO4s1iZt80roeDwG/HKtYu7xZmvtbL9BvPl8O7Mcly9LSWNkJ7mB
uqgKrbZE3/5A/SQ2K9Hr3rk+rZYZMsr+wBvv76zVjM+DFEXotFQ0rKF2sDPs3v7825NWwO9Zng54
l1HM4Ojjk0OUC8bAWYY7FhJbPW+iDV4dNXYdCc7Mabw0HDkJIz0Gt1LajwW+dfdJ70DH49PW7xJL
6mbWEDTRpzKhYqkscgd5q8P3jfQBTB5FXeAa10hBHxLdjXfWND3NHxGjXddqwgUqjF7n6qvaMNVE
hLrIqIvWD+9SdcB79+qMdFU/RH2lT6il9RkbCmkhQ+cEGAmb79UnHU9DMEbID82RPeovgnYlP5MO
ujSXMzPtRFZqKziY1BcNMi9GdVG62XqIp++F330nURcbAG16IJTaDR0BP92z9GjlM1DNx3GyGyRU
TlixAMo2bM0LUpPt83+P4aU9GxU19IfWBIKfJ0LqS46gKo9NpRcHMfz5/ouHfOwl0KcmF+38gsf1
RpSxEtg+ydXkxl9qoPicnGfNXOSQK0WtlUCQk1YhnQ3E2ZG4SIuhe28eyhAFpGC+19Ucfdqp2fNE
1Dq2rmmUU2Z6SdBgXoXL/rTl68KrpCnM4YJK4emaPLc7eK1jlx9bwX4VTq7Htptlh9+FNdLifFJk
+2dvRoC061jby/n9gz3y8TMo7IQlZGEtQnXi8PX4M6Pc9n9COIl2PklzahxY1dM+2zeLlW3WmNal
O8wl/x1fKoK5WVgnvNhDJuvSy2DiB9U3Fh11fu+nbobK8nG3jpoELPU8eC1MLJ+wTCQw6htpHPpC
RGIax3RRjebWTiHViVJKrTfSLjUNk09lNSN2v9Rf3XPtZSVGBGbN2iipkEFZKjocONxwPNJE3+G4
9BJoebrh30stCsM5iCzaT4AhjL+DH4mMjznwiO04WD3PurW29uvF7rgNORu7X9NxJsebIdvZYSyl
TgTZWlZ/hDAHEg6EQu5bgeJlMVL8WOChVZZXU+lUxpPXLuHRbY+/IPxFppTQXbGGuOPpO1Gsytiw
uEavLPs9bRCcD/Kz+fVRxRsCGeLlgNLbZtuR43v2hNSQP3NaE1VZjl/n+pw/QF0ojmBfrsQuegiX
Ry/gExIqNXwTsb+a3djT+ZqgUgPTTSrL6GKUZLoLfxI6lQp0lBFwqbHqPjY5uuk8PjNwBC0P7H1J
+jvdduC0Wp8xt6f7Ek+binIRFn/IxVHNE1kRAFxZyA3tBDWv/nXTdsc6gDmnsYU+bKJsfA/HUj6Y
rnGkoOaJDnfRDakWs0vWHhc+IcamEUR6o5TVRTFOC9gJjZxEL5CxwcHHVIzMFo5+r6WRbnrI1Ytt
OA2Dep/dsL49lfVau/gg+mhkInhFqHw03njaqFN9MO+febXZ7N/o3fwLJ4Gx32PCOpC5jrZ4s9ra
bnMIkYDZ6qT9TQGn05ylUm0yjl85mdqHWL1nhoRPSFOnec2y1/REyukzn/7HKr9OBfWZvqv0hIln
OwcS/J+/LMSbg6uuXlJvbE4fcXNnqmrLsYVwWQSYLqBH1prqndbptyqx0m+WbDfxtIk2BOsd6gPB
weMx0ctPuYYaWydksH1RjYmSbUrlOI72GVn9oBMVtsiTw4CfVxGbszw3Q4z/Lods4Di+qgS1L7s8
OdtK5q0u9zvAy8MxOUxqDXekymxMtgsEvH5L9FRXA/PsdkiNUYusSQthtfUDBJPchO5RfNgJNZGL
AmN4rDkRimVJDN7P1+n9Yxjo4vvRFMLtrzQ+oj7PRcI5MHyGhQ8qcXIuH/Fuf0xbw+uplxmVRx2C
UNKMmvqgd9RaakaCI+D3ovm3CCF/DseS3FpIVGfD3P9EdLfx/S2l4Qk13Hnc4MpMULEWPOF88V7G
bFDU+kRd3aGrpTK2oXkigFukGMRY3cTWgNFiOQQ260A93ulTOOcPlCqemowFKw0gZEpL2drEutXh
PhMXIwXGcPSzJPanjMK7bzTYqiHVkURhM7Whmn93dAsLzWXVRELbgv/BoMzluKa88/TQOs03lmHW
DfMKUlYkrNseuuCT/vFmVddoGXjOrpxLntwmfZyu++B4dPK8Tk51M1BjqaRDgmedkyIFeRclxIaS
zDXs2PxOtSmHgAQJaABL6FIT2RYr+JXrfYnTIG78NOjR02aF3Fyt1tjh7WN+r4zJVmfhayPPLdPA
jKHpgjL2E5eEp0I4tbBogqxpZ+JzXb4k5a4fKTg3NI4L8J5BXI46BV4oK9PbSy2KlH0saj5jkyLC
HR9pvbayvrs0WEmCNySXjfBgCEhN3xCOLEZfqLn4MU+SEYdyWz3KU7VK43GiVwfhLJhT2yov11UW
eD/Kbw1z/sD1j6M4zLUd5jR4kt1oP7hmY9T5j6rCqcIbSRHlJcY+VCKeFwgLftjtL8PpU4ofSNnA
jdxE+zz82U01h7ceqB7WWM6Ol+I9qY3mDPXaIVEHOzHhiVRTplm7A54OaZNswyM0bw7DWNywc8l+
YRC4/sA9U9zrAMLMbFv6E5WIRcs5ei5gMt11d+mzvlb3l1rzRGNOdwGhSZoo8iT391JGSc95tfDK
8v/K2NFXuwazEZKaewyG15n0t6JsiMlDyDOQYazXmdVmt6jktbg8sYRlQ4lS98mtNsekWTIh+5Iu
Cf/psZpTGkHjwYwOVzr3Vlke/E8wR/kYTfs9pLQsFlPw2uLsB92xolrU1Dz+tu8r0PLWQ+WsNy27
HxD5HH62YiFlKd5gBoUqNC5Zk5URVbQ+pWHnPOcdDlg7hb6E6YjtYu0MAUUuomR0pFbyarBwBma3
jEAudYcFiCLLRf1g/eWDECZF4PGv7WcjdY/td1Mgbz+8rY+YrtZiJJGZ74+B7Xg83Y95mohaNiy+
ucGWtcIMA+adWRf9PEmjEzNY6gmEjHbTkcef60b0vexKs5+AEA3cM1bSuFyc6scDRlJLSkLAS03z
KAkaNxCMcQWUpBsHSXoACe0wn9V5OhsoNd7VLcb/QUZALW2hfDReozB0uHfYwsXoxVmslxCk0hZb
Jhe/nPuN3ETAz+6Hhmb/lu1GnWReF3wBysTx5d2jph+qbGG6zm5jjgG2ezZKpIRagdu5e+pxydQ3
lPHZGFslVOVcz6TlqRO1bG00P1FcFB7w826GfwUYS2Ni2xSEWoX07xEtG2UWgLNn5tjOZXO3l1gx
rElDs0Is3S8X6nBjCMyvm7UHtDdy8iwLVhDH98pHKfDbVTHTBOS/P2lh43iv50Pfl9C2ItJt7HC4
KPGjBhV5TQr4nq6+CahMwBQ1l+pHQDkK6EKBVIpfc/BRrj9itE1T7P4DMuzXMSCXUq+mj75cjqnt
OSPlDhSf0+ZZ+5nEqbwk0sEdAYvX4yFEByQuMvnM7xyw4aLtOlM5gW1NMnP3mTnk+LsAzb24g/i8
mFgMA/alz7FK5vY0moyjoIWSSLnapUUMJPFn5P43LN+NeVWyGgT9/MF2KVO5u9OSNmCPCcNUHz9e
0rGNojMbkjXpVD9HOc6zBO/9KRKrQRQBZvox20zAl98qp2K4URDpj6TPU7fxceqvKw4sgzzXptU9
rrQroxBzX4qAa5MzvWt/SObgsGdYNKODV5ESDfH4lobFG4GvpJpSVDnE9YCH4l3yvpsQb3uWwNDZ
X7D7JH9SSTMAm59YGUUZrYKZdQAoKzMerOm4p/Kylo0+26EptOZhV6jKeB4GmQpxqISGm5Ctdpc2
D4+7nk8tnlalGcoSEdd0W/PwS45ml6d6L+KZUW9ZMg3vEUYUACLLvw8fp6WLDRG3eJNaQiuW0F9O
QJ7MAeqiI+LaVGes0xYxGNvnzfWLpBcF2atcdfo1YpqW4Vg4kXFcFR7NhJDrdpGBv5GoV+u/Ehsa
nix4DBrIpqJKB9ORGNfOVdbRshZe0PVwzKrfJqWy9IL6e+vh4NHzfjRMaM324bd66MhZVs+0o7J7
ZjYVVfTOhJngSnF5Lw5lX+KcFVLld0aentPfNxiOYVhPW5n7pX8Sjek8yd5XbrbAoldb4GGPxhsa
SGywKw3qdfVhz/fmGoS/e2lBiC9Bxnw0xifYyovIurAXI1cj6/a/IB06wMSjNei/LDrx1TOHRRtI
0QdCo2oOglC2Kyyn7eOkYDZ8O9TpvJz7DoF9+AQBXBi06NCdh7SgILQA3IAT/fFe1+jftrcYQVl/
SJybte7R1tvCrrbY9LUyHAvdYm8SHYtKsuQpvvdOIPPYLER5QJTfyrb+DmXj1yScVavwbVvd/Wds
YO0U74NsRpAvkivRJRXdAKgzIIseSwEMKZz9FpmznsYRmo96zM4s3Hc2NgUbiKXaIBxpqx5F//tp
RTwsYoQ62ee3s/9iM9l+18LOJzVM0tcQZqX4tEDsAXrGljVzTTYem0nqUPo6we1WhbIm6fQufpA1
rfKzC50S3AT37dVHFpe2Zi5cquKissJd7LfGNfJElBzxhhtXEatAuv7LCQKipa6mewju7IWid2E0
eqG4/0QEu9VUgCIhUP2xgKonmrCW4Jobn4Q+XOGaEN4fTHIb+kEK7T4FQ2CK6JMehzxNVRcMtA3a
ERojZC/kumRJS1r1weGBLI1/c37/XtaKH1g337nTfx5iIKp738SNty2uVXLO+VtCG5K6cp0IYWhS
BdyFsypFdEQBcmst2LvzkE8kJhrh8rGuOPitpynD/N9GKWudrTVevGr54RPoknoYlMIfjrFD90N1
KGWgCReqT4Zc79WGy9ajqPFtnrWGDAwS70wD83NDogqN7UuRtJKVisAHSJDIS5idVHoQKu+xZik3
pvm67jlt6oZi+a9iUre3XsZPws3YLyYZ7c66nSAC2+3SZ8aAdLJ/z2EFCfncz/Yy5VKAkDRat8ly
sBdeaG6tTsgz+YlMvVqk9uaAAAsEMCQ2HfFm0XKjyxBnZLO8a3PFyDj9fKPyVU1ldVJqBgEYXmYm
TG5Bx4mcPV4kzPXio+8cOmj6uPkaVE8PLhhi+fAvqG2mCpa9npDcqB8/210H89AT9WjLfMayGQy9
6R05XHN2AFSqbGI4Or6r6CmsEREHtextMqV/aLarEcpSeAatYyOU3rcU7vNwdWJxH2E+bOlXbM50
lChwXu4542UvgJEiMinSL98lgsDJV03CI+8b6JugmPc9R3gGnGbDjhzvIfoViKz19o2lKFaHXBE5
wEoMeeFD7WIH9S2DpI2Qb5/Bw6MPqq8j+lvhNJtXpFforwPqRqFLjF6Q1gHmJoPPLG3OCB33qmYk
wG6JYblyFoolJc+GgmoDP4Nl8YOSu+OOe8gP+JOVsWvzEPIOLQkJP+ukFwbjCpAD3LtXUaU8ykWX
3OA8We4M/CF3HYJcuePDqI/TykJdeFllHLxB8RbuRCt6dluPQJnDpnPGILYLR028dNSpiOeWGlEa
iY1UKzmHdr5M1zq1l3M5M2G3tC6THAV93MElcfZT90XGiXnkZKojr18I0/MbB11cZS+92EA7jCh6
hYO7a4JdTstpfXsoaL37JPj4PNKzeuR7XUaBaveJpNqPEhBYoXvLy0D6HKYRapH464X84DxmLvDC
rgHJe6x8335qU8qGkEn/UM90a38o8A/6MHeQu2ebPzYDTrBxG6KewWQsnGBo4ONfskuNy5gZ7cIZ
qBvQbGohIePFBeQKrI0Skr6sYmldeAymMcYqw4Vcc7IXL1ULgFZRYay4uU8yYRx+1VMisNmbxnQC
V5yoL/k7d/vLtGROmcugU/uqdt3royR82jGPMxVtZMuWST0OEKG+Rt8MC8K5w+63uNdyHkDBOGWb
hfJ7jb9UUlmBnljkrmKMdvXlEtwa4RmBJiBbIS6KKYt0Ip0W0yfhJMhxzhSygW0pob6PiEWw2xOx
XOkKh/z5SMNOKqRxT43SVOVg+j8sFMoxrmmg4/i2ecd9h4GnYAI39afnbXjmZZogtXs2/3uIPglx
LWxFxqWEpRM+rtNS3ZF7rArgtWBxhOwxktKNIto0A5nDeuGLTDLyX4vGGiPsNkzLxg4SVQqqTTxU
QC62MwH9B5yAZlSX9ByCK6Kq6+hYnf/3Kk0a4iWeea1yYoush44V3bqDd89QcBTnEXGfT6grQYvn
/L46a2bBbPghW8HGeTyoonS1DlPOUYTAbZR36wAacSzmL49FwwtfKAbZRY71CfKqpMPLHbpCsZzg
NimjfPfDQctNhfUh99CTmwZnPT5P5LV/mIq61F4wqwKo/ewduiJWBYUEw/mZoOPdvAn3yUJky6K0
P0r4AYYs0Py7l5mNmuTD9/NDzMy9JDru8XXZY+SAZjVGvXa/wIe+a/GtIT5RuHYj47cbEIUmJWPK
Eu6qfP+OPGigZDtglLV7IJo5mIsylJWnNRxcd87KSMpR1MfkcKL5SkUbLtfZWvusBYuGNA7ec4Lg
Swtm5VS2UpMo2y/Y7rlgmHccJK7WKcIdCYMeSGsEqSXCjXSr1ygC6Gl7ZNns4z8lupvs3+k4wL/i
GLIUO/LqH/gQ/9j/WweFcNvevbkPoIQS/W5fgZ5nitzBrXQJLKD0otr6UCD78Bs7wgdvtIdSLY2W
P6NjgXOmwqbT2kYwQnfD7/DLWRBOxK7oWbEJZoVHiLGPcjBAQwQecDyFyccr++N4lQqBRBMLYooY
Rxbga0HYrRXP7YW/qLafDE1UTOVIR6wxu5oD5v4iO6HCuZFFW2aa9bQYRA5s6VXKLuhJ3W4zYKP8
gwIJ3Z+SSHpYHLwujf9+aoNBqvIyPjhJfhRwJC7550mpPnPO5xKkjKmF13T/sYRQUBP7d3PpPtHp
nI3HIfHq90IdmZ0m2dSwszbTCteWO/etn2uo+Ej1wNUdj1BxEVkADF/MxA+zOc0v1q/uxLBUf07u
8fz8gwBsHOBVYsmxpTl2rQI2Jp/SHiykHMsI3lhUdgPdA7UuAc/wU2UxDh1dDUzAhCjotlyI6pyc
aymwNx+lMRdMcbSoeP3mQxT/HyvQfyI5Bd3KD406ef+w//7fCMEmOcy2al944Bx0SuwgaDrThuZ4
Jd7SaEaPXwfY/sCb+gKn6IUb30pn9Yzh0mx3y1X64ueaAvL7dfUB7opgTejtwXD8ggo90GJwUldf
ZK8RUf+rOM8tudQNt0xy/aUKm6ZOQSqiDnHte5dT6lmtiQNJOHGa39jj0MgIbzNvcCd3NulJxSK+
Dx18v9y/G138ckaqikEd6xLlrqrDyDWMd4RuBwvH8ULaaRi7BFflFcbb4fYRWsemkaP8OIrhlzoo
uyo+5mYHRh7wwndn0qVDFbHPtJPYuQ+WcxKVGM8WZajgVUCan4lH5mXKLmxqHZ2FwBWSgeqSliTf
zI3B3A9R5EaFPRxL/OqlMwL6PrSnqhG6GKyg1U6UWRZqeGU4afAEPQCOGA0h/vTCNMtdA63xnA0k
tGY1sPcAxcmPqiksNH45zq2C3iB0nq14uaBtQy0z2mLHbIsnDBWvHtypPGyYdE3/ZJiJPaJUKtHK
JqBF0NOdCPEqzPW5F/jlnXQTaEM9V79Y5SOXsNrU7aev91SxOFZEt/SO0z3Fw8QrQtU/8RYGRvOu
NaqmPsbTX2j4lXVILaIUUcb6CgNhv1R/13qK3t+PfjL+PbsLC1KFX4w4AjWbvIzzhMPPn1/C3AhQ
gLjCJviXgKeNZym/3D5VLZ2vfyRXoMIaytGi+gDzXC6EG5xZY3jmjBWDbWugbRxtLm/pzowg8+cW
4K1ABw8g2M1V/PZJLJkiT1rsvXi3hEyAxmcocan19EmlOTIbUr69lmFI8b34fPNZsQYsSdr54BNw
9btZBuHSMcHiZ3KYhos9KI0EUsr4aCxez/0Quh4WjOJylSeXhP4BAYALpmDw8p9Ra7YKjs+53W2o
KyZm85+3eBW8x/wD96MdVi4ILRlNJq9yGcnt7yjHCDQQLzw6b4lEZKxv6G8R3dCglFG19tL120bb
tGA0B+2MhL7wYSZp/Fo697+KESdCWCaH4uze24/s2OT8w2XPIgYGi3e4TC418AUjOXHh89G3dSEp
LsHL2Q3BzDaiHYVgNCc/DPZ2U2BZ1bdwm/MaX5hjLMKXEJBLD1pYYN4Rf6D12MbGQhXOJHOCRToQ
aMPxtGFICcCPLqqyeK9/IXN+QJZXGNwgW5vASuRBwK9AvEArf5mg1HErmDu2jpVvrO1Jtdq+nn4r
UOhWR2J3qbc24ujodBFO3WKSrx93SxJmuuW2V3mEPGQKpzCIvo9ZDSoK58ldNNEqM0PmUL2B+6u9
20DOW0TI7neVeyOU3NvQ0MEpulqPLKGR/5BovKRftJR2ClejvwswMF0Ac9Rl2r0LWZvBPz4jZigG
QMn/RAmy+A+URJPmsm5su4pvKPRxHDyk2p+rBOpoufk+kz1TXALfCVokJx/agvhkng+E8NgTwiEu
7SaiR9z+mmN49hnteVB7D+RrxzCLjT71eCl8htl6zUAwNYLlhIHbj77SoYgcM2QJrzUGoTT8+T91
+S7pE084abL+SekIeQeud6UR2x8OFNRDmG2t4yqOMVn0s2rrzomDE3eDBp4tdxW1cUuBm7Rkarzx
PkqOL5yIhOOKUkLfwrSyESDlga+axpzbCKS7j+QeD++gLwcDEJ+e0AZj9d9HNwtO4omZgMg9AOee
jYvj3ZEif83C6vP6H+cw4p0Jr5SXllwSyvC+AuovUi2aloW7x0+MFxzV+0od1vAJB5bP0FwCjfZZ
LH3SHMYlopZaY3hdFHrgJpWTHMFnD74/miw9dvCdIJu5LRzhnHhZ/eiJXtLloAGqJLs8Z/VIHfP7
Dv6jfgBgVmG4c/9mOX4IlrTBhmucBkBm6oRTx9m7WYn68KMW30s7tJCbt9FTXTXXGVi7QzoM6SsC
5YPV4kyx3tX/dcrxn1tl2mGs+vEHHfH6oUXNG34pPkkB+RJ5razkywuqQIprzyIn+XuYhnsfHceM
gQZjSTUFWPy62ksTQipQY3tH9T2JNPkwvVzhsPZdfHvQc3obmJSxa5HRjej9HDsIlY9k+oTtFLS6
diw044C+qPBK17+uRBpBTDXU2ld+gw2/pGhNHLSPHCC8+oRfzZBaW0QxH1KKNxqUddYS3i8zCVuX
FQ75YWoetJArteYIM0aPFLc2VhxRpaCzoyGF8dvd3bjawd22BDridZ5vKEz68xKOLcPZQCVLPDWU
2+mVs3eg6ryGmkUqCXcsBzs9OT11aME04q2dEY8OtQq4Peo7N56Go3vYNpl9zhp1m4S+ZsLzP1SH
ibhX2r6OHObDTxXLqC69RW6odEGHDWWa9Ev6WWnfv2OJxKhJWDDJQDtUHV7VnOx3pzj3JgRpGgAf
+wx5iW3OMT0Q4SiJ7Y2uxHFWErvGejeUCJcS0+w8/pEG+69UiRcgD56QUVwZ0mhw7tWe9/UXXyq1
KHQzKQUFiSI8RKH8j72T6iVCOcWo99YxLkTcSatJAz8+fVw3nvrvhMib1x8pF8QnDwA85DxiFrfa
RC1x/L3OXzurHL1Qh/Dx5I6LWoVYOpYELaAChbWZl5oPRHh//cfGnrQiOBorOcDaH6EgCek1xACz
BxC24OaqeyzWOSEG2nX/oLQ4GUwHcv8Ve5t/vmbq27tTMpdzRTtUUAY9TwcWARZFZQMhyUQOCiYO
oB0+kw5t4VCif2lfhX6RCcdSiSx/7+q+2vN3xbC0Irb97BDcd5oZydgfZd7cRBEAvzhqvHuNlUz8
/NMThkpvfEoP58U1SU/gfXfvpMBtqtU3R0+l9ihxHBei8aYoDlu0rvKQVyB9VVfuWrecDQilLn7e
TVB1719Gudx3H2hugL5uIJJFWHyfISIZJFuaN8CoRPlb9TIYt9qUtuXLu7tYJzRyIGmCkoJOgD2o
bwDJi1UF+E/bI3qz6kzAksAQ1inixKqOqKWIImQzqfs89ySshMUZodjAMvXidUpr3J1oeSLSk/QT
LVVlUvQzgMHc6q1Uoa6TxBSYS8A02JGxSsDzR62KjcWrzEPGhhfM59G+eqYWkmOvI0yHjNLGXGgO
pZ2Wkhivz3KSgZo6+jhO75ekojPtasAMKj1v862SNpdnd3zfCmX9JmJTVvsBWJ9B9sjF4tqAxu+k
qFRozuGmU/1+/Zcgwo62HfFAxjJDtpaKvq8qhx02RYd3XSSPa1xCEbt8pfR95BJDKUliwrwaTH+g
5hL8zblhRZB9szfUMl1FUviavY8Lg9Y9JJwTruxP+GBgzoAooIShdjb9wE60MOEQ7AEqKnzTs9lk
588XqJgcB3Lf1yNM9dU/unY/vKkHAvmpfaDA4BSTAONVBYAWdnce3RNXGQmkpbPV04A6h2SK6GF0
lDBXtXO+bPc5uz+9cwm9bGM+JjYzPIFHCzQ5hdfv9SNVtXfnrCehc/FF7jI8OvxFVrmxBH9eWv2M
8m+1jY4DS63bBKH2hizGcLC7Rvnejf8bLTU23S2NoGTeSXfJNPRhOEkxz69u/QDuliyP4agb8pQu
lejsY69H8ktQGtj1jPrAKXKfjzT8XxuPAhVqDVL0AoZWDaxcPxi1vE7ivuSfhDh/eU2yefNod1hA
VmV41gKsYKvXqhDgkdXGK2qgujQ7/F8JnDCPSQqfZ4xq3FMaQ4XSB5nrgn2C2gnW1NNmeopJUvJp
a5mKtUuntS5v8piMny0jc316YzqXucLYwr88uYmaNNcZal06do9QMSgYEfq1YyQrJrmPjYlBw5PF
oFCGbNkTTtMF2olWD9zGwSb3TrhCowC7ipULLZko4i8dSwqGc1L63VdDm5pAL0SL/hi3/TP2Qz4J
oPqLbrkeNlHkJ+4MY6cArdzwWY1RY+WSvzb//RGi8LxXUJTeiMjOd0zWoQrWy2chLRxZ93fk9Y4u
l1kyKQIgSm9A6hEzbLdLfcR5vp+vRfQOUG/9boptp5raqE0PgrfuLw5H3D+nGWVHEjQoWZITHChE
vucmnqktSake5E5KmxfcwRH409JsxyPWimXuPFygfQEZA2mKIIZe8AgDMRtmdvuVcgqt0bD2i1sD
sWeUh8gzHcJKkDV2T94cNXX5FpwVBvSVkvgOONpJMN+AhLztVceyt1LZq9cvQKH74oA9dBqjUqb0
P4/NvqVobplwmc1rvXrvOjWWOpQHHGq2NE8wZJ91Z4mmy2KONrQuuhg0FAwx0PQYowkizD2Z+85C
CAZVcg6SATfJ+/pgcymnEN8afDMes85EX11Y8bQf4L7E7dtweUH+tSkCPIcO22p22kHpGtxD+MMd
Edq9j1TeV+1UPH0UMdCzUn9VT7YD2gfuCF1DKGAj6xOlMFossHSdGUx+Inx697aZChEujJXE3lC9
dyQwsNxdrhz90ai78OAumL1BuFuG954xon9MwKx3xRNkJOZLIKCMmd4Jk56I35Lgjn52TR/PdUtL
1R498XfYXOSx0o7wj74lXvOixh7a9mBRvSE4UTYS/XwGtfL35Vk5o1gxLywprw057fqKZDoPqM3Z
1vc9W3w9dnylpnfJBD8ZQ3n2uCLIHo6GK7yGYVpRSdBia8jibLgq6MLbd+nSqcXIgTh6Ly+HUP02
Gf/dzw2HPmXLoauznE2n38fjZTiYMj7jDziPvLNBHvw2lCquhSRIRnYF1Yvfoq+iS6AKDyPwaryH
Hv84NTkMLEFM40hz3+Imup2Zx45bhRzgTFlNuo1VGB6RcZJL6DrIDedFoLaRhuSXDKB3WzxaBszZ
fum24yMYTasl+NkyYu9uJPrCecZvMD3YScEl3OQeDCVL+bsatRazSE/zqzZaZsr22ygRZD4Eay0v
lMTO4QAMM4VUI8MTS+JATTrLMR2PPWj/+0FqByJZvFz+nFfWnvo9EvY13l5M+ExHjF9SLeDt7Oxi
0h+4rKQmLkZpkDhA3PMhOeYVMFqZpzzeJbPdAmyjwkly6M2OlG4tfj5kL6+UyfgQ11rlh5pAih/h
Xm1G6a8fWiRxT+SnVtVbujuV5jiKv4BbAYIpNTRqfVwJwfxlwtGmy6auyEWxAnDpSyw/Zpcs7mPg
t3aL+EhQiUGcLCG9pHONYf4DtjNe7ZofcrDdNZWtgquwBnD+FxWYbJhHvBqghlo8X4Jb85FHReYY
lYUrb5E5PKocBad5vFTC+VwafnHmDHR0nJP9OIweUVUASoQWTuagv9cMnXdwPlE2eYBouvH3QgQu
pXeIC8kH+Od6JiXTekc+dQJXvBsWn8n7/4Av3vyM1WPL0ARMb69VfHSKVzQkePWuW4BitkZ/3gyl
5dT6Q+HN6XmmBGA3nruwIrfhXoWgdzoBf4gEx9P/kmR2AnKiFqPg5T8e6Qv2K3w8n6NBCcbdJy8d
AUWA//5DEBAuedEpfEq2HMScyzHtr4kmtSNUlRP/j0SYku2y+Ty4Gib/0fWVP/K8lNokcpqvUuzx
330xcTicCD58b3QK3DDWk/FUBK5Ok/chC0h1cXyzb3KiGXXvacGsY7k9idu6d9OdxyfREbzMmJRf
ZzXIAUJX8MPf5ifrO18uT8RjeYARUEjA05lO8fYrnQhsE13XtDohrYaCumlvycqbEetL/z7OIKlo
RXiFdfHDlZcgsvVddVnLGrJ6s6al5oc3WHEPcLB7KhJ2vCy5gflqetBZ2sz8qgGPjYJc7KE/8Foa
DfK5WsztsqBBmlNyo87KGapPBRbjONMNJE4a+JkuW/yqeGRoy3mdUsqxllVGM8fkzWKM5waY7EfA
TIy+U6tjDK1bA68vTDTYqI61M3I1kIhoo2Kto3B0ApEIQScvu8dHXxO+W5CqJBD5DXyj0Q5DReEo
P26Wb6wSIR/VcZgDPufoKhag3zXMZjBR1JSDYCGK7KJWgewalwyjskCT9qlr3haj1ZzU+bdJFCPE
NfVxOUgC31aNGke2crRLcZQNRICyzL4MH8xr5gnROJqVuqUSUCAU3cXt+EBjdl6B/kCFdh4bI5Y0
6azXSML2vQWH3KxohTMOejnFJBcqyi+U0JMAwTQAiteC6zLf6hWcd6kOIH37jcexcpT1Z9nnIxAR
9e2xorWCiiKxXCvhI2Pi2hHFspLhU0BTQT6v79EB5J6ZsECjIIpoTWFhi260bhpaHUIx9C1IDV1L
GtEZh/Ue6YRVI41u4KCHOFii5wUztf6kPzOxCYT4+OPXg6uhivsmd/yrO2/lp++db/6Q0/Il+FRn
LYssqqFzmIHmOewzcaspDbrIFvIhB1r2hLANBNMoGLrih2mhg830/qF3bhK25PgYRj2u4kxM+we9
d6s00u+SS3bV/TOErlfKmjbXp0ZhwZW6wIX7LnO4G8W2DdjDMdaomlGkG2HkexpAyJiYdO3ApCTf
ACyy4x0F4xT636Ojo4CMV/v2gJ31msB9LwqDaBGU5YDG/Y6OJg0qf38OHQR6hqTzoAIDjLW2mA+Q
4tK5ZH1dyPZKdSVAWvu6hFPbmQLMK5pP8MbLoYlOahkaDKh2k8DwGYlpeROcMTTPNvQlvbW4P3kx
6YWeiE2WaQVZVFMnzbi0mjGx83V+AzQ7wNcJowynGYGG+FOriYoX6JaKRHw46QPpOs98dwxFqdrq
GO41cM9G7juxSViGTEWkuyxWLWCmrX7x6CxNY+BP6qt87szKhBDGiuAHaIeajRh/gzOasoQI4ZTv
nrzyIA5NQHUMizyQkZVO0Wp3iKB27DaFuOZ/oSgEi+x5W/C7OZT1pPR9R9RnI2Ah2WU9wdrIQgZ4
ukDAWbgKGuBChcvTGibFZbHRMCFmINsdtcRcyzNae6KCuQdxgARbhOx1foZUQo+UXlgv0MxCVWlh
BqJjchZbAuJkf5NEm0G6XS42vCHtIodtuaxApNTwc9c0/kQL65DmFdwklG26gKE1jMNxYI94jG1q
+oPjVB5wZ0I7ouYA5N+LrHmY8bcIQ5dZ/nCHdn8lYDbWxA6YLJxXkdKO4AAStGdLgNeVeyD5Ie8d
eLtzSN6LH5MmEx1Fl6Ybz0DKlR9LwL/oOH0I2/YHexufLSAPE9bHgwySz4H9wq9lfNTol36Pbz8e
ZgYLGUdOum/NodyorjoRFs68vmLv8sMdeMtTPkDPKTAX0sTVtsHjMfrtVMzojD1kFIheuYL2fz8Y
i93ONDnP5qdRTFucChn3AhbPRoViySr/LYRMc/qsnxtuzvet9J0JElsPQRyFd50nljdQ9A+7cdYc
IwG33Qy8waUOiKTrjSoTEME+cGo3+bRyxOx37xoTZeuCyUWxXGoBgjxf4eNF57K2S/ZVTAeqHqSC
GK44Xp9SwHnLq2LUi/FGKjvo1hrshOjCILNxLNmQRckaYx8HVQjDIW+6SNjiIuu0g1IC5bZ9pPua
mwlS3voiQSJlEo/klH+9eRMaPfWOj8PTSI8Seu2/7GFGo6yhpybSTXjg5QlydJGtCum5Y2IUrjmZ
2cyGWNQnx4HMSSsLrjpcPkf9rxsMdF5TillOQhmRU/YEugjfk6G8rqX9hSQHa/q7/jMJasxd7z3y
icbVCCa0O1MJLdM3kUJgonzjSbbA9YIyclrHBvBvSnfYbAE6o8ocbPONVCIloQvq83/xnTfVarKi
qaVoOrdS30nsIwWq9xjg/DxohKEoHFIIilU2sVeifjN54RRbmFZqHuLecfwBLpQatDruqws4IOBU
P1OmifQK082NKXoSsvl31ffbRu2GebLcjF7l0ZFe1qFcOXY+0nNDmJa7Q/2/KaPqgJ3+VuUvIfUh
woY1cOh85eWPuDKdNZIRObpZ9b51GDYLsQSAYjJ4nfxpf/JxB28km/lR8CnYYvbfCglu3brax5mY
mfpMhNb3crtWuc/WKrK2SCy47BIekjBTap07AKCHO0e0GeTVdfQQjpYgRcvHS9wtOyqMisUXvNR8
AsnLB2Ri1a99GUj4MzdiUwZSCqA/it3Pa2Z2tUnQsioKoH361nEwgXCMooEJTJQPY5IaHB9aXDQf
PXp/YEx8HmuUigI4zBInIdGNLUJKJS3gOtOKaO9CYJlMP/yqeCNstG97/VG44L5jSICd2sQqNf+Y
1QLgGWCDQhDcR+ILhNyXCIOhyl9sWWg4uCUbjULXhgcagPBzGHI9SDRLPkTxEqxDzKUlZ4AaB0cp
sU90rG+M7pRkX6TcRiGvu/uECYZqTmphL8sGXjJNWNSLWab49TmJ6OmaMseUKpppzhVyKZvpSBLv
gC38VWyHD9+6UyEyoaDJiL3Cu8ZM4y1fKw3XNCff9yo1Bc5CGlMaMsHkg16vUjt0SaNgVIVjxx66
sjqv0PpsoieEUb5NRf64fftwMFpni6JvHFOilL3tFCDjq+PqyrxkCsO2uxc9KEUUivvfy8fQh9vi
x3/2b+cdAdNQH7LQw0KyhsJSzaHd23BzWqjFMF+mGl3gTioQBLbPIMQoypNzjRoF/HYUFD6pwx/U
EXKxVhUWvCtYCQ416s1eEF7FaInFQXlBuoq9B4Qn3Cz+FS7Vs5p5Sht67jRH4/da5cdJDW9vO1lP
DzLOPc8JQuYd/4KXTpIhMxVqXSgf1PO6oS3Av3ucxYWO9Dd5IQSV/o40TxuugeSH/q0ZkmRHB4/x
E/hdvs8104yDs4HaAHdRLb0h0WQUlQNssFiUYPBbM8rs+PN3HgI2iXikrTwf80UjjZiaQnd2BDZS
NJOGagIbnUsJrxCvlc+WmLuSSkL+HkzAtBvogn3L12e1AZpSYchqO0bzNEWwF6l9rhD1je22H1/l
9ApzBCnn2XVSSKNDXibuSzQv393wKPG2azz8/z8ak6ucSLEIqll2UE2G2MAnzwJA9SMOXRnOxw1Y
FMK7/vtrKj5ORSRk63DuGbKKCjKE2McyuqQm4XUey3T33xX7Z44PT6enRAWionloeVzUBJrWdXtH
HbInI29MsODNN2fIrzXyi73A0vMsA+Sj+LHSDdMT5jTNNhWOB5XaX3Mj8AYfIsPpjceRel7fLQY9
KA1XvJi83Mn9AAzm/CP4wJ0wyED542sASY8Yw7ucOy9kJ12ZulwIcP/5T+WDBK0s8eLhUuU+6lNr
nRoAnxocfmc1HneNUNPZl6P66mbOUHlxoNMldHgs31QMt9MZmWGwUzleD47vgQVW7maS5uZ0VAP9
nS2XNfIxGZ5oOlw6NcJta/N18iLmqRk29e8/lFNJtYysd9MNAlPDdLpHd14YhWSBTvA3GcVE54zi
3n6PCjahfwKIRWbtmEoZg8Rd19iO0nsSaIo1oHW6zr+eUwKNgKiSQkr/qen8wAN9bT6NtxDtJnwV
+xezM6xEebe+VZ6oL3M6kIjqgORMwTLueqAtwRJbkhideWfyWK2F9+DwLOF16PeWmFN/WBCwNuCV
AfayHFeNQAqIc25ymCpmeC3BKmUOupnJGd/C8Utf4iV3RatI2fBH2WEXqcO0xdI8H9ReCZ6eyBbL
nmHi43y2qPK/YMLyB5NMQ7o9d9M/M31EjoW3pXzinPkDXkG0NRcInlJcv7zv1g78V1NZ86BZngd/
JXDWntYa4mDwhHNWO0WCD9uEMqaAhXvRI2IcMGNPM/fPIlwGIMKWrqiqrE9gXYB1VuOZYfh7e5Kl
L+7Mn8EwsB2X6EQL3LNWT/Vgq2kCh0d6W/GIUVsXrrG0+X4oLohpILUuvLyOm9TImTOkn3XEuzQ7
ePd8kYHo7QaB4i+e6XaDe6wVQRBytm8XqodSLQTHb6wBns1K/WoHYscJ7CEdJqixUWaI6kxp7rKE
4OQwe5GvFn11NdB5zSUCDK+0h+oQnbuyYX89rA+zYO9cR0+7PbMwVMhnIhdOpKUAc3UYF2bKffUl
V+CNV2MMdX8ludYVYCA7Yk/qDD3l7MJZDs1CsUqL7SvsHGVHRHj+zJsS88zC5Dckv3ilEfbAo23u
1woQAKdy4nq+4g6vcGQ8sD7TW6sf/eCwH837WbswtHLx+NnapuaPSMSdo0WQ2T2bggCUQ9eXh1/i
UvqjUEdKcQizaxy9m3YGRJ+haL5YvVeHUmf3gZ3p659bygx4+hf+SqDjYgfDH37oNAOSdQbH1OaE
399LwtF2uYwzQf8BUYivZQN/bm8nRVdZTQ5CnnPnFGny4SzXnXZM09nlFcgQcFJtHuLKw96sRIVg
/ODCH5HVYv9g2JxZT79Qiqf3nhdo9GiJsBpFdZlSaMsd1X9x/Hu7EhnnX/jv7J2YbnGI3Ln19jqa
+LU3qgWmlYnlschpz7okzz86TrZJh7I4kiLLz5vCJJbv5lAe7/IOFYcM8/9LKjZGteMluBBhPJ3h
kk+c0e4cTHhlJiB1nIkTaOapwu06/mMvS7nlwY6zTf8wP3WcijqZVEeelVgXpHpyT0zPbko6CP/k
otY1Yen1oS8XK1o5AVrtOpe8Fb4HOVEtThCWf1fKERKbbxOfnrPu7+/hSydLWIx2ls1LxNA0Lip2
h6+Fd6EzUm8HAVuU/AyImWKnNa6Jo8drJk+22ztzz2bKHJge1cAwGnr6KWOoCpk14m/ijUYbuAvU
M7nqd05bV751Wr1dh54d4ZaVkfHhz3+czqswEExlc6wl3CGTO/jpsGfnWk+7ImsSscCqONFB8DHv
n1uxjRf1+a6Xwtqo0q6QJNE4STCIHiDMUULZQUHhBB+EOLDGU9CvVcQw3OBE+iWuAaCbIaJxnYXx
ZqVkMfEReXG6RggADO4e4TrN4ROK1bF+sJzXQFpYQcSntW9mPGquqOdQPN5ukfSBgU2Uv/xUoec1
kArHxUgHZDNQksOsThnPapoUGqYtZXOnIOoi5myJK5YLcV+AKoO1dIGy90s1YhrijwZ8rccllmpu
A/Lc2e5Jw1eUVTvaEXJOlCnVZE85yb6S9bwZCRN1698xWqw8idEqUNc4RJSywd/1REO0+VqHfQS8
BBp52XiRniE+L9EbLl8WHEOmXKF3NJcKUEe75Xkmcr3YdgpeMTTl6eB3T/FDiGYzFQg5H56fQ2IQ
3z4USmRZU8YIkQcbfwlFsjwcQkYGSPklVylzZ372NzF3fyPqQbmo0jgZghgzoJiwx/jARpcTNifN
Jt6XZpYtqVcagS/fzjGLz6D5yq/CWiwgoRlSsxU6i/vkEMy6HFkdKNI8BJJNbQwNrvSbiDfsZ4co
u8RgLh4rS+MpMZ/u7k3SwIuoYfYIkwEX4AmbUJpW8TWiDzM9BYnip6uEGGkPuh0nWiWB7ktITf0S
IpAhz0hheYzvOrduXxR3l0oZ+82EwZLJaoq7Zvmgfp6+h5q7S9K3OYwfkZNavEDnhRidiZD+uRcQ
SRrCjOFvtA/8ozCt0dcnbXq2Ae7wm3XBk0kK6bieVOK0pAub2/YsfL1C4lmysBMxuQB5zhG17Vln
MrScjxUhnByfVVHvo2EMYvmDpU1du9VpQqIWkb0joRlkfa5ZC/eLrrTDIzT8mSDmNM3UcFksmlBv
M/54vt0r+5ed+HmQ55ovnxLqui5gj29Broh9SGIFqbd+T2TU0FSum6ffqcm1HIYNv1SwZNqLPUbq
uN2aESl88+EjltRjWA8zupJtyJzJAlz8wuXi9PfBGSi2E1lxd+3HzA1DcazP8DEzUnwEAYCOf+Jo
Cd+ddVNZzwVs3E5AAJYvEPvGZzs5zY7dfUHJY4u/l5L712dKs9mlvXDDEidUG/12EQmsFGQMQbU0
ru8Aw8Wa0pvaM+hEsMesWHnIE9/5Rcug6AEJN4XBOPdK7S17lzlV3bQwbnUp0iRJlzoEejhiccCy
8WILnu8VocwIUOBiPx63p/5drT5NSOuvUUuoH8Xq3AjcpWZ3rwCb4eFbMzDPe88Sn7JnrIUE2Wdo
ar52+PILnOR5RKsbM5oZ+SesCY+tpmn/jsKw1mggzXshp/owiMQr3qekIF830yEzA2gzS5xpx5lz
dl8h3+b6dvyRPkgiqcHRF4d92OPIb9N9Fzcvrkm5+XNEvW0L77j9iomX+26QLtSc+0W/E0hI5Kn5
sQEflv9o+FS9I9/lrGpAdsstI/EMPMAYNsBgfzuRAfzARgKOQ5A91YoIbNkINolEqDbnPiIXucwR
ds059LLQt4hCy+OyP04Tyb/DxlwcG/Xvvs2jdKhc58VH4a5RqQF1o227lOpG8gS9MnrG9AKfJAV9
yqeTq2OEh6cs8M9QEM28TqN9eWv+M0tb/VDR5iWQh5qMAhM6LBpIvCX53hjiFlLiQo5YMIvi7BQ9
N7sXo1QYpHl8CYqD9frfr/cQ8p+La75D9jNcCgaYLgU5f9SijTtXqbCLA09dO5voT8FInfFya6h5
rq2bC+l4c87FiLtThi1mz0xFHYqmcvxteGE2yNaQk7+mmxeNctAbYfTcD++cIFhLykFPU7jcGo1Q
frmQPdcl4hSOMIZ52wGUaKjZHNESL/Te5NDmaWpeZtJ2pW9pqwVm5Va88+IP7xOTop+8nJpt+jhm
82c5bg8mC+lyf+rewnKkFSeqRAElVl65HsASSy9MhBpiaABbmHE1Ri4BNpF095ecr+8OIEhkkEOs
vc01yY6F1DkBqPeFoqp3jE1wxgphun5zMUhEvxJpOLR5DC1kGPbwuJwxvq//u9CcNQL0E44osZhW
LMYlKBiLeeZClJQmHgmYbSV0ujyxGnl+wC0YAAFdeYg0wdvS4b7BijcN53LGlyRlKuzrOg6X6GQ5
TgM2CmrtTAnRiucvJVxv0nEx7Cy2YELjzvawxMDfL2LwQNeirVd27UrDL5LOUX7j2P1SwIIFzqx7
j8gpJaRnbsnVinQe3CBIeMarFD7UC2tE6WNNQt8LdZMPWMCtwAdi0SRmyMXAO+tYjfZxz+80kUhg
XzXq9KUaYJdpg+yYklZ+0jmzWyhW0NuLBoeG3fEjlxfsMzuM0GMPQf6g7JOOxRzt4NrXH8iAJDjm
QaOk+dKVDPpiy0XsT+QYzL/NIxeGxICelcblCXEgGZ6SOd3F2oeUsUn7UbVqiwd2L4OcEdKuse59
0rSdyRllOzaZclCmgBTenFnr1nFQtKNNj8g60W29Dr7+2qNVNmTefxUprIg4AJxG4C+tCLoWs3dK
E31pVZHCYas1PR/DFa7vU7aAB+AayJoKQDht9pSgczzZoniXWID9f0IP1Yg0B0q+HnHQa7YfoF3Q
W+8AyUkNWzpQGJN6rjIBbTp8MyJZcepyTBXI5UCzB15hmfQGl1cmJ31BdkDV3t9KblPBK04RySx6
gLeBTyrVDbC9ua++RZfevEvs6pT44zwafG3qHC1nBlM/6Mn+tu6+vGHets7GRBH3F49/QQ0XGDgP
dB2sT3uDsx8g1RB3/+noJdYC+2kAM7CCJ8ZVrx12WydZK7rVMAZ8GAiS4BOzAcJamzeIiL8at5bY
AvGI/x6c0M/+Msx2oZXDHtZL/Z4aHCtqa3zXv7eB203mbihzAswldyajKeMVz7eFYwWSVPEa8NCc
RlPiiypmjUD9cHhNrss7hdhPDrVdM8U3TaW9d9lsabVX8Txc0BxyBqbnYq4UqDiPVr3nBqauu0Cs
ahoHaVPhXzt9/yjiXiREc2b+VLjVqsAYVbEhpN6SBvPbZhFr9PmkMq66Ve/vOTRlm0v7xPWPNESs
wJojyykyZT+PYeKyhxx24Y8c2wTy9N3FLAj/8A+L0oY8b92KUamt7ZZfnJwIWtWYOMSNZaswWPzD
kUsMocK/+v02fzCSYQKMo1aLEb1v0EO9iM8y4nDXQXxQczLKvDnBHswa0F38klUOukSYzm2C5Khd
FxMe9ohgbDOCFYF3JZANYwj5og0TQakQOPwOHJtpH4/N18fEe8dDzUa/VNgLjBty7xZls5Nuq1in
i8jQPSg8EVYB0q4ok7PWeXowntOG4zHP9gmoC6L8HweIN65AWPMZde3wvr+eaOp8BtQ6X2Fbj0S0
zd0WoR2RAN1zKX0uM28787MWoi7e4LIMJHSH1JpipbcDOEPypGDCOGtzrcLFbT3nHamafIhSAWFr
pmSYHG4eSpuZyRtX7gFJl9UvLjKpQBGC9/7btjt3JqQLslWLk/IiGjyFpD+Zun8MdfqA5mjoxZSv
k6KSZrwXsq9RMkxg6BMd+LVER0r1uKcB5g76TeEuTmWTrkWGxyAnJgVZ5e2xxPBI9xVcF/0rttWm
qEx4uZeO6ZxFTgQc82rE4/ftDJNXUVVrPDDH/3IFjaze5WER5c57K+rjOi698O6IdQtKY0dPin89
uTyITywg8QqHemhOeylSXvA/7ZYjPsc5q1XVrESsSFaQ8ro0AXk9fntN4RJkUzGP5zsos6Fq8XGS
v5aZVgT9jNwVNBua2TsCggNWnaf/6/hrZPNynZBnEpzpePDy8Z36CI+rJCcx09BpyffNfqx2iFs3
gyWpSNc0jSTm6AiotazJujY5WRz86cqI7WGqLeCPRq3ijNIdqlFchQBuLSFEyi+YbiUjLIsCDuj5
fVPzsvA7iSNQkrEUukkGSVcFc8ldV6mIg6IQOtsFoC6FG+eKXzRR4J9qerYmUJqp/PNS7GYZn0Qg
TkC6eW4aL0iDdSmyLD94p9+hIypymG7vYRAH53j0FmfLb2/nMjg6pGvwBZ2jImhGQu6MK8t8zarI
IQoZwNrdIiQaGaHrazGvzJ6cI3yqgUjQPqvYfc4r6xm7Zt45fC9Hp5OJBcVrnNL+OtQjEGXs/vmC
JoS9lJkt+SRcH0t2XwaQstpP9IxN93rnOJdMmR4kLcgHQBhXY27M+d3gz+Ib7k2fq9G9QeE93ouA
X5beQMxpBZn7WLfhGTWbSjhvlon3FSwfRV2xMsbOSEszIKS65571rImWbV1qvj8VtWZdV/Nd2ZDf
NvdSOHbH9aLy/2yJNlnWQioC5nNujVuqzCAx2LPU1PLNdPrmTyd/iZQNdCo4zZOujI8DOE4YoXF6
fcbR5uq7ANU4eVbHNHtmuZFUOpYQbNQTtEMqWa9YrhYq3HCEvq9MUmdRsM8CRjCZBnsQ93EEvSYa
F8IqX4vwr60k7a2de5W8Y5/CZKbN8CZv8xqCPRFUVs8wswzMJusxEMLSSIz4+UkrQpGJKwjVQZqs
+zInag5+n/hzDd6T05pEDbKnuYtuZE4SGwm6JVFHVZHk3YZVkxpsKXbTShIcFianN96pEofL1DLZ
Jfn+hwdYUq36QvEQ/IU05e16gzHROBvyFUADSB7mRwLGGIA4X3WNhz3ziE2uLrLg8WbjRclS7ic7
1vMwZIBQdJRgRC7/YIlskfPHADh+tcgb4IxHs6nvaW4373pD/qN2TbNLFY2lESEfdmbrCWq0qRRS
LDN+qGkOjbJvd49g+FQ06KPc/X1eMc8yP3EnWWR6Mu7/BKilSe5Ih9xOwi35yPOVN+mwt8Mc6sEw
R5wSLvQX27LPHa0uJsjbJCwH1LML12SzZH2lN/Ma1B32wWJQSmbF9+6TIN8jY+FvYEj+uxj1VDjK
ViyHKk8cupGQuZl5lLPOtd6Du3bNJXZIZr0rMrUyCG0gywL7ZMv77K/F5uT/rLalBX+zbtC2nxMe
WUosfsUVQ5AqwO/Q6Nb9guqwp0wWywOUdp0OvdsCjpuVm3P6xU9kPSJh32xz3bTDULnZpDtpbiHf
UfOm7EmeoEqtZDnzgbOJR7dzqyhIx6q7fSM1OxeyOp4YGhPzFUx02lBEjz4R0sIVnohGIqr+2ObZ
CzZa2WubgNxXBzAeTljVFUt0rT33TEFYE0ot3LWLeZapwU7ZHBpIhMAfp8tohpNzI4IYoQbpF2zx
L8HikK96MpgV6bdaNF3V/iaqQbx0F2MAy+sDPPWjykAc2Wkix5EWRbim+VfIBVNLJJpjAtU3uQvA
0v9OTFKh/po5Kxp12FsoEB6iFDBtIEtX25q3LFSV3+Gm4Ao6uxKjKm83CieDkwn2JYap0BoGdEVS
mwcDHxL4A8ffmE/+4wR2wyaha7tIYNjwMPeTtiJ7ZEtgwyKNTl9xtQ2uxbVVMelqCuZEGAc2qNAO
LDFxCaXbyxn4mtBMyUsqOrC0H6YdWqYkqME91a8Vz2LdM4OHbGqrcJTdcLyBJWL9HhJlQyFWp5gS
KhvDmSzqKtFYaf9jPUG9/y+vjRYzB2Wmt88m+iMZmTmNFv6vwjVq3CS3CLIa7u5b3JbQHJhZO69A
mk8mUCJttoYV43y2yd7S2JAu+q2nov3FCce3CRyr3JWngbtFlVnfZFF1HWGBak1ruLAw+DO8iu2Y
b+2rrWLqyYDBBySwvcfWr3RTj1xxeHxt2b3PQ6bBuJxS5sKEMxTFgTWqDV0fF/F/bLdr3r5nrdYU
4ESeDU2mGLZSeT3M0z8ZkqoxIgxEto0G2YFdKfKi/h66zYZX7Iwky1hiBBUk8mtbnCxE/Vsp2DEO
swGaCPz8anzVHeePrdBcc2eZjTu7DsYxZKoBIJjZAY1bIQ6GE4Njw+doCR/klumCC2BkAWDeymCB
akMDkXwboSa+bHvSMcPrv3kVkMYPjMRcdZwIKBXu972UatQA3iW75UALrewgp+C9DgyYrQcPW0Fr
ishj3PTzDjcwYP7hgoTwT6f2GhMAf1okvjFGrUwcEvLCRlaUshEc5o6CHE2KV//bvZwzWGO+8nlx
3wIDX7lR6q9HnAe7AXrXo4qQeO/RXzhtNsS2y2keVFKmVKRyGzpVATyZRszoqjtmdGspdVNG2B9R
jWChhd/V2KNlsMKBk941PR9sAsf+R3/k+wBWMSkKA2sl2RlaETUkGj3KGT8NdKr2rSpjA7hUcukG
A2cjL855fbMbreaLOgt45XZ0QGKdY5Xio7J2QB9J6tIXHcIsKtEsbarN9iiy+dibRGT/hqXXG1bp
cx9w9Y6qH9L3w8iGSxbxlRanErEvT9e2JbBARYmR6GzdJ4fvFel+Opo4dutTYb/gxQQn+K5Nuyft
Ifi01cREl4j9NvfOn2ne3p8uX+UtwAN9FgcjfXs9WbBw14jjYC7ZsSGJ32BHP/KA3+tV+JEG/WqE
ukK6qE01u5wkd2cBEvEwYYrdAmplYpbr6YyU8iugrvYUMBrYsD7heAFbEL35Wad/bbz5+ywM7zf1
8Pg28zhvOjGJTM4cQDGDdKfcg+lejtqbo+D1KhjY01FFOMAVgjV0dBD3v2OwMdCi9N0RSseY+4sN
cigS+JikcNoApziKbE3XggwAUvCLP6H+gxRD2ayojaoA2NSEE+VrkV+xqk/+jwj+L3sx+Y/vTGgn
afcMY/L5KdItTDfu+ZuzG11xZzWJgwI6cO0sHdc2+lQYXnRkVaXd6QTyo+DYVtgUcnNoFLia66DH
UGokUEzt3xDnUoKITzUFQvugUshQ4qNUg7N9EFYzjnXsnkg37TYK4MRFzyS9B6x/r73Vd9Oh3feZ
HYMPRFy7ZTn4GLuR6izpoU6Dnr3Ho5tpQtjBZ/TiL847KDeiXxhy3ANtvWI2HQNyslQVU5K393jB
CHrFpkFZkjG6VKEMceMRoM+34LlaWfqYx0BsjRLhHcE+yQSOCf8NXDxRxUWq24tSJVbyf1bH/+kP
kIa0UOYJvmOlMaOGAW8yeFNYLICandksv5tDLmSqOtdoz5gLH6tIIZb+MHATVufJBXsMRBR7ojgb
HNZMjjeJG2bF14XQJkQumd9tL6urCOqpQUTNvSrU2+8YqqUfjfDUCas4gOhh7usGIE5pVbtswZ/a
pkGsyAW9xRxj750qZ24lQ5D8M9XcrutKHxBnCzkJWjIzzWrTXQ9tmCgIWrbVSo7M33aZzhkxY7M3
dlbjUUAf+EVCfWIHryurZlGDA/D+gfqXr83iXBSce/za8/dy4qYjAB4HmhRB8Kn8Hue9r6Is48jy
YsxjyFSDXnJIeluIWO3+vJ7iMKFFKSu+IzFsyhbjqbXdDetjZ9hfhNbJZEttYNZSxqXngDOH+jrK
qP6GXre6G+d9yTloYtOSr6gfYI7nfXJLzRPRJC8LL8cL5AMi83OnFRYHDvR1mIOjw8VRDdwhLlgn
rJq9WZrKESyqQFpfLIu4t3mmoxHTUR8o6bUnNmCtNuBXAX46oOAKHYgNx6gsKoBMK0prv2Hc9EIH
79s2Ubr9fntoPo7Hs3fJWsi+1QFUo3R9mS5CWTWzXUTaZh8bTNC3zsuSD8iycxhGseTX/6mA90hP
sT9TRri0T2vvQK4TKKLw/WJ9pNn407PBpUvN0cY8oXRyRG/GNNkj1DTZH78qJz8smSkNtTUJ5KL2
pqTL5Vw/eqQ/0arzKxYCWXHjYcADxtub3C7XDPDXjVLzAYwSb5ArD0u841RJ5dXlDnOXUvxqKZhF
wCdc+tlcM6ivUQo9XsBHN7IYs2bcAC8pMF+ScBW5eOZTDTUTWYLpYz0RmKKyhuqjo4yDVyW5omTU
UGd5LpRC5tDR8M7qdNtJaCx6qVDYeWWo5HbuUa7Noz2Uw9Wc4DtpjJkOGyi8GFqI4GCgDB39bBqm
Z2Jvw56mNZiYDp7mlXpgC6iRWXQjwuaT8c4449dHUSc1GhxGneS0eOwAMvxC0LisXChh/kOaR8YR
p2aIIIF8TBTSGN6J7eOxVNj9A2V4P9tRDnupXJ5o9fIz2k4BXOXgG0UyQ/GNVz1+6Zn2KIkRLvp5
Ei7sHWAmqLQ97ZDX0vpSdpqdCcsrtitMUgMbFw9hfOB2KDcPDtsU2F2cHAUZ7izd5axm5OGwnjwS
xTZrhCGopSGERy81bxF7AiTVuko6LnCfcNxcZr1w+24GaQU2CVVGRa/raB0XmPWGBO/D4+jQPCTc
7PauHT/E3tO9BVZ/UMfCio0PuGfO2fwMmXK4YwfKVhM+7LsEV4nFfySUb5Nk+tZ4lqH/T/vlN7qr
b1bpq5sy175tX3A1cNojLbU+vX7qP5z3z0bjOu4DZCeFYILsUkMrgEaqEzyQLde7tKHdJQb5gzwx
O5fSLTTPCY/H9/T9/SS2VgDg/zMgFyd5Ci3YU6YrAJfL1+GwS7145HlBcsCQH2DVmXuuJgP8mZgh
olL00B8G46GUSoE3DC/rfDU4TtBm30EE2rMW6HooOj0WAI72mXqgbWMkpybLf2ygR35xGtszx4jB
DkRvPQmhtakBX/smjMtSVwkSneR0cdqUWk6gsIf4qSyh/jNi1lafWayoOFf0mpqxsi46mjI8TtTo
VkZYKNE/JBUvX9HQ9bt10tbTZslrDl7qLOKfhqZCakxV52oEzNjWO86mYXhdbJ1e11U60pzN3Rf5
vCfN2MeANOrI5a68AludhDIZJofCIxeLoKPQOAu62XSRp1LiRthc2ma5fUDh7AdA0Lt3M/BQEDAS
VOqmcQLFPPpBvykCwmzDFZjL+7Utcxbjcj32YMdIqvG1MacMdKwiZI63lOQDGsyzQItNTXIJqhB1
sVnzivk8fnDiGTxTDciNDAkZfe+tRHKcdhjY774hyNmKwJ2cLShforJpXWEfLwf66zFkZJRAW+ic
QGACdG4fYGL9b6qiX6BWCFX4VmEIKPh2wRpD1b2UGUbwwJqHsKod8Dt0q1IWd4IVHaSvqMsYoLPy
at1+V6XCZqj4ZwYJcP7E8f+JlCbDx4+gxoPE0qXmR4ihKw1JHJjzQS9fxqjxEkrYJFWGTZ35qkEn
aDWlJ9B5RbyMQaHqlPa4tavFAxOtXiTbpuSHr2Oo+qYUxDwHwg16nMQOTcQOsKG7lbaEaKcylHWQ
Rd0K6+sWKLvxbxBM4tBysWWmS7Iyt02Th19bq588XKEb890Zzee/exvDdf+rvvz3o2ZLvxaLpmba
zacs59w+CwwdkkUb1imY4W4NolrQ1tncHiR3gRMYQG28vNsf0/KcR0baqhDSyHncbDine4ay0FXm
5OtJeZh96f3z+iOivwzhK5B9mOoXLOROmJpxSNPlCFVTOF9JjKYEOkjvnTNULS7YOfQuKtzbHqIo
YPDbCY0YE2tl/bbrio/RyOfNA79FKx/WzbrpbVlrOEyDywYM72A94wSIfqhCNirDhl3Ab7DygPsm
l1teysxSiEBHWL/3GV5J1pT4Q82C7J5/f0jHnZH6bSztbJJ5d0iav8Vh9qp2169TNq1mK28LJXWz
5YoBqG4WlvwzPLvghokcseeFTE+MzoX/EgYb+sryZpc0FIAkRVa8D2f1VSVbyu/tZwooQYnMzRz0
kNYZ+isyX+xK/pUwPiCfWDYSlhifJKRsOnC4nEs/ITt2i9bDC8ncsfW68N2mAgRKdp3SSTibjDVU
RJYDTYdH5zXbizBG+HsMA8CYBalnL+gO67qVrKiIRYLnsWt5DtgoRdRSeU2vk0upNxrYd98GAkd4
34jcK68c+Vtc/X3D31CMvpupCuPgLmCHEbnQp3nxLKx6CLUF2224GcrKdexF6t+2Dwo7s3FhYoui
FVQbDKhRHkykuHe+a9EL+6U+DydjMT2OOTQY9rlgGxeE9k1YXJsK9SOXN7+TYxs37o4jasJyErZn
5shIdP4YuBkvhwwfXUfxaxdM861MCRCWIlJNXcRr0SPYzMDukKfUXj0qp7VQBvZsHKwKxvWtqk6S
IdjZku2BBd+I8jxfGQtIFPRJgzLfyUPaUo8ziNnOeKST9xmAn3hj9CCj9l0vBR3v8qUcGc8tEIK9
QjTUsS0NmaQoaJLPSx3B3yYlQoad/3IrdP3+WIZDI8Q09AOkUhmDBs4sylb4Rkz+iBe5vYs7jTgW
flq8LM6jWSxzx6KAi17y12yjhjmK8UponA4ZDUX+MhoyipyWuEFUU3xp87FDoqo8dZ2GIylV35lp
8mh1zaU+/F39wEst55frU9Q73IdFD0ilXSAu3gj+xjN0Ex1fqsTK+BlK7j00j6FkK6n5Gz0WgW4S
d7dp++i1T00VPohXRBgGBOsFx1ZCA3iLUj+CbbPWe+wkDAGiz8nGnpj853Z9kg7gudVnXfZex/fF
XxMRGp6UASNiOgV+A/UEOvFgLJd/jGaC5fEDpeH/5jkVNCbd/TaafhHb5v/SZV0zlfJro+csj4Qz
2YDH87B5mJAKZwsWVqk+8QgoL8CD2M7Evkc+0xIIViG4wbbnZWdwfELT4y134XxQZAE6l39mabuu
F5E3+Aq6A0DOzBNomxpUeGyUj+oybtFmloA/0XAoP3xAaPwuYdhEBUNrWk/yWEBMnoJsejiO17D9
ARvfZ1vyU0Ux+mWg9K4oHKqS0ufYEQ3BlDHtuJn42beUc0ycvbvyb7efl9DNl3dcmfkkhFGvqB8n
vxPFLUV31MfKQlnM3J+h5UsPhzNDyHkekZEQwpYSnOMrCT5mrLQyx3f276UuufVFbxPRkylJg821
LUT+P0ZPWkxoGY12kszdMsGtuDFo+YLHPXqhAFVU5cEdMxnki5ibSSQG2loJX1p0sKvJNH40ezee
0IGfaqxxpZ3CdCsaS2KSa2q4hVO3lpVE2vC1W3GNUi7Ty8cbBDd1sUu2iZSB7jmoPedg9LI39zeX
7j9mnDQdeauv+gFU9hDn0UhGQMUw+uL2EexhOU0cntGIa84YlGh6cE1uw6iYP0ARuDrT6Yn/MuEQ
qOgv5Qvo16+gtQ+k5YLA94ImIR1GgIku49sfZg5N5cKB6VPHtAR1ARwHZRUmZv1ZajX7l7W+xdrt
JbFcpt1B+HgSKKXGpPzbFPco4P1YeNDWHZU39qAj8+ZBD+GxSQnHaQixSPzIzqKC+OO3KjA73+VL
EIRB2UwxmzmVL2dK48NoHXldUmYcZH3XQjvRoDsKLIZ40GXqaaKNYQ0A47jRWFm0p9AMWTuJcnUt
WqNpNbjWvVAuECY+SnknkR9ce6PcXjIHG4u26z+gDQgHsYLuwtMYHz3VywjaLuetTPF5ftdMYVb0
88d8E4f8SUE6bxQw+26rRPv7dYP16w1yfpOWTg/cvld6ZR+QkQNasxQObzF5fB/v/9zaedTiWKf7
/sBbDbVwo4+BzHb/VpGYutdFZLabemmqoxWbfoo+GKsvNHNpVecr2fSOq7uJ1T7zs0mdOgTwmsoY
SVWHJ/GHSNzxiWVSSGQMiBDG/0untsevIPLRDXuS5rZK93rKnOovavSqYrFtJ7ZKGvvPAgcOiGve
Gr/YgC8+7itcW4bRocR/j9o+A1HJVfcD/FIkX2QXdqShMQQqtNY41lCyyRQUaeYWdVtWMGV0Ja7T
g8NyEyOm5jD5pHrWcL+/6HGYiLKhFoeEhEtVKIxeyuakap+5sZLhJuqlhO+wW81pmLrZUjZrU7Py
qTrt10XriFEona99iWwAqEGPuSKqGDcnrUzjhcpDilz6Ywot5M61xIRxU24pOqengCdSgLw6Ycat
PRCNCa3aIJeRekiqgAebW5k7jVOkznpvlkfBx/2fEkr5fBIyYECf/Ycy1JvJcrkE0YspiCru/9cH
nd/P0Qe3bHhCCbHjQ0BogMlroPGCXbQjo3ooizFdkMVOx/dxUpG/70ozBewJixDqsj73fGxmqvlW
H1OiyuFSf8c5IardXXoI0FCvDP1/U5k6E8Zm24R8YmH/tMRCN/ql67stL/xCiqzR+AZ6le6ZzkBr
lP1BnLtps/iN70CkXdY1OBaPRsG+tvQpCvodQulOI7CYFQ6XBLS3nbBo2Vmn9BpXm7m1K4JKfKbT
whs7wLzME3DnpDLrEDlwP3ZddmmaQ1kJ8HYu3U9Y+SRDz12Oe86t2T9B9bPPqWxTtwz5infRWVe/
lAYHShLMWG3TMKUJyt4w0aiysM7hKNQbkHZEUf9iK/uYbalBMEJXPfCkUblRpZak9UzohaH/wNII
WDb5m47DffYSkMF09TUlT9E0QBsGIK2WDHjhvfE9CexoXPvTt85H6EB/BkIdVKR4SwiyqtvLdV2d
Ll+bUqeyPeh+ocJcQ//BMVoqEXezzslCpISzuRbmt6dTCD/aK2SQPfFR2yp4egdJfZ4L5J8uH+nz
ZM+JENVOrs36rHW+j2oRukrAqN7R9RW761e6xutwBn+zLUBzZSm+OmgvIUCkZiGKzBe/xUZBfqj3
kkoZLCTVPBZuPFHqNzdmQ+bvJlGZkVstjLUMkHlMbCe33iBXxk/61vPkUsX0HppiP7pRFaRZQQJS
UuzseAzOcM8kAd/eHwEHJGRu/hTBh19If+fz2c+EHrUN0N9DUR3sJYGtjrKzFbcyI+2GkVvZNNHk
RIxhR4wCicr0k9heTDw/jWEdAFH3ol7VJkPbXgYY+we5Lg5ECALBDYJXlAtOYoyznybgYfd7UW1C
o1U2ABdOk5bYzVmbTa94S8dk+4Y7k1vlLJxZ9PwkKu1aJv9pEtstwQ9CRvg5nW45cIc1J814pAXp
20bj2i0Du7ymrPq4Lwn4DPzV3TFK51PdwITpYkpGusvgZnVogOT98UoY8zRyQabmlPxoM3Btj3BX
UlU67pRxMFCu2FNnFCAmUVF3L0ZggGzM4POlGs/sTsKwia+V4PPERMWCGr/p7010p7kkpN5E9PTv
xrmMDb4ujZFNH7dfvwIJYNIvPd7ScxI+tV2PZFg602m8nXiSa2YKa+mXNyEvqJsYXhobNDMBO70n
eA5cpMMhLpjd1XCWuD/qeSti+ssL8v3jVNsElor+HMu8LiFMaANDQ/QAvRrAZMuwKhbETpqHmI2c
/bezA1YwtQmxK0M4/2/eQAjXQbG/sInkK+zkMaSccJAixFuyPjHi4VuJmT3au2JMrL5BA7TrAGNM
qoYZ2CULWMnSKx1L2yjtlzm8+LEruXmcI+JX7GMuWaE9+P92opOv1Nn1LQTf7AbEzO9/kGODLgp2
g5FD+3MyCEOvL12tKFs7mv0Y49tbFrzZzPY5KBwIheqRTghIszm51vDf1CBGBvKc77pxAgvypkst
zkcRaQClJLs+/QpMn58sLNMpo8TaCFNr7NcLIa5R90hz+r+k5phKtYTZ0xj2YfNZBVjA+Tn8lsFH
vFYhmPA9d8fqP3y4xAJ6ZJNItXadhJJbuyZdhbRIcSqN23AtJ42Iq+7+61tdNnWfZTuOcDp4hrZZ
RXEzgiorcQuFQE81295b6yTYbYgTkSqkeVyWxhxURoD4FbH/Q6OMcVDsBGnZ6j+n3FmmpU66U4h7
4t9AN6tUzmTT5iC0wsjjgeqMPsdVCzj5t4CIJSRUiJ8rwwofEmOvMAWu+hAUaqi7ijItY2YyEnik
ByEubIBwBj3hu2GcChwj0hJHPwAdKLzwGWF+dVNt4tO0PCph852NldVD4e7MAE2V82w2kDZCUnL1
CisNZeGLo/motsM7BlgLzaKuHhGs8FwXxkp9hUcOD1D6kTHC1UzCZG9Iwy/R3MXa/YKpQfgDKJAg
fFO0AtLtzsyk/sHlIksjsIAUWslt3ZmVh4ZAxpQsf2Q9TgdBdJfB8qK+RKnwCT6PvW82I/UzeAHB
gBFyjtikL82R5tstZG8aKk0dt5GaITrm9m5Y3p8WFJfPvs49kI6cTrOd4CdX40jtF/6tyOyz5wMs
UgjAbyS6jt5SaYd/PNjIil/NydgwkgszI5dTr9+MLmKi9zZGoKSNgjAuulVg2HOeaRrP+6PHBNSw
XsgQCMSEgP98lL8dhf/HJekcAs9gWQoBE04fEjjyeAVrMJJFcDR7uwsU2g6t0+cdfra88rZFCRoJ
IfBC6NGgd8nNolqwqAtvKBMglzsSsyY/j5I0zdi70OVRLdat7vu3SrvafgImbkmlhV8vDy9OAtDT
8bX/aJqi5YcZkIIKlQh2whq30f7V+sXYX2ivbvrmUrOdMVGww9tLfTkpHFpvWGQK9IBopOHJOb7N
rRc53x5eyTLxoLotY9XmVnkz/cI7dF3NemKni3vG5ti6RG6PWuc0GUR9xZDz+/HbfXvlc+VLQAQp
kuGqVA928Ae38aRvaIUOpt9554BV39LUb7MHAfl2lYGnCdbJSIEUWfOG1IERYAP2I/W+bWaIij9x
cGCIX16izxblGHCxfuQ979ik6Q3qVzEezHXK5dKQ8X1X+unimgCryHYyihVhOO2rnOyEApLpVKX7
Ho1SiqV58si1zDzJQqNn9n+mu7+ACE3+sc9ujjRCjDg8qTZp5c2Z5JTx6da8V7Vcr6behxr+Ffrd
s+YZwwnAHgFPzxsqRcK8GlFtdEQysAWTeLetSWB5nTP75y4Kv4w98NfdespfUQROlr60TLSuAKnp
RANCvGT0Xh/9EoZpOugKrredJIUYTXaKMzB6OhDEtYkbbIvF8TTsY/aGQ4ecML0hHl6wjbW6uQBX
cG8Oe3spkAmNt5sxNAZhAJ9CtXAFOKBzG57c83dGXW3+Z3N7zSyMvSC1dydbcmcepnLwwrxzL/SA
HO8bW8Ibz25/Tdb/awn6qX2/BiYlL9AbKvH4Al5xqwNj7sgXAiUQ57SEQGvlzqHm0aBsU7/9PwxF
FP93yES27vlQtrIXurntzlKojsH4SkZD6ud+H78IrCe/z7rtnwNd8FJ6wnw6GJCKU5ulEelOHXcw
c0m7S6dTUntML6MFkKb+E/wr6OsWvC16ac9nGp3hfoM0wQPEeuij1r1u3LP85rvjJfx4IYPd2O3f
U8CXc9iIclID3c6cPeKE5Rr8vK+bzwAFFCaDYOnY5bSAwKKGRqgnZ9Q+yujIAYIZEOj/cgIwAG/m
+vFjgH9dB2KIEO+YfNXoXFvlgVcArCmmpeWZ3N7b9Qm1pTu4JcicFTZ04S2cGCG69oA5pwoDKrIl
KQer3Ki5/79ay9u3+z5imbutMdzc2TaQgSuCPO71+iZPwt1reB45R+xx6a1dWwvMLI7WmsKTnyVc
+RZr1KheJkijX4eQhxi1B1CgEizo8sKvCoW5ZO9GXudK2nOS8kgYLWFe9IBt7ypXXpIhho/4WSIJ
SpMdH2gjffjlkFNw2pgeOIeztTvDnHEiePt8fI71ShoIytEr7GHjW3+WAmUKYEfmWoVsihr39TAC
Y+tb9faQT1Bx4wyaSh3YG3FT5Rjxr56dMZ0JpdL+PpW0Xl7+eB8MUN30ZlJ7HpeEYwMpt/rEHMUZ
1JmgvxW2bTUNce25bDbOJO5crK346xhX6QK3waZYwrlt3fduQiNq+TyWO667zllwOsQ9wE6/dR0d
NhRKCDn3R7TdwDUrXkOq5JrC126VXPkzLGVewHr5thqcchalsjnecPq0Mc9XP9DQHHQFbqLBkOB6
INSD0qkeNgyp/8XcbwztgMyh9M4gdQzGSBbvi+ZnzIQR2vqGdN81/eIDS9VC8/v189zh3KsGz96y
bcYELRQ5Uaora7VWJLS4exOJuxwfZZxQ+LWqenah9DNV/UT6XYTviFTOsbEcr5WNNggXb6JaMPWX
0pIT1SUR6FV75Gsfl7nOhRbO8TyJbEWp4fGQ1Fzhquuw9D7pN8VqjCzgvRJ5Cmb6vedfHbaGdTwA
ZYbGJ1pr6e+J3Rb5sW/CMr+wem61nGX+QhxYMD3dToCTrx7fSCpIY/FAdlOvHMxUtvOUgji/+rJU
sr38KNXFisahZqptSm2hMfgxU4L3vtcdip91JqRoKhNUF0MzoD8g5NUIJqzg11JblqGceCupXTU6
NlW8R24qqeGhrKqSqYnzdoVBx1247jSudeOOOdZcCa6nUuiu5iiS7AMcl703yJUupzQxd64lfs3r
897k+NweDIYBfelPpyte5xb/eqNCQNMtky8rd6rlDoaZuSqeeiApfARgQl9kbrsNnbBM5F3i4DuV
xtmC7BbNf0Bm4cNIAIKZFSVzXPPKYYMIghI+HdXEfda14EIoyJ1PW/O6h8uVUnZGumjCQUuZjQqL
Vm0eaK5saYqDgyKz4lE/U+EfBDhpTt+Ne4yM+sFRy5V90nJCVlFE+VHRP/KhDEsstp6S7wkaAqPY
YeJtOzxya7zrL0PXs7zecRnHWkGP3f4XQnRprp0Ta8Zdg07UzH8jUk0+eRZr0t9j8u9gMjF9Inyc
B0WVqJkh7zXcv/Rbs0djJyGmD2ol6Pd56yzcx4vn+E1RlvL6MtdSfYBWFbW2LwDmWVoyR7bWFHqA
qxXZQS2ItM6uzlktUgY+Nk7NTm5S8f+LzTEW38RoPRKaQyjSeCb0xk79gXJQR6ltSKJVdjVsUbio
FdFh+aS7gWd2Q/NaJIHgH5DPG59b00RFee11FzQ6f66YZ8FrERG4u9jXm3DPm/661XCqELopU9Zy
XuuXOiTjdayS3iV41Pvv/glNqKFWJGB64FWG4gv8jVlXxzovRiX8uHK0byrOUvY5Fvr5msCkPF2c
5XgbltP6PcnK9TqfrDE6LwKzpzeN1ZiiIXTLAO69ZPr4Fpd8sHWHhDWJDYcAQ5OxOR8zwd8mGROe
73zV8QKSh+OQM6YhCmLEfGyZIQr+bRWhqjQr3+vtMOulE8ajfmvLzc4qCyr6WK5afze3VFvpARWS
MArloeakbKR5PVF88lfU0/1KO5D2E1f+/4scm8528JsSVuToOu1URcxXK2rDUX1XgJhppEWQQzgF
v18WYtUDOp5m1J1HQ6qjgwglRuotC4zSxwVGoinlRywWZ1sakwaJGC6wswLxFsEec2MmrP6bQHez
wOtvd72PYlwZlQsadFigZ28SYwJmoKk8q0kBiwWd5xif1lL9TlIJLmTYg8S7+R/QggT7l9uXruj3
0wwbFIMMsCoNLSyn30oNxQG0Et9R5dBo2WFwdPOe64xrCySMxX2LeqzxPhKS9oniFxVRo9CCyz36
gXcKASpotsRL/MDwj2XQEg3oXEhxNBL5RzvIexdTHqrtf+yRsdl4vYruPGtwzY2bDBQGsWdIn6Ic
cfktEJrTEXdJKK5zLFBfiIGwQcl6rEmOGO6zXZ/LxA1iUVnQVO5O9m4tzOCdro3W/8IslBKXbe5M
NA7YO94gMdXA0hB2iv3iJ/ecTpU6BZ0tPvBrQ+QaAayteaamWpW0QIAlOZcSMY1c449EtMZtKPLE
crRf9/Ptv+ShNJKEklnLlcsxLUblkQNjW0djH4s7ZWP4ztrH9BljS1SXC1v7sPZ+zgq7eIKK5j2v
QCeeLZ6xd+Mq5Vf494ntNfd/ZNBVpGmTSRHQ/sA0P/eg8M0lMNIc9fLBwSjtXGds1R7GWYN+KD22
CbkAqCV36OaefSJPlcDzy8AWn2ItKqZUnm0GncJ2gykon+ReJQMN/YHcEX86tbWHAYwhRfBkBVWu
JsuKizLMWwmMQ8/w2XmaWWx/WEWJrRcs6otANWQFoEtmy4j8SEzy7Y9g++D+yCAxG9t9+dU1cCKz
XZeS5vAXPjn6SSFfMOkL82dTQWfeerP/ijDKPgATjDmEYqZSc73zD8fQv5fMIN0WBMLtkRvaZOex
dMcXm2rxpDQLO1uX+VBWIT0s9OZN+oFrbdv9e3E6GIyhx94A6qatVe7l2Sth2MScykgAwUVvAZoE
jFSFPW8LL4i+bHN39aaO0KgLH4hS9UCFYicd+4nsnRC8/nCMES0EVl0sLQ+J1kH8pjC4KSsVqMgT
2ZMYC9uAIyeaRaBJaLC1/+Zgt58HYtB81TPYO1lEo+d+Cnqim5wUIXcA5kbkQPbW58oHylXZpI8H
nWBWrsHmX5T7oRarUKC2J6U4Mtt6Xi6/PK2ULFMzMztyjmUnikw8j6YHl6hk8DSRhh39JzWGMHGO
MMbtXnoAHzqx+PYuOIdJNrlGXBqHGiwLbthQs0ijZOC0IjPJQabaU9AlgOMJPfz2e7J3w3gVgqeb
QiggvaCMU2XuEkkS9rYxKTl2wOQaMnylbel7NwarHhuTvu6gM6R35UqKAwo40iFraZ5TQpZEnsYj
1ChtduItXRdR71SxBcETQ5ff7mQni69ZKezmTBRynlhjMTIpz1cEUxwNTGZwOcwJLEwGq3yFbDlA
xxmp1rDlFF+JHiuDhYqIP+RzOPMNLjhEkymXVrBnrO3WV0mE5mkD9bpOFUCt0TzeeJKQjpUjGnE7
Tv4sdvI4fFuznYOVnUD7owJ0Gcm5tcL+lfe8bApaVXSZMg0qFSBANtos7osdN7PMH7HPKT/fncPc
qK95UEVAsiQny6TvDQDcGtQ8OO+pAE3qCRz4lg0LBNx3Cog/VjFnoged0f9lvfAp9vvQ6W9+EGfn
cIcDYCU7sqzqLoSvdYHJf59dgT8WqBRRJ/2PayjW4o8QXP8UwMPGibecTpXfBM25KdHt1vMYWF4m
w9zJ0Dy2o3jf0E1aGeNChRJ8Y//tVuGDXtMWqXhtRtcwLUhEtkZxLdsioROR6LW1mZbSj/BlNL9u
XTP3tT9f7BTQqqeX0oNcfnODkUdUbNSzO7VjyvEM7QlPw06Lk49I+ar8uuy3L3HNy6lid/BZ8QQB
g+2gbZXxvUZYpdbymiroICrvhzqm2rQbNjrcYZqJ0b0k8DBPmBQ04ypKl2LUCYmfCr5UqrJzqRsB
xQwf8vtACcxDE4XKjJ1I6R8gxalczGY7t3TqNoIY0UXZeGM6v5r/puPpEBji4F9dsbnHhvVteU6V
IMhGTbOw490FNHVauwxhWY4s0TbWLWhjLmD+2xCSFGZ98KVoI2pWsIYEF2ogsinQ2bnfBzT2od49
69IKtqZNr/xicEwNjiSuo/gmbWXCD3afp8M6KIjpHvv/EGCpchTN4CvAXRoNG1QkYLpJFOrML5BP
VY7LAamW+3uSA+0O2nPeFJIpJi/b4TYPy++CdxPCTiwZmjyLKx4V55UIjGzOa1QYYg8NkRWmqeWz
G+mIh3K/qsDVU2RCndwliePsEC9TSTXBDZ8XoTXZYJuPNFeWw4c+W/7czTc47VVVwtvs1t/zEfuM
niDucdY6DdkoMpwEcqygtOHxakkmw1YwFdQDN3Pg0UwnLWP1bjYWDVzP2YbmF1Er4ZTdRjVGQPhc
EZ+p41gmgamVgAZ37We/Vj7W9IZhEYKjtlrTo+y/NgrgaEtpY+FMk38nenB6A4j8i80W0Y/A6I72
er3JeTU5qmqsRIpqoYshjFfCo99XdsaJYPxKqYRIp13GxMlPSpT0zDenjQdMvhHsKVVhyVw4VOFI
m63F/vS0oiJqXKmQfP5uBsYKjWgxhDNJ9jj5yWU14qesA8+11pSBar8lm+yR9hnepDSE9RFYwBVJ
Wt+HBnbPJEDt+dkazTtVFM/+UpUPyBHJXJAKW30hmVp4n0YFvl648Kyu021uG0pxs4V24+3QzsEO
deIJv15T0bQiBbyOCcirpRUiuG+Z2PYcl1jef1uoB1JG/RR+aJBnhsvYsnLXoZW1CpecdWr/wE1t
6e5IB7t4Spt2Jx/+9mkVh327+3UmMJQMdulIkAsm0oAda3Lw51tEz+nsAjXBTfPYVtDclFtdSOt7
N6RVmH1bN+Rwi8naEe5952G45iz9PMe58reft2mk+hhGXGMVUZxh35fuQz+xBbHyAvGxr4D2q7ZP
tQ+cvy4yofpVR63auyKuPmlpXa2QryPu9lgJYAiPxry6MB432x2hC4kDa4XGCqSZdckFCqhr1dj+
rUb8iz9wKjY6uYMEOO03EZmytDahEI8EFUu5unGBIMTFVLxoG+Jz3sgdHm1yJ4QDaZbNjRa83T+9
DD6BhEtj/cWHNeRlRSnIDf9UEWbMQk8yoggSvkNLyAJDpb0pQO1bmL0YhU2ilOB3l9ldwXtuLhfD
q3jwoFrPI5d5XDqTY6ZGq0cPkhNqnG2mtFN7Ete+Qeb5AED5mpQXaghUzVvxb2zEsrKyUk1av62x
GlbNDFhnlfUK1ldVL/yVnxWfXoKFR66sn7ZsB7Cq76S7mgWkzMevw2Ng8oZ+BCLRNgxVGUw4QPEC
l71Le5v0UV4uC/bg7aeQrJYGK88aVwv8sU3CHE9f9wUlDbGQJD58KchI8CEeS9KJEF51jdkk9TZG
/hvdDZQA4L/67By8VPo13//D8uxlu6y3qCft+x+F6QKFDClBlr0l7ZpK8bLNSyFzEaN71GncFEwC
JMETAhD4xp95oWEqqjcAv8TM7JpeZEgm2M0tHpEXlrKMzUtF50WNTIc2LMuaqSTfZhKYN4x4tVLs
XWRrhYEdP7bQVesAqCKutED4+DIsqYFKtk9M4Zvskii25CkC3p/EiAqYcKj6I623ZPTEiZcNyZRo
bVbPLyykCWJUpQpiAuoQk+hcH8230G/BWTSi3ePwsXUrHYL5gjTwW5ue4fYBt12RFZ7aY1tY4/nm
YsGSXGSxFVpGcMHoLaGZ+EVrIfKy95DHA3DeUSGjbTfO8BEcuBz2amDldYjxUqRDzhsM2xtwLXWI
7U/H1NOLh763ZtEBYE6CMGRNH//fM+ZrhxIwEQ2nkwRc+e5qJZXyRKMaR4oH4L9bGhcIkIGwTgsw
69fhm6MVFcmB2M12Pc8jtKrmbLO+13PC7utzex4Hw3rPC63UTR5y2JSuwtj8QnDzBOcyyc6c0Edj
uGjwQUCHDm2UCBN+LATyOpuhSc2dfOIiURAge9BkFI2W2F7XKvXLcGedWg/eQrexv0BDZCdGDZF5
lR7nTDPb8956auJJeucgRfw0M4JRLySv0wDIdypvXRIYMhpUEysFDmgpo3bIpakk3Av8eBlB3VVW
iAejtI2iNPvwu09PqlDNNhp1d+5M4/v2s/c3xyqcsbUNJG/qs2uydWTZ2kop0PhZFzK/G1VknIP0
0L+Roas7DszVKEpi/v2r40Mowti+oje9wcN4ft+C5jXMqrPUkRL0XaUn0kwiY1x9gG1QN4aGx7xi
SLoNnCOuvVkPXSV6kK09lJCuViDSFTOrNmXHjinLcNVo3vT0uzsUQITzphUy0oEJVNwY5n5TxpGH
dUqTaJxuG7b/oF9xwta79dhwUNDt6C3vw6WOQweCU+a55C7BCP2nRMMjj/Mba3pcvFOjUNpUDWcC
J82/eavRegPib8sxBGCPUBokMt3J+uhRctU4HiVNPYNB74Xd3iEzkO1dIQ5l6H13soo/Qn23Lkvk
/OmIVfa5cOAPwkuncrZVKq9y0Y01tT9KvWb6eXFh1ZIEt0PHQg9M/L3EHX+BJSpvYbD2pRVDS/6a
x+BviOxoQDbStd5wKBpquMDLXH7velEBxnm0xMmK4rAaUM+iSILjYcdzpf/Q/2j07YzKssFLdvWw
/ZGuexLsgnIoXcNr8wzvDEHXbtWN2OpK0GfPw9FDgcQDUJKoMNuyBQj3o/GGMSvzYTd5bakCteAt
n6b9KP6ITFTqrc+HJnFVoUCE9G2YVjIcWYmpn9CWOBuvQ6baVy37y6OzDfcfaBYU51E1SHwLk6gd
Auxmb4N3vEGEXHi304PfxnDa/uN/YG9QQTfMFBIVpOQI/7oVNOffpZEIm0lx8nzfAMFk/EkdGucH
SCQIB8wbuxaonDtLjAywua2XZ4ceFrhDqTLoU3aJg2Xy4JWZE+hfsQ36lHNci4TJrJe1w+5KmjPR
fHHSIxDdUSTkHc+JpYrQDNI+/C4SM5ZPd1t3LP8ikNjE6xyqwfj6SHJmqQS+RCHYaVdyraozAs3m
NSA/kMm4GIwO2gApTTVohtGkOcIPeXNbqqXJ6FKdnEsspf7m3nahYnJyhixbP02NxqmkX9iJhVBZ
WcLX90zzb2P1Xon5p+Mbg0heuay1nn0Wxg/VM1nPwhOE+Jo6SGyIZQHcEBwnC7dmmAWv85M3bdId
6KkBq7Ym0axwtN/PRzj7qEsnpFIu0qKOUphffXU/VXj+sAWtFJJvXaBhFGhX1Ouy8hJT0XexMkap
EkqJ0jpaKNTVsxzFXWpqK9Xn8K5hIVwiRTzXrKqScUr5Sodu8R9QH91BqEHw3VzI3b1CBMUipGHU
e6zxdlsqoKTZqxEnJizKrFsWq9PbYhJRweoDDpGkjbiD82MYQ1Nb3NKue84mJsLaxw0RnxhduLkj
URmv9/exemG+1a2W39msms3CHpADgcgDK4xay4QdLI4crJl1qQHrPn7Qz4eNykCNXMV+0o1WPcul
l+NR2zLUfzJ1yoHiaSztEffoXAT7NPPytrTVlTLiG1O9actX09AxyB+E9BU26YxNOUngBZYSSEIQ
PRvb3+fduyqTl508swJVgZiJybPhhPtXVhmiespoLyAkGT2l3RhsVqJ3OMHjGv36v8h32gMOdWsK
Vgsc20CAJQRGsiI+wJ407Ua07UUieqDvXB/OhrIssTCa1+HwyzeXh5v2z94AxpHviOeXmYZPzeSn
9n9Aovi9KmMxHVAKAW3XfC1XqoJBuTA/Zl+UAqmHNMJaJqi9OP8s9P/AT5J/g1Wp/P/p9Qg8nlLm
T5KTS4WWXqEr+FR9FsWBpZELGSkhZelhcglAlq1Sq7vzJAe1GuUuxR71IzVtEQJ51ZUtQl9pcNCY
3l6OB+lX7E2uegDy49hiz5WNA1w6om6ZFzkKPHFVDR4Msu220BHLNX9RlBnEzOYRWjan25Mjkf/u
B+mUKESktemY8Ullqv4FqmPejtUp2ZjZuNMj9T2JQl/nSSRyyKoJo7I1gjugIbNmXP5pJpQSz1aD
Qtv3aBV40dgDIZ3NHzek8rk/9m9jnCasClN4iFu64rEbAOcnnYOoVSQrRB2HT/JQZXEHtEf1B8Pb
Tom/3NpfUxv8DDzlKk0EeeCCNAaSP+WHeguxNpcniNCJchPJTnU8N3AvSzjOMGoPjf2T+FZYgHYr
hj7s4w3xUrm0f9sS2vvZAB7WDJsDS5MZ28XuS54HzHPq9c4oFYMdub9ggCPM6/mK0Uo/ik7kMpBM
gABT7r9hoTW7ubZMDM86c3Pi5STcZo1ewKutp6yCsad75pKudI/kJ+216BNL5fuEW4/yZwCR3YaR
s+bY4NfVbgvnhURqD0qwh0mEPqsi4QoArH1QsAMtObg6wwlzSLwx/+wnQdzHRDEwMLgbR0bqjEDB
whydiv+KMtvsAzKWUzURZsz6NJkozmzf9WLp2hzNVgwcSh6oZ2EOdsslRzS31EuYF89vP9J09cV6
SLynRkOyia1IlhWTDuDCcsEj5ekFMg2RvgkG60UgEGVtjir5Q55badzTBuuNzPAPb3/KU62HH6tY
zB3y9tLibDNpqTyPV+GZvtSq+ujedzyb5dR32vHoUlX0Pzszg1o8tMrm/VFLvs4wvDfevx6BGJ9u
3Q4nac1X/8Whh60GiWhlwTECWdpc2XG4ujteMeKIs562Kf+7Vkx5hKn44i+FA8kVqzONkXfaoSh/
0A96RXtZw+2F2gk603P5RRijHgFQDl4ikvlEPg/zsySIyHdBSYTieLMHC05sTzaAHp6CxoDySP5z
LEcd7w/7gdgAtBQ6qKgHjD8HYGszFLCHt4qbNivcslWQtu31XmqVeYwr+gSXMjfnd55sx/UL9c+H
wgWnXQYPyZax6gKfoCHrh59Aas9DYorVo5qZQxuYwhVrEItQFFU4yhnRFcCxj0xkcBXhdXefOKbW
TGaEOkgPwJ1QBZ47wIizmqp1d0oFAEsyiBPHjS0k4bfGqZzMTkbskdEqerCg4p7qepbxQOWbmJN6
YTVGMSHD9r8VEP+qh+PgfM6Bz2RzrQfuey/n2iMOUM32nn6tvw+Yn7txrWfRYFyUPCjruTpbIAfb
ZhZMUrWumtcwcB4xr+pzAR8rRVgsgh+vRq3xdAqmhcf7D0HLCOq66OLPwTTo/omfuHTNSU+ISlYR
6Cxnl/J82GDcAUqJE4XwADmC0riRMDUpfgaSxWiswLDEBZI4JtpZDBbMrpk46PY7EUkMddTnr3Lz
pvWVAqmEyBa5bNaXdrxonyeGEgxLpOZvwGgO1ozGjPshA+kbjWQeAEXi3qs5pZEBeL4Swak3V42q
GUG46ZTjLRr+ifOfaWvCMpeCWWTKCXsbjc00V3MpFZ0jJeYdxcg/DnScZ837wvUbOVKyY/fKKiD/
kESndRjV0dInxjmiBHvbsQxDrTeNgjsY7L4NiI29q2ncSlQzY9pyfYAgyOZzqrYttzBcKaU8Vozd
NELMgRCL6fccV4+S4OqDASnkjMWhltqYv5wKrrKrJyGpguffFtOjcfrbWrGyDwPSQxhnISTzJnEy
ocf73kcq9PNkKzNwBp6sc619La+/n/W5ZTUaQtmMW1R9oGtA9vzfxZqi3AKNhK5LqvoX8iexYlRc
oLPOAhk6TKZfKgFU+74jLHrwavY0nCNYG8bmSIthDt1V5DJETTzDSD7um+/RqYUuM6qfuBDQTFby
iRG1Oei62KL/CWhdpWNN88V4WsvrEi0OZwn9/VTV7zjT3U7LZ/exK43aPTkEpGNfEeCjeY800D5X
1I/NTsyjApNoQvcPWotUkXHmjHyF7a3jarsw3svyUIrKHbRNVTDfjQblCNkRLL9Lpy1uqmnZc+QI
BwyRLbjmoI1iqF6gou2gFuXut8V28elLWX7ZPkHvKOJnSeiGbYmzEzhWYEMXpd/pMp2YCxnFesCH
rUrONXCOr0vbLGRYlVJYp4d1WZ0C6EfbxWTmAu7X3nzgwkKR478xFJqcp7iiQPAkK7CAbsL61tQZ
jn9cVDovSDNrA0gMJeafkQoFDXUMhFGgWE7nt+/R3vk/PsvoKMdQjIAH9OUpnX8/rywnHg49W3xN
Dwvwemgs+KMnrzynhmFq0Vuw5NPzfXGs4QU4/06Gcl7ZH+GayevjwlNePcp02lR3TPl5E14E5TtU
mT+QdxBTZ5JkLZXoanXtYWVEeIpwzc5M+qLVD1lHWgGBKs6vxTBLNfy+EpE3kR9zADAPCKUq8/iK
2Io6jMM+5BSP2AONnfe2Ku8YCNbcViReKveL3DP8pIt7EVEge9a56Jx+D5FXMNnyZMzjBFh5zcFZ
pN8KOK7koWzrRO7pu5bvRaU+iuhCKOoJLEVHBNKBX4ZAjL55YBw+iuF5wxqvOnEfuOQcxlVrVZ2F
SPFBnReQv4RgDO7szNP933mNzZ2glOQynvGY4UGw0XiBq2IoHxO+Xgc5WG95CNlQHynhL+QIcpAb
Q3ma7rIIBShCqhTm6bURZRgazzOYOJAucKBwT8ISVTb2xA/qcPAIjSDxngMtEhsrWc8Dop85WC0H
vM/0oQzug4caFlNrPXGa91PB4X53scJOq4IvVwkUjZ9B3vnQ0G7P7BT7tqz8RBS+d7GZRdAEkXyW
6vjml5ICBinmnSFAXInnz6338oh42XJnMCxd/fJIOY5blCEzekAXqW97AKWZffJ/+n+UoSD3ToA9
rq6vXhgv9jY3JNF9AGy9ojyJ78BfmDfv9r8di/1U2W1PT1GbkOjWbwrW771FcRTxeZYUoi4efdr6
vrGzYHKbz0sBpicmguTdNEdDW7erPOCRtSsuryaVNIqWyFQkh0WPpHRkgdVEJOMKG0bD8iZz/Hha
oBUmDUUJPiS5xW3RRXN/WJFj2u5beR+HHM6mxtfER8ybx3AyT0rHORxK0YOifDyVPsCjb/j/vTOZ
fzwGVnIscPhV+VT9hv9pspIeFIqJqIJnAvWC8SthgVYsp5n1yecR8YHe0v2Xywxlu0xYyd96ThJM
8TtMLozLPnPLT+VE2NdCc8fTYgkEOgnMZorfHIq5bGtwExzMYpVnJW1AzTAYQzSPYHVIW4owU9B7
GTEwZvdIFTCvctOigD28iCwDfYDvAqRJrFCrrvZBuV4xWPa3hqFQzriy8fj860wGXyQTIIsNRg6i
uHvy3eW5FnkiPa3kDqJRC9Da4nZanxl4DXS1OepDaJwFXl5TZ36qaqwbkXW9cOHXRP5RX2Xy/5q1
dyxVcllhqxO88bWbkJzOL8Dsuipi/PdzkL7/rWc+EEDv10/qLLFk3hLA59iVl41nzwdczRgf6Sxb
lcc6HZxEr5r8Eck+oE6tZFgZerUOtEdEjZlrphO9wILPS7h2PVUKeAW48IqJme8n67f1SurGIkNh
cou6yyA0ILNi3i9+XjABXD7oJXRjru4j7Gy7M5OvNsR6AN1hpwJ3EWdIuHL+0u4CzSi0l+zZZu5/
O5U4/mdNBqPpZAhgRBA3PLC9vdySCvQU/7NCfcIcP8QteS+ZFW4TDx3vkfHhMwNf/in6tgvdmEo0
XfwXifC9CkpsnKfdlroJia7IVB53BfPw5BjBeWFWqSoYC3R2dDi1VdEcT3gqG6gH/3F77Xhrg25D
gnElKjGb2OctaELcjaqosswNfZICCLcsqFeN30YRv7JBWMT3caEiRfIruqrD7B9VyUfRLrEUzwCi
Pej7nooH7p/aCBXn949WgtYe1AvA1MuimpZN4SGSvBK63GEXtCKs28nlTUg5zU+c1w1xvcxB4U+/
aVeG3nKX57RlQxY5WWaTHd6L5/e2AxK9Wj+larPbV3jLb8fU/ANyWm2fQOWSPCc3i+fwLWd5Fzb5
6wJPA9RVI0I+k3kFYU7NZgQ/QoNTlmE72Z3vDn7j7Z0xDblwPU1JjvgZgj0VDOVI55MefIYF+X7X
c+ooJXxoWe0zUZzNZZXxebi4UNLoNKMRr3U3lgGX+Be+WJ1hrnvdI1fhjGlOsPoQXCJjKdIyeVNk
WOkMQQY5UVaduKpySM2UMkFP7w1KPqrLixFwT1iFgC+mYcOL8dSAWtYEghj0kic7rUFSGIVstQjW
E9AtnScTityadVTTcmjdGo1ThMtHfVwNSVHY69IwWNdC8619DzTq7Dp+WwD3SlKB8WoGc5jJiY/P
cnFdQMUd25uj5uMEcOfAhHEcMVX5vNvM9NrK4xx2s0pomg4aBkzoH5clnQVy3IrNh1hdm3fCq7Qh
5RyzhBP7d10FkwYO6mW1/7jXCQ/uoyOlA9d8sB8y4Oz4fH3SMzjtaBT7othwr70ihbizKdDjy3b1
DRzMpivVGFNXSsjCvuCqOIMVd0+PCj8H9tNrFIlxDPzuIjWPNe94FKVMGQD+wN+y3A9u/6JasIVI
9/5BpxkOIPn+Sg9MlQKMpcs54q09t+A8PKUcHGQMfa4xu/iXFzU/f8cBllCD9khZm4A/Fdk/b8k+
gupzC+TlN2pHF0PcJFoagiO7MlrDfwOxfIec8LOCd/kszfAOGsfMxc9pSXnq7E+drCJ7JBu6l/S1
1KjTMrIPyaBbKkfx7tO2dNfPwDpTdXvwoMyjNS6SsG55DM73ieNNc4Bk/ShO4luhFJ79g9gnAcKp
89k05lc5PHmPYu+9VAsgcpp6w8QqP0KdA0qIXyO44sRvA1/0q/wLN11ymjjjcdkgoY6egKFPLEfZ
3LV4E6be975SRkabBuR64l6eR/un5zo673cFS5fRcWERJOTwUDZHIMMtMMdQq1+GSYBhp61I4akx
6RA15hiQe/acoAZLKjUiuMY/2YX2Fb2MEH6mkuQ+C5CMR2dUrhqUKUSOOGuY/1Dwrbt7HTsw1Omp
tTdtpyhYxL74OWdU7uOQCuS7xRawcbdM6VnAcRUS8Q1XU3MQq/qvlEyBEsGGe+r0aMoit13NGS4k
8UaailguwxdYobhJiCaXSkfNpyvsB3nnL1HfRNn4nEIeR6A+JOzmCwlLcMd4u+ZVm5gKQ1VCRZCC
mhKTafFpdtqxSc9XnFWK99UV46kX8IvLxOfDPxwDclh35v0kE3eXnBFNVoh25Y1yx/gPdw0iQ9N+
nq4X/ydSvVQKqGiiHAmUgT9A0PTlOeFq6ArhhaKs3haFCru2ZyX32oQynng+Sa7SWNLn3asENMeq
XQfsFTBcPOo2tV+kGU240QAeWvMnb+lTuYCtk7zN5G9n6Y1BGp6Y55n4m/d7gz3opRr0Wbz34ijR
dESDMLk0yZN9yOoN9IEeNbw+kLSHNWCBhcCxMd7idOOfYRw6nlzPhpBzDH77F6JaLf8Akhz+CTNO
g2kSJH66VgdRhiIsLJX8a6ZAEvBn9QmUXikHkJqoEr2cOklkDYm+jZkQQPHHcBhW80yOviwLWHE3
0DtCIHpFQCxnwYv9KjUYJKgriCld3FSH1PhbHxDudKdoyVRPcqGvU4abgxG0P+VSwLluEdysCLwp
ZxwQ6nI6MpgBfsvPXN1aEItueaybeMLj0nKVvZUTvmqn14cQCRkd4+4b8lLCN3MN8ZurVGWjyRa4
1gcWnm5Pc1RTi0vcEBPcWdwEFWq20hzw6T8+s2l6l3y3Rv9vb99Ss74r+9FVYt5vFAssX7GmM7GA
HrsxgRG4ITF2GbswOU+/xcHwKMrF+QEHX/z7U3+1OP6IUvPy0/i17iNvaA7w3JVnjOo/f88TG3Xt
I2Ic6xk3MzJ0Hiyg6i4J+6l7RREj+1tXOA7poCB43QTfNJ1WNaCstFN30VHV8JDa8ZagDdHqIT/H
dM0kVFlXafNhqSLjcBnfqMKsPCdbvWqfCvt2YGg2p0E4BLzHYxVzqemuvaAMSPa0cO8A7r1JaJpF
IMF86x3o8Ul3VT7vKxp5zatTC1AnV/jdmrs2kP6itWzq1qwa/6CFn/M46snfS84eVGM7ujASDr3I
ZgjmHnIicGdMjUOZOdW0n23laJMz3NH+e11JNyHnKNEI00/A4JRb25fEfKaU/ItY31TCnGnywYip
uNeDLQt0KJwKrkWeMWeOhjIzxVewqJo+NOJ/ovu5OfYaR1I6KP4n2GzcigFmY61LzXXpersigVzz
nEaaMpwW+cMSgjxQxC+GLrj7ACwTF9EyFO+2bd/2KmtN8t5XSXxDa5AgKu9VUbKiOPXzbDEzwyJD
o4ACCWcaPdhlV3vuMSK4ueJ6TlDGHYgbTv5sDZoHBpSUEe1gZtg+jjLyKofDJd48Gq6j9T0ciDiQ
CmR5NpiTXfMIvtqG7ljVvg6DV/1MT+VIpPNVGxA7aHF33v7WkTbvbkaGAc23HqPD5Z3Lsm1aSPeU
m7LMKFNejYTSa/A0zgbNrT9o0ASVjnDHWEizTQfvYGpYo3bvpE0d/AJHVxp9I3DeBbXtoLbfdWWY
28EUbWf2ONudEmC836kwJ5KmRvlG1fJdgjCeJTTLDC6vJNrzdtbYmBH1bEpXq7wnYN8ad7t5qcZy
y+RWusn9AdBNuw9iGxctZ7EzJ1lghSNuD/AaJ3QnSfNAGmdP7zBlsuaCABt4zBkmUqK5/GRaWiPG
8oSDKrNUaEpwRi/XkN/8OnHgUoHbfH58XPcvEP0vnoVlw1qLocl+SZcM9V1BFTRWx4GxRhuc6GmX
jaCUKVv+TlZYurvLTeliJSXkogLZDFYIx0siWf/aTjRArWvNLOY1gTqWAJepJ4PpJuc9EM3K3KHj
EmLQTDnmZ870DqAn76iS1w+wTCP716rigStQTJ6s+/ubshOWh0fOfMcYnm0wFLNhgBCywrC9Y8QO
r1txEykLaTwfCFbFdkSn/3JONhnER5fXpb57yUXNZ0Mu1ezGChhRngNnlmnrML3YwmBKu8YwTI5v
4qvJhQUiNeo6e1rBpfritHY6C1UyzEHsMS7DMTteKSHh0pLyUAJ2whrDeNsfTiOu518+VFFG7wLt
kLoNkVDA20P1wKtwXNvZsE8k7bp4//G1sFcmPTab7cvF+IzoWpB46HxAX9KS4DjAav6I93MNWa7m
2Ba8DfWTm3WnAtNI1jlateyJT0T37TG7/laIw+D1hLtszk33Zx98HCcFaU6i1sTDa4DEZgZKc7zP
m4NUDO4iqd8RxpMLVRO7YkWWwuyGknMCkFOmQga27IhCR9j0zucNmPiPbqctxJ+Fqm4ATB4XjKAL
BSX9Cmch6iOpIWvBC0Jh0+bfhIb0CXeEzLjHhL3Bl4TwoUvoOZLR6KclqXy3qZFMDdbZYz65NKYy
fuRZWDrJETp23cKi7SNDcTkD127mGz57NzpHUONrYzff3gejmA2qnMVeru/6SLp45IlHzfjbCk33
Jh7vHhyOzZsyUIZjwP0oxcI9sXQmVOtNwA5CTWnBPbXvcbLlr3a0PzIfPrVCspP5UnfxDL1rGkUh
xirWdoA6ivqRUE0ExNAMVzOvoUNIU4ADESC3sjlpvmXYj73ZwuMfL4sXqC4j7Ovf4QJL1G1uhEh5
BEPI/BdDg9xtGI7f4fl5i2CyJEKyvjDXy0Ch5SxoKsytBl4Z43TDECSnj4bPMBb483zH8q8hGgO0
FLDqU6TTAUqOkrFKSYsAyl6mxcgeiJ6GEWY22joaXSLNmVPA96NBj4a5/qhwmN4oqmAIs+/QnLpt
vsAGM7rLD732iYOY5TDveVmxGYfQNHxHx61OpelB+Jb3lypIx2OkDr8tVaj11Ucvo7Tj6cZMnSse
dp7EAwrDsSOlWqO6+e2PoWoh7Ze863wzFOvSTaCZAgUQPwYzP2FAqPJCp1DgiWVltPATpXtqiXvC
CBwplsGgKTdN51D53txL978KFVMO6/wtqbBlZzBHI3DyzTdodF0DSzXTtfUSKtD+mxdSfKaMpjxu
8yj+5NAJNRWZt1mSHog4eYOyAxfeUM6+xDxZpAUkz7ApJbiKlV2WddiB5HADiiTwZtKWQ1Ug8E7T
mgFzPO/MqsqoONur4uxtucQjKVJi+S/1Lcglo3DAknfWnxqpO/FpweW7HwT+CnjRd4dlA+padeQQ
6NPffmex8lXRuPmebGBaJLFTBBL3yWlmcU0TDZ/TktU0CzpYPjsUFRD/0AJOLgzO5eDARFEguhLb
YHP+VGdX/uYA25ZKMWQriU/doMX70tgyPD2ipTTCqeMKlFNvnBurwl9XI+AtRRciifyj/ecQ/wDc
bfG09yK4Mxe5b2dHi1OJ1o9IPdYphAA/zAS5KM1fbqlrNoZ+B1QtSFf2fg61Qrjn/q421IqCxnFV
CW5WWUe/0Cl51aFysrqGqlg5snk+cuYI0+/Xi7iZvach3I+511A0LuI3CIMPhy6FUZXRpolZNgPD
fLPfmNb/IvsnyLUGwGFIedmlf1myAoR4d8xDmlsIapcKLkmul3xjHJQPCu8qJTmTY5x+esd5qrVl
kR2ML9kJHP9H9wvE7afrDb6RhappIZ2KkoKwXceq+8gnTaIQ2nHmGXLHoZ5BoP7C1Zc6Q1SPtDr8
8WwQnPpnIHCXq8RCZ8CNbIqZWF8TKPGHm1+uS96ZxcvZB5LpQpxzNntdd/Kd0Tj9rhc4oX8q1Li/
80zEt8Nu+xv41GYGMZdsfqCGzK+Dlcr1NEfwImTYwTEAXsFyWJx2MVIvfoh9niCDLmqhXFc2Q8q3
E5KJxTqb/HiYMyQnChLxyVBfNQQAIxL2McWcW4SbTC2snj/PVZ67r4emqDJYFZpoAZrOkMnP7i5t
xt1DWG+NtBjfz9Q0sraasmuJxJX8fdcHKgrj3Xs8Gl9YziH8BOdspwo7RtOd49b7mRrK6Bk2PS5/
vfrmuqPHamsQNO1DWzl/wCUDqXdU4wTUhHyNvQh3eOJL6LDVf+dfsJFc008GMkZ69SrFGuiDUekz
VfaxXs4RGH9IzYyeubfz6jAsF3HEty5oXtQcBKLPUXzK/O+6Z0JHAH4nx9bb8Vz8hl3OOhJlzWpX
Sei9JxeYZ6KlLcU2iBTLy00oAdBoUpoHObLYk6GoK1eZwgL8MbpBuE2hV3W3MrVyTGfgSH20/0sb
HnmB9XlXhRQe1ZobZ2qwjt8tIJf2EwXyAd1Ebhfjv8HcyHWP72+csiFA8c2oV8x+h+qdHyXofYrC
d0cBp+nbkxdMa+1K0jSUnRQhVvh99U7cEp9IKsj8Ef7iZtlg45XEbeP/07pcUiuFW5I5QkIArapO
qAqFfqXx7xWjuzlFZ0vycPIJPeBHdX9s3cuenkidJZS09gcnhSmG5XHdAwDfN0UjHn6JFyLl028j
yIn+onKCvnlY7qwtAsdgt2oikAXY6XzHwx+GFL98HH5hl3cfjJ8Y/g8+cE346EFWshvSa0QFEKG2
DwV84LjgqABGaiuC0bPp5nGT7DGoFLnT19WghKN3QeuIBlC6kuwmTbEl4wdlvUsUM3RsqgPYV/UT
1q0+RnVMn1vBASbNNfQwZjQUMEMm02AOP2b/crvNauFZvmE9PjGUDoCTHZi4Q3j4B+XSEY28vBPP
59RBP2brvTk8v6kYZtBfe2sFtNnnVmp843JBnkTvllW8yy5NfrqU0oJrx5YlZ1Fr5vLju0VNwRLu
WP4bY5h3PX7iMtwIHPA9W1pyzqsi8SxaBGrLpu+Xdloyt/uH0vduDwZXkHyLenhWNpBFaIFhaHXg
NUUGgQ0PKLI0/gCsGzXD/I6STFaLJMqmkOwNYpCknwX2ILyBRBBCLz88LqiLe3lktdvf4ZVH5dvC
B9hF9Dax0PV8oh2Y5/MxMQc7abHTiJDeou9uVop58S7w7YsSJNct7b9RNfPrv1pr7qyu4RfU06kt
NU5ncmHgHZZEuJn8LVS17nNqzy/QFAb0hbxJrfDQHGCIv3DEvY8nEwpRXSUX0yaNpXWHNz5w5/yb
gvjQOwKUROfVdRl+AQ+z1yT2asbQdRJFXH2NDugbMN+oGs8PUlITlSB6VeLEaAbLMnDM083KzIC3
EF7AuxcUIjXDCLZ/N4J2vEtiYKnRLPTZImecKXUkzz1uxbj0N8PcVQUBIFK0LRKyAe0MHK74/Ifx
7i4f/SPXaDEdYv4gc0eKVf2Qb5UOgZAprwvIzPWAi/7iTaxb2Q1oJVEti9iWyXUpHnkDfZpvkd89
7W1yijQU1bJLALw+5DKkqY3DyyFSZ7eJ2gOMIXeg4xEF6TsRnfv9MkqP4MPvkxXGyXZ5KxFsXtP9
cIrYrvzuHzI8a++zMFsTTAIiUTIK4FW2km6C1KbJXeMIfap8GOtrYlmKWRMzWA2kqjSpI8UYwI7H
cS/j71aGI5uMcpR5kBw28l0H9wCF+fCauTIikk4AsIgFELbtXmhISjWt1YZY8AkYWeXFITjILCP/
d8kTh2jD91uc8tj0Xfmrxk/FrErLAacXLDdgCnufDHNmUDqGS1F2S7UYYtgMu/A8ZNJ7wAkieCau
jn76iKH9mPIUw2I5ZilsLjLa+VZhSi1dtDmyxEyhju7fNIF3jGpRJKEBp4TKhtiBAT6l929bISl9
jR6+F+dFrOlwghOai+PD94tVe1bb42QcoiFKNhSaSeIgzBpoNQYCS4VuMpjJ3oLG1pY+TZn8Gvhv
wIMQ+yItxTd0Der29dhOiuhA701hu6GZsldy5aRiC+Ftbvahl8HF1w5XyM43wHX2KOtA/fl4uImL
AWmwZYQVKtsca6U9gp8d9W89xhPL0yqqGJJaTC50K9tG1Xky7YpIITUc15Kjnr5BmWRi5NMv6noo
/wp8xc7NwuF1BnVRSkh5brUBkyEW2pV9V3wnXYPnnV4EB0hJiajCmmnrIbx2hIdyHSSeD/VHAmX2
HE1ARQuQlrHEOTdIR6Dyr3QpdnTRrejdVnq+r2UbegWBsbkfL1KVT82XMvRiYNnUVw0EgptFl40Q
xOIUbM+AhXTpDvWYwDCTTyAlCXPMRv0D9PvHlrens0IdwBX4GyV/tYVu492ql5kdNEJJarw3WSYr
IQLPOCKMfvvRtm8ePbio1t7tsvUiTBAIgych5FQyNUgRCWZEl3PRYkA7bZGtetqkPobcczNypc4E
JzsNXojL74SNuj6cKxEbZRprGbNYM9vuYeTGhLtRXiFZy3AKOGycwdMbqzvgMBOSYlfLcEPUbBjA
QY5gl3QnQdOeTptE3TC9ErZzrfVJYRT5Rn+hejIoq24uYgp3YQ7YcXeBCYihQDmcrWLoh9JR9Or7
v+kKEsQRkA9d+Ba9JcFZBiE+0wsdY6mFGw3qk3FGdQmKIwevL1Gv0UZ4uIelqCOMo7AHeOgeldus
xetKcaFLd6Kw0/qKZ6hD/OmnPEL9tzlSCCfYSUC7ZqMhkwjJnuLKB+paUY1lYo4kls/RUkLDZgKo
Nt9j1MOzJRWskFC7P9T5JMsokWGCv4pjVzwnEtFZcJpBAiVe4EvTYCtn9OdBx0A2zgH4WB3ZlYlG
GiQRZisbgxK/VzYP3FZM/zP9VFktLqtjFwlG/NpeB/TYm8vyNleqlt8UHVn+cqqfo9hsAXr5lxfe
U6Nslvd6GKVYabycTuoM9i6tfgQqhYN1n0ewmbMfMqjjedW4rz8ZpqzwfGrXwWjS7LItsym2wSsn
cawEiGThQlFcQzj86vEb4XDyGKuSyHR2AieqoSwebtqcaKJ72pu2ZX/SI9SM73niNcWyMsaltUsu
+TCra5KuLPOL8Jg/Tvk4T3xApKDG3m+MTGj85FyOjBSo5IXK9xcmLzf5ozbWdbTiYkwB6acS6DPq
da0DCeG+q8lU7U6xW9fUEa3mChNKzfYo/UIpWq7xtyJmJl3+/fId3gnvFk6tYPQL2pEtQ9hPsFqJ
IbKQiB5Vv4EjMDex6H1QVzDpElf9RX+CQI7PguaKwM+Ev2kA48/S7Bf6h/RwYgD/Ba9gLoBBBhlW
n7lN9bg4mo+BypjKCiamY9vkeuitAmrhHnH37jbqghSbDdr9ELaKtDAbtz1BoCUpGKrDylD2VLHm
LRmKWm8ugix2flECwZMMmPjwbaMmGX4zWbx9V/XSrFf4X4CMfbXDZpwOHmzTLSUJGlBLTWd/pI3F
zmguZOOiYcllhONdG6JlLo9jbqneX8syJjtHPZdr539CDJP2k/zUwpt8PYxccmXJ6HhrG6/n+70t
Tcxo46gt+5PWpY5pMsqv/onpfjUmrghJvuhvqKxcJ0J8TMarRtvGPzTVRynRw/vbzaDWHDzgwBiA
BT1ldkbWUgQ3bEfThwB+iusFQnvHM4u0wgbZg/E6qmNSUsUZAPH+8MunkRm/GMyCeJa7DmcPdDtE
QRa8l/wMO6h1bg5iKpQbHDcsdhiFlWcV+64ZmYTJX6vehwTFa7mMndFWRBUAAAzWRg9lzPZ8wAIZ
Atn3b+w+XM5QE7cQPQSju0fHUBSdUxPJMmmMZMekhubnDMJ/amlS+gjTkkXoEqTgmbkrZfBQoxnv
D1EIk7sbqSgDYpGW+sQazFh3hTvQFsSMSSicj7yTsz2S2uH6Ya1gSmcItJ5UiCyRcKzFgMw7ZJe4
mbb3S2m34mOhp7vEbLgLluJORgvQPD8Z5/E9ArJd8WXd40ur4oBqA3KhC7IVnShHL3zCTTAPIm51
OmB0nLfLJi6sfN9lqg4QTz8w03yAx/8HzmzfzoH1v9nWLYy2QHfVpPiWjnUCLLzCAmk6y0PCFDhe
U99sXbvEziJHHunZluC+eFxBPDDO/kOzBNSWM6hY7Rvi5PtrX07L4BR7Tr6TJ2Tmr7IgDebZqGbf
mUtRGYFUMaaYBr532EVB2kMU/il1J63n1jl8JL8qGGJPpMEY1CYtH654QRX3rTqZMOgQfBHSISb3
WTFcPv7K1+whloA7PYAxXp75EYcxgz9xjNx1ypITeWW902Th1lTCellW2sygkaOpMoRY+PisUA9j
5lq4X3np3Hga76W9m0h50b9hoP14C1u5EmIM/ieX5qilkhAZfgcGhHIiKQnB09LuDUDYEcBEW4SV
Zdo1qD9t0TTAPgJtsU1ytAUxHu33cm3QhPH9piKzq/9vjl/HIok2eNyDlzXVytOFm2l4DPmz2g9L
LzznRgqHHuVZM5bxLlw9VrNhqheSxzcq9T6S2OxnZeJn2aL82JMuYppfNl0nyxbVSDJp9B7lA/zZ
TOEMzFyJmCFqUkbWd2CuZUn8PEYJ6X5GxmJbshtc99sYTKqkFudIMFszgwwhGy/QmJ12YfepZd54
W4winFbAZ8d9Nh+tNgXmiaUB3bJTHnM3MhdX2bWV0JlYWRsVwi/W6fq9tz5oV2kHFI89cECsGbyp
C6RnDQn4hsQFu2uhK8KpeFEtbbe0/mL7wyDUEdajTCQh0DTHWfaS3bfpYyAZd+5BkIQuVQdQb1vn
AflbCBmHUN+mWzKN8gctNx4raDKNMezYoalJKaoxz2RB47zIRlKB8OBwvn2ovNbGpOBUAnXgrDXg
pojh9kvf+SRAjG62N/VtUZjjRbfTuEqckyONZQzUCF2icKipFR1n2EMo45gjWhQxrYHPg8j/rWfv
l6mVQuq7LOg9DPWpHYAzCJ3A9kx5HunDb/Tvpoji20zCkokMrbvztSewtSd4+/RU1p4IeLO6Bd7H
i6bwDdtjMx9BXm3xatqwHpJLEUiTpRsgp0tTdyrptcbD5Oqs90uN5TXJ5+qHTFSG1FiTh1muv90x
Oxtl/LWYDbZg5HRinz495Y2GCVM78SaILbPkw+/ztHoiJEXgqv/Wk7Xa8oQw8wC345OAyA0yqj8l
llQ1wdSJV2OwpCSDAq1WUd1ZOJiu0Le+iahJO8vTC3mZiH6mvxFGXkEIJT2Mb1MzdygJub0qjgEp
n+jF8PFwnr+mGWZrjgxxfb+cjAqfon4Zk/fCXKgKtCyqjWgUp6kht3+SGZs/2kg4eJJiGZOxFuV+
T7j060bOBkDEtJ0dssPZt8bVgdubirteZdvJNAmETHsilQYqlceD+CfTnP7VDZdg8UP/jYLClJ5+
rlkL3/3VaApKU/ByCmdMCYUaCIjnrkgbsfCSyRIFZMA/6oF+dV9CZlszzytMDQwgY3yW8GU0HHa0
azS2faACUcP7u2xnhKtWiKvq+mQ6KVOEioiRackGBXHOwoFQ4eWJmgrCI6eTJQCDpJl24MpRAihb
UMXz1wtZrf9qARvNHifK1Wc0h9m8DxYd1H0cq9A4b2A6SPoIhnuC7JoRWfFzO9KEP2gFKp6GpnR5
YmLwQ+yQMoEEAnlqM8OgmCNt1D9VUHNLANTT84nMZconT2Iq7Z3qJ1NXYkRfttDeZV6eIva0f76q
8dFvpH/myE/tqu7ZDas8HJ3tvUvTOysjVThLQAVBO5JWjt0zRzSxCS0b+X0ucUMjDTSmeCfatas5
9tUwwcLZIZnOs0NqqhyKIzTCTUq7Sb6Wdm13az0fJevsM2m97ZHcYGYK1dwgKgimOUG6/+2ajSA2
ST8zhuVatiIQbUZ7fn+DIl1CI3B+n/rM0zVF5Nbuqamady8CwVOPo8+xmCMxnKLzMlh9+uGAaL7r
lQFlYbE05SZv/5eR5GfGHuNSgk8BPYOjVbKRoRMNLnINjLWoFnwr6+ETYHYrfsw6xRsns/Cw1/8d
19qIOPZViMZc48tvCkv5QZTrJn0B0JJsPM/VUnkCJkIfHPMfoKY4IZcReltd9kbF6EDYSY1a+XuC
QG7nH//Xiu+zXOQ4oyHieNy2lE5sXezSIp1y4a+Br7hswKrqqIxUGgvqX38PIiHAZC8VXBkfY/iz
mktKH3O8dFctSPuOnhALqwzvUYyj6h/DA9BZuos7PpBxmwPQSHEWF6Q3qztsWGeanPVtzUjSkbHN
F1zk3pQw7D2TmaHOs5LZBoYFaqH1KprajJW9A/DKA1O3USDDpfLuE666nCOg9sdVcgjQwBAm20mV
t/q1t2uxwijY59ow3apeT4h5XmZHgzuCcVMA5viCAU8kCHJyGIkoobWOjcDATn8YoCnIm6CxQGwb
GCnDo4pndzg3fZYIsFyFD8Di/dJCd7+Rxe76luvKfpuOhavISaHDz9RwbMHNJjzNN74KdAjOpEj4
QdNyjPb1ZnA0ou8W8XYndN0u68DK6VIDBbVb057aNprm+Eh49/WSrP9EpN6fv0FsJBHg8i0sercI
Fd6xkQ5ILP9GLXghmsaIVGx4iBQuPBHypd96ASUL3LVCKnbPZYO0a8cYJ0iQLHDiO66pAfCICp2V
TDIujDN28/As2q9uwztgsWN4EWQ6TTr/YAe/Auk8TOZAEYkifsZBQ17cisft0xi5bHPyOg4hPkIx
gQXWptkxGkgl0NSM1iUEAlBZ6PqUQLElVQlRSiU/RUC0qV2NUciVktteMKc5NlWeoBqGeno/AZdw
qzS7w4mq+EYSZfIHPo6ScQ3Pm+BlOzgwmxJDEO0YbCq9NrjpcFxtXmJtyCQp3bkncW9VAZRB7aPA
2XMH94k8G3Vr1V2MwnTmvj+o6SwVHeG1WaLtCuSAG2DW/5elbsUPyDa4NnUBf0vmwlqN4er4f7xP
6/Vnf9RkbUoy9n4KeOnBd4DmbuB/32UVCt5yrThK7S3scZkeVSq3mXtiNjGcObcl7sJNwcvVqNya
OP1EQhVZFVOLE69o2Mjgprnfqh5wH8ToaWP6fhrqeH57u2qIgGe5XlpLSHicTQURai7PadrTIuLw
oc8kQwxM9uFgF1sdnMETeTELyCtogE1Q4Ibinx2cDNPSn5cyk0NMm0ixjkw4k7jHNvV2Zv9SlUAs
K6ad39bwii5Fyf99TclxP/cUem0f80/WwJiaHCWcx/UxK0F3kwdxcw1tSPUs3O+cHZ1+nKi7K0/b
h164PC5tFGx+EVdtUoMMGjAEMQBG496q9tXnyx73FbHzlSqJC0isdErOPYRPBku5j38EaYx/TYEM
m6nPQQx+L057zUzeP1BPd9W4UDcnQuRqT7Qj/k43ZoyakKQCFFLa48flFpTPdQVibZQ4kf10l+YA
3tohHeRTLgW+uoi5BWZmnQNCjGo1vAB7Na8+9hGcBDBo+thrwxo9FSoY/0Dpg62wOydnVVbI1XBi
TnU5AKQcS1Frl/5eT+YP6+Jd4h5VCBVbuXKUE3lLbUbVFAaW5qXhGRjEWK2bdMH6hVK8XMWM3v3Q
pjI2AT8FjHOejAse/jza0acf9siqfPiNt/Ilf0y/PimTJeiqVew1Ygvym0vFY3QubMWzI7P5/0Nc
JlRec5ulfBxCW6PQOpW5ASWNK1ZDLX/PrscVKyJswFBy8QiIXKnnppu8Xp7siC4moWVvgKxKzDh/
Kf5XrY92oYl87NK1xxtO7bgoqmrtChypv9ggrSURKvV9kEwJejlPM4N8Vu0yaFgd2amuhW+vBGE9
101/FVsfEnJXq5pMcewM9dTZ3pW76Et+gfDWVsxoDUdUWro4odESeGZyIAuGCLM0tXyxTPUbotpQ
R+SJIDglzEgnKXyewI5hXoZ9qKfheg8vQ1ZjpGvAo+46RS2/rR3rqKclxgCU/EtaqM2hgKn82BXd
SYtn/v5OkJYti4sWdYL0vgRv8bCZqZMHmhcBtKHStEYUx8qh0Yf3lyUIpVl6Ba7I6Dq7XX6uI9pt
X4fc+BnuSAqnUax7Yt0JWwqqYS+KzRxr4TKg2TBx6pnsDj9ME0//8t5p8wao05Rk2rTV5UtlZM2m
pRkwZepNaHHRjHmI3TwcvCwWtCu1Itb8SMTpqfX9u7T8Z0lf/+4qlUyX0YKe/iyoWDTmU295ghQa
SRn5wI23oUbYhVTHxOY0tjtojY5GHJGCSUHylk2C4PB0T9fxRf49RYzuTwuIVRKf0oFE7HfLl5e0
iK1jhFsnhSD2Dm7V8MZYidVYxrrGn6ZXlw2T63ddu1kzIFlWZ4Yd8C7khFCNuqY7YA7aqTueDxqO
SLUlKOV1qnlT55u62dYlR+PzswGZsRC4k3CcJbuaGltFDKMcGXdeFen3M93fmD6KGoQmzNQH1Bv7
/BL5AcmbRgNv7V6rqiqK80VJdVWueZERZRJd6BeuoBLOQpWROdqOgeIV2oW0mXZvcSa+ZpYfEupm
NkxHrZU6LWzW30DWcL2Ep9+EyBD6kE1Do3EeA4J6277AdBKyVQXscGzXHOmdhdXkV1Z/PgxBP/gc
i02XeFI15r3m9wW/8NSeipSeGr2+L53zJsPjT58dBbg81hIn0s9llGgc7LzYlitGyQUd+SA4YeOS
T6GQcy85b4raKvND0aL5jVLM6+5LSTG2nzQzhArQf8uQty8Keg39EsCEMVUlw9LwM+O+7HDAPLUM
leXQpb995hcIg3WwJfrgbzKNy33twWdyDJVcKSS2b1NvQ4SLDPLug/s+Tnaltp/fWcO6bkjkUmWD
W6Fnmtb8qhKFhNKOb0O/eq8JeCVvn5bsjxwEq7z19vd5kp31nOhy9iMp6Xv1yb8vUm0DfCzm1Ekr
pqn/gFh6G+/phXINIMv3zsnDahI4EVCxntbuQVD8YbcFhhTaAsA02Z6YR1czXIgTDn5q0UV2X2ja
tw1Rai9QR/kUuU6nlIa8cLXqbFNLRpNkE843m10UaS8kIOi2Byb1xQ5HHZzjDxCLGnpp/ZVoLjrT
Ug/o/ZU2v2/A2guPIa2HTUmISP8+lu00u9yj5k3kmomeAw/LHALY/rnvYDRw7m4EF3adcnb+yQfm
Fyg0gVjk+LkDMIhHuX1+6MopU54f4xL5AcOc+sMgtZAOAvA72C9+AUsyjq6fZtt8BwYDztPJZqV+
OqgiL44frnNpPKBC7UYQH7WgtIdRdYbV+avWch7imJAdxHTP3Af/Tl8nIZEFX/hkxVWQgO0OqU6c
mGrx5CB4xi5Iqo6O7SzFNnDDrcakMnX3B1W/3prZ2/Sz7qUYnbljSPRpWbHn+UW1Ct6NFN6QF6em
nrspIeXQpSoxxdkKC6vk35n5zNApVZ5IiZPRa/NEbk/PTxyiOrPaxCWx41oFTEKphru1Qw8iHOX3
jzqaJOEVMzB5QpPKFB+xCunBHMRGLhREsijUnofLbHD7YVaK+7LoDJVRQReXVFpSUXnVKg0Xi5OU
HbXAn64wE4ftzIe9t2VIZjHmfEfWvWay4yFsvfX+1M+d8fKjfndRf5025IeDBIw+fgEDTfx74ZVc
sANvZ7VKd8hYCWDTIFapXYd4fR/Cw0zgHDC4o03R4YlW60ElQT+t5L4cBxtTwSR1BKgZfag+POAZ
OXFQ8WzGmrMqdi9uLTl7iqF0AtSKzbZmQT+MjEftJhjRrGGHSXna5g3d6TCB2Xd2WIMSE8NKXjND
QxklJW5sd9/656AxBB8Snu3LpKAsdzfkCs3AilWugDp9FfKrf2Pu3AKJbMHbJafu61O2PT1qRQhy
dh2At3j3FP65cTG1j7eCO8M2GfImaEp0KJgHhb5VFbiJ6sU4wVNLdDUNgvWlqHt37ppB+dEaT0wL
6suuO8iu1r3nLGqj0D15uSn2T8bG8s+scQGXTR6HGjsXe6meUb9VIRfqcqJizDW7HGuDg+/0E7LF
tfJB2WtqzNwdj1JiZl7GGL7y4WarOLXy3lh4vy2J3o9kyk1Xyqslr0aFmMKx0eyI9nJV5Sg+St8c
uF6NdTj4mUsd67cGCm/aTGO9PFSTk/4vWz+JtixRJcOq/MjkVbXUbl13FK4YccL6qpn3wR1tfz6C
DlkLKyg2EnMYAj5w5nQ4IPcD0cuSdAfanNgFalC9x2nisdk+0YDrb97CZENxGSXHbthj6MIzK5G+
6+lzCXkSNuve7x8QqlJRKaw0Xh6w1ZjlnEEacEC3mZSNVDJk1remwkSRWI0uwVJUdoeWNXmdyxkY
Qb3BUgib0b5n/TVaG7Ojv+KoPuryGQ1sSchMS/frhyQZjK7t7xhquUudcnk3xeo3PL6sX/Ge+bJv
O5Rg6lhRwTjix+HAYR10o/Fa8XgrQ2wdWl+ehZZQHa4kn/puKwPJY3fFpcjIjr9+69v4dJNLxCgs
G4z92n0mrRkVZvPhde4dWoWt9jblpTLkdFq0XNwfcIpD/k2nsgXQIYwnyWaVX0DSxPcZUJYvnbm+
w1N8lZv8zmFSoUkFYcAQlln0gl1zGiuUZw/IYz0tUrQ77bYRXXg0ykbMU8LrlQ9AzxY/uyi+4d+U
zsDLSzfHJ1afmCzLyzyFlG8GcycyQShoRq98f1MGoakXEwJKS5pvLGSUEEoM0SgM+LCFFJNoKdGF
q18Z6sX2wkCHEG+BptYgRZUGmT7YkxFA9zldSOWXP8LR7pY1a45n1wSZ5EYnX5XESjZzsjBkvmhR
UuNGSkqJ8yeEk4Ywy66gY2K5/+ktTGrvGSQvFIolsEAgqcg+cNB+aqxLusmzrEoz50xrDcFC5LxM
1UsLAlxlIVa20s5paGmchUKOsdHB+X+KFX2Ozs2axfv9JmmiKBQEsJyMsKX2TPPNUrO+2bDlbQvb
R4NXs5Jpe3tXaU0fS0lIwJecvS46EYdz9cH/FoIJvbFwRyy7/znwGSnllDWJtB+16ZtJ9VU/N+ZS
dHpXtJlWDO5ki+zRfKMyknGTD/u6PPFvZQlD3QUuBEuYGxcJg5g63c5jyEocFMCo/3Tf9OR3bWok
pjP7dINOcgG4/jaj1ciyXr6U3DVFnzF4d8P8DCGU63Y2o4kYyrLnWa8omrqXJlLTa37qOjjVHRHd
GXfw12d7kc/ZiiSzduO34wsFvgjhemaGi1JlrEH6pGRr4WG+GpV2wmd6AP3gHl8UP0lT/8gEGfCf
2/x0bOYSTwIB33i8lohXLAlsow2wnO3GOjzVZ/SK0vDRK/9Cl5N1iHZwT/7RS5dFdVA011kqejL2
LS8LHzPJzejJQoa1+W6vNEAnMCgyT7JZODleEixQyrvpM05XIr5q8QzNB1CE/qmj6i9mvPuU26s0
2yDiM7aoX3pXiqSUzx/pU6o1zZp2C5Yb50uI5b3uu84cyii02u/XeMmdAbENVcmeF49vY8iem/Xl
3HRtaDam042QTuZ6MOfMhysU0qO8nOx5NyCOnEBWrOIuzh613DXVF+yAUKqPNgApGdCRzAK9NwWy
0iLEo57GEDi+qDd0+ImwgQytDG/tKQAlSYZnR9jFZxZ9Zc2mC6h3qVbf+AsMbm/n9dGNFFHCwFN0
zwEwOPPWMtknLS2raCVxofSduB/eoJfHjOADKttWNFUJONrm1Ufwrskw36C1K9QF+hwXdzEnlXc+
aZsSlksVfTu5mn1VPImaVXqvjobhrT08EU3y9FWS4nbBRow7YjgeXceibgdZVdBZQXfy8r4pHJqK
NJTiPV7Ke+2LwGm8hhxgmY8dorvHqygVagnb7umoyeThEOXG/eLiqUyNCQvD/7zpFQjTjIsIdp5I
ZbLaeAC3YZwAI1XzaAczXToTek3vN3dqJGwMinyHN5pucppEo3y3kYyb6UiK9fZFXLlb1hxdLI/P
OIzsYsRMGjI/JZN4NVP/mHDHylvZH4W2hi2Zhf8UujmrhvRLSJif29RlOTRn2CfbUBhsRiDSE6EG
bwflfzItIsjj2W+t84tozIGQWu/v7jzqYWTQfLfRsDp4E2frnIy44EMiytjnfg9sAZI74sJCjELa
K4jfRE6mj2rLsg95QSwrV7Woh1CxYtRV4roTnoqy6pOp0Pw9nyb0bcv8mKW0BNF71MNyYLwYGhB2
IYvg3LI2CMZzEc9NtD+oPXAKeNQtMianTP1OzfTcGJ7LmHptps8q03/rh+VUMVV6GGT7rjwCv6xC
joq4AF0xY+3hjin0952li2pQiRSfKJ3zCnv2dZDKrwmoCjoZ5iSb6to+xC5+qbAFZx2SxjdeUtyX
A/vIWzey7AU5zO71TrUabtl9FT9NrUgmxox9/Khv2rxjUV8Kjt84vApb1l7mAFpGvZi2JA34zycQ
Gg2FDmfodb0kX+MBYAyr0Bely+T7j4xVXaLLrL26qMf60b44+gCUW5YTGyyPlmpZQFjkZj+4onuL
Rv56ycfYabmum1JLZrmBVjWQvlrgp6m2ZIWSNaJOtCs9tECCAcRNdnMEG+gSch/AdwD5ZTRfn7eO
E44voJfmMeApSxfevZzRUCWbiyrUX/fk6clq8x2BmY5Vxpqg+atGbkaagd7JJgs7bl1Z3B215iLg
E84LrZDaEDjdZvoo44KgyEJHujHLRTeNUgYAkl5PS8h8NC7HMjuA85NKUSSB7+tPOHvFGijox0X7
ZCLEn6xRieRD9bGG/y7mXnOjpiMQG9TCvyfoR5yp/cxOiE9GuRRkcXBe3x47D3m2azDsp6CDfDZx
UJ6MbGX7JU/mt2n9Ynrz4JxPBB/++S/c1pkwulgpx7rhaoXr8xDmlHsD2+EULJ3neOn/J3j3Pi5B
LZmivdBHdwbdi6XL7rB8lDzXHbw4d+G28IAB7V+BoHntpX1pKhqfkN+1e20lWgDfWRUcc72M1M1M
4QCVXNiXvSIqBUfZfKO4xUP1bkDRwAHTxdXGeUrVil7jl5hacGYM54a6Zyg1KacF83M9mrwOVjHC
yUj+nIpqbNjOFKk7rWKtq2io3TpIzNQWu4U4CqopnW7unT0UPtSFjJP95D9yOAe8oULqBe6/WZg4
S99AfyHQ1ul8cfG72uSjfVInxbJfM+4i6QHMRDwJ0xy6oNQOvx0v9FgH8gF3DFXRyDdtFaNymqmY
ThVl25MfLvm8oWNxW5rvjD/J8JO6Ck0KdxOkQeb/G/1fsuK8N4HNH3zEYOgDrP235zk/BiEMhURF
sc2siIPec1xczmSf2Sc32LfEkC8t93UXJVWuswlTsajlhCzXwDS5v5ddkMDCM0nWi2NsDyP4iWJR
f6S+FOwQIYQhh2RAYlJvR2R4rXkgfWUbnTHzH7dtv+lPuSsr3r8lk6JTXdEpBx/ok6EDflfsr5i8
urNlBxO+3sxl/llVMsiBkMWYhcz1f6i6Cx7LFdNj9bUYZg0GrT8jjwiOf68hp5c11RB1RSMqAmFf
Shopkt6+CFG0eSqDvkvvqCyTfr9vOfTLiyv0PICXQ+xSlMy73RTWVV7QKJome3fOTCjwrR9+bJs5
AfWbuhxkV2QHe0gHZdodgLoYCHSir2WdC8NUY+h+7tgrXuMOOgj7rQ4A55Ae8tF8zBZfzx4U3XVo
9hA0mx+H2lf9DlMKgQfMnBCrtEMk6cf0qcZ4UKP9DeqnjZL1dOY9N+cuZYOETc7c2ovEoDlUWXrH
EpHa4HHcoDUnaV9dN1648OBwnxvhY1tUGPWnfkL7vfH3lcDHDvmTrYJfPqq9Q844NB3FdcIuoE/0
+oVP/6n94qH7zjc/C7pk+5wYeWTcNh8vz2rzB6TMFsBLsQvGbVF4IdBnnYglEZC+ZKAdMOyqRisD
Oz9lOnCld7MR94c8M4+ha0qSjrYIPFpjSJiGxDJ5Kmr88Z7NmIbAcr/vHT0ExsEHIXPXymI8NmRh
1UPdOkqXPyDnYaGyMYBkFPnRPycJPFsD4gDLkE3AfGfXiSIDQcFlOJurDL3fUJqqkETNLjbJffaF
lQs75qvYAuX/WbeDhGubsdMrAT5XEQ7YqjzYZmC9xJ8HGaYsCySXc/b97NhPhhyba5ErxpRQu4v/
849xEzpwKpq1w6aeXZyp9HRjBbbTmI03b3crelM/Y71qaASpNk8jVEsNYqujzRSRU/VxtIYoPpyB
uMpNQ4dazIGjrdGP88++ph1KgCTWouSNETR6a/XuTKnAhBLM8lp90CJ5lM5OxNfrrkYr4E/t4Hs5
DziRzK3D+I+8qhdte8U3aGz9MwCIUhFJC4it1SBUUDO0Mf0WHPFS/anhCTLtYNQb98WH6SOZwkz6
OphIlOgRM2a3LHnLJBhzBayyBCkzpyfpz4fN2U+PC05+KsiXFjFmTXsi5kxA/PXF4MIJ/4MILPrK
R4RjxuB3R5kCNOahx+DgUA+wGJ5K41J1QhsoAAML8zlNHFID2CbiFwtGNEmjaRO5/AcMAFUJDba9
IhRg+b+ViEjWQQawmxU8LDw5DnEybhLZCJA6x3906JPT6K1JsKmxesamUQ59KZdUkfIqRHbXLWlu
4AMhCQ+GgaDkI2KP5Y/1dguRRJZSHNFbKF63ckstQnau+DXquQONSF3zOBlB7/vhXE4kyXhrhVUA
xj+7j3rvmT/hnyMnCsomHXNGzDzAuk+o4zcBxIKRAeXdOfDxc4A8699tpns1g3gJMqR7hrHsbJBg
fRk9InSBDVUye93P/DdWN1+S6XC/lgruiLcb26zOMxWKjKl2miLPmQLpmwQ72DpjxetZpBX+tAWS
EnDFLFHkhW25C0vWHfeIAwcwc4P71qaHV+Xy/wopedwlqFLUl8KAl5pwfJts1wvKcnVKCwFkkYG3
M9xmSiYxWN0hTZAHLGbTk9OFjuPIfAexC7EwB0dkTaNO/iohL2jjb8Ovb+JclFcphIQyWoSAVYeh
4wFnWD4MFo2OcqZVgVp4yciHXK7PiVuYclEnJ0znC8GhfmM7jzSIACmm9QUoYRiPD6LTRlFEhewh
OE5CMll750CoTChp0np36lP2xBHButNPQHt5uHXNWBeTvxeXfcoYgIQmNQWTr3BbKaD83v11WRy/
NuE0OfwBsUZ0vM/KEdUnX900Sr4mqbCUw42ZaJ1mLEhDydd1wBlTZekYXgfSC6/sEhTAVtwLZIyQ
/M91g2jItnPIjZrH9dEkPLPwqtL05+ecodcjBVXyIZURqPqr/0/rbzcSGiCAoFhFBGY+XZxIAkbH
I6PG136eGTADvOkwdiB1KmD8WbGIl7LnaqrGTkDMZUHe0zikCSn86IwqI/JWmWqLRMkTUhC4lKbY
pIa13F5kk6ck8+lIyyqw8AUmb6zMCxa5eu8Wmf32jtOXFny2yJJKE//nzJRWUQ4nRlBZeqLd5DAj
afOTXqLdv097wEGAlKPoDYCoGhzgxSUu29l3oyWDPAK+yXGXfaLiQDc5jzT8LIA8abSJusu0NUh5
OXsT0G5uaxc3f2LkDvd16YDBWZpK0wjcHMvQmNyhuBTJBZx9xcqq0ihI4dhJ0u3ZIABVG11I2wvO
Z0FE6+h+cUQLKViOTJZvGosK/tj0KvMI3HKvPRiMU2Q6YRHRVMiOI05OpsOFct+h/1oR/3aO9xmq
nbQlZTBFRhR769LfiY26wI4+J7lWRacUHmZ+4NCrq3ObD2ftdiNurg+iA9rU3BJO+eLhHHAIxQVy
ymVzlRzBM84sjJ/jZ3TiIGwhJpFhasHIgBv1/njUEHeu/W+lEnePZjftsDuxAxBnDKBMmUZopWvE
j7aYoJMGZLVZ0ojpuIkdGwkXQVX+j0u4HZ7qUJ4OAfifTw4DLbpIRMLUjZHqhjVfvG4Hh0NEb0ER
N247Z6PXbrWM5+2T2kX51cJNBEdj4SJGpT3o+iStJttdglxtBkRpN8PaWGRukOCXd3MDAu99mygK
K8TTMBkR/5UFVcnutEpUX01dE8fW1UPE6ZIdvgTk9yoWpChs0NnFFrw22afRNR0EBSi3TQI+fa8S
+yLkYi9IGQRlwuopRbPt88kCIGrvfNsvuenyLSZGRcDN640uPCe9MUmB3fEWrEzJkyQopTBKk0xM
4z5B28RhYoiUd8J+J4aB4JdYpsEfnopPpG0Jlocir/u6GY3nH0gzcTTQRtaV11ynAc+g0KIpdc6q
LkCXvbCwBi/3wyainE3dDTLxGv5AstXxDhZf4jKy2GSmd83Kof043Iqp6ngYjBCdReddvD3HTHyJ
isVhlMy1C3y7Kog3HQOKWHCCQMQVdllhLz3SofEummgNhvVGnfUQgr8qEIU49h5U2KF/O+s8f6wg
lIIL+RONWnI6OqQozEr+5vfOy3CwpfJkTVIK6pRuc1KrgdnjVFmNfWrnLQeTx3XqezQSa5jSds3e
nMMjD5IJQ+OfkNAmBZ52rGhmHeAcBMvFq/HuKZcakMGuRk3JDPulZRb9RGP5LUbisbvLr2SBo7PM
Grfmuj6mz7DPdh8AbccSz9EzaGkZwpYVvlrFx0cDVxXEVtPxQZcbMR1p4lMZwc4S3vePMQ+UhcHl
Fml6g1XiZL0rIhO5z4i0Har50dG7WutUT7tJPJ7VFuStEwvXMFQHjQbXXL0vS+LlfaiX70J9PpQZ
//VMzFoI3HVyvkiJIpqe86z76MavOC886ZujMEixAlCE2gJ3Y4AId5B9lY2OQ2/JdPtFGXkuzfLl
amL5OVsk1svCHSV/TMLGltDy8wZL3iyMcQB4QH8tPvN5emuFJ7IX4eHuOOdvht5+8eVgiJjPbRFJ
jYrhrPbRQ0Hv8NhBKvnnUq8ZrkrGNLaVJsATYkoySv6pUtq2nvefLAdsPAg2gH6Q4ty6B4hIv+3B
xFDv4CvWZ4hagn0ESVR4qVw630pEZEIr3MWEn3gG4rMLMn7d5UC+s2Lhy4l0FgB1EUupJF5OK+G6
fwloZOAbCXZaoa+qL8ALUJzVO+SZzGLqSxZBULIRKb7mSWpm78XbFzCiUHzjLUYf7OZRkRH9xkJp
X4ZeA0sAfvSiNRHT6/zVEINWfr5zOG92svzFHaScpthuiVsQfe7mQz647/H9KyaVBTdxQZTt0ixY
Wca3gtgCKGunB4jaJhgIIJgQNoA6yfhcoyCTpSjec+RkyNdeU1nvf8NddOA3ijxOD/0mwoBSstog
GLTfaX1kUYpQJyhOx1p8K8HN/1ZqwaEcZj/61cgqt7SqpEek+XKBUuasf7m8v1GYXxyrFOsUMThN
2PaXgX9U4BinmWXrPewB5msjK5defUapg44OoJHON4gpSnAHeqsLpAHyRwRD3KVhBIk/jEC8QOHS
jANKcGCPSk3u2GrGSef9MKD94lat41Pjn2oiyAN6s/hvAxLAH+DtNhbRJ2NnwYliIwpzOlRIUeWr
kK2rGRwaYsR64Pg6oq3+0qnGevoix/yBY9ZyUNBdgQrXAsMrG1psLvEO/nrF4jfmFnlmesoWYowF
koVCe0qvzJVf3HJ9D65ULmvBzEVJ/exbBhOU4DCW6eMb7+U77DB1iVzktMUs0wc+XniTSm5iQPQz
uIKMsa4g7tvfD2yy7XtZTggp3uOjk3wZPF2W2psShF34g6gXlIsXy0lzbCNeeVMMZgor8vyFjK7a
KHECJJMZsD302wynSxqBAdBxjqHnzlOMshxis9bi/za1qW17ZJUA3MrwLBBz/jORiQwNOK4W87G7
gnwd5gAY3n4qDE5LyrX/nXmfunW+tYtA0OrcrqhQLEhsuhVabefm6xBFsW8Lm7yU/cDcYAKFqmI9
MlRvxJ2KsJa7IqcAOBgN4Tf8efBq9+m9Qti2E7vZKvY+zXTXW2a1mpYWFc2pIztgWzqxFz+yte8s
eHEdyEw1d3sJ7+52SiK2jOmvgXJulBAGv4HKo7Kr5RN89B0lBLedPfCCUctNaJIECFJjM9R8dzvX
/J669clmcGpFBrkpkaqDgepkSdMncS2059cJKzpYZy9W7n/XXi4DhGoh2CmQliGviIjJ+mogyLIZ
wTqTYx7weqCjhtoTKEk5dfrsTzmbUBpibjyRpvz9xBsEiQEWaSe7bbKEq9rEeJYIg8ZxPpsnOSSk
9RKiEzg9fh22P0h+f4wWXqm9dI/7Mp9jcZSFg7ZnXh5sKpcgCa50qxoqkmadCd1v0TETt29b5ZoD
HOcfqIHfnK3bV4qSHZ97uVE03lLDNXyzRdaHBzMkAhh1B2xV55fBQgV6jWZYe71JIT4/JrdbuutU
Ibg3kmlHMCnU5ev1Inrva5rFEiZZMUInSHDOc7Ub53iHNnqka03S/0ARrMM+c/oRwZftFqDb2CTC
x89dRnPfB8nEX/p24DONYFqDhzYejGEGb1RTpxf3R908zzaqct/ICc5yDvewntap7W/BsNCnKWUM
nJxIexOQdT1rycHP2f2IwwcxAU03nExHu9R7OGQjmxvKVytoTU4DBA/1k2Hxfv1kfJLE3oIk4nFy
+EKfF7DCgPUEHLASlRPkJXaAMXLMZR8r3QKF4VZeUk7TpturGhjM9QVoDxmidJ9m0KLH8m2lb6ko
pxWqWPJwSx5zhNRbKkcVyqDGElKW4u7fR2aPbwkGYHZyj+Bvdvjr6fgCIN1Np8wvkzjr4zbgqtB3
G9B0X+QX9nExxa5Plwtb+xEVb345REgyKC6PbFosPIiZcpJZSjM9hZ+TtDA7K9bxV+i94MgNinFm
BoPNV8PgHwnOzZkaHS3I3copZYZMtQySd7EuvROccl+oypG8NzIUsrJH8HaR9QUe5LZNXQp5FWGP
OD4tM2lRzCGnuZgZTJBMrrLQEs8P9sXgHadINp2VOJs4lk1beggGoGob0r3HMJ5NlzyniNB5176W
pkoujDaXe/CMZB6WVcHRAHBxBLQ9ScFi1IG5BvnbF2a6PaDdPrqv3Mii4z8ZUOrhB/uyWXWAOY+q
80k5VXII7pmiOSg/QlnN+cAcbj8+NcOuZ5GY9TuIQ180FGzIe6+MofCZfIjQhL+CtbR+Sp5Nxlby
ISjYsgTxpcDfb01WxxQ9ULIyt9RTQdTYasjx2n4crnTqGUeGBcxqZ09eiLZHoKMzDjqpVEavnI//
R4nnP19QTTwFhtN9+25f6PxlffhzJY6s6lGSzj2VjVsa/qj677uLVOz3+gqi2Poa8l1mzAJjML4l
YBfpnn/YQjxleStHl5I2oi5P/kDL/Lp/yDbHsdYTEFuTnTYsoO/mAHYqwKT2KyQcohBbPvQpWz4n
l7otxbmpzawd4OX8B1PoA8lM/TKBf7+WgQykBbClWgb8SPOa8wEofCPDTXtgXrBjMmlr94x3KC2z
ipftqsViHbfSJ9ey9Erljs0GvEDlXHiIiHfHWC17q9NdRxdkHNJyscPVjfSenRonhwuLUa5ZLJNY
AMUBnDI+jc5lc3RaKq8VhBUaQtzt/4+KmT7yi+g97C6YsBlYC5rrmRUVdUm+HOMfYy+Vf3DokdRH
mp+irvgWJidIwGOdz/5lzPdMEA7NK7RVMk88HI/l4e7ab/QagDjB63HaGRwpIAKKpLaeFfFeH7Oc
zZK6OstAimxUqt5pVcXncYwo9OswUaP+BgDAeJHwnCUOG8LtwyYjhbO/YKmexo2J/lYI3YVlL8RI
wNLd3YtbkUlO5KuVYgRsG8bUgj3tC4nUhC/ZO685YRz+YqdCA3YY3QIjext9FSvGBYOBw8s/EZYf
dnskG5kVOrtuCQm2TQTB/nO3moxRYnDh852qmBsSXBpguT3sttKrh3NUXZYrjZJmM4U0ge0sspZV
eSqJdtJUzsqgUY0n4UockogoNpMdCx5fDCyKrcAy2yFNX5sTFXVoKMR03WPQ5CXconPzIOKXKfpV
6jAa8w0DLxj+TAAGc8nyjHmPgBPcxSs6B6yLYADpuyhLCId/6R5ny/wmIlRb7OuSNgci7YcFZi5e
Zg4W2KZCex3aoy+yj6v/xPj3mCMmlW3odTrzxUxtwDNoWECru/Nfyh5oPheftrKgoEuH4upxBG2o
AteQSP5tlp2SUcRmwBCRnqUmnBV25D+agkXie+MOJwxL1NmzFoqOMuOZaUBSK/3oY+MY4OAZbH0g
lHSjdh6XIh2m+nUnrW6JfGw7gkldBDPb4iv+QArVVYZ7rmjTehyJg71hFZX3ljdu1gnDYdCXZuCE
8ulP4bjGd/zmGI0NEcP1M3W+ct3UYgi0NxoY8jAsKubumM+Do7/FQ6jtqBSHvwyEFa6GnsVPKfMT
pic9qsUJbmC1Qf9fgczw07pY/3Ab2MgMFppZj1HwSEEYAdkvEUT1MBv0Lph7AUQ1Kl4BV+Ek3wjm
DCaYemW71Ou0sXwr9mj2CmEoWOL4NlFDPLBHu5UdPoENVwyV0TV5OqsBguNTjbcNx4LMDXJV2a+E
fyAGIwaWxXs4t0tr3rxxIXwnV0N/mQGNY+N+qBbuf280PMWXRFlGSuwIhgN2NmVhTfO1BOqGAxEJ
+XJytHGMdKYI+Cyz1vtXRIeQUy3Lygit8woA9/NOK8oFBUI9tTsulpMrVisHfP8uI+IWPXd9/TrO
UWbB/JNNbk0IgEalRjuBFvkH7DXZgvGDGNb0fTcb9ldcWeQjKK+NULqTw0eC0wDMa8DT+8y45Pzn
As81S8rOvEJitleZ1x+8JIqseJuoMF6s/svtgOlHuPdJwIcnOC/UYK6ECplXA1N6NaSeO0LmJhul
xBviUK2MEv2lUnQO2b/dadBtuvDPT8CV0dQNgCF/wwuSAJYJnzWOmLOTakbOI/qTFxbEG50ZVSW4
eQ5MS/QpbSZrjKdRDnDLdV8d5EiUyqQ6pi6xsReSkL4nk3Qj2pidwAAq/WsEoJBLiaLgKCQ8a3FK
D++DEv8Lahg7szuIP0NeynYn2g/S5zQG7PK5cOut2apUx3CDVFrds1Vgy0unCKb7xWKXJybUzLPg
13+SIhJc1n84sKqxX2I/ri+2JjzOB3nZPh1pxsC1ePphMDCO6xa3wy8GEtHiXR816MsuhK3ZPHbe
K8VKaWqiUK+aMh+j1TmzQy47hY/4nH6hm/dYBYQitvDayyD6W/OKyx1pSz1eUxrNEw+9wSBkwui3
wkQr331xvmTueUZseLppVapmqKbl/+wlkOH8zeP8TsxnmLpDHJU7N1DcpMNJXu3XrAi9F0vz4QE9
5trfmMkBza4LZQeiOcs4I4EDP2ujmVAcVN0IBNnSYql7KIScvpZWkUFya2U04Tm0S/EbaAOW+XBP
eABpvKAUWbuhyYtr3CG0XqZ6Opp8cBKM/VmEpc465J1nnsfJnq28S3SZECVMfiAeEiAS62NoknqO
4jWxzYLY086syIUikcsn9yXuirMS2LQKsVnorA7G/8hknWeUzmY82IhwRi0IwUgOcWki6aYZPUEu
EPY0QcMa3JO1qngnmghCPc2WgfUXr5GfzXYdcrVjSioKpRxug1zgsTiZJSSkoImAY/QazLOUu59Z
kqxXN9lpi4T7DO3Lb7BDqZ4Cot4c+qnhREgd5RPk4LJ+YxICibwYUL0fUdSmSleIXd2yRuvgu3MU
4RFnh6okYi/3xJ4jzIRFhsE9f3Nvl+aSrELOdDecz1ly/k7STUQU0wHK1coqzm1Rc5aJ+GYIfAgU
bRMGtrLMo5teyz8WzH1lo1Y9yN9UiW1HRgHNp98twBSbMdgUSXlHhgLgPtUvuwP6/cQkDgehhzvt
Xy4Llyo48pZmfv7RVfxiESLi/0xaR+fmJbxJrXr1SoocdoAe0tB1N8xxMliXxlE2b8pEThHrUIpm
6xRtWA7uFL+ee7jtuS7ToSIq8M6GHlvF0oqBzFW7k3WeULwuuTO59CH3PF1aUW21fhZNhZiNmiQZ
h2JFQtmATbfnbXri1zoh2n5mZ6F4Oodn86Nt4DR088vk/MWLhHL4V1FvzZcwbnX/gDdpsFWE1LLM
HJyP7rfx6EIP4ZYwLWtZccXizSP+eR/yDrfYw8n6tbXU0ayD1g5wNZJTfIWD3hL19+ncuE8zMbHG
oA2PTvPPWjnmmjRLwRJ1jCiG6r3F+gg1jyODvZ6cCUmaSYd9hqF9Lt/i1VfTegoKJQDGdZjP1sDs
QjPWxMHhKKeyPX6/f6E++DiFhZ6+ZW9XuKPAn6pTjFje3rbzXIpSdWkUgSrmOlshIh6TVs6MmEog
TjAqNOD9Ksy6CdsgZzInxeY54I21XV1/6WuMBTtWGDIX+SO+hIVy9Qrr1Oyi2lZtXsk+eEoxzPuQ
Z8GFdUiyo7BmhLLlU7OdygOpU91IZGr+tmvPCPgfmOxwbxH39uzQg8jAkRwYk4dK7LsZIvCGcU7Q
5TWaWzH4/Pt0WJT2P3wb/0OKi0BUegwlMiswiSQ+MDoxKzs5t9KU/uVPXdQw2AL84D5KmD0NB18/
oH59UMMgufmX21idgwXTjd3lqF1ZvC5QupnwgiojP7GUAww2l/oWa9eWAcg5NNfb078YawDcTcI4
3o7XIxclek6VClVrnYv1Moa/jHTDVnzMMiDOHMtHr1Fqd+LRa5EQM6R5QlVIFHK9O0KahACLwGN8
aL2tmSNLBTiazW/6R/0S46yt2hXZ4o1QBnj0mOmFHSK95+hI3HJQIT8U9ofyNVa4FWOupCcIJwJp
PECRkNLfFWtfztPnMcEjdMWaEGxSH1PM4mrkVqnsFBzO2Yd0B59ZEYNbLn/UdaXll3LOMYCYW5/x
wYnCo3qsVVmdbLUyWSEpuh7IyGXwE0hO9OFWmpYnGKZzok79zoDpyj2x+fm9O5wklAyyZEeAkM3p
kWx5TmHUy4WJwFXGRmnniXuf39uvHlbVYHlftNC5FLWa55h7QQpmtvuM9uvSuUnRw/rkfzYLsrj+
k+ZejSmob42sRuzuRbNSqWlETh0Gm39PkqQ1rEZO2/Y5E8H5QIkMFepRsGG118uCprt1mO7jWU7w
XGL1TP3MUwYugtK0cU1zixiGQJeenLk1w6LY2NhECd4HnhRnqXi276QLT+7nVTs20x88T5ur+vkw
OmVEAS8REa3DlnHjKphqRydQalzMurMb9C7AIaG+EVyvOyHmipzOmqnnHWhv/vzZKovIkTuPl3NC
buqyBCeTh+OVcTK2pFS6gEoCnz+ECGPBaE/M5gyR59sl7KONRI+ugxCzmJPzo9Yg64OM1LW/Klve
HGt7SXY5LNJ9TgJNA9IoQ3zroyULS5l6G26lNfTJlQe8nwZbJ8eUAHxTVt43XfKY9Ua97w7TCQwA
20t+VV9lOz3QUbOxYw9fmjOk9AJ677MCVVqHWq56P3F8TicLsa5lBN+wdceaTTvr4Mdd5wDtvusi
u/nwZ9l6VGyp2DcOyd+YVdUzGHuYHdIy8HiipB8ggeCjGUnuhl9VxztPYPahHYpdSiIAdOJjmmL1
tRY0qPo7sOgybf+Hb/f963qnEKaVuwoy2+UQDETPvjLU/7kgtdE3uZ89j5LwQdIbUFuQ117/RKZx
iDEsf2zen2/EI1NSz08k1STDmm01ylwSvvtZQy0DDg3G4fZRYGDYMLfmJR0igYU41cLCd/uXvz82
jcDxZD0X5Awi7Ig3Ezm0i0qT4+mKyWdSXkqUtL9sNKo/Lnb3BNA6pDzeRJNwpppMU/6A8wpo6HC3
8cRPgWUk5TQg433yp+ccFPz0qDFVO7Sfx8Sr9qsMaz/A+VLQDiMigkW2hNGwteA0Ik8VsE4iL1ij
YIceJ3wEyIlB9xJ7HAOMXi0O67+vIRGK6JNQSxZ3xnkzB4NICaSjYFrgFEIu5jHnYzzTDgpZJnhs
rBoDf0XdQ5nTGAeqyHZUUAeMURWnwlQ/Ru8YlxIBjFenN8aB/XuyLSwyD8/MebAt280GxG13ft6S
UuvQdmLhUnFFxMztKlurQRbB1GyqFm00v7YjzOCINlKMN4HLO8fjjcs+4HPRnyttWzzWIby7q/nL
XRdp8FEsngx4eCvSZdqf2+ouCQgzjO29gb98x2HrsU9oORof61Jjm6rW1u7g4SaFUSu4QCtbjmsV
7uRshDl5d8hy69birfLInHAA9nDSPMU7ls746aFul6KiskUsUyJ+i0YOD2cWqXrgQac5+MhJzo9t
4c9UFuWrK7ubLOX3rqDknmdRgQvlXhOwMO6J30EBHnoAcSeNY0XRcD8BAKXxmxng/yar3DOHjGlI
HOxad6e9ZFMHY2QNYIFer5c3ZVDqGS6806T0xCbP1o/6VN6tIPbFKuvaEFSJTtu2wLnLOIWDTLJI
zr4sQCjJF0Qt3tbiKqJFMK9KRwl1J3UfhE2KBJ7pVv7MfpLRPfyjA7IF1rHqhe4Wz1MzG+O2D7pK
vbY7zI6XAE/jWuoa1sMB05BwqgmDAQgqKJWceutlm5qNzSel84ESXyWlSK++lm89OoJlfDo2qKEs
8Hhz2WbyP2xuaF2SKcS1s6KMGZ6HkAXQNlfMPcaBPCd+5iO1Ud17EtkOb+/9pKc01pKkSrcNIEGd
OBgkg+bxOQdXbmRtk2m15K5J9fM/ECahRohcUzyOlY35/fyxCbMsDoX+AEe694XOUEGUvXkXpWMp
EcYGrcAbiz8btpWmoHKrRfXrXfmwbX1E6ySAFDMAJSn2KQXWcPE30l6ZFC/T1ZqqyCfDrSLOjH8+
gASRMeScPl6SWbbxbwTLep0rjBOYU1Axd9DfBu8mW0kAmZAqEiUbECxKT76li9rS8Y6eROzBtU9H
1yx+5dUFsCFy22mcmqDgJqN3NBGyydBwadn9gxUQnrz/DgSXVPhc4X6P3f4ktxRdtqMP8Wp7M+jT
v469pJhsbcugAXOvjrzCGXPu7JW2f5xeFDqxMy/2mlDYJTvvyg/N9p2by/tWz3qCLJPuG7NJ28aj
PdwHq6gpeatkGmY65A4ZGnk5UCILewr9An5rVCmzqBAeC+IZuT3o/yQ9WFnbY81izP0GOMh09+m/
8x8Y+AD8K6BUmTaAwT9KDrEyp8k9CSHm7enUkb2wqiscfif7xza3MGXdAca8nAEsZaxmDLPfzqMW
eNlihFWRPuVz/xGHjK+n9om/Tz+KgdZD1G6hgFCsX3/GfW0xeE4enTLMDvlwMyjnAREsf4rhflcc
6sxQTiUDaU55Zo60YavaC9EtMao1W+k77dQIFc2/1R2awQkFs9Fj30uElW9YxAY8f7ppTyDAWr8N
BMSh9N7s+WSufqAELdOJ6Bx22S9surm/psYmMMm/kuwkrqoXLcXakTSEEO1JmIQldBjeMgg6DRlM
Dp4MY65H16BMz6jNSViSVn9HpOaK7VUjflhiMCLkDbwlB0fDWgRxJfm/0B1zRs2oOx0Sv2K+gWPQ
aOla1IkMfGmRVUXobHbXF4EtjuUk+zFR/I4QMQh5IW1V3gLtaRlR96uQste8TRBYKMNoJp+YSkh5
O7qA86n7KRLQ+hbWK4ogXnyY5H+F78YP8jh7x/NnQcCL8vWOtaJcquXF8aNosKsGQGLEVmw+k9gN
V8cDgdajq3Dy/Ts4OtpJ3pHINAI729zreibCVVBUkJuBE1Nu8oOsbytOUdJyRm56bcjMSI3dkszw
mND40HG8mY8GXLf0ZJ+7ZFh6FzOybcR+OhuSjJ3hMwW7rO1KCpvcW1TkNg/HqBrio0tDI/k1ZopE
mfuBxkrVvsV0u8auXUd1G8Ps3aHFPjj0wjn9Vgwd3ZNEFD5i2MspHsJ/gNhvgG9AOrJOGu3bniV+
xMkWS3Mi+DSdIGvciE8RrLLqJjM0XB3qVDwYoZiKc2yBjnnvnGRXots6Rbg0xIF01uS81aDwlz8b
Eb3sxL/AFXO8+kJXSX6on/z9IHzbNNXjM1Q8HSyaR13hlgX8dwHFksDTCrkoIngTeoYbhWjYfxDJ
InSF+dZ0vLIoS+1JDEaxsWpg1u/cG10THlawyRZEn91NY+8Eb3Nfx+xvI4/cspRCt5j6tV+YwFlc
I0iHf17sJfEtKxnY+QLNaKR8/t7ib+tHdN9/GHLPt2mwN8O39RhHDSvoMBvDvh52KG1T5O883X3/
yHrrSG7MzBP6Kf6kgYZOAGqQLROJSMiYGDSWGRgazLssRd8O3O4kLqy2i0vEocacrd+RaHl32Nzd
sTnXsIJZMQopc8skHyYfdA/SWGAjOlbRSm8LuGR10uNsQNXygXok1cLN0jAXv3DV2EsMXb+LaGcW
4rOBVQRdsdLiV4qmX3P9H5Dq2gj+v2erBktVvI1lovaSKwp/TSZDqV6oTVGrbgZaktz/I+E+HXnK
IAo0XdtfKfb75zGZsm30r6HSVutMIW+NcsX4QPmh0vxb1pw/gSkA6yLGYHZ/lhK5GLXwUXOxRbwu
HfbDSPde2MuPvBgq0NF/Mrg4AXZjECBULUwJsVN9xle/im8QOzxJW0HPBcnGN6eJ2AEMLPng25SF
F5cTQzUY70uWhl6yPNpxWLNoL7AWpkFGhd9j8UBMgdaASBXOyaxjs0TY70MJcSCyqkQ9+78mzOzH
jYa2yAqpt1iZaR68dCEzcZQd1uYbYmH+eyAI0O4d4PgW+O1/t1614hMNTLpMrpT+5VG/70akNSkd
O/DEhuROBLQqe/910qgkEYOLYuEc+sVf2sA0cJbWnMgafgcPRPE9EZQIaLbIcXkzespXbVuugwtk
Ied5V2jRvmxrzhbKx5NCkcL4zcvRk6K6U73HmLsxt3+9yK4PI8Vo6lRTD4HumaTDcl6rW6/uo0uL
z1IRMaD+l1tviVj5JMlnfHp2fxaTFAnfNXadIr+vEwJiim4x7cAITXtGwWkipaCrPuXwAR+itI3b
cWsrLZfkxrRQVg20LEiu5AaCd1yT2WBaFvnfqc7uI7C173Z9WhMzQ/lvouIJEYR3NBwotzbQuTmZ
xrKOhyOkAYIG8Q4wzXxd2v9QHXHWk8KJjsZvvs04FOkFZoT6r3e1zAzUeEeZUUfPve1Ddww/LwKY
W7DmeVlyTevflMeo4yeiCZrzhqTYtLM2V4yJ2wkPCpFb+aP2qV3JYDfDDQqkdL5HYR8RhoyINRy6
LBi2sp7LxLm5pyPT+OCxEP11Uq3gxfxtjxLtCzyAtox3Qk5IoOVhyij/UVLm5fS44p2wZdTjX6TR
4WpuAUSzXkVlWOuw2G6C65js55yne8QzxeocEsQCs0oYruOvc/OM4dkoNjOmbUK5w61fzPPSUrha
ynHrrtlj6+Te6tSrAj9ZmEt9TRHxyq+yCfTqP80MFe+MFvIqeWO7LoLkfVRPuu623yiDjKSue3QQ
l6mggPe+bMpM6pJopzWZUGavw11llkJUSC8PuTSek9nnr1R0zKv/U8pHR566tyWoiG9jUFP6oPsz
wiYQz58qsJaO0KJgXPGUcous845NhATEhDFyEVyKYqGp8dLMYQpjDNAQX31CvWtQp/fRv8uIvL0J
ZvZzX6hK3cFQXC5LDFzMDmZqb5prPql1VWlu90ZRFR/6zBNXXR0Xdnb2d8kmm6ku0+Cl7bzfTwB0
WJx9dkMCt02jUf7QounPfZoSz8OrYBZyQGu1TEIfJGQOuYfcE4H2otpENxg44Tbbc3E8fRTbXk6k
n11BbD1G4gHi3JD/5QNNjdBmsdcIRj5qXuHtwG5VyEDfB8KcP8FRrZX4/1+VUQd047xt6LOyPdcM
S965Jp8xPdCXAYEa6ZABi8R/Eug6CsZ8x1FflEYpqxbQ42lIYwT01UmXQL4iLsdw/ZS1UZ9PMFEZ
1TtZ2GfSWUwYN0umVhOvFXmttkLu2eJDFz9049KemzEAxnShof0b0FgCX9w+re8YqJ3o+FGFfm8b
XqwfmzXYIUbozRi1dTDhpbBXxLVrSPZJhTJ8zZAfwuf7RgvqdqS0dGE8bP4zAj7yxpEe9kJbVNq4
dVqD7EZweN6thWAVOCkICNKg9Ztf1qrIN1AS6BNFsw0s4+AqCcCUoRBmBJgm67V0OBFhWFflLRNs
FHPIEamOUg5ae3XBNRJ+K9bx4XOlvvzDPSN9OC5+TiTD4axmjqwXsc7TYqv38WVNQfgljHxLjDxn
JjkEYw5DfC01RO0b/DscYPWQ84k6PUugYhBL/nAGZG6wLDoEXATB+LKvWe127gYCAKowBjB54AAY
TmRnhwmvKlFUL7vXmPzI12YuRWtLhYbyEtEpDBvEuh3C+9slAe0bwdclJD8LB00rL2pvYhNywk97
osubbB2NbHuD9Xoo1FXSGEg077O9VPAtVTdxkMNJjptwPcd1ubcJsc+2MUth4IeiH83rSkfGX7iU
Xp2aNrFIRUCnD33Os2ORtSZHr6WNB5aAYAL2n89KMSrWr9NkjTLYVPZisrSD6F51+VxzZCiXvuB/
YAzja3i80ErQS7fJaVKcYOCgtZr7wMEi9kcU36UfJRS8mPfgNRSH0HGYkI0X7hk9XHEqmC6psuDm
bvdOzI0BZaMzRSA8oHjw3YxltiiK1FtJNzmeR4EEfIOcv0VDvkk9LFIpTnJI/GhNbcXBMoD7C8Jd
MfzUjR/iOpojibjMD71tyaAn+dZdLVyPXHBcQxfS0gOeuJ0IPzF9MRVDbVG/ciR/51luHpMC5neg
flYbKMVVMD8mSt/Hkq3qt9nMbeRykYew07eHRfpblXgvB8Ec6O6s5C8z5QDn79rsZUwKQaUaj58y
bxPV7UJIi4ZKWD/5OaO4WN1KjMmkrEZnhYpytk/sn//eAA4lqR0xk5AchY/DHHnMaEED5KokOkZq
DCnvcHSdBEvlaVgQBbw7QFqdnHRTY//ibcth3vqb3cuBqoykyJBjwj3sYOH4hjZQk9EmzkfLuzlI
ab7THqpadYVO81UjneilHTmqfspRDN0SL4ZQCqZOA89wOi8hHRIutCfhz2p4fuG3rgLYOC817EV6
MYQb84pEOd9GhegmMFmiGB3eLHa50pi/VFDQpxbOGkIZzRl0NNlbAiUsB4boSJ600Zy/oDV5EsNI
3FgL1wuL8L3/+uSKuGPkf25CIaDw0IYLf6B3i0fgVHcwENS0a64sDszaEJKJvFy5yBuKB12NRSVl
33bUlnxi/wG/Rbe3gAYyFNgsFpsZ2GHWv2BtQp9TEhsnD+cGmDfBDkodnLUIP183mwwT0ZxIvRhm
FVmG3ArDeasNkghxe4Qxh3lZNTup5RZoATE3yXh9YPIZ6HDJ+taJCp6YZOeRzyiZnGlk9ZuxwwBM
O+uCiI2X+IZajjOHohClgkkd6/niwvxTswc6i4IV9MQsPAV+0mKDQJ41o/lCE03xyJp4VVwHyEQ8
YWoswFZbxGfns9mPxeCSlc0rtG5FwzMBatliJ1LyTvhLpkFO4i7No0cJ2VwxYnjOx4IZz0UoCPTE
tQhDjOVCaasaCtlk2D+zG1pyyvHsnzG/j5eKYF211T3ZFsSJRq4gk0rSWBuEnM60oTs72E2i9TEG
UHSutt6aNLaX0c1S0ozb7rKf7IHzNEMjEFHVytchzaEH0MUSYTAerVmPPHBY7ywqAmUudFixLE2u
HxsCvvAmYgF2ew6qGTaiwR+erb8Og3U54KIYqBQBjSmbr8chc6Rghp95vUNWuNkn0mbh7LDCwX3w
0rditRicsqLaeXPfvHWstvjaQpQ1qPkcJvobUiTzwSm3EY0mRGICtXdUD0CeIRAe5NyOvmLFWdK7
2Cqt+EnK3hAN2sKbysDReXsmlC8hlX17H1WAFXBdMy0gGGJKUiufJJOsfc76iWCsnyYHPqgKpqbR
kuDooh87UNACbZGnPrTxTWVbEA7ToSStzWFiXfdEzm7q+zIlN708lVsKriSrEnRpe/3HRaZw8obA
xlHsx+khVGKcPJYdFoYkQkkItFmOcD1jo+bYKQhkgYqgJ+YTbgPSoQFJSkRGYUVGlfnBjyZrzmbF
pbpCCNVg+rn+MfBeyf5aYiFXGCvFGof2UssQeFJZGLxQdeuXMFW4TYVlT3pM+h60zQAy+cCcljCL
dcHRjsw8VpdA4g9LeircGePIYLI516xP/HL+Ha9eJyHa8NtuDCRYfTTCXw8oxfB3lSw33O+dURBw
3ftaImWt4XIp8QXwN6W6fl1bYEGdhjFZp2i3h2A61DEWlHKWRRUVvhScafbHwWhIW1zJ7q9O4KXk
wIzYxAvMBPe2vv8rMdEJ74KDKxo/iZ+FnBTh3uuq/3c8QDP8vTcU+ev+A6SF9a1MN/kQ0CMD1xVw
rdd1WoZ3CNeqfyzX6qp2M2NEd/mdEQnro17Y5f8AEFy77rReewG4ZWILXQoBOs15QrAHP49jKORX
h3e2SOFUqEGog87pUlLaORUpYBerju9W6x20co4cEDPf+shw+zeOEsGYOeH8AqMdfudl7ciLTuFU
gMhDyatXPrGZeefiF/TSjuVarwyDGxgAkwwfrdb9CYMrbRMzkZt5qtgJd3NFWLOFa5ewSQeQKIYR
oPfR7BGgdejhYUpkEmafguavYx7qH7NS7T0LoHrBiMpiCXDDACZ30POWl4DUsJ3vXEnIxLqL6K9K
4SIeJyQWyn4QRk8g47smfpIsPNgJQVcbT3O3SqbIkV/34zRpPYphzgi/wsOgTS6R0QcT7SMFI7W+
BAOfHWHtyfF9bFbvfSRA6xrvHzRSCE4dHiqmwUPdC5RCqDGi4tDUn8rP5xcLZL43yMX/QW+IpVJ5
MbEqSvtcGxA6W1Pb3LCAafHKGXvFAn7Qo4P4own+OCxzTkGKJvWu7H4xEgPaf8j9SEL5bV++yY0g
X/Fng7vj2lBFwNqQJCQPZioID389LfcsXfS5+AofTJyOmr9a2BSNzVdRMrBV6fTzWaYDL4JbWL53
rl+vmM6PiCeO6CM4sHsGEsuxpdtYrRnerzTVXELthqW7mZ+L+0VgvCDpPzfxcOIObSULcvh1wq5H
4lIB48eztRTMarSi9ni+kAX1Z/PU+o7RUnxueJ0N1nYWEf/tpmTWHh9BW8m76RxLXotQPv8oSvZz
4A1Wz6/cwyHiLZMPiIOje80uR3JmAamRhB5nkdH4vBhMDNR67flSdlh2MQ68thvZl/D3BdL2kFK4
A6eDTvLOvRlh3ddJ1Xsuh/Q7/BOJYQyIbC/qLdsf8m34qhb3tfTkzIpe8OuALuroBswo4qqKjkZm
QZt5be8lukxDDe/mvq97bcMIPhhHnK/iIVYwvZcsMWapObKPjbt/ARhaEh2/YrHVVoLmnL3RHnSp
uMEByyevgrN1jQwGgujA7lAuWvi79mOjkbeVS8Hr5fAsdJsviV9Zgv5ZlHz7Gr5aD/RdMGagfpBi
qnrXCOyOzIDeG/ULnEtpFforq7Ac3yYGLBnWjE4cA+5DHeSWVfZdfh6sdFU1kp1zg9c6EnMHxOR7
VZ2/O2W3xxS7mYa+Fp1ToUs44J56PYlLJozKAnGNXzdcY0O/y5tI0c2IXbP8jfS/lg3OLJLV8QAf
Q9G0V/7dT4xVbd7HvkgRmCUT8xMwSmlzd8MyHUGlogc0XRSvVZEZMX3K6cOunP2g6jcr2uuIxVCf
ygSTRzZSTN6JEwRqmZ4XPgF8nohTqGLRexMArrKcQKGC7XAdwK6itG0FqtfkOheWGJDAXJEgB/jk
+GcpWNQgtr8rs6F2SwFa+/wk/DzirVvDMgEtGE5J7PljywFb4WdMghVKDwYXK8HoGdpixeI+H4ZT
RuYpcNDl9Fri3ST7ds1j4Lf5vAGjd8rxEft9TY/X400AzKOrT+9qKh/QSvlc6P0MKaso0OB5zKI3
SL/q4WOVEgF62ymvUV1PBkx90jnc/RJ1JFmekxfhdjqsGm4DhnPJ89xbLwumZthxlLMvDcFKgT4r
GUvmo2idBxlXW9BH8hrqrfzgjJQPT7nzM8k1EZmoja34U+N+DsrrTKjSPfYYoPt80gRyGx75N7+v
82Aw7f3HjFcKHLKdZiNrBoOLB7G35hJX8QVfCXA2GvQ5/ylU6g3u+lHkksqeiXWrYIOsgVpU6Szy
yFj9A4Pp0UFXx8EYIzQcOdjhOhB7KTKNkUin4PpyPoFa7T5Bp/q76v9mt3zyqKuk4wogBpSZSPi/
aAaSYrc/sV0Eubch0MzRZZvb5BaZOR04R7U8AG8B2bFVtcDTeTt1zxmbypgsTuqWd48eY8uYgdgP
BAAk8+83MtW4uQNmWtoQmcxUM0BeOufn37ICnP1cmCjAnpHGOlUAQs9mKdGgKbQsF3BksaSKNAyb
A2yP7zzV9ybgiPksAJaXpdqe9/BBHMOrF+ROgxuMsJde5zQ6E+su+u3/+9JEvUfvft/NFeJgpSq8
K/V/VHDrREYW4dBB2X2dfxBOJlXUm/WrEhSy2HV6G0UGQpMrZpYHKZDuWlINUlliZfP++1R1KB6n
2RQVScrgyLyrNCc9HGZK94OXeg1h0kG5TTpUxerGpSeW+Cy0oeuD0RocTjpkpdhfsahSLZwONrX2
xBzwetQYD9ltlqh3FOWsLyPKAE37RtY3ttQ+iwxGT0lvrmA6MUIM/90uNOrr7mSv4s2shrOYQM/a
QHHDc2nrse6vANDXkIcYVC2zRIiPrZHkCDtt3F+DspsMfAqWTTKhQsez6WhWD1yRcGBb5dB6/HkW
Q5JsCetg9aDXstLmUHdBn+wH10VvVRQYNHBMZ32VdnSFQQo6DmG1Fixtt1HvUDSw20ynbbc5G+8W
0gZxwAfRDX+4PMeoH562vAqChxDYKI6Yb6d2czaJXI64+h7no55TDhl/axTFDIS1kFF6qF1o2Ykj
rhJOdkWoqkisspYL7emw07+I75J9AxixNKLDoq9RnkizZVE0kxnKRdk1nYFrFlee1913Eoyp9Qe4
HsHuLXmLUzpCVKN+6/deq1f8nlanoGKRO96gskPtwpwZkmtLaLPkR+NmKnybJN3DpUP2xKR/KR3s
+3323cQCPZPsMdiBzT0EtkDtzr1LGK/uiiM8YDao04cHRw8ErXg4BKb3Nnk2KkIMNI/4YwNrzXCP
gh1aBF4oAJKYqkAN2aBP+EQXdfUZf4ywMItEKbJGGy+2HAfwPxTgqyi4hWd38RXK+ZijBaKRqK3S
wEsMVwKlEaoChF8KJAzno29IFv588ng3beP2f5seWWTWaQ3bj6DvSaVVfpO0WGvVaZiFicVjC/Ep
6mbztfy5Otg3SMtSMevrSw0CPKxQMB1fsC81WS8gI7SG2gthuZ7c3KwN2+VdjIz76WLgevpGizQy
iWU04SYj6+wSYfXkhpeP/Au1JGkb5fNfgyQdtLRbEVKkUjIUEvHxeJRViDQHSK8b2OLlmgk1+OYu
U3TNesBsQlo3+4/jC97bRIQLDI86cmWqhbtL6ZNF23vJy0GrcorGcpGBlTOqas0Bf6yVWiQmbSBF
+V6N1bfRZ7d+oerAiuWZ9WtP4p9Z9Z+VkRqlN/+BUaMxPwSopJ74XTZ9vDSXxxK4KYcdvclgNzDU
cGAam29CnSEttt40bYnCvmhhLO9GzPDcQS5HOVss0HqacsGZ8lFj3WEqYzEdl7wsJBm88oeyEzK8
POT3yQ3fT/lyBsqj3Dl/hzQW7N/ohMiPsrNQJRPU/3uJchVAritc+OxcPmonv/5DAh2ZpXTV2dBt
vMVTX1VN7sMvQxxBYhwhahfZ1peB45rVMm/bdjDSWpodsp/4ZuHqXWR50bNZmpDht3QQKsm7PG0X
pUgMtsB1foAH110UQl89YVupqqn8GqdNMkoR+xPlPYWFFyKZIeVZMpYg7qmCvP45910Jf6SPJ8kI
//gOpRaIzPdtRAinOM+YDuz5HXeQ53I1eozEc8MFLJKDVEi1TBxltuhdgjTBhg3QlvTjBfdY1jwU
aDvqulkO1oVBY2a1OIr+GQGkEW0Y1cINTavhSFKg5o6j0T5M2JRymu8EGTZI7E+ZHwTDkFkYNJXz
zF2IcAD37V2wtGHljKAWoO52GVTctC5W6HE+F4f2TTIlw80H55nyw9pDY11Nb6f3kE2YFbWDQkZy
EqlWniC+FkWVkokagsoVg1PItBEc203NCuFBrva3w0LrAj+r+K5tbRF/bMDIuhT9nxbsgpyPO3n0
/XJVAMd1DSoktxD5oHBZU9i+4n7DBCeQ4kNQmWa4Gn6Y1AQVTpU6EERf7kFtvTuxi30mCQSw/XmR
Dmxk88QCcFTV5BUQ0DBjMOV677ukhu4Hb5M6ybdGyGGuFjn75OLjFkKKZxEbuYpGzyn/6HaS83Oz
++Seo5k23RmJlh8AxyKWrv9UGFCHmQQRgJGAI6RcnbNQrzGV4mmkTar0lNyYbK7G7kI5nLqdlAg7
Dq0ANtNDee2xNBrzw0/ZTIZSZwj7htDDtIvHvZxE//I6WnuXpy1Lea/anpC2UU6DYfvptu+S6Yo2
QXVDDYGyUGJU4fBLt7fNjbyyvtUajtQSBGWpNOUh3qK9XctLkBOyWNPUVcGWHa1wHruonKgGyOw7
RpIB059aUf+ylB6i6FGZJMldtgX9hNpvadcmvpZJlp4AENqWmn9/B88kM8402dj+OvAkt5Jo+w6+
zMp/XUopS41Vfm3Zg6CpHAxfZvsaAA8mPfJuLwsvOkfmXXTwtfjJ/Jda4l++I4OyC4u+TNZ3b8nb
6TuAnzfZQ/QBVIM2nxChft/rCiKyJjlC7kEhSkP+RCz3EfhQnF8A9ihJi4F5lA42abDFFyejIJgW
Jbm+5qKC3gRBDrTAqlX8DXzpggPgT/E8PyM7R+mbdmDodg1PC8ONX7LnswJbiExaVqxIL8wvTJYJ
gTLoSQKKTqjWtXiMs1ksOQFVJgICB49MaDKZlF7/gvy0otRTY1si2TvQr061UIQrhJr44XHVfON0
vzk27K1RrvnIB1hs76PzUQ25iLmD53Z6LhPM6wrLORJuJlUQBtjRfcQN7nczxa6kSlGrrI3Rz5O9
Qwyjio21g3XCFl8wHezYz5WwFqC0C8mhraL3FuTKlpN93G3DxUToiGgyusvVQc3uzzajPuFobKe3
E/17cVhuSfxa4+ukV7S9Pa3k+R8Fdi39ZvATxfq2zDb70TUg6rophvlYhHQgcUSZFHNYVaBPMpKZ
KNnGDo49JpJQ+EnwAH1uwDG2tYQDescMI22e7hAVGTBZHV90RWW0o6v9VfloGjfB85m7Ahzk78j8
Yvg3LlXtsxLoS1347vE4JKbGQIhIPr2RH2y9lmhJGMBERo4ghlxHZMMFBrCdBZYixSPYV6SFZKBF
RnKoSJIiFfjXuRqYJ5EtnHy+WHhPxm6N/QMJwb1igDEK2dWFksAa7HYZg+HsVAxdmGHBAff3gpCi
AaDKdLpirDkUT0bU6ntRwvTuVMk0FfXL8lcPVaRs9+AuAUnSRae9IXW02jK7wcyY4BB0CH8bb2y/
Bg7qzezJOB2bMaMYpJ9+/H/L+lnOk8plXW8v8mcLN2UPjJ59dotZStNtsZDzGJzXdYd9AyxG+3Jz
387ROHjcY17Oo9cxriIey2XyAplx4DxP8bcp3fj18Tb61eODcXBzebWeMc/TMzeTdriyMoS14d0P
2EsnR/g9CMbvmnentRCW8mZoIIz3Ghrp5ipONDmkUrM9f5C5TLcTUD+pQRv7pJx2UvRI4q/CRTJy
+dYY9z43kWJCdRGCQ5wGib1Rr9lv7f1ASoNO18sCNstUtIrjQOIXoLfvWoir3QDGYMfojgigO2RJ
27I9EUQwEEtyP8UrJjNIcSYWljYkAszbC1EdT/YgPX1VJIuSqJoKBO3Zho5IyTeQonzWSpRp577T
EgJg5tHdBACY28Gq1ISNQmt2PXourIdVMaDpVyknerteT22euOtpX0nFYY+HFiUNb4BCia4cjH9Y
5Il/5DmcmTsgUYKZFNy7E5uHGEWIqCmNL0u0DyKLANgb1zxzizxoV49iVsNGIdtAPyhlD+fdVGDy
rTSIoOkIudQbEQGQZ/wIyIzFMkOlOCqTF1NHoLnTXZCVr61qUr+lTAwJZAD6FMd4rVBdIbk0vGzy
yDQpdhKNBHSfMgLetmy9AdmtHP5E1tSTbPnqWUv7UqdCftPEoljDsmfIfh5Zw7u/YBoBXOznnc7k
MgPBl3hbU0sBz7xI1hzyUjQNXad2fyJ+rO9PGh5kVbN0m8jV2MemWq2MLpiaFEWD+UhKCCR+o/PK
W6Qrj/uhn+jmb1cAKMFAX1reV7fFxll29UYGeuE6AFg0UzyLdiK3a+Rt0OBrO5ajSp1GHGarHaEP
hPWN0WWkIym7o/3r+MePvlXJoockG7lWpH+PThyjn+oryGtX5dWj0OhSSMogBmu/RcY386m9dgVt
CU1Ju5dvMlDgctJZwOKHgDeMcLeDC0t2JjlogEpxX1maMO+/D9KWA2pSMcCzF+SXf6xu/XmHEEMm
raMES0OgEYz/8xhL/6mOo5A3zcFXv3LvWLoafVv0QdAJ4QuyNr/2v0zd78uDwezd/xjozM//dNYf
BkmKHD0Fk2z0IC/odE4pNrdJvYd5YZpBsOZ7KKV5OiMjsBXIVys0ZqJtYISkzjiuCy3F3EGKFDI0
JGmWAEY81TTgs/W8I9Cro/QtP/fC+1j/to8Z+c0xlKLOUSBDU9aJgL5db0UTjGnD8X+6uV+niNQn
n3d3JIngPMMtgFOMkkm+VxI/TmN2AETKfp0mi54Lu8Oife4jf4HY7u11Y2NsM7vKiutmsk0RNppE
0rWN01DxULXaL1eg8p7LLd3SGbLT0EDXNGNKCLf1vjqLynxy4ZvAqTtw775XAatCmSVxlagHYaPC
kmfQDe3jHzIVAd1PSm3dxx63oCpXs6cKg4SUB/289GYUioa+/0rv6FsIGh6dcZ9lzD3YCi5Ny7aD
uGgVnlAsN5Q7xXsMPqyv5YRtBlsmPTz6cScY0oQ/l/gon/tyT2DZ/BNcR1zJp66K/H6t94rPeaLO
EfJbkdzKrTv5VAeaKn6inVuwmjtuRb9PCBNwusiF6u49QXe7z3JHBzfq4te9FvJqyP8/IgxifaYV
nXRb2i9keONkjYYSz9LSGdwwDOc9MnN2qJZq9oTWd3gGYrovuaCRjUNoeUGhgEJPo9K0H4ajw5W1
46V1+PvVXJI2v9Fgk8NOA8HF586wZN55ZcGOcca/qatWdvlq4plNv3rGL5q10VOIaEzSPm6bWRJF
wW1Sy32ezi4h87bUZkLYaBSQcGpf4YNzNS9e5OaD44GwIMOknxrqLQ69yQqFFxWMmErus9/FeOVI
Q0LcLZBzDBpmow31ltYtCYHdZXp4ckxFDvIykn1/hSJuNfcE+gWMsEdi/fyBTqfd0M+qIiHHZTTg
YVUMuzjV0X+Sb3PU+wyfNnwzduawfx/GkPDpWce6WSrrSTfFunmjXyC0fltvVfv1TvjhhJgBrS+P
eQXm5WbktG4rutHKWUGuVKaypDHVco/wWzpCr+XHZdLSvskPFBi/Jb4XdYhi2n7uHqIbz/UoWX5c
9Y7412NoLDhENGr/Ijs/9fLLXy5mG6Eg7XSsOleHrLEtBHroptyi5H6UyjqHvNFwXlzBUeQknEEI
RbBebJB5GuK5fqsdoRO45vagCQu3pg7Q+QOo5tpaiffQhsFTcZTZ3Rf4A+eeuVPyYU0weMh6ogPH
eHwLyIa+94ft7va6un4cXIGh1B9vKo16+psZvgkEb44v1cAyNiGaJtrQWRVuzHO/g3Obi6+QppH3
OPyXU0mywrax+fW5yqqmZbPb3hgJytlm7g2RGwDCO3g850r2prdFOA6PCLuExjNtNa+wvEE3QTvP
MCtewdD7ENcRzqDInJXSPXFlQWwfA0g98rIGVx9syG0VGb5yCMycLeT/QgGUHd+yR7LQTqvoBv8H
yBXFmXJxETsJFYEEX3bwb9GWqeOIV2vOp/0pr35bR6g2vym1jDSMiXEP3kAjVzr0Q9GQblkCyXsK
RxaYpSIXukyeKGlwCR39Md7+XcuOg+ER0aVs26sYyu1tXiYsEUpyzMd2SKDVNpLmiUC15f5o8u4x
CgJgvfwQo3n4qAiokVkh0LICRD/In4FtWm6cY7dQERxT73+kGOrrPGXJFF+SfQCUv+/9CukOGnWQ
iyHUHBHZ54Dp2LBJja8+x4gYNOn1oNAQPxkpzBNDVyFWhOuxNBYfOsE6YwdTBPUL6qEoY5mJG39M
2DjPDWS6WaaygsDUDAXvry+Akdd3xMyLZGwss56hQZRdS0Le/OGggJzskvaXtztaIyHZKaeOVR2t
UYAGyqU4xgg9WXenyL3QS41oXtdApk25hBzQnFrYQC8AyMtHYrKpJLElVnEflwWYGWQXlx+uw6KY
i0tqDstINOGqRIKKFGW0kaTeyAdoruIvpEuZ3ApxY3h6Mt8mujr7IzbJR6ZkshC53OACS0bhAW7d
STdNhVbvv3Bq46TYWfx8bbF/kTN3w8pGR7Uzz4XYd7kTLjoOXW6qFiZ48Kdz46rkPajhqy7X/dHi
WOyRyxLSMV9o5AbibdXooRDj1pvr2JMa8kTVZNiDy6L4S5PR2bSfK5Tkt73MUMiN+mnm/hGc/OTR
MJ+On3WxUhfO160UgvIOvGcepUjvE1hZgZGjGGzTQYpyTrfvzN61yBjaEBY7SXPsBCNZtgyl3UPc
59eBlj85a8tVO0QR1aRP9nKCKLe/dNxzHqGnNIm098ktQacogJl92ViduwZsKC+palf5TMQAus2k
gBs27n+kSAp1e47/Bx94spY54jh4X1FcB3DNtWuLOjT5l3OQXFVuosGfP0dSROxay/+GahokOHEM
TwoEDpBkoLTolv3hq/JOKVJwA36RpezVj0MWlSJ/qzjcmM5B21rLUjr1Ch2DcyyxenZwz0o4uJAP
ChNuVSzo5zbgG7mjhTLXUpApaFa/Nv97+fSN1hkcjarLWSQ++5yAty09AbGCmWIYFxEfwEriuGy1
Bo2Z+S7jWrRxfXmm5eeUhDvHXO5h5ABvbIzZNH2qhaOUMIaVWul8fXRj35xhRd7AjZ75VAa3Bukr
VuB5cBSUgnYyWiW7Afq3hZ//pizEiu+F0S97FW54uWUP41rW0uWjYEqD2lLs9badporvekckryYw
VrpDabd2CosdZ51x971vzI8rws4pJt1VED8jfRCqcG1LWPf3QHpKd3J2a7GMQiUIkScpahkbQh1y
SdUqrDA/qWPEYW34vH0Mhg3Z+YM0gOyo8mPY8iDDnhc+OtTH/+u4nogHpq8LfGSUck+Bp3Pq6+aN
lojnHiZ+dRiS06U5PV0UIgqJEtcIQXPNBQ3R+wD5yZjaF6C1rqqS1k1OVUNRqSjFcmXe0su3AOpY
7G3VYAn0yV1eaU4TJoRx0zHXO+4wr+tCGfG3l57Zm1eCSlzVQHUORyWGXSk/DW46k4C6mpZTKwA6
y1+whfWNntjWzNnz0izH4IaQmXGKB4i7SQQlebIXcsoJvCYZqu/8QP3B2ANHgzWXtOUOLQHKEpbk
CZREs2wP/fdagyfTCHmPmLSCAqrGbJLdT/BMPFKpQRh3uO83vEAfslysl9LbijdowgRfbfyyrw8f
42J6zWXio7jgWXZ9634fctGKQY/cn81JqJWxWZ7RxLAtkLl4ZTX1whkHylf/C4mrL6FlLgtT8kfR
W+GK3j5AqeICuylni8dhLUvdn5+60HxJPvW9h38k2f8SAOnMSjjp2q6abdApW3dIgKcKgwU04baA
iHkshMZd/AxG6Tal7G0D6Lqx50ve4SFKG8G10aAVKyWmDEi/rj9PxeIiuGqM9fL9GCN5uq2bWScb
GJ+nHtmMwLgQLaefn3wPQdJJi5x2XtZfTrs8S56Ykp9AwaG6VlbDEPAjD0P2wPUuC8OmKp4BrI4f
Xf1g/Snf4ukC3NG3KhpDmlYMuP21HcnPySvu0F1TeUqrLNPSiZmBL9dsuQz8sxis1Q3oHnZh8FcG
qThFw45B2mANyrIQBnDJHvMQpMl4mRJF6380kHvJQx0IkUX8As8f1w8AYZ3VgCTODWtKd7aQN1bl
fLBf8xov36spdFp5v3RDzhdFqKi/iUwwS1HBPsxz9oA5z+1xlaUq4TIgAg71J4c+7rdfPRI/mCqt
KKG+Zupi36DW99v2fsDMpvlt/xjtGVo2d0HZMaY2Z6+ZQyM2AE0/zk4v+8X4s4PEdrO1qGlidLNo
J1nSeae3o/D7PqnSNMPuW50K/sNOJmLtMHGKIM9sLz5GbTMJfOCox8sfwud6VXoirvBa2/zma7kp
f4/osR2jZyrQIh1on7xysFbqv2sdGaz7XYWEiSjZCTdKT+oqHKQLM8yBfZX7jfffGkIhTJHajgLg
t0ro8fViMCRGn91fQPmIuoTNKYAcTTDSV8VAckYFLCn8ggd3zd/OZKKcG2tMR4qYmyIHPeqjvsqi
nS0a6mFR1eZLj9dpjzVIBOU+cji4Tocb2/mIR0m1VJQrtuXTru7JafbZcKGoQZiljG0scX+gOl6T
1HAIIH/5aV/k+IBa677lOSQkINjoUhAfexNuY3BQxiM/8mjr3lKHJYEMFsDvs0PoF+/4elz4JQMp
3/XZrFGQBLbnz5wp48xZCboPY3+PwdWkx6TCKGtUSgoctN9Yijd4R2bBUpXZty+sHgzIMjYIte6U
0YIgJcXcdMcQr94SrL5L7HukrZHvpaQfJlXSiG5fRMFqApGLqsLAkU4dtzdnYmBymYDQUTzfs+Ev
vXEEoL2CTx2ODcxzAePnTPVbIw8iqFeM/RPzCO1r+pwI5hgSzi0k6CbR19B922cfRBHuO+NF5fI+
VEnAN8pEgRfNH4oEE9gH8uVV8hpr9lHhO1XNqj88rJ6vDtcxV5M5JGT+p56F4nsHjj6lIGVAR8sX
d0Ul6mYdfNSKA8KfaOSs/st6SSXNc+7Ss2mjPzN7qwu8dpcCqrokanM8lvS3FteaNL5plahC4SPx
Gwi7V92bexjFi68YVa8i645RIdKIAUKm1qzU8YtHcfr/1Io9FDhQe8Iphv6Fv8AZJPdPU6ca8B/e
FD/IcNoAOzJLCOoBQXdDKPEGZohpxUqJy9ngWEgu0Ds4gLaRBtVS4FxsDOxTN/aV12MNQHm3LnxC
50ctgKdcVSmcVThC94xI1ZePXm6hObDEJ5vM/Md/W3xKJaSpSgE57+Tu1e0CD/LocDbFL+2+kTKl
Tn1eKSH0zg0U4vzpoMhpsZOJ/6Tlpo/nYpjq2X670lJT/yf6TFqNAAIJBkJ7eLPw36UlUV7fgc7e
vOKjk9ZOZPY9QRTuI0uqxPW2hHyymtcTCQjiQViPFu4WZRIlhnpPyEKmydR1v6D1ex8MRkTsu1b9
rc61VCm5S9VXvXHnGivC3Vg7jg+7zlcZChvIJ5FZdJQPJy53Kf9emTL8NWpF/R2dv4BRFQ19NSbQ
tAVqkqs1wVUMnAlxLZWTc+jiP02oaIzIzclYzChA6dG8Es+4tPs15hSVYZ2Z5LxjThT3jVhPp+6e
ybEDhwByGhDh9GLH7EBS8CicxFt87JJgml/TF0Jj3DHZfHd4KihV21HodibnO5Ly7tgMU1sxYaIA
bzzZle9ubSmnrvlsvrEQRWNVc0ye34OC1edsuH3K1ZHec42wwupw5C3Fpp3XP1UdNStgxuzMwTDs
SkLTga6yb/lqjOQTxEAfj4A+uj1ei1DiAFoYAEw/pRJmJMYsynX3YFASbIGiCr5kFnR3/VneLRNF
QJF78bAceLaDz5RwG3RLXIkwzRcrbtbiFQYNlM65XhW8fu8cbA/l3/9miI+imADehDLRpTWRa5Nz
gAOqRkJH41IZhMafJ/S7AZuN9h+tNx+4Uj+etcy77/o3Kn9uGaHShkhtn9nAtKsGG98QniRBgB+j
HsMrhHANazPflGTTnk6yoUDjyi9PLYYg2YpdlmzbKbBJAbnpewfiKjEk6p3kLsoYo90z0aFNiZ5j
N+P623cut3ERcF20doTFwvrubSLyBuzou6gj7tsFDsaw3OFFg6jTN6NdOJvi5Fxvvfb+53ZwYlqC
Xa+oKbgZXCsF1XKSIKk17heS/TwOOk/VNCA+x2AlFc1pT/CkZWSOlg1mM0vHfV9pSzdWJlA8CtFX
OwK00YEPGHPNHkigfMuzD79/etEaphJj1DIy64uJDa2lJk5+Mldin0HBi9GmXAa6KnNywyYkMRcH
cjkRJZ6x+k70ejUZQF42viwZkVdgfli/nQSTclbMn7QlOivPeK5O9l+aLtKpgpzYiNgnaMXoRs1Y
0yypMxjtcMoQuIzTdlPTShQG9S+U1CIMzdV4YvvWRrv2kAoEq2H7R7Sy7INwMHQS8G85HfHrhEKo
bkIb7iq+4497f+wILZEIVdQUsiHBaZuWusbnUFZbtC9Nt+J2I7EqurpE3o5xvgoS5+FW01scsWkq
CwrLkQzQu4/znxDXvub/ZtEFRLbDwNmR64XHpqq5U01I/XL1kuGCRzp9cG/1lhMqAADFfxZ31WrN
+iLYtPZcIOeZdM48uatpfGHNkVIIdy/L2uZ3C3INCbQ2DUZaIxMnyk7Q4f+44oa/kyM4i7BefIfo
mwUOqdGm6FmE1tH3Sg5X4Z2oCPFDebq1X2KFwH0mKRF3Vi6i56WbwcyRskDq6kQs/M69XWbgiVaF
0fczfsYJxdxO0FFnqoj2ZHoYMmYVwLOIBvDWKI5S8z1q8jjGJ/8D6Nn3FqbfqNJFZyrRkQHUU1ru
X9CbjZHlNaoXYzBie27RUqtcqKGzo+aIbUY9c8RSahzSNdWMZ6X1wvBfnuS375GMgdKfMHIvBQv+
YwcGxh//hgAfC1JLTl49BVG1j9Bi9VVHmhyDznYg+xVeoPH79VqJU9DpBKr3klYkQXMEgUuB/AE1
DHKJsqRF6L5SbI10jfzquFLnBqLuMm66fPZFKlkBuPIxJVNq5iVSWIOICXpSpeLT+rAnXeprZ/gr
/CjrRIP35mEDBIzjtYSeIu/H0gH+wjW2LNhbI5IwuJDMhtKGj8PDl0df7QhLfy28UULs8wiat4Ph
KG73aNaJpidNK3E9AtNvrlHo+kgYpMRbVSpcOe5P3MnZHCrGja1YFKIezhBR003Umg+EkMwHc/Aj
My5MF1w25DJHF1hGSb3qUe6MHG4nzZvKwq/FCP1LDrEwfF06qhSw40DLMEMxdXCYJqceBrv4nLRP
MIPtCEmNy1GqfwRQh3+4fhtud1NlfNgNbvg5AiSussSdIgjUpdOP0iexNPTib+WifBbX13T49Xj7
gA+Id1HWSEFmHD3NTo1pnkZ0rRA2whfM0elRTydzTQT/xHBOCHtLFUD6XU/FWDIP90l631WF07xV
2CVe7WnbkATdfIcnq2VOIsgKiQeZEhOcgXBbDr+sXlVY8T4+vds/CEb1aVxL0wJObZWIpp0kpmTd
AsYtYEPVpeDuKy97pwwaTzBMJvpVIkRGOV8Up9/CoCRkr2yeZDrC8UkQOrL0zhxKa+kkBZnAvPLW
DKCduybJva3ElTHT1rqjoHlszN8U2GB0xLTNp0dIipN0nv6Y+ItCCPths7CCRFvR0oD0HnEK25wm
Tt1Q03rC7ofMXfrlc6W18vteTdfEHOZqV1MLnCP6baQ8Oy8kiQVpYSFi79xqy72uyeQadOHK0/Fd
3T4Nb8E0Vhwq/ex6qioY1y//j5BJgqOfhDxRBp3lOh2S5xIJxCYzgqDUJH1kctdTob4fRCWxG2Wc
ZRhlxQDrmlvw0oF1w63QILhDqq0S/Q6NYlzhRz9iZroZd8tIGybpa9l/Dl3SFKOHJJobmLF9BUEn
r6UJZ1UM37+aVNcFA6NW7ez2Kd+HE4aZktPZ+ww+jM8XT8498Z8DMly8Madr9MEzj8Njow1SOon9
S77s2tsWfTTXT73EsAW8UzezgouN1neiMpk17/juj92m90wlG0L50Dl5OFE8yoMaYVH+L0dDrtma
pYfkZN0XpyTSw/gMwInDgpoAew4F3nWAFDrmzvfoSN19boV2a3dDXeirdob9uasGBuaJj0MO9wSz
doNbiTuUTUWFDKPxeqssd0pq18pjl51uSosGhuYKcF/OhDLRi+GwWKYtGLYxZL5bRYjesDTpj8J7
75PZ0V0qtatim1ezgPBKisDggcYJMGYdwwcOc97aIjG1KZ5ImsHz/t4iDLtDWBPjoVvq2xgqxBtU
T/+qw3DXDuHu0E1j+gNBWNd8JpT4mEztQe9m+RcMshZHhxalsDOfQ6SC1cS48ZlgHl7uNbkJmO+9
/tFx9O26tlXM/ghOizPGn5L4xr+zdUELkHSb+AvPZnzxr0k0o7FUuVSXgpRotXWAxCCpJomEglYb
0VoxNI4t8ZjS7F4FIi7dcl/8qH7+TXs2S0I/QqtzxY36W3Irem3fCTaZP67PM2ZYQbYd4wk0QUmj
E4FJs6FN8x7SaCUJqBbhsS0MfJ4pR0iiHnCfMSCwEqidqyyHw6aTNmGRRcgqrtrhuZLQxoVdf9Vh
zJ9aIAgUCXDFFRkTIcVQYUWk1CAEVkbRvTU89UDTgYPk62dkGQU5MjTZR1FqDB5RBvNsVcpPb9m4
SPuH+Ssfyu3IbNT8CG0CdXYtxUpB/MYRZW4nMmFAFNrKWSKGo+eR1TsA0Fj/Vt4dkYoRMwvBl09G
IC8Cs2uzWvbpXPvF5IIquu6QxkrTN5kWtBfMQvfeE4fgII7kf7Nx5Ru43fcoRlRBdy7AwcG/yg4s
MVCmbjh21K8/FjolgDg+q621EBK/Bgx4Lkn3AB3BE/chHOCQkkoF9PZQ8XsTE7UjDHZ6VLQEw/17
rPsiDeM+nBf0/uk54M60puq9/SV8D1hAqkGW+ABNGThbg8BlagBQekNKxIoxfYotL+ItC9xM959y
EUv9su/C4srRnDdK3yc5XGsKZhGEJPkPbrynYxkm6ahSQfym/kbExbpFJZ/kX2uf4PUFvatGJlMS
Gtjqot4kUvLrgz3SKDMLI7rnSTf+6fi66orDdT16qc29FqHzstE3sfEU0u6YI0TOhiaaz1d6C/4U
t1li9FVGSkAKyW1QyznND+GGzyQbBQXwPK74cAsRfmRqLGzze/XSHG2H6y6ulM0Jg8NGI8f/F+2H
lXDMmiSeiIqM6bIXm+E+7JTV0YwmOMAmYk+hF+tImTC42nGJue3WpyYL52fnMmGs01QiU2zU4vSW
zfY6ay3t7KujKrK4iXZ9cohhZnmyPEWF9HPCh/fB/0dFHeMi7uHt84uSLuTeP/gG/ehyFvDuncho
Ry2iPeUJypZ4UaMU/ooc+Ylib98hV1O19mq4av1hynvv2/dLrZm/xvb6q7HUN+kanFQjDdB1nu35
axrYRzH032jbR5KmXr/AIfHpqtt4d9iedHqwABIHSbOLoqoHaqGt0SKXfpbAUH/HoWoUkLzTsVCn
xUIYvHfewjgQrgaTh+aOotS4qCIHtiU83ByIi4evWaGN3pqeNwugkuiefYwLeRC52/oLHLG+H2UL
baaNo/zTHyVRVj3BRwKLTXD8gUEGsSOOg///8g628YBYqsV2l0+HdANphjfNkSkeh7PYo+0LZPRn
rYTSLuWTlK4Bi0XzHdUR2JavXAXIdIInUMNmG0FhNjMBGrhTx+qJmc3WdwaS2hrfnGVcqWYZ4icx
og6DqpdrQZRocCT+tgLoq4X0uWVfpAfYpddH/+LN0iLwScIbLYdO7qWRBRZ4u7xZI46dCQt1wULp
Eect84vyMrBCGUWH1WmmeZlrsbl/PxCXja9D8BViHRaEV0o1SOrDNJIUnIq+K7fCJ9U7o7tlfpb9
zZUhUQyiW/5oWn8qfmEP7NwMfcp/Z7QVyDuXnvHI3V+KbRZb081YA2BOKA89MdhjdSSUsRli3J8M
YcUlqsNwGOuyroaos62IaFLC+xV31TY/JUB4HIlfoaEd0lEjmcIPZS91yhRwJ50fvBZewwn29i7T
UNBZRZI4NKYeZqQ2H0G+baijnSKEBiHGO6PQfLEkUIfHZoOslb21wp7oSLjJMHnW18gi2oSpzZp5
sQVRm52CKhSUvQpxa8/3wlPwNIodosMFGqvMPk7UQjiLNAXFiXCCafCtjt9R3s864i/VtH1XBa4K
A8gpYLJ1H78u6ChP/Qd5QFsi/brvF6ZgCHCticPXmcMntUCF4xYEZd7yfcN4K6+xZ8I5QErRW37Y
NclnXkikoGoQPge8UHTyj/UubrzkleuIQ67tp4lnH356qI/dSvOTBuuWoiDZBk2tG+XNyxisGO70
+OICf/9sYs6FnJfJLV9n8o07d5y4TltPmdMuFhysIeHU//N4FXu4AcVEs891FTg917JZjpkfPYDw
i0ZmxZ4lRLn8HdKJu/8d31Zy0ALuOIQ/dOLcRllnO110fFi1/1Wc4Aup4MGByyVW/pDTl1o3tpzm
Xm6AC9YnsnxrLRiaxJ5sVVEIROJ4l6pHh7aoUWlhJjnqwtcktpMznyYqwv0UH+kzBpMuW/KuDIQa
98ztHmF/5nboFbrigS4/h8beos/64v5mg7P0a/A6yd694RKQrtu5tOPw75V2Sw65HEToLDrWaFw+
OOBxiLIWHANZmOOUBjUpBNoJSTTCqJ6cLR3uAY6MWvrYCo2tEFO4Ad1M5/l4TZLiZZeYnCDS44n8
98blVAlpd+QENFSraEDlvkAQm7GJ0BLIwJW2wY0FbkT1mDmuwjNC8kfl/+u71BsE8n4C4Qfz1+B8
YuOGhFxSRpuakXliX9bZWLi5CYUQVpg8kGVOTRvJsKeZkXygFnM+Kkqaj4mABOR/NOmViD2KmuIf
8bl6MtyxIKBpLgihwLbYPdakzbdx3SJQweEZVsXw9B/tMlTASIf+a8lq623P4fO/HyuvZxjURHpX
CkOrWfrJiJILBmyszHK8SIh/GYVqrwu9ZWtHUX+FV9ZuJY2kyups70VT8t0Ns+H2ZcrtJpj0n2lj
hDHXuE0/8dCUaDhs/veXOcpkx+1L7rOfgorw+qlFajBzABxsLNs9EwTf1GmL3FfTeJTPO/KY+95X
9XfsxJv8V7A7Py9GW3yu3mcBy1KGIXdzXvLZHHHpeI6WACl73gzygugdfkoaH29PIwefgS3EqzAS
hs+P1hBZDZxcD6jZZa+ahN3AmsQ82t1LTcLYOvjQJEU2K9S/T0nzoJCZ2kowzEFjeC7ZQuVlRlx2
DdyroDU/nQZfOfuJuTMk7Ilr2sZ2bK9H6FRJcrHJkUasE47X7V13zQpiTX4IHyMQoIycZHhbieVt
R2Cpqauy+S/b8RmsTL1zy7kaWZONp6xxaY9dMPQp60hEXqXyu+Zs6/PiTKJnBF9RaAYvRugrleRR
HlDL+n3QKiPXYvX2NJatQ9/7np2Nn6u9UTFk2CfpgDAGl3mMXOse9NNnQF+kfvYyti0y7NYj075G
urQusTH17qB6YnXucBaAo3N7pJwyKnCu6js8M6UWE23mNZ0AjoA4MWOGNsvVGLIsdw9ie7CpmM99
qBRWnjM2cs7O5XrVhsQy/WWSygCEsSoyIk4X2zSyBQuViIsC5UJhQun4gvFEmEdJqTh5y+gSW73s
fSm3TXz/LayAWBGj/K6XFnwQJL+1dphQmspjqd8MNWJhu/ZtLIv5lMb1OQSyjSDbPbcKz0f1QRLo
laujF5kMtPnZQ6KDWuL4PWPnPQ7WC8qd9uGsZnDSlT8roQJ+xJ2mQ9H3uot2Qq/JWuEqnccER3Wr
8QIAlTeVDRcghDozsalE4cFNi5jfN8rbNbRpEojHJF0TY7Djmw2beickzpx0C9nJP8j433zFq+ie
TVcYUWdgSL2IfMRQLWbh4isTmEUACDKn17PROg+yU75awurCOtHkD3J709FtYhmYk4RJTPVTyRtd
PunjkLi6203pQtrxQ/hDMV+Far53HK2vYWV0NHGDGteSGn1FyQo9f5EPm+JuPbKKhr9+SJ7ljjHT
xPbMWmvjVOQn9tZHz7hwpnLWiGy43zsRjUlX8AmsBTBezNGW8JvskUlHsi8kUyFo0lYd99rpFJf2
4SR+OLO63oihsL8hSPV+PX1+U4lFkU+CjMNSNp8zKBDFNsn2ZjefYpWNin3mOjujr434duFwXxSe
qPKKrm49nSTRbsZmOw6XN9mJne36J00DNpeM8JtaO++FI0rl1ChDqZbOCHP+jDyVV7LIYixrpsc1
J/SSSXBArWPDcszT0oekkFJNgKZYJgd7IkHPoh3Na3xavl5f0KUHXmnlCKU4jOQilVT2zJouUL4K
JCzjsL3Oz0/SQ4Dlptd7YjSe8iFRdTa2dYGWTdPV+fGWcmf9BIWofS1X3ax1bB5Kv18/F3Oz7QrM
LOqPpeW+JM1vZH21tbm4YAzlTUKI521tUH2HsCLcoh7qge20zE0isZLgeUidpoMX6ZLNxCjJ0yrV
NT14G0UMesSA7URBGNL655630+56KzeYQOyMaJ4fEaPk9CJ0KC+3XAeqcuP5jiePC7+2sB+UChvk
2AOS55zrPB5rkeia+gcYfJnZro+a50G9qoySnHcDnV3W9HxMyME6fkalgVvq4GWoZ/irtDdxHk+6
K1seaAucJYQ/b6vGskT36tQZXVD3rnSgOh6t2nuS5yOz7mUOVfaQL5sQAzbqPSLrRVLBvJuwdpj7
bYNhsbh6g2taFlnwtDAOtoMBnjwJQ4gTftSLTgX2q92//nu7ZPtqjI8vNwEOREzUvOM9oK2iEcXo
MCmHkUfXI3smSktAWGnICCfIu4ZColIWe9SXCQVMiMNb63oxs3mf4KawQbiJeU3ybaA5Jc587LHc
7SAn4RVXnra98JXI9caGMpYeJYYF9BJvUOR/Fx89JP3Paj++UdyGfmajUxyAwD6dEY0ybY2OufYM
BNnauUPeQNM8Ax3/mSGSRXp2tsqLwZW5bEbLrZSEcrQU66peRDDTqNsVzi0sGoHkyLqbMaLSyKEk
MabmV9jnDsgE8gJLcn2BZipjIA/OoRogKRpVYydETXjN9JhfMBXV85gLZ6rvbMyrmJFOugKILfB+
SV56kM7oe/u4f898s3iKb451gUm7sNjv9DEGEjguIvSiXrKb1XLnpwKdxHIe9S2hMn5Xkrfmjsme
Lkqp0MTOexx1GKSoJKFIzyscKSRXD9Z8iLFDHU7KFExaWmI5ZJxtXE81ZoE0Inq/dU2cCyRHBy8i
8tXOXXwGVf9Z67I73KQUAsNVBPdfUeN35KnA98fhHAcqXh6rnrSz/b+a7st8Jn/LJkf8EoVPfpyN
UU6DOdxMDO8At7q0CSRx/9GRLmrUWQQCpsBjTMTPy7pXG5qyM8tRfZ79egKc8Hg2XU0nDF1Bt/HB
5RyvJisR2E9CpelpFaKAIgEySevdMaN/QO7qj4kIOQ64uQwd4W4OsihW3zD90ztDGKUCcWJnQBqe
QUi1j7cteVgGTLeomzD7oCa7VzWftMJ3t6RvzI2HYEYEsYA2//SIqvyjEz6FLih9wW/qA5/W1rNj
Pr/4xkksUvpIe4EpV5B+lEVjHlqAFVXoXxZJx7xz4TNDRC5VczICUrrAVX4gHN37K9p4x9uvCCOm
Q6eK7IJv6mHqGRAd3y9ir96aSQoPfDtbHS5pdRUD3U/IbHDvOtYkfv1DsrnaQ4ZtAPSw4NsudA1O
UQFM7G2dSY1dNXlCthQHvgOhsyEbNvH0+AJ10fYya3GyFwlxeDePzAFPV1du7+WcGUuGfhTJZ9JR
HgpwGhPsKcqvSfz5IqVbJ8sL8oMZ0VPN75je34iE6GEO+9DAGTS3LHHJn4IDubXfRShBZWj1lmlU
YZ2qS+AHz79ALah2e6fMBj5vFgkzOxBAp2XvaWTFo+9ZmUXmNdMmkzAQ/ViK829RUqgLzqPLFKJk
6bPjp8OJGwlZiw3NdX1pF2WXg9cAdtZ2tluUwKLtZ1b3geCjmnuOgvVo0rRXJGlIUOFbspOFT+LR
UlHKufL7wz4wMifd5MB86MH0n8XR9S/TNGwi7aLmTOLfyGeyRVjWu8CXg0xYhI88p3hsoiGr+xE2
80IN/46I8AeWauM01KodQtWWna7fNa3vHqHagBH5vBEIzj1epJY3W5eiLuNCueFMpJ0ybPIv3LpR
iGCfaOFYKzVTxC7WhDiSLkTIDxDgSq87Ya7abZo+1zJ30xnEKb2F09aZXcT5OJpNkETk1rsC1/uk
SxUDuf8ZKkE54XFESRF1kzqvFINLJyQAGBCbd4D8o+BlNbFTppYcWNj1c3A+G6xCPcdmyr8aLEpP
LDX1b1iNJIBWWOKv1OyvEi5s0op6HnnZxsfjOmyXES/pN2f/cFq0rJhoMOJF4NRTe5h7exgIJhq5
EY12jUWtcanMBo+BTES+wxoVXSpWoG6p/2lUF3vi08j0HLZ9U8UI4hjVaVS46Amcxcco3QQpLP5X
uEYpDiLeib6UzOjx6PqmvBr0XusQz2VXvLUV6U4/qaKR7EFM+xIOQax0dQVJgVtn63V8aNeVCpbo
lhfXo75kmNQ7YfMRyonUGhdY6Fm+JfH3A3a5b8B7Vv2dNMiLQ6kqW8TDWH9EBQQ7+9DhRbVZpdgT
LW0fd4G/SC01YiNgw5yuylHJYorpY0r/e+cxWE9GLA60XU2gXBTWo2p0LuWeK4tjsxfuO1WlzAnm
6+ERh7dYxRVDAY9dOkqQh6v3wsWn14XgS/cW+v4AdIWKGR38/jMLpgMTHKoq/fD1F58iifX6CmsT
fdqOW42au+CtZajH3GQPwuGNCrNw6vXJa8SazFAWdSgq+yVs1uDhV9+6WvORBj5bn+SZXRJ4FTsm
fUC08wR6yI+ifq3ULsp/SHyH17D5AMEcWrCsL31EdawQuShVzWCmNub1AA2ic8jj+OYZWvQWuR9O
DgDNy/c/DUeatkwsJgp9Qv9r1OGh0FIk/chNQ3qWbcJ1+rqwiEroO8rr69fs+/FuZ8qm/6m0VLQm
yjtlu5K2FnjPimBgHpvlNDjQP1BuJBfvprpy+XRRTNtv5H4IKTovh7EJphs8SigGhnobz8JNiwhw
P5iO7UtZBFmEIdJ+Jtz7++favex/EBUwXT77B1OlepFg9m6nbHtbuU2ZVLYuwMD0EeTaw5h9SjC5
Y8AxI2o1NKVatIZTfGxn08ZGmC90SP26FEAe+5PaKiE2nIw3NZO0lYzUgSNlgzvprNLnBRSomJu+
mOeyJsTDBr1p1HQPO4HmN91ncpyDkBFXEwk+n8cCD+ius5O8VEerQ8bziWf8+EbUiTyECxSNDTBR
NKAkHjQu41iyTLFt//GF7FvqCTcEErGdW+Jeh+0UBZcpRiPXvcxvtAkeQOSGtdJonPaOg2/PmfOJ
PsKwaqeXsW/XpH04aBzIaNq7jGr2plvvjsmS3qp7OPL+SGDVsD+Mw5gW2qJHW02AybjG6tHAFwZP
royAqB9Qe5lHYRa1cHmlsGGY1IPuBTFwwa81Cl5Nby7DBoPjrYygZKKZQVbZQVHVFgcoj4LpYse9
9cXuTBJYMDOGlC6UV2j8+YoO8L0NA0v+FH5C3iSV8E7sahnLQtznZWA9SpK4nwqzg9SzAcB3Dad+
MowuPydcDLWyCg8dQ5dxU+bcvvAiv/4SrCgrDtZ9RCw8y0+fTxi6t+0fixDXXcwwMJdWMofDXZ1l
3YRxv3t7ojvjNL1zHUsNEMT/sT00441r3AFGef5FQeODDcrhIynrzQtbAA+Qj13mRMCAW96Uos+E
v46lj/ZDsTAJTG7Eu/jr/JLb0438Bbalr2YRuZgdgSlUkshglCpuTPp73Y32zX/vz1m6Nhyc/e5s
kEi5vCasAUgcdMMSqUXjz20JD/OWN21WVaQhw+70GRqnENW4zNdXBjmWdHcYYrD+glJmdFPbqSkM
nfw9MzXHVyKD+Edd0NVTK2AY48x2LdO2p+NBWXvoKweLLdVu3dVs0DtLN13OU/aViWrCatxXyJbZ
em7rYva7BTRaTifIUKwtXozi7jH6C1/XyBe8hQS4XB41NesYgpp8mYcPVLLZ1GBZzwpXlgQpz13K
dFjzdOfEQMQYp9jSqajEly7gKJIu3Se5J2Y3IUcwlxzjY4th66yMMymilCs7dR2h67WiuX9jHBWt
u4S80zDmeSBGnCPQvdXBCbQCsZm4TkOziLEayd/gfzFss7EMn7TxV3pkYAhYPqxW5Z8NeV+Agyud
HFLSwewuV0u4KZfZwzfqF8bYY5LGYI9oa549EX8O00UlPcaTQlha8KKkUagUCugCon1X9Jw2cnFt
aXmSKE+ohnQxTtiJX9q4ge2ZdekFGB4t8AEuo6+HDZGqyw5O+X0DCaoAWRBALO9QwiycD/83LSm4
yKJPDK5QMIUdfhncTWd4bf1KmNRNKOq/WIh7yHBdXpjf/TC34dLdiDSQse7IFOXFI2ZMfOetI28J
Z5O3V9VCZ2ubcRrtpQbapG6t0cYkgzuh7tvnWYuJ6ah3fefVV13qhuim8tqCszOX8nydQ+CTjxeK
EM769BJ5bWcMvx0S95bwvg1fEyHHU5OLsJgNaKxnSDRnVHIoX8v2ZJviA6cQ6xYhZuH7iK3ILeBW
mTbECxEcrqfqGwKW40SqpstF5f4XDIdQbaf1tqigHrVUwmHTtCuJinucos2HYBnZRBnCmshWl2Oj
iBIYysNlYPtq/4Ouf0UAAVrOZjbodYHxUTFo3moFEbZ1dS6rHjN5ncDL0N+Zj5VKUM5RbU9wdppD
BT2QtCEJCFoHxULZzy6uzLlorqg7MSJ9/c4LDZ7xA/N4eZKH045s/xhRB41OXotHZInrxJfjTII3
NyH6A0yLKX5pZ1fL+NsFrzkwVRSsrzYCx2SE1ESkAnaA4ZoLRTic8/PCMCcWXF+q0W9mcNymDlD1
LV6JDz8cfz/v7LaJgAgcDRwaWS3QW2fLqBwwBOeGdio6ZInAbVPhg9cHJmGektDzKoONPPbeghmy
SSg/bbFrT96yktoKpcfPjs7b71Ssdr/SLU9HNzsuxO+/Lg3PjZNqDjRqFKX4269lyugytedp26iA
KBB7LKjGwMA/o92sqw3lthOJlKDeKI9AbM1xiGU3rsdp+QvLPtYVIH0CAfQvLmawj5BHclZ2l6sG
ZAS9iXAss0qF3/s6Ga31XiRlAhlPij6iGyGBjU1tydtqaVQY+v3BxbdYZICTCUokdCvzTYIXztDM
WDn9GXNfMUZItpEo1QvL/y9q9W2Mc7eyQGOKkg07k9vfAGcz4kWZkC8GEUwGRI3gxU7PLarWtLCV
HRaTIIFtlSNzYy1KKb8qgz42spAPFwenpZ5A1exdhGRiyeJ4hUS7WpVLarx2odRfv1eWUJKtvolN
CPB/4+9iDyImHUoJzZHTKvcT7WDZmWj+GapETSC6u0EwW3B44eixrQBzvMVsFxE8cKMQ7ywXkNRc
l88luTLYFTJpQyWUu879iiOiAmIirf8ECsu34rfRf6xfa56J7XJ0Xk1ZWG4i9VhKjnSOrqiicTls
KdCfe7SYyWJoBxCDD/No5sTowQ95PF6dXg8ezUOYUnzLL2G+Sryb3yHibdxDh0gQ9HBdPyy9Nwxw
4mLtBzGOT8DodMJmuKOaE4JbOwh20KYhfXZva4BNFkYjZFQyA2GZsXs1O0ZF68yvT3T6HVK8nFuk
nXbsByEfteUxFvgz6E4qBKTTwYOKQnZoa9gKtnYZ6bxbsk8+CqJmmvLgDLQKlbxhWBlBqUgxIxjA
6dqs71BGXCgWEEjt3GdXAnr44osxrxVC4+517tYFxaKPJ6eAhbStCCsCW/SPohrKoA4gSArhIUtQ
SFPhMqbHyQXbJDJ3UtfgP/hY0QT9dAb9WjDy0PeVujWFQ9woAjSVpGX/NrLwg/gWaeupJbYwVE/I
w5fGJRRx0zL8oZ5zc2NVsgwBiKcuW1MQqpbey2kUtH4nt3laVMr+bk6F0IwQOVVQzogCZHvJPDWn
Z9iTAmh9o/0lEFNGjKEqFx+qgDGU+cNQLAyFXrTHbxns+30FLh15Ifg+yaxZIc1weZWh5NFLn7sM
/0/bztqSnSh8AIC+/0WjLJK19KQcmJ93VPZlHpIgkTOyxmgGsLxP28feNT9iR3/X2E0+5FzxHR+s
2wpOKvqik//JEm/RbX8CPoUElDPZwblPbF8GTQzGDpX7t55Ku7otAZ6B4jC4Fss7pXVydCOkovaS
jiN1iP/i1cSTosqDnw+HOFtVfs7FgP9l3Ax9BiFb0QhvASqnacpJblN40JTivTCchieQRYCdpnoL
+8LTV2DquXhYoCtIOhY0D3NLYS3M3ZLtSSyqxi51zYx1FF/By0IuBt/KOE+skpiRP6BhRWF74KBB
nYkZPtL1TDd9yxJTgeoUf12Wex+qjpheovTYnaO6w6KtX0gycsMvpewuh9iXK2PfjyshAvwbokM1
prdgixJmbTJVgIePMw0JVog2BD75iraGBo4K1iEmXmOvftu3tHFWUx5p3D90U6mqBIdXO4vVKKDZ
ws8IcEqFKbX+/LiulPh7UkcBN5wePkUCSYwsXPZ5uh/8epLPE4feltAQmNAVIIanPbQwGEON/jZ0
ytyWDv7ztEpxriX3CQm1hYcadQ4qrszAYhu/u37qH0WfCaEqU+MZAjd36A9gLtf1HYl9GI4TJvPH
8wMyGXW3gji+eDIEVNn+nWHMnKRQms9t0eVxsZPI10kv5fvOkoKUXObwFe94Opwi1G/jH1cUcaS0
deG3ExSYNwAqLCYhsNuSY2kWU4cE9xKqAesfWtt99J95QW94IqNDyD+0XwV/mfmt+4Z7pvVO0YXy
yz19D1mc5RI5brt/exNco+guy8J1MkJ9Br49GO9JqkdKroYJmISqZxMZoTQOzY2aYyqihLBnwTcX
hRTA5lo4HOLSmZpuPDbmGpEjuJpobmcoWVwxc9p6dFTcSdw3umPldP4kPbYUuJ43vyjv1EKeC78B
K308s0leQNTqpzv1o1cOfH0TmsfABm8bh5LSd+9Z24OX/Tu4oVlmAYA/Kt4QhhWLKrWT5suJr8my
8AlFto6KkpleUoZmYiSa1yzdUlLlSMKOvjCdy8mzL8COsvlTQxLEWwkGBFxaN1GuYMYAdXj2NO4l
flDFTvh7dhCvSMWNAYRyGBTNjwbj1rcbT6RdK6Y9wxFikoYHZ9boDyvkQBQD6VCDGU/IpUe3lnVX
M8mPeZx895HMj5sSfvXwM8QPtXqYzIG2xtIc/P6mm0T7Vxp8PaUtEOgzLuFb+vIXdJVR1KWZvqWV
fZiMjDb1JtgiUl7emPEswvi1oRfnDhha+/MsKOYjDa9FUhcFkodgxPMh3ttMZEnQXXy7obNw2WKP
F29RO3uCuB+mZav64Z0y7lKvGIbLDpqCgNJPq7br1N/Geexczq/bdWBmQ0W3DRWoDh+0jbKfcxIb
xHyfpr2zu+E45LAwIoTCBVpX//ey9Dm04Y40eYv8Tv+3xaYf1z1BKhB6xL2uK7A2WOc/0sJZQEVy
h6IfkFWgbO36cdmoDt0Cy9Hqhf7CDcoXHpKh8j1y1RjFVU5xOaqfDoxzRjhenRopFPKIPQAD+B1V
eCPWXufmsK4QXOU11xB6BkKW7zCpyJN8ZoBXhxIx1rl+4K9OtkBzEvYQKetaTjJYJN8FtPINMlBI
GZ5jRNZgG0nBvtcnRTF9hoVk/PhtbfBOhcKp24qvWa8FyHGp2h6pVVBJtyEhGCQOk41kLEhm4GiX
dtirfNF4IwuSWcPix6jw3Vx5Q1DoUXnWta1sBbve/jOhppBVGwKKxXYxdcHdJb+k6FJqcTtxVKkV
KGcxW5jk7XXTmfNvV1Fy2xryo1dxQaOJdRVymCZJDJArj6wO3xmp7zMi3KL/EoYbOC1JTszONPtV
NWrdnU7InWGpd1FHli8RYvxkAOpCr5uUih0Ic0boKTPj0+6+staykvxQ7jvlIIQlh93FcDw+LVkX
t/DBOFB6wKklaOR7OGPqj+/X+wVr/8rGZpaSZMxXS8TPR+DggPht2E83seDHXcLkMX3jgFo0FEr3
Ct1bSUqvK38KAe7oFwlnJKVuqVlpP7b6VAiuR5rz9KWmClc+7AlCJUPgGiDeLy+vBnUulbPBGIAk
ttLJYnanZ5TRBX9cfFhKanXj6oGIhIVhnRQZEYdw9drB9FnDsKxh6E7L9UCXKDfV868sVT5bBpAb
wjMrzJCS4fwk0xi3f9q6eRo5grHIF30Zkf6/1265gkwBIUn3nY6PvkocmepTAq0PEV6QaFcc254E
UxO4MFn9aESYe0HunL7/IzgkqvsWXL+LGrcwQI+LkXFzUvQmrK6HIZSgOI5CiHp8+YaQlR81xTf+
IPjoWY86Dw2LdthqEHjOMElZB547k8h4Q0aLWzFXYt//NuvX+qC2q+2UJg4VWkDgBzBYcwXFiCHO
MFv2loRuUStdM3qwnbM5to4cVjQ5fXcVYwZUxZM0DiTKlPUISUZrsFVXbD1VjVL13vaWgyxVhOlM
Kv4Ee8f4JuYNWVmDoTo/PYsm1QYPkVS9JHC2QrvzJOBxsNzyldUUvFGBnbgDEa0JWnOoskpBz0hi
UvybFh15TixulDZPmqMMVD6U28PmU55FOw0+AXkvRYznGpuaNhcGQQtuvzi/HUF42Q6Jq2VYfGRT
qT77ljyt+K/ND8s7DnXpos5jSlGOKc8Jt9UHutBXWhSAN4S45H0L2L0a6IcSIOdXVigO6S8ujGqp
KAnRqL+RE4rbEcuxB3y+AQ0g2VM+YdyQSjRqmnuHQGtdH25qnWLjxOIrpzqQzOnZOm+VlkHpa61q
JEasnUCsoiMlVhzrHxkoalp+dvj7Lmf5RXkgsjWc+MOPpX+tAKqC5sR4wcRBdniVWmmYKHlzLFgM
Kzwb9+3R/WfKysV8hhnpbjv9DPDzBJFjUKXGhkmCZRWNNpYLJ0UjsbyBpaSm8HnsNExa3gKspLx7
2fBHMjaPdGtq1AEUs2sm3k7jjR8qHVh33f/kE1cYNYpYsqC2J3wRCoaTLaGVQFzTlczo3LGyI2X4
etyjNuAFOMxb4kWsLi8LNMivdeHP0xfc5B3PmGD+ocn+BgxcdfiSYWmUfvL8DH9kzrUC3EMTPWxj
bsESKLPUZqy/0Ydr2pHAtf9vr4diD/ctIU0sqwp8nVPtQnGa+7Fswg1hSX88PQ5OigH8YmM6z0af
ida3OY0oUwxQD7stRczgP/tgcUOhDstDxbeWxAujJJfvyry4VGijTUxaImGmIAcqYSDlKo1CCk97
NdMO40ZSR2VtrSjsc1LcqTpR4qVIS4kpTcAxYcNzF2rrc76bR5eWsdLVlbDiBsONmIiCqWxy8kVY
uJnwpqQLvcmqfr9KOr7nju0FWAEgCuYHgDdjeX9FJbXO70HtVkigZ40PmPiqlL1OMYGWbg98oCPr
mF2SRkyyJwYFKC3DscwxE/PsKbThYUr+WjC//i+ZOftb52szqogTsQHIi6XObrXzEElk8WHet+ve
E9+PdjWtdv2tkapMOjxPNXGj6K4uJND8n3UnypUV0p2Qlk0MGOSor66tEuZ46Wp0/s+35rCUGcJF
HyNh2sY/V+xhH7sTKPRGHqJzIWXIjNIyAYhXPA4Hwo8BH+HpZhZ5vMpLo2YLusxeZexeYtcPITJd
6oq9LHeokpVhokckHbaYmGG1KMwojeQzAA5duRFbvTQ6vS2iY/6+ygPiNYpB3PY+JNALty4m662X
owwICB4WFYW7zgP8vtDX4tvmQM/RcOWAaop8ge/FGTK7Yffcji/htyNgzyylJxvV14AIzu1zaUzB
FcNOFHk1SYzHi2Ak27AHUX21FSRZ5B91RTyZI7eOB2qXQXkAJZvz7nB1me2YI56nh2zOYhfEZaKD
X5NInHORVK8caEQJa38ZTxDgTwcia15KwjF2Kz1cW845RtoepL1HQsLU3NEDZmeuHGkQoFA5cIqg
aPh5RH/eiEm19QW8q2rpjBS9S+qMtNxTlkjcDGPmwNv7Sr2t242kg8H01h2pm0E8c4ZTK/us0e1j
bYsVkP10wPxaI8MFJ7CEwfcfGyopegVQl4YZeBW/fnSFS7Ec+tarKYzxrD3bSA+j4tSXSLRxa4+t
XcStdG0aHEnj90w/mHNjAlFQTFjeScldyyiZ253sUQ/halpHgWWCLdeSUf8AvVJhX8DIh/IhIaj5
/UEBSQuV/MPdODiq+VpYt4ZC5pjXq0h0P4M1g+n2C4yMz7AUsgtX21X8lnp+2tGH4r3PuBNGdkHU
zuL/APdxNx8+pycJpHMAGihxkBrvUJ86HPrUSgahXjO8Rpcx7maRSuzpUFnJGudpAta/NV3oG//h
CmWLnOM6OxWoEOwAPZKEtfSqf6NeEfMkTNOPaix7JmFdWsI4OMXjRxoX0hzeJCpRKEGH0yvI3xls
E7btW8NyQzonEjvknZZhlwVkDtC+XhZKOhdwCVmBXGBlbsmFO4dcKDaJCPvdwQyWdcz31lLRDvix
GpJ+A/Le+BfrEaFFIWsFPcIEX2/JfyYI/M6oWdosQkjf5ev67COCOFvu1q0jIAlA3DkqelByKzew
j6RYdobqACOco7RoxVAR6Z1ywWGuw4XLVBaYmvyVqOVNQEjveW9YL1oCZml0ARsC5u44Ja456uld
sejQJuarPsBm9RdWS+6fKZ6/32OTWPILYQQ9urCsg8KTXSp/vi8dNvrJGAvTfW7dnfdqKP9awzMq
nP7OIE7175wM6vxD5BMIdNcuD2QKzrm6Px7/TfCGvg/mX9ycpzCUZjmP4l7IdG8lkk+kpIxvQYgq
Pmc0oKNm4lCiJJrSyGIpiBJ6fRQVp0Dc6nwU2zw6dpIJTK72QJPzB/g0Yhb1wFUhJ5C4JgwBkVII
idINSxu6w+VRqG90SpC4wTHOwU4n+PEVVcpC3KKRIOQb7XeBejfbZ1UFig1jNLpabAG0VEbf4QPf
3t1is2hRkUEcHlrOahl2jF9ZisskKxZB5E6B+o9p91G3gMbk2S74qpw3GoEkmhNqVkly61XSbEAn
U8cjlHbClkf9vSF55jESpnHxciDwIVbmWD/lG8jdyaWJxYpYQui0/12jAn/UYeO6AqotsnY0zWUc
d5VjR/vPLrwbgwaKscmc1RL+52U8KpWuCzzOPEN9wNhs7yWQgfdtrFtmN0ycczr5wNNzpKGovKHq
U5WRFU3HGN5vslFNPv/VTNsGsNoQBSj2K7O0wR6u3GYvwmbgph1ECsz4SSLvJvSHfbbG5y1aKIK0
uAO5EV1xtljMeQK4RbosN5rwSjuook9vQ83wCTIold94fHVPOROhciWH4hmNLdFRGimWDFeKr4DT
XwNbEDnuzgfaD1PvC3sAvGI+CxWn4NLWWQbN+LDED0GrOvDcBSQu67jziNHvyiF4FUboD9qJpaiI
wsxftSug/Rmdb5MRdKQRx9ppMkFl+U4qjevxji5/HkXaq2x53vVyH+VqwrXoGlSZ1TnvqQTND4Nt
jI7gGmshqh6wZo6f9IZXhMFGRhQ1w+wdYt4J6E7ysvo1RIl9kVbyd4+JkEKii2c6E0sNa6dmytG1
+RXS7no7F4Gn+j4LTY0cokJH7xpg7L4i7D5hfLUQ97wZWlnxBEaLnjv6dbcki3uyXNLmixYMpeRk
lqZKJsqoqXoUaZhJFlmNlUpcA3H+f6JeIn63qTMKds660Wd3EDTxGY6pJbgFdKzw83hl5/b067I/
C5GNSa9yWZhjRkI1KLGxRO9Kb8mvrR0P+FHc4xizaTGbSe8go9EXxH/vD3Vm5DIxe2U7tVcldx4I
V3ahkp/KchgHPdy4b40xGRDhgyTK8xxRp7iRBzN06M/UhW9gOu+hesdA8qoHPp5+0axgCgRl89iL
l3DjUKAdGfFxH2Fqa2CBhjkD6ufu00lXu11d+SJtCxsx+KKmisWCGBUm8tYBN8MqzP71m501T/gi
i1MEafvAhAEUeyzNuvDxn5CHHb0Vw46Mm1XCQWd+hZ3v+99lVcmA/HaIZeedBiVAq4W2v+/TKhPz
nyXNxCzLebxL1GoqKA68S3hZ9WnFot6uVhLO1u5d4qeBhxu/iIeTLLMCwqIS5xg+8s0O6MfPlC42
r6tHFS+pIF+ahLdO717JhiFXr2Rjf0jX70k955MfJH1Vdrolv/Ig6Ri6zRSc5BWFOTopsNXEW1Fv
CA4IX6fhxb2HpIpK4PPMgd+3zDpnbKiBofeBbgqx3cka9sLL7GHcYwaoteaM5fm5Ff2TvJMIPq5F
M0ozttUIYXAtZ4zc4k98ZlQjMh5xB25U1OmgwITEpzxMV5lEj7YhrGiTCWwijwmtTuTDI1fhcxwj
jQY+W4dKFyiL6ef6jYJPLikg6YOb50znQuNL0DzuwusHNSTRfKEi0TbImEqpNUxlkDccHtxwDSew
SJtbs3zUe9ZTjZ9pmMk4aaRARVkbeWDMPfX/xLZhCQYkdmeY4yiySjm2A2xgPd62+ZEE0BXa5aWb
SjzUq9fOaPnWVBhNHu8bHuK6decC9xPcor0zFiawJ+s/rgvgxsjH1LSjS9GYuGgW1GhKBVJtP3iH
SrzYnjmVBE0wfqR02n9Z3mA3gpVn/skpen3yuPI4orPVhA3bgzYzvOuZzSkBA1gAd0ObATEGZfAO
nWdywMcnZaCOJW9o3fYt/SnZrrPpdPpt1lUvCLB5wZ/pxKvBaJoUn4IkvhohnbSvZ5nmQRtgwKq1
o968RHtME2T3VuZ8ChNufeQN8buh099Vx4SCo4ZY6lrt/ufaZ1gD2oyMZ/03rma5FgrEkeZfwFhY
JUnR2cCRIyCse1tYBqb/q02Elf33X0nQkuxWIsEmGk6mEBfpkEBmW7Jwhl9v4w4mTH5xm0bikEoB
b2WjpWZdD5qMyihKUYh3F9yiHCFYjldiuTLsZYv4Dle6+Zc32dVScuTegyYxPj7RydICqoWiJEet
C5auzPWcyFoQMCsxRkrBJaTn+B+2M9xfSKYNBTyNC0PVu61y/s6EbSVYqb4yjMoXyv1SZsz2Yyr1
gYdkBfth92+Y2Puv2t/nnBPOC2wwyHG8I4o4MMDO2aRAKk+VXdL5erdwzxAJvj7EAJj0uw5V+0CA
acw8+M6LymFDni1sRSN+CHwFKaldoh1M667+VObk/28T/jl2wOUYgZPdKAUAzEAglfCkgE9tNt8L
VVLkEPU3mf9V7gBzj9Wr9FNKWqVV9RWvNDmHZLCweH1gencyfqEkVTEXddTO8a18qPyPTVbrJH93
CTKCkLgopzM2p4dWq+2ie5tjO5V0nG+5MCzV0CLbbwLoV8fJSuoNpsvKJBV1OmXZBP+5JHiZJJ9y
hcUQpIL5EcGIa1uMG9CIE+d7Cy9plMZ4drjzPAFF1GmihYtOgGMj0DF469Rf7G3LaNmxauLvWYOK
541z4LtBATGepl6+BLsfCz9OEGektLNrQdS+Ih5JUNDfCVSZGziEeLd3DGpD9BcxemAgTWhWLtId
k7a0/vH8ZCaTVp2YwJsvdgWlC8U3OWvNtichD4x4kzTOztYE6B0eCH6LmLW+TEQt9K6PcDRiMVwL
4sDOpOWAiYPJoi6qrpwd8TJNLXwFsPTxmgQQjkx1/RMF3MjTPpoGJMlMWPgU8ErQHRKN7M+Toxiq
PWBnLhOs6bntkFezNmLcXKXBq8vtmFIGf/8a8wiqPc4So4GB9OY5DYau+DgA6tgqAHXDPB9kvwdd
oSO6b9Lj+SdsL7oDwjr9LM6imcMN0tvRaEqXDZNUj4oUgdZpbHnb3Y3j4KHJiOj+Voux1bsvFozL
qNA9knENfkVM1ZsMf6do0oQyeJzPbOZFUdBoWU6ZPXpDaLwf+LooC7T2LWDRzTH0iZfZ4ij3umPa
YO84a5kVgswc61bOIeXLmObQzuS2bprmNocS0ebafFFZ6DxKxt9eTLE05JR1Q1BI5Qqf4Gu9xOgK
BY8sdmy1i5GObrikENtRSp6zvB5ybzPFvTsS7v9B/QZJS3fJ0kSVr8CsQBH4qLgOLmWCcxxTz3La
Cg4o4gXL8He2QOvAnmemPpGzNBgnrAgtE72VIyHd+PxNcmXNoFWeDUeaRRoUxvMNOgk0hSJrXPR1
YnEBqrgFCHuIAzNCxTKEwMurryUfbaZ48cNG0/EBwV2HQ0MpSO8XNhgaqlha25Slb+5pmLpXYQSX
Wm/O210IjAWvmg2RW3VkCVkXy7IeHOpLjGlEuNK5w3BZpOYek+QQWWDmgM02oyczQ5Kr3u9YrWHe
CpyvOlZrgTeAI7wCl5dk5URwQBX9sV/DZ10bAupIlgo1PWNG3j2d2y9qP8uQm4dYoFKSXjt6rsvL
WXVj4Y4DmhIVW8gDPY2oZjHx5ytViR6SLl6SEwDqMz5I90myPSHgB/a3N62afuQjlLiFVgVQ9CEe
aWoPrQgOXPLhaOg0J66hKeJ80RPePpneRJGWDdQPT3av2yPMcqeyNXE+B6Gz7Ckz/3fyKm1IoRdz
KVZC1OSqyO7D9Lj/QR/F5MiyX/U25qq+DYMPaOXMhJXzwWyf68ZvLRWdknP12ycegBDa9upmvvTz
aMvudnL4of6+Ji+egLH/q6+J7c5ZW3PZokX0Z9yh9mgHiyZO4fcsQKqeIx/tfSdpOg4JGzPbx5ir
Iu5b1+kIWLRUXQw/JVAr851pIOPwE+vzrcgXNshRIlZaampiFqB4YYCZZygGzJbbSomA6lCDSNoF
AuTrUa4BTWB8YMZD6+stpACP8E/EW6bkIftaPZpPS0f576EWUL4uevu1IYm6FtZ3tdaF6RLYe69/
tn30tY+HPfrMSSdxtnyud36mA2eSTS4x+ltRPJvP7loB4/mBYIpn5Ae+eWsi0VEKc+uo6VteEVwS
Pj1K8JrnFotEu9hWe93dMulHmCDc5yZ5EVBB3W+vR8sxGIBZUaZZM0vP5zhxiAcLOIAkG+TW0bsR
YEdAQDtVvkL5DT7pyZ24pavHFbssob4KFUMr4w7OVIHzhVmXTRMdBbhDGhalVWENoYR2Hw9k5rFD
+zgBtsaioN69wRFrQ+sCLtRsoMryepVlnPYGs/QUWDSWC3ilt16N66f7OAdAsi6s/vqOGQp1t1bo
Iw2ZgF86PX4G586DfPDbUwqbZwBP0uC0jhYaQfVMBouND8MH4u4pF0AMDn4LMmR1lbSpfPwP6lgx
KnT/xGNsPdbAKOCzc28POmNwQ+PJp18oSOGetMpsrHdJp31vGJ16zx1kIR92p+Q1UMOSN+VpJ3Re
7ftNkbpgPRo58ua1jQnCrCzi3aF7Bla0rDW1wesItlPUsm4u9l+rfYcHlzACgKEtL68yf7V8JttS
VZsFqNEiztv9Ni+9P1/ynvP7TBv0NJqspJkINCSoKLhdwDwL/ANTks1lEQuuW7/50bVU175u9CUE
jE8t0qc6Q/c1l+jTV8GkGQn1FF6WeeTndJ4iAUvpnkNxjW2J9am0YCOKFEJzD/+ada3eTOSpJfDW
lM142DrcpBQvay2+Zns2sMZroxWU+w7flFXb6q3AXBFlgi7UXHZYjEyzweVa7PEvcIh3Pm8IhmaI
lj8H1OYGKMM6jllaP/l+xzieQ3tHgkH1Ph+FdpmgJvwa4zrmfpHDSdkQECTC93VwdSEkmAdM88WI
I1AOqRuXTkDQbbtuNIHx4I0P+Doe5od7SFTVBuDJs6RSuXxElar9VnbcCwtoiKGXhi/wIDmFtCRV
D/wCbVPNRtNcaq1BZM79c2quqJF37d6TXEAbMidlCBWCQgZfzSmv1XOkGSE1YhlIRH0AAgI3HDnf
fmP829cEBWvHf+fI8EbaSyd5fgW1/YbYHfGqZMcNPgSc0Fv1cw6vbmyPQqfsfWDV7qnb33QOWPev
AS5pC7kuvqT42Gj1KiBTwvnhUIOAGEmD/AKAEV+ZkEtmTnOUZs8YinfDDJF3biaoz77gcnAsXoLj
pPJap7ssNf/NEM4kzxfE0rfXAy/fZk9irngH9+wTFE4WzIBeU9UJfQG0f262pOTdDgP7U3o4+T2y
KsA9YZx2p4Ri98BSD58WL5Qbv5ZHlzLZ0X6nSddQoWgJ9okTm/4wL/gSO37d0UjnJGYjm/W685O6
RRSvHRScUpIlV8p7nIpMQqCEydYDXIkzrmfy1FIIzRlKncBD+GWGjbDNJ71cpAi+WmuelxtOv9Vm
09HvCEybQiHsScaNuqHorUBQwxNaaMG0xuLLsviz3lbfRjq1nm3KBfNWv+5ggve1gle92SBinmVq
dalXDurQ+9BEyx7ZB4tNfbZifkNrM5PSZDAvufouyN8aeiMRaJQtW4oBK9n426TxD/iQg9WKfVuR
x3sr2eCpLjc3jI2uACVW2SwzA02nDjGiNQa6JFkQs1NFcSnM/+YY/d5mRA+sdX3CCstMUJgjqr6t
SrYsrmZS1FQ7xdZ06q+4R2aIidXeASsfEn6XUFStH9P18gGL185Oi6h4CGeDRZSNYqPYJIavcKTO
bSlLN7C8wRijdkf2KLAa4tFH73Gbxxb9Jr2b8SNFNw9eR1jlM1xjLuesZB3ebAA754HsN8UiE+RK
TCt+JnuKZsnuL43rjH87+4iriBGFqAdTRiv9Eo4uE2NTkCUcSATfseH4YqpxFKHPMuCUTp8P8uBR
IsS/T6v5YjgRRHtpCM97bE/dOi9f6i63Z5xveQyZczGycvOuC4Tjrz1Q8lYxa22O/9P/NIuY3snd
dm15Ewc++/ZFbyha/CTQjOMU7i7TOfpMFR37jDXSRBDRYhv48ahoQDGAWo7zSjs0P+b9oizA6ocr
Ekz1IeFJZWUf8DEjufzcp6W9/kRct31QxwZjQKm/aqsvX4ZQuUTFqpES2+VL+s2U2fYZB+iTL85G
tGulJBBbcVoEXuOP8E3iWtaZc3QDdk4Oi3l5rU6N7Iis9hhP3vpIM7kovDm00QdjjnEvurznVLus
RmCMU4mghNFZX1fB80DVcvv0xFdNwXhiuRxMtWR2zvRh6vNaPKLxQ9s914aNEc8nmcT0tEdm6uaA
0oF/ZVIcI6o0WyiVXpQNGP2/Ft4jN1TJFwPvWQwf23E2ifRz0tbLZkyPDIQVSgqW/+O78wRXqKj/
F0TSsnbVHNeUKnHBWRZqgqFUVdzeDS7972zNRPBpajhmg99AhKutlshfDeBqgbl+lLjv2OLwXZIe
BbRVMFTbpONe9xyP+dtnaovN8IHsCXapohW8B7VoyezRP9zLXBrdiuBw4TwtcreXwrJvOwD/mGIX
LziTWJ0u0J6NL8h8ORsZYOC7es0DbA65IaT5jfNV36TAu+tnFo03Akuv2LIZjO/O7oLJcZ3IGF54
i5hVSO3KQyRZHeppAMfvOBj3zQO587HvxfJ/qaYkhSshPnKhyQGeeao/9c/IPW52zc35j0PoeqSR
2NZGGluPdbNVQLf+bm0mGbDTfpXXxCLRFMaz14ogYXVES74lBQlRHevSPHTdAOgdY/b3tnMe+AB3
qBA39oal/IL7gC1BfUTvKQMl9tzvDSxjkk+PNvghpA02PwQyrIaMBnxiAm2BDaDARiLdCSuGMN8J
mP6LumfOdV/EkKMoJucjZK4UKIvZhFk8GoswIBFOd12F4tbrAKLnyRfRXQHYH2YNeYah8njvvj+p
j9ytrn+X/ID9qmJaXjUxy6P0qw/k3Bpo3qP7GusxBxPegUcb/AsRQQeF0bPAMxlxSad2LSM92Xyz
o2OF9Vt/ek/W6AIfeFQDhAu21zh6cVUSsugL2TnOXv2b3jKVVtbqE+uxoG+zMMAglIzXsEgaH7bT
7mEPPc0TXl25i8khGLyF+c4FQ1hyNO0ckDGmr7W3vFF4RmEf3dP0mifTwr0SOtguFq/f+oD/TWQR
zZxgizhSNm2xI6uOCWsluXomZVZeVrugLc/pp0a1loVXfvMoTLapHc8zeAJshIGze3Cw3ADZaI+2
9u/xQu/LwNBaTk/z1/nPHA3liYAqmnBrkrHZRAPausA+1lF1wWIc4xlbS/fdGBYvC1rU4A9bPEd9
EB90Ve72V0m67W6Jr9h+jDiRdgJxCNgdu/i+2HmF2S6kmk3ynDifXL1CpRJCbcxTD3tyVOz7oCsu
PqcWxXlzPxfhnmnSv8gyB4SPSrjk7ZZfZbkK/bfXhBQ2toK8DL6DAHpkeUMIVtPFfwg8vRBLxik+
ulLrcin7z5OQT5WwDVPNRphTOTSFHpPRGQpOu+NNbQhJeBSp8k1OJXEQUrdlY3NsOWz1nYWwIPDq
kiUYML7pTand50of7NM2V4MPWfyiuhhDvX6cDjLGD0Lh6SCyG6q15fB0psjnNc5Aam6gbtgCCa2q
QFWIVgZiT/MXn8I97qzYmgDdUt2uCIZ8275vRmwpqStlQLnZKE1J2veYHlNi7FhD1WbqRDkd5d5+
GoBs92XkcmLu4vYWaIZdJC/Xg4jeFil9z6EYx8Zpwwm/uvQyy3HrhmOlZovn4neEJFuJeiyRwTTd
wgjtbpyLVfeYzIbPYPH2OihX4fxDE0R5ABd7PRRzDNAtXweeo7jOeo/KYcsG0sCiNI4axdi8S5Pq
q8UIeMUV3Os/fAz5DZ9zVvZWFs24W8rfwMMPLOGRK5kq2uyOgKBym6fIUVDeiXczy6QEy9zTQB7G
dAjBKa6bxL3BDTj6u35dJEq9jOWo7zxaVhI9KOo3W5np787isIvtDkjNai93gL803xYnXr10pDQU
x4zR3Aawy1AguzEL1kkaJJoO/xe7zSvPvycmMD9/fqTB5uP/hMnCixFB4JHlLbstQ//x5a1KxReb
1FSAr+IBwEGuWin+DcfUIoUZ6pVVDaLTtnoM9AQ6Mfh8Bjtryr62sk5EMg/DdSryxVLkhce3inzH
JG0H/z3i4RIypWUV2fpumwVOci95N0B242cQkekdoKIaSuCf0egkmAo3Lbo4jFrO9gLRWdZXcY+k
jAomVlTHyfOVGzZS1MWZaW1Xokm5cHURPdAtJvxg4Q/dqi+NLB6rZWPKTDe/DHlewFHH2/cBvHVD
LvHs5w/w9NLo14pb6mY1OlwHoNeqRFEQI50svdLKq6Scw87AYXKnuotl+dF0CO48GtY3MMRW1qzO
wLGUWVhqlIlj3gpMDuporMPikbTLxBaDlSiyNA02A2BJUcuEV38bXxpaszvc0s33ZcenO4XFJQ/Z
MyPEigiJQ7ap615pSBjkNZcv8EW24vLVEE5ncGFtBctFezFJLnXg5CdTcuW6lLoNkYmX6ZY5zo+M
w4PL0x9rBRkcddbUhkMV5ShrGFuez/Wxm53bFycwg3LXQhrruMVnZ4YPtRH6aq/7pIjfrpepsEsm
kjz1Gcx04c8ppaPdBCLuzRmmvzzcWzxSB1fHIMsyBDL0XGT0uxBVH5qgCOWwmrMptNCpacm/XoSg
7/nDZ6h1s4Wm5MwgikS+pefbMa24R11tgams/OsxlfGq6+LChJNQSPD8kr4gutETkCQz2n0C3VDI
ZZzASDY22y7hLuYygxEb2tO7eMxO5yVlFrt8Cp6+hGhaBKmVOaii3hy03CcDWngU53PzOunxsOOt
cDnjLMy+J2KqHmv5ty2i1pRU6edaP1iMdw1zaidmlPCocrEMUDYXXKOPfz7/VASdE6k7R7SqFetn
O9S83Sn2ATrNS7WpYecH+2au8l5wWaOXJgnVBOG0T5cWScX0a96BrF+bl/51IzwYwAATkW9ZMlCq
l/D30hUI5whdMBQu0dChPdeiEIgIdXwtestgTEuZUNEXZtcupvHL6B/rN8piXigHjb4N2OBgC5s7
SGCiL99joQEaiwV9XexiNEubsu2gszbB9idEPoEG6J0JvulKmOwfzLiF10ymNyXGdWBQLf2WAX8f
9XX2mL/qv0SGYmM0UjudjSV9og1y5ei8mBfXf/A3hn9EBS4J6uyTPPWX5Q6cY80jd9SnQL/KV9cU
rVO4nTpMOtcpJhg0yAGiWVelMs8E1vBgX2JEeMfYkDtgo9G4xMBu4hGabufS41VvAP8mFYCOAD/O
D2ZedcIah3OyNqeLvamVAVczsvfewldy2M5E3nZD8xjGE2S4oxy3ou58Gyzics1nz2HFIEMPAAra
6WgwSnJyXefLvnMJxJ6NoqQDkpqH1xTJLDuPuf2PTOXjkuphvRMJtSA0cjYn7tGzszeqNrtZwuF9
FOJbhupafpn5Zo7y7F43zbYjuYldGHoq3KQWOrKyP6dRhR0KOJt4Kl7Y7rPn6VgJYNofDFW5I8pO
Tyx1TFdIeg1PUT1ChzOaJZJrmTdB1vlsKXrDoXvaAUrI31bnf5rSUr5feYZ/dVE81JD8+9osDjEC
hdDAzc9+n3/mBaTgTCKu/3vZ+mR1bkWrsHmeOrwIIMNwtWjhQk55mDj+Ts8D9RrowB1zOxla2wJP
MGlcXkPqxzw+if/pFh1nkOfhRmvjs6Rv1G7yLzE/ATERAmHo7GsSqZnXMatUg9OuPM97n/YHZOBe
wGo1IlPGeZZWubr+W6o6zOVJYsbwENagu34P8D9cFQZJG8Aeaevd2dR4b0AJPa3p5mOZQmDnr6w3
so6fi9VcWus075fOKYW4eKgmrJ10YgHWtVwc2P78Xqu8WZi/5T8O6ZBkNC1DH6IJT2yK3nExYtKk
VLzV4L9cOW7K3aNJNBTvQtx7mhwYHg5sfcP04eGNrnvDdac6v1Tfkkcmc57ywwuxlIywtCvSpSj4
QMdXfyrETs7mojmg3+r56e9SOA8yTKa06fgDGRZDriDlK5SFK9kV5FIY6YheSEROg4DeFd3HiIyj
f+tsfx84qpEPpBJQyiHzRIqmXPI1H9oCbAJuWpsMC7e3gv1O4AKlo4ZYGsXYVVl1DDGDjBNJXJ+V
2nCQLFlZivr/JCHV6RZch1SdRqyF65A5MPzGpzj9/1dI5NcANGEWynYnfD4xz2oTS71vJYHr4r2W
53nQhGQoYv/uA1bhp3qE/5xOJcc3V8RrL1AgviNS+bull1jB9fGVeg8v5GnRTZ55u3/d5xp5f369
ZdvuA1CC97qUsQPquqsUTF+b69Hsxr5bOL6h10dU1Jc73xNJALrz1NMJpPUZhpB7aH+y5LPEbLll
fKdaMr1ckiTUrimbElVPu/LC5JHFh4IanNM0dw5E2pgfCODV0U6N8W7R6/DB1WYRpVkO3iaBAMdX
XZmexX+IUpk57Q0xc/S3bcWE3QM/w6ZRlefqF7YeEfAO4vabK/Irigtsq2Ecll+EHFtpsGM5nSFi
eG5KMzkRHgySPNl6ybZA5IvvxCvzBem17yGUX5HcQ5DUkBTRyj3CsDCyDo64hFhunDZkTyt/MH+T
erSBdqo7q9rhOIMA84xDfWTTjfXyuzZIqTYl+1Ca67LHl0T7a5p7+gQ+6lfX2Ldx3VWbZP/fUMPT
7FP6fp3/t7o7F5N7IqmNBrjsmy292Ii230pZd93lLFb14Z8o5LD3aYmDvbREhXDAv0MUX8aFcfCP
Do0WS9FnNLPoFlrmtn9ofguo6JjyuRe7GZGPcZcYJRudt1eEjuSiF+rCII9gx+bugBaRafk/dMgJ
uqCdZWeXk5gMp5C2gMyllVDk4TreWXvuoMdm9T36cq9O/blRfd7IYOc2v4JgKVHzojXGZd5Bbf1w
EpgJ4h+SALMLzZRZQbV7EJg1YgBxBc2WR9t3TrmGCtyfTdr6E88n1FlVhj7iB7dtiYGgCoFwzrni
223tMWy0OJem6/WVYFSXvJESeYKi2bW4lh4pSWgwEcigU4I0Z349IIdz/k3pIhau5IKp5NbZ/UH7
633bccdd/6gpYaKNJMLUodPVoMpM0q7K+PTGvM38U74GN2jv/jo0/y2WDZ9ggkNO6+XvLVKSE5pM
jaTzz56A7Z9Jscgls75o/Ok/h7M9S2dZuSoIsKyH46ycnBsdKRdAF1dJDMUFWx2otLc55we9COI7
C+SWtl8FmOhT/w6FAA5V+/gU86hDWl//sZkGZ1TVpwDzDd28pBQYworzs4uB1FbCZtxYyn/iUMnz
/UJxlJN7qW4bFKRT6X521644UZYOyr4JDPuqaex5pqhlAWXqSNGtqOSfSfjHahwiCgsypKfQA2q/
l0MKrN4axMJ8zouvIslzRXBSjFvOQ+r61whmftBRY9h7oUQPS6XesIYyle4i9g+XcdObXVrerogH
93eX7nPFEXbqNY2svHbVDTn3tm22Zc4B0iBWiVEkgshNCnxe6hOtECCQKrmIgK3igR29YjmoblRt
pIaxm8gyF+fxfJMa510wlAgl0rv1M5V1bdQ1kb36CoSQ9SXPLA86nxUogC3LXtZa6rpJDz+Zvn2b
Wq/EHtXxmOEoWI1JensvI9IECFTrTP1YUSUVcCzgpQKOAV00zUAABN4a5P/U8opCaL97s9J8fGyg
pFOuXerRMYEJ5Myr5wkQK/RcbSgNfYngv5luGTkEHJg9pcxgRz/xHBqHFNz1bAzFUXFy3Guhf9GT
4B4+8rR+6t9SJ+HNDDMCyAQWWdFKqb42cqM4qwXhS++XdHNlOW2taxNiojBXdjJ9bxNUhf1iL2bn
4IraHYGNyDxDrv0MqeEGiXTRSA13r94sv+z4Bn34m67rYggymWGFMvjABCGgIAxEeVe19BofZDhV
qgiRNU2KY8z9hmmu2LiJYUP/cdolRhkzbzh5Msphi5g+D1CXhm8bcB0ZOBop5NP8CvFZIEF8YncS
e3Hoc9E2ixrcVwx1Be9yPtPgVic9aKb2gkJsGd9wMxLQMbB2JwgtxqAabSe1zMwlY31gXhXr3Y7/
ON9bAXlHM2QNBFVs8gcvCUJ5RPfwkBa6wR7zrcaZNmaPzJcqZ2LCm30l0QchEW7UK/pzCK3m+SHy
vkfNcSizkk5GaLcuA0M0dXYuuQ0hoOfoSaAqAIpZCM5wWxS+ZF6AtfGtzPGQBkvAEJqDHXZCIYwu
06WBjFgFpKNO+Ejd5z+x8PqwxWb3Eyyod7BX+l0b2AMfIxno6EOMEZAVLuygW7ejIb+41dYqoOVx
sIkqhjCyLl/DxmY+VuK/ZSviYsm6Mk3eEkWinuKk1+Ykefy31YPcrKvgVMjIYXHqoGSPWBZqUd/E
sV3UJpcP9memtI5Xbff97zkZ0UtkEjiFK+2usOSX7RV52AvRXXDVmsCxcFhah1vvo+f4egf4INkr
KzG4QUC02l51gSmHpLlgGHGgJ67SjUVEq6Jaz/20g+0aHppy5vCmBC5Gf5V2niYB4c69L+igqUN+
S9algvC+LPGAvE6imqDTBEPk3FKx2+9I7q/R6s0Kkye6jqahUtKhHULrGMXMyHnBEzNiJeeSTFND
5P9MDbdwxWAD1fbXxaDhHgfUF/xj04nZaGLQWjVSXM0jT92ARKtwCy7WvbDyonN7Q8uMJ1qkWES3
p4SN4sgX3AcgJQtv4cX4NTzL6vxyrvWndcdMDyltt+UbcaI40raoqPzofep717ICuGQv+ehSp9IG
dkaosz/B/AVsAzVbuwo039IsLsGV8S2qxiPcjQK53g2guk1jTalY4EGkpZAto7MzRIQHvDjDUWDw
y0FQRHMq2F8axdAVTZWWa3FjdsDOsYylcJ4wFDk4cPhfzYiRdN5D7hGyXa4mRZkel2VUBb+a8XuN
Hsloe39/toZeadH+PR+GU1mRZ5qwtt6OcU4vYCupxzXCiAk1e1BOSoFSmni4pGsV9+Zl8I5mBcxj
K8/ZLBZnAPVxIsljsKyW0cNcF5+dbm3t5BE57FtmRwZZqnEujHS/paFGo/6MIsJNdJThcYgejotR
7NEqpcEKEFJ33JozJKD9bFyDg8eSTlWQFqqE1ZpOP0cM6W/F1eSCRDiXhm3VmsmL0v1lKLH4gf7u
mzHU8nd8CA0GTJZLMs9f2LzTluwFu6tmvG3HQDk75Y/ddamoEQlo6h2CFLg3Co8g8dCWy/fGL0s8
Dink2nSxZKDwreDUcEtLWvpzHxqQpi6K9vy4EvcnqCT2EHpOBNnZKgmq5uMe0FasmaJ29aGWYTVy
XWEssp5iUsRAstSLReJpAmfgIYTnhp4uW2k0eLDg2IXZMMe7w8BKY6Xfuaxs7ptvTO2avnpt9ppD
jM2X3UBp+Ac3CZzJv4JYEOikH+BgXAZSsJQDTJkZbbchY8+e/wpXqoEP+MmDHZYg/3c/mqJcvoBO
0JF0GkMZjlAF/QaD6RCnAFsq4HCqm2EzLH+F30Y+VM+PJ8JNHaRPv08PMMxI0eilqsxo5OqPTknU
egSKAn+vPQXqMNFcpueeDOyN9Xv/xnUA/sHkVtD/axdeYsT3bRPMXGjNHJp6Tv8DkrwuNloMdCDA
hGX4FwHPIICaTDVegukOWD5xt+jYtgNsP58Q4cDQ2wHQdC6npNfolSdz0XQN+7s20Gwf6QsNm7kO
NZNcMSxw/Wn4j1NxSWVnH18U0hJq9WSL16Se6dWOvg9Q7OEhSYpQjsh8JkJPseQqEncy9Dab0jzH
WLq/jMiJnR1mjdA7Pr3PvoXVbAIjnfyMDPkJlNSP/Gtn6WV7EdURsw0TqAyhO3iKCdcns4zVIzTi
XRyxysaPdqOfYzprbnT8+YpukOZeEC5MT86xFQcvzeyGdFX3DsNo3vI4N871S9Ez7pTXS2hC9Qj5
BfklHa5VSDtpXTXbNuhYRirA6F0gZmsRp6PD/A1dL3GcUux1bZvi7ZupuvjNjWjEm6twzCS9iQay
WwuTLc/AUfSEjdC4dSe/5zhWlBd685TX50OSI/7pDXHv4TLq87m2hb50MVDP/COOvWUxAxSTsSzt
zUyEBUBc+jmc0Cg5kkwIAmE5NBtyUZxj1L6+r+3lmP/sazv7oGmj2zMyIxAX8oLLCG0jyz0RSTOa
MIB/fpJsUsfPCI0XP3VC3DbaxyDp+LD5SMlmIbTbwAea4FZ56LtTdny/dMu49wzoVR0bXmqWytlC
RaF9FrBkCuPAoTiDU7EIvlmifiuOAEHNzidNl9XJ92mOCFXIQGxcx9AI/PxSKoruqlWtcUq0nUCv
jF2p7JvMrZf5+KNt1zjU7jvvxYl/OmUWeuEUpYUcD8QmCag6EEoXgAatYi6GvCPrnDNuzeHLpvSR
GDkTphGlTl9b/iYIgkmUjDtxBaEAZ/t2Cq+LiuUeWV24Ia+6uAxVPjef5zKRdrcncoHHBVISin+2
LJdAm7NXkI93lGHd6PyArJkmjcnxxe3NcQNyb/u5n9gfgLyl5JtrTVhxCeIA4Agb8n7nU1b1PMQ/
j9tLAs952uO1Xd6cMxtVpdd3PEBRhkLMp0JiEWrfNhUVElsk34m251lsJsy9RGuMOSy48/Xt6M2w
xspothfU1JbAaeo/uFnz0OTATySyWeY78hTddytMnHTup/wq/ZmgYuptHIEhwiB9DEXP7WETQEAO
SiQU/ZvEvGnL6Hm1czs6FdD6QMbzJtdALvYDM8ra1t1HuUz5uGmhgkG6po6aPOoDrqJJQ2XW9XJR
fjh0ql6BlFsqmOcfRrmEsiduPoEiAGCdI57gbw4CY7Z5Q8RpBmHquGDBSFiJjM5l127j6MZDoLph
vS3q4im7D/JbaRqWeo5677U5FTlDl6Pnsz50DQfrzgRcySfLKw+B2NVPgdFbhlID29EIGGX1igAC
QUBv7TxiQ79Mxkk7xBBgTjxLs69KQnnT6whwWfIUD+t17CRtZv8R9n+/EriWRw46t+yavKkRRyv/
WLad3PKO2iREC6EsyGa4iI9aB2Vf67W+qGxbfE4cidAKigU7gt4RqkDDPbklN25/XgsaxHhSKXaP
6fEuVN2JKKZb8+dKvsLw5G7ysw4JB87OBo7dPDwdS3tsSRrAIb6hSxPghGOLVR79Sv2s9I0WvVO7
hco+rYwUqovorA2+mwCvsECGsUqZSl4vfuYZR8eFB3FjL0syg0VtT5xyPC4up9Jn7u80WLUkHTes
NvVC5rKCkUTuYDcOo8zDjnnGkRRM+1XsADPp5Ngc7ILqLUI5vsPE5lLCTC1/ZEz0i4h/NZHjRVBZ
E+lex4KWpD4bj9kW+NVaDpD+FJfICh7pAYt/95AwgUa+aywwus2BkeTO64PM7kHjFDY2wkemnAic
iX9hVqI43rs/oS5pIVsBq9Rw81YNxkN7eKeOL6bgUU6Uo0kndOv1pboAVu+HqWHPGBMipi2kaO/O
NAps4jkQTu1oCAtK9ZwNK5aBgaq38j6JM2RhMndd5vYSYqQvpfTEs89PTfMRL9Zi43nxQyz/7VYs
gErc+FwRf7lIsfC9HEtyLMYwagM5IuBjETUMDCSxYM5B1BLNyipcwoi8ExOkV7QykIiWTkqQjINR
7TNBNAsKPUamolaCur+56Q0Hl+x7c3Ugr/LoPxGzHGeVrQOtaQxgdM2nMKuF11SZ8BVW6z79cZlX
LSlhfe9Tjfimc9+D0bMffzbpvHS1/uGI4HZXIWqwWN6l/kX/oiPBvMj2CEB+SIbsimd7ERz0uBcp
qTW9Ysp+UxTWiN9ByWsFiyrY0ynHhBaEgvawLTn2NMDXzsKvrLXLKl6Dfqt04+tIOL8VIBS2Pm3I
/pF2Bl/lIkRg5AaeLnKrSJjQn1rtkO97U4bxND0gRj2wRXdzviaJzP9HoqzDbnuS3g52Hd8i2+oh
2zN6SHrOjaCjDFfOz3fhQj9cxfK5fPm8e4WcsyNfIAf0TQEeSG+FwzoduMiRM/RLhCP6FP0/Zuvx
nnoQF+bwdEMQiEvOwujyA8pcb1Mgas/ivMlkdU7e1M/Kk8PxDPgr7zO5Y73hOonzWKAU8KmtRw0x
T/VecSg4gDKMBSRC5OKeRy2tPLxqDvkPuH9TKG8mZXdtirkN/HvxYPjXsdhNXmma44qZa1HclYYZ
r0drAcLrN9+kuD2vbxuQsV1HuChVAEdIMhoiYTk6WEZKoKo6aD0pNgeANOh1we+nBnFPzo9rcibC
fpEU8B6jF0el1xrMdScWskPotcayHeANvst+B2s5WG9AWo5npKQSEzX6kL4AXsai2a90XSZltc53
5P0hNv/chgR1DFmYyWbti4hWtVjgdsZFEqUNOWv12sxs3ny9Aim6yNR2jSiJdXdxpTj7+kWbK1yf
BRWQiAFsQOqBWwkZ3GAvIiHqO95ehah0uiTlOg3ZZNJgfEomeoyfIo2MPt/WDjmulzmhU2dia4iB
c/21IwpSQBZlDbrbWUlbskFLEvhiGjrmDUhQXsJxYWFfDBay3Q6CeZVYUWbO+5EBKPuyYS28voPT
jYgFTqTJnzjVCby0fcuggqogikrahzGYV0pMWGgPYCbP20mAs7d2suDJEBaoLEAmjAK5icH1uewF
GKAKY6OkG92C3I1U8A3FG4V5iBtbTnNpMfJ7aCcahLOXymvz+DLViZ4b2iEvmnhr470PWN+HVZyw
jEK+s/InCLxebARXQMSarxlgP+YUrnIjQDR2i2UMU4YalOeRqxgNddJW8Fn3Xu7HUm2K1iWKjZwc
WYmZOH6CFnGy8WZnAYYHQYIXU9p53xmeWcDyUMigEePkwqZrdU5JROo19HOZX8rjRKfcEY0zXhm4
GF1MI3BQecqoqr+9OcxI9qHsvSkHPnxfTJll/fLtl1RM91DOPeeMfOF/RKrvuRarlhkJNGBwrwbZ
KIgAiQDnqV+UAsYq8hXyC3pHiT/DYNClnoEPpqCR1fDg4uklhZV2B2F7D/HtoVBAoyHqAHuG+Fts
vqk2bXBo80QZB7pGhSz7Sgk1AKsuyul6rHVfHfuEVvBT93Q2DhKpAgIePN74E3lEHKtIAdrvbJSK
hFpuafZFqoCelA5MER2fU7BPWO2oHhXtb8G3Ztx0/hpqt13Kn1t8bwI87UBiecWflvQ0mnzLpv3S
QV1AJdLgIGRMNPk+OR5qlflwUQMBLc2OtY5gIgYiDAx5bcVkjvv65H68vKym4pn9JKpxxvycAUD/
umucRDZuHv7JkVjYOdm55kKF2L6N9nhCJHQ2bFnnajKpaOqFVEHZV8W6P52XUCzVzzV5EF49GS4w
xllA+5l8xBDg6SHqeESHJmC4HZmROsbageNF/pvkIq7mdtCXYXpj7fi75NxhtuFyhxpxLRYA1gYz
ojiLhDpiFkYe8bId95YZzT7ZGdDEjSFG0q1BjYxwlbRWjLbSwFWOR3PUux+f8O2DKpZ20Mr39OZQ
+1Snvtc5kkpECdNvZIF2ikJbJk1e+JIVVOQMErjVvqugmhFR22dmULK2DWoNWGOqxTQomggij+7V
947e2QSXhwhYeHrCEmhDoE9LSAderikc9GioiRBllhpqeBSGA+H9G/xu+xiw0WQeJgXUaBkpMo9A
X1o2EvaTVmkdg7/4oP18NCU+DshxQZv5tz4nsMq05kJ0XXtVNRhLLnjB/Q9ygVumwP1Vhs/otEza
MjRQk8mzo+KEYTZFzlbXlXu5LW4M6j9UArcnUhmRBkFO0CsWPilUb8jM3w1b9sCj1jJC+8T74GCX
Iiozvdt9xUuO9InSKFSYE0Sgqlzb1m90HJjvr0B5MV0K2t8x+Rbz9Ti2GUPukQEVlJ23fYXuXeB2
/RuOuyocO6oGyFs77jsL5cdEWUarZK0zeJwpjMNs/bG97NjoaiJO3NUcpitVC/Qf2qbK4BLPdM7/
EPwsqluSjazP7L1Ug9bCMirvfX1qlmfE5zuKpCcJUpO2ycbWKZBmDLg+CWGlGpbmL0wpfUeVkFxh
mWpuMcf3jxMR9bpOvKAdM/GhgYgTiKJUOJ1KG3ibLoexHW1YrSefJ9lOkxGfmQUUs47wVeiblgJh
ey24978+bwpMhtoTwj9DY8st1n5wR51e8ndQ8fx6xCiC/V+3yvEvorw0ZVmxWDOcVivHMkE/rt+Y
gfbMNs0wNwqiVIOePiDsQvzjJPxcIiBGTBC+IcSwLg0LFpeSzTjGqvRm72Lw/pkfIhL0zwNHLcQG
2N7mQ8UMLUhjSrwr8jnZVUXoTfm18yV3MssYcaTbdh998JYUdA0MLsjIkQcYnE7iIvW6oSViaynz
LOibtWtA7cBSapElt0cfOC6pJeWaPALCgmj4pdD4Ph7FL8c/ypl0vZhC7cH8w1wVl5lSzXeXJiLf
OnCaEiQ3Mwbo/avVfyVtAsr3uHqqgy5Jzq4AAKueQjOWF7B5wZzJmDE03XN/TfEe7WhxLAJaupCu
qCqC0uKNo0emZqJKrqboiIo/CDldoTs4Gm/FYGchBzGA7W8x2s/vO6Qghr+hOnDm+abFh0hU/kHL
CA5fhlr/PvCTvKf/g/Q7IZJWm9jRN+9D4EfkLT/aA+LYySYpGaMGNUeP/bubqr1w9A///kE2R4dc
BP9RVI//ZvMLTsPoVPYggt78B/cv4tQAPNW1sjUOZWgFmH3DqXtAHKSkGCt4PKl+maw/uAR/MG7V
lLS/qMCHAgU3pK1HKqJJ6Fj1J6smsJ+iVLCBuR8n6VW2HL+CypeLNrQJ+MfjW4p94LN23n0d72M5
HHxmzC8bBlrTtvrTCxR7oMYbkLcW5T84sKrhTlSZSSDFvdGlL711shRvIg2BT7fyC4K6lPLJ2C4S
74B0NT2knu46aG94g2X3XN1UCQ/gGYdzE1gYw2ChBmnR3DpB2ConwfxqNVsnS05KrgHzEtX6SpMB
HDtGC9scH1dZABRVPyrupHzadMLIHlRekKn7E2nfGoXDh84Vvq4MiE4Jpo5vD84IAG+VJ9O67IN8
mtILJcyUubIf/TKgAeq6AjGZsfXuiLshYpLz8eVZ/A+STJPoD3kX0KBzlI+b72N64JlncJGBCfGW
udfzTVQgc3esCJuBGBS7+FD9dwotRLh/JeBkAx4EuWH3gkr6Jv6lO3yjnCH9QTNRf2krQogZEo5E
UzfT6PcK1L14+J1+TLHwMQ6NBHv6s/vascS0sIhaKZYvnyrB1JCB/iJUF9960T8X12+4NGSu6HJr
nuZX1xD+B13/MEgxHERdlnBT8Swkaa6PNDKCd/wgCNuZ+LGTrCzGlAj53AtY9fSIUxxJThaPwd7U
4Kg++oJzgTveD5nu/iD/VNS2QbJGejioZcb8ziD4PEHwWXuU6nF02P+xrMLYIoNDonUAppm4wATY
gdUmQ6iYa/LQwhYA334h0CIJxWwsn+xLaS9GGMTzGBLp0t7yGuwARaTAE8Y2kXBy3amz4hqVLIHQ
kHoH8Y/v8f6ZKroa7A4OriPJv940r5Zqd8TS1wD2Fusfv/VwIxoNq7zOf7zxBmbyD/phbm/bgl51
DYf1FTSz8vdej+h+lxwlagojtnJ+geB1JBVm2jFtwsgdP1U+q3xYwkmX2okgRzWYi1a9YGaDPksi
BZ5bkBz90CWvz0L97Ylai3TwpgkSIORNQuR1xpURN1yHZB2/W7PesfW5mjxN3km9XvUChmLuBdYR
kGOF34FKd8WcZbs1rTRU9Kedt4rKTkYJwkQKvFPRRnwTjOY/hgtr0hSrP1pv292xm+zv2lwpaZKL
aBjiJ6RE25qYlxU14tyADXm6091xYyonfeLK5/erra1OPa7XQG1glADE+DDPlANlLu7aGjYpotUN
i3fY/LpyQcSVxXc5zERbwdbFnJd9D9sTrk94ir3JzSYcAR4NZb796wSxXgn1LvFPZ0rbFEifbn9z
XgS0YR+4zHhSy9qmgY/j0k3EZZqiP1pPcF/Y7HlZ1G+3t+Bsb/277QGDHKX3uiC4/13mlBMiJz0w
c5OnBTofDo8FEH8OPRLhEhxo5pUx1/fXxLTvtf8RCkk7rimypgPY2m3vlmVh0TgLpkuPaCItyZgc
SNMOlo4unWGWAGg7vqW2WOuhxEE17P39X6yzcWx+MuchmVKPcl4+ZfwiWw/gCkg51KJaIXzkwg7Q
mU7dgdin/4sOKlblpBv/YPzF7JYa5RveMOFPlxWNerxcgSec5K9+amRCst6lrEWNlqOEqCf77yRN
KeybRn3AJBeUPagnN8UtlLuDeLTlRg4V/G2LRmgXKniPfS40Aw9ylsSfA++f1cJeQyTvnVmSSjnx
bZNoyqoOk7lNHlnZZN41LQnje7ycECsnJfqt8ElRJrskA8kQlA97yzoIj1XEtNRIHH7mBNPLFhoT
kkR0ncjiog9qX+ldByKxStP184660IaRzKMOwJAdkmFQLkXhVLFrftKgzWUiuX7yFoQhtrvGq7nF
Du3dscPyNHV2P6otKoBPmW6UPrCFNS9lNqU0T4DxwwrWyt9iri4NNTU+ExCJo86QZz4eY3ZSg6NR
vD5H3QyfZXxZUajygyaS8psmNnmRNgu5bx5OCIDeZ3uqA2nF0kQ6ddqZbGGB/fgZ06dx2wlhTB84
ArT/8X8TD1wqDaJNJbkWpkvg6pzRaHLFAsoQrlD/gc38SQpbXiws5mqTKx/cDAzpr/MjCPkPuil3
w0iU6maiQc9WXDSJwKOtQXXS/k3RKLChPVsZiJR2hATLzs3Iu5bb4dHIuO7jZyJqEKtsE/A/wAHV
2QMOetoy4pIEcJoQ/eIK5bP2Deq/H1fBNMzAu4phr58IPET+sQPu1cn7ef7TDEaxocREmgrU8oR4
kd9/wBjQe9Ao9BiKhIWBgC3TdGyiUNKCIF484a3DmLL/2w7XytnTPpXHHSn+rTjC5iSdTrP5VORU
HTvIav+MIBcsUZefHh6+rFYJSGhUVddHAl/4ytvp8s9KbX1gyaRSuE6w2CFdPZDZpX1C4fvbJXxr
lFePw4eE11SbQXkcCFiShPDlFHh0b0wRIRdM0cmio/N+QvUnQcfDd7lzVzrVmeoCgydAXDQswFbj
WO7+KwJZ+rZtUR8YZB1imVQEHBxjiJQK8vLrZgmFtrJ8xHmV60r6iGVL3odYLmhAiKIkYWNHAg7F
fTJFgZRGL47pcnSDah/3wejBt5Ug+bEI3RPLJT8XKb2JQeEOc4iHjiiZ9paGgd3ecPRfzCvkKrrF
1LEaJdtD0e0TjdTzXLsWuZ35ypm0ZOX+nl+JkMmmQ4m+YaUC/SRAQ23O6wguU4DXaH6mNO6Id18o
qS7jgkEAF1reYIDeB/a2/Ytv+l6WNhra/AVZwZQ+1U6OWog9okuAdI/nAY405KHT6s4UenW2DWR3
kWR1nq5+Rp1jW6PbTQU/N5gLgdjmnRn5vBrImQoEkXonvTdv1mxH/+cPwtXw28impOs9X5qT8kAG
GWE7lZQNRhf+uBT6CM2dosWSAE50axhDdqatlcdPdN/YBf3At1EGPjof+JFpC9ydspsfYmo1Quy9
0oOmudjU286ckDAKbL/694+79DpoA/itVxXlQh5xozGCefrDctFGJ9fgUfQpE4NRp7gMO79ApQqk
vmL+kxE8OOaK2t6LOoLX90hfv/ziiExqsej4u4Vy/LQAIZ2zL6n+T6mWu3jQGH40luZ99TDvZZTd
uVp/ggMLR1fzBM9oJjsmaqzlvHOUShr3jOaqSWjpu9nHnHlHn8uTlMq4mMf0F9Qtyib02Zfo8WYP
n8+JASetijyioVZWwsSwrMEcwOYfZ4SxLoQx83HT9ukV+PfgF77DZ3WIV4ElzNdx/hjrEw08JUpa
RpSGqNELStjzqCcm8C4MYXdffAP2AEWVsxIY6OVqSwzc3WPOAT6BGra12InUGnw4GVm+nKlw4+Lf
OloBh+wnhH73ZinpsqiFtyaYUiXg0x+3AIW90M+VZel0XUMz25+wInJhWQVcz/jK0gf+3to+w2/u
zwddpAJq5P2lF8+xJi+n2EUDt9MQhQ/52kUofLZd2guVPCdnTW5R4yYuG4P1z0X1oWqmPqc/A/R0
hh4U+HeAk64/TM+/lce/StpliYOI7t282lRIVMUG1Jy1kn+UGXkyLNp02ANbdTW9GcfxcXAJb9Db
niuqv08QJ7iulXWXN5OHBEsqDoz+HelTvvAKZR75M8kQglqhZSnk/VqzhSPxjkAkHdxIXO5GyXzS
XB/CK3W4IRiWW1tVkIWKgD2wxqB9+jUlvWJ4PxZ24atX/sTSPzC/6kjBlAYzhTxOBuFVuYx6zL/Y
dxS3YPBpoGvJjDl/wVSkcstDki5qvJ8xJfqY4V0B2wNaO21mt10Z3AcogwSNTxEYNKgRu4zsva6m
ZcUmfP/mBA84qWn+doMnIGXnbZTxpF966BGPRFuV5vXNHPzTXrIkN0zaZnkLsoxpuxaO2r5gav3J
zy9EYuoSfRv+FPxLBLVW/KygqHsW9faF4cYJlYvs/5i6Oa1Giz0sVd904zWmvhmj/SQyTZmFGPXf
gHbwB/Ibcz9i7/Dy7TRRlgN4tAHN2T7znSE2KhVIrYio1h/ZeT8vJ8Ppw7WN37BRKcdYqO7WSk0q
sG2TnbMK67xues1SmFWIqxalKo45BLI+l99abHMD5jIoea1511cpRii3lfF7lDpbxfUU4Ca3TqFD
k55lfdssGy993Z4FpcdfyjR/pLnwTXJva1PG4JJN6+g4FhF29xDo/QPVzqqV3L4SsqEo7PELX15i
zmEHX8DOXU79v3MI5KxP5L5RWlRqBZ5686p5HjqkK7BwSLh4D7jYWeXrNucmD7qfg3kF7i2/JkZe
YY39UudvxALicHl7nEFQ11f+CF7eJwLXN3NOwyE6J/3lugcJhLEqslLmcCroxvVSFWkUYAslSoHg
ReXG53S6o3yY3gRwxWDdYmvHR7NBkcrtSHnXyd1C6IUiyZrZtHBdFcocP26jeuspSj1IgDHHizcD
jBA79YDt1jxOKGuWB7bDoLZ+cZEJYwwPThiZ5pPorK5MY3RbpKSzN8HdEL7W2oxKz+wwZt5M33uc
5kwjvyZhzHlCT0seZ0Zz8Vs8E9gvvoogRwNB2l1ibCFlMagZV1XYab4sox7ZQOgKTTe1dy7wBfQO
68MVvnVpqoYMjbsFhzs+n+j/ewq1p2QkcJ2D2+yUwZ5fW59ssajU14hMOnvDZyRYirbphhDdQu6N
2ip91mKOx5hqrIsdIhi/XuosJ9Tnl/1NwRx5GMgBljaWwIrZxE7tVYrhr8mMXKMtJw5uWeyIOHJd
7sFQMulMni2SZfv2dAUe7vyY1Jd585rO3p+2fawHNLUEQYmwi1WmNC7aBU2KHQ+i0R6S3DzHjwz3
S24YxcaleZ6OGs7Hga1hChA1y+WtrzXGyAoTz9dEkS5FYnMh/J3Nrl4U69PRXDqVIS3w0bwMhdst
0JTUvia1m/fOGrd8R1h5fRCxJ7Podk/hREmNQpbqme5VT/mrfjvhlXQC0DzKFXaCvwiJXoRpSZ1r
J3inb1kVepaHfrXhLBHhTFV2NzH0C3RIRvTQAnhcmD0h2DJOyWd9u48XUY7ZfCBuY6mwPlDSVfeV
DqabBH/l7oEvZQm0HRwbnGKlhT92ChcHsBIULbHylohSLy5B5Ene6mk57DXG/FKwIIhdOPBg+h9g
tEgGSAk2LUc0LDiqD+qLtm5rP2ZmIzz9uJADFuASLcPbZeusx5s+l/X9JWGPTFNLiuI76T1Q1g5U
om0UCL4zJYzRG/OB/SCiUjMp7DV0NHUhDc7XDfJX3zH6a5rFsu9zTD/k+zH2CkiyZebIL0spCQ/M
g3l7jeUKI+ch0t0nVTzaopO5e9k/FWoZz09zJz58IRkWDd+m8ADAO14kegxq/NEJHyPe12DLv2xr
U92oDRWmcBopb+4Et5mvM8ew5Q8bCG8km3yeka42P5Wg9uyotn6wTJbrJLqzv98Vv1WQHR40RRE4
qoHs7xHdqIjmU+7nM2RsJ49L/5WQsSOexpzsiQ1+XaYQ7Tt4mEVFg24G6eOWMx/8jn3knYWlgT+C
khCDGBAmCZlogzNVGmNFS7T2tl58TXmGwOl3lCgOb+KHoA0l3NtKnI6dy9BQ9mb+3TEyhwmoP9qo
aIho9mQ1iQJpgocVNL6voHzQf9nNV2wPg8cphS4GvLU6YkfJtmMHWRgHzaDx8+NJb1YDBcR7zqHU
6vjZIbwwkB5YRdTclaSg6LgBHtNSEhoasv+ONzzSsX0+ZgIRWhbhhi6BbQm47vBjbFL6nfzRCjzU
R+9QHsRVt/b05G/4J3gJp8iVMYaM/hP9eRMgYxYNG4JQ8BkHL/GQu/SiIfq+YrSIsVLmty/X7i47
/iyT1Er9K+5DGlnKcVjWBPVS302pnVQ1EA24PsIoSGRWv2lIVNbJTMwsf+9anjgKk/TsYp6/peGB
iqw9p9AfmzW1xLXfO90PA+76/nc1f4WLOuAWnN+n4MNNLzLOkYP3NPkOLzZG/rOpy7c42ummd5Qn
14CHsQhkOzqCS11PeodHoMZ02rLp1P66U5vHfoZOKFfge60J8tJ0M3WI9HbBtwaHsvPg/I3tD/qk
SdlnYcgNrRMZPNBNR1gfVRcAG9da1TnupLIYDx2DWk7WCy8ugH2SCy9cnHE0pSqD5KcVSPUjpS8S
mpJummNfhcemg9TFenK21S78SENlk6T4IofJaKur/WVoH9y7HOj44n65TIVMSE5se5fKVI3mw8WV
ovyvUC6G2mzFeVSj69PVK8tiTVedeSwJ3vxEvT9MOaAFxz9SRrugZK99czxbr1zW4w49gJ6mGB2G
7k6pzr2Q56tDojrKYE9aTzBdFObyCUWEqqVd6PGriOc92uFxp4WLrCCeDpbCw6MceiWuqoBSi2wh
6CW3UMau7IpjWYwNBNeoEQxwr+p/3lIlfMI+8C4lxK5XDcduNPBZKqZYtX6RpquzqngjmawXtwmm
VsG7TQGCbyeqWkJ15iLM+o/wh4b0RaCcPqUSoZHSZ9u1aAy72wUgGehhxgkCGH+iTx+GYRCcX4Ub
SkWoG72J/z2vVdHaONiMwmWg91vHJoQgaoXRyq5DayRgms89XL7gth5kB49S1dTbr1QS198r22X5
hgNlkWx8EvRn59Wx/S9ZMnnRZwqyDgrKCRG3HiFBcuA69GcXsMAkgZNDO7RQPmVrT0hABXd883RS
2x2lYizLDqBqPASs4tYJ1ifFjGAWsdzEN5neU1CJBSrS9dVS735JE1pVvTSugFTFxs2XwCwj+jUT
z0I/RSqHRQbaFKNaA7ItYm0sKNJ8TE6qqXumeKLHpE/pPTAjfk0dZQIFryCpHNCV+dQIlRCx/7kG
g8Jzf8lIwv3azg+lXvuV4z86Bbh4MYN7M/biUwKtVlYj5oakD6LdV3y3Eij6e/eMXF2oDVrG2IBS
aq2BDqmMSgivIVK4E3LswXmWBgUtCIQLdwjGZ9OcEead689ITZ1pHAHqmG/gYT/5AtSlhnHA5zXe
hI3uN8h9+lbmFTlyuYRFMASQJ3r3s2LUWoZXNGKUx2BdaNyAQTB43RAb24+PYbwhkq711uf/u5Cr
AjqbS19HRR60gkDL68o/69rs5PfLHZ+JR28/aI68oLzMyl4EXjpvuTNFG7VLlsAw5jPS7gswKZlb
6So0DWRfwUBHRkxI9i7ZIKcH4XB9Dw5dT5AQJ1ES+SyiDSmEWF/4rFN5E7c/VHAuBmEd2tD3bqJf
UVVwROdJNIwiaQSuLaIyUxxHMjytdkHnoGGtW4r67gDDHQCZ97gID8eJhDel6NIHKOHoHosc+A/Y
2jgYcuImE6XTnVVmlFL4Xm9GSDOiCJ8qwtWrE5pU+brgXC6HzkJHTRgpuJy+YfKJKW/Fb8yY89Ul
JpqNJP6gebfXvi9ZmQlXALVN1Hq3Z34TnMoPd3nROKUWnpFHYfOCIwipSDSj/+eP0JCT0EUykk+W
xC45OvoJEvt8MnV7RC2euIUjQytI+kbAnJfFw4WTXwdZuoPxDO2vYAr+F02xV6CZ5Mi7tiaU5a0t
hlzFKtDlXtO7L9xmo1rn0MK8QtA9+GYHmyWdLs0hYtKtF2RUwDpVaITVZ8LWe8ra7MK8WjcdqXVI
X/RcnU/u/MdQwEkp3OyBDRccAxQjTlhjrYMCIeCSxa5x6CVwm1H4OUf+XnYegdelftc3zoy44HdF
NqRl9qQPLI1f6aIloPr0kA1tuZvLxurPrKkDcjW9e16aL+XB05DdK8UgtWqrtew3dtiuhVRgHssD
v00rAZyywiQ8NpJZej9TrJFYclzrLlxmSAfjlmCa0OwgyWwLTHm6WePyIx/XyBzxkUyKRcd2288W
o59H56FRZ3Eg0Rf0SksjdmGfYJfkwqhJ5YZgN9e1cIfIwiAsvbkE+w58kPlNN6seOpyw2TRhk/4s
SnfsT0SavGbS3aNmIh/9TJlA3omNNO/HG8RCpPz9KhPV0ge2dpl/DB//oNvdTYwYiQAMz6iF/8qn
Yi3G1g6Vx8yMxqfqJK8BWjdpqqzAr7aC0/Jiv6IpVT1cgJ/NwyrVMXH17O5ubQnArtgQ+3nkC2JA
xdKThjYk6FtUQAHZVpfXqpAF9Hwzuvviv9jnHwXLUQ9h5+0jZJvKD4pOm9bT8P5fxiv5zysiwA00
RDLjLArx8yQmymYOWN2ZbzW6MqIRL1QUgfa2LDjz5guv51h2xmSZoVL6dxy4iTQbiw/MXH3q0rEJ
wGn3lyRrUQWzOBDXFaoJQ4SiGQP51UKWKqdY9hMvuA8lvR8fWNydBzJ1jv9K41+sf3GTkFCfz6Q1
DGXYIqS2FMmEtWaz2t4H7UqgQKa/ddv8WVdX6Vw/wzZ6RAi2Iz4Au/4twDJni+CyLLNGnbd4eb8P
kCjW8dlPTPVs/KmwmImUvedQpw9OjJe7QNj2+zF+80efJTMtR7zr2nN3Ud94F0js4shAB5E09JpK
O4WUA20+z28Ku/juynk4sDMFRLEfxdUx2GmvCj3Y19lVR0oXkEu3CeNv2GoXNZHsHKUACO/VEN4G
kpUHD7JpxkHCzB1aaYq3+jYIT+07k3iBsUWVjR6oSUFcLTeveKu7eOzPIcuhsjP2t3snx++HPZJ/
H2hrwbARbJL0tP62P2/nwUf7f669MpDBQUkj20feWMg2dEOsczCZWiFtaAClA+4gezW/vbrZHbOp
gYlvlA6l46G/5HVnL62waTb6qJFTQEmB/QTaAf9sgPdE8PLxlBC0G6OCHScnldN61mXt5meHebjy
vov0/BvnZPEI+MFcAKEPh/nCTG33aYN+/KaNeTgrtcKN1+Av9HU7t9lmbtB1ujxkS9ytf5JieTA4
rtBRalZX3Kmlz/x9peDn7UxoSkJ4FaWRJDMEPRVDvtMPxuxYtGLjiM09Cl+dbAInKE2kRQfM5Ki9
CgQ9+sI8t8p4K53e+DaaKtoiOQVDzZgZuS+cnwGXDXWQHCnZEkmpbSPbEma7jIH0HdDybtnICkLt
87FBqrLUbKeQ+3BtzIobG6YR3/ruH/0Sygq4KB7c1G6bjqPVSDhvp2N2S/tCS1f2EmmdxIZBEO+5
Ozc2PtrcmeUqcxhidhYpyXF2y2apQmb0GBtt+MkxYEJaYP/41Hnb5yVEEaE7VVdNh1seXW6+eT+A
mktLsSrlpiEMaI5SI/rBCPgFyhhN/lnM2HhV32qcYdVEeBzJPzLjJIgm/B4NSscFH0UW1jDKFwH2
q4hV2k8DkymRkqQim/Ur2Jt/WKbjZygkOwWiXoTfP/65/bKLE8b4+1BMNQ4ZohGU4aMxSTe+7JQ8
IfELRpyNQg5sSAWkBuWLHzgQ8HMTj/JZ5+8I8od2RlYnUymDflDAOGu0hoZSBmXG2FpzjsAXsE8i
s05kp0HZ+0M0M2O4nuZGnbEu25Jmp5NzijX1XBpPIDNzFZ94CiqLBfdU1V7VWdJdRnNdwH5aX+rw
7P1qZvkraKSUCUffNPabx6KgRuuWpRggoyvKBHlTTsmEdybQoQYTn1e8hJK/437L8G8tz/BOPNZS
TLyJTW3NjstVcU6lqSs8av/75xPNsrIJJYi6hhtXowOlNQxVV4BvBmCWv6VdfS6wjwbkdVZrh+aB
aRsstleIW+Vth9pn1tx5h97lovCazVaO097VH/6C6pR1kdDupOJ5CNjj/pTc7YlCYVLJzLTLXff6
3Oa/bjy1iPzuH7VfHYdWVkDNtJoMDhzAzvPmLqUR0v30yfCV7CiG0zCmGrFnEyooUCip+pWNrdbr
XgpdFqx4KN89F2azeIKlH/0xEIj/t1lrwRiLfxDGzS2dMJUvjabk7TOTp9rTEsaPoQmqVa2kHxAS
EdkJi21DwyrPRH+ytCOl7c9ZImdYEDZ9c+9ehDnKNX/OkBiLuP9PXUuHmuCb5y3lKg3Q/o/kMcDC
KFI0FIFmEcN01RsL5Q9XTHUMoutnou1g72OM5EvPRyasvfU37JWARAZ+Bhiq9+ZcpJ3IHAcPwjwY
GQ3FwXcFUBRQnpnat7cKoVPaTGLZzhBcz33fB0HjT+TdTc4SDpBBqPDBja0Cd0I8suZ7Fx3umeeu
ELGdy3+pzGiaC3jAl6w+lx9m2yTEwH8sUz3hSwn9+/Nw//Uag78n08oQ4L/MjTd8UG9Cb1/ykhN6
60Xlb9ruEohtS8XT5C9Ul0nsq1QkeLlpTfxLwFGpGLB3L/VKjdrKIbTmwwCBaNUBoYjLkt7EdHwb
P5AaAgZMk+8eDvCS59mIAmpVTEN5s1xaDX4mzNHr5MltucfvBAWCVKHLYnScQpjveromp52DSj9K
Qa6pAqf5wD6nzvUqTwj3h43Cn0ZeTs/wDV1uvz33db4B/J/Ep0C2I9y9y8a4erlrWpEnKNzNk6wT
8p6qydWNE56D/wEzL6HDHKsQUR/a9Py8TlMh7HkVeLR22H27ZzLTolxypOY55+idWqZK4gcmj5vJ
M6AUJJQTrRk0c0KEhIb2V2o/L6+EZhJKChgiGFmg3tubQkBB/nxRTcncUvjeYxgJzSEa5Ds9E07g
KJF5eHsvTKHeUoSROEoWLD/3ZU7g/b8ILj4Qd2HupAwdOL/T5GvVbw29/ggqpGLCHxIyP6vFxQoX
UzGSpiZico0Lo2IMkddg0RG7KQK2p8tvbSs10wN2mHUv7yDJdqi0l80hUbfp8BiZkaVsneEymynD
B7/0BYo17Cught4XuxqpTljJo9cS48g9koh/7qzhlj3i+NgdDwqme+RAbmnMyRxJQ01mrJtHezjU
WtfnX3RAjHmkCxzD6KSUsug8ZIgIndxlyFTFug6isBeycDgU5ANfYwMFJRM3E+5MaEBN1xAovUje
fzrqt4dKgkdylGMn7/diVrvECn+vR1/F2DwjSbXo4xJWoPum9M5RdV/EYYdwmMnuKxnn1+0D5V12
2r3kzvNTToGHk0FjF2w0l1UDIjF65vPwIcIlUtDwXHgfA+l1HhuyL1qJMMiFC8HXP28djxeGnrGp
U0DHjZNdRFusTgotBHHYxCtPnq3NP+i0VSyW8hKMiqcmGKVMmJELnvnhtrBOYRsmu6lF/4+K9/5Y
f7oDY8IbPCKNqPsyx1M7xTgnAMlzaMgNtc7VkQuhqNpkgmpkzd8zmUWbaIHCuw12Eqy8rjqdbO4S
AaR6hsonLISGmCcVkWt/0gYGRUfV4vhFPkTFf9IegbAt0jXwcSf1Kj8DiK6ERQEloLg2pJ5/3S2s
FasqdJPHen1h7MkmPEeyw62Vhe0wMnpQXCHmPx5MuJsvIJGGe89OV4kGinygqqiQ3FnrBG8FctPq
RHH728KYcxRAY2MJf+NXcqhhPZ/zs2tpWOuvKHHgttTxUGX4gZskkeSJtet8/BFEMvKON9b6aMQl
1Rk2iyGiXBtIT4gA8c6CXJ7xVtUtxFw0dVT5wfbIYa277Jbg3ViqH4aFZNdt9IPIjyO9AvQ7h/oY
Nb9daQGfngPVAlzpBJXo2tvh2u/0NRcOvHN5yFbDd5g0yAiZw0nEo/1wwWa0pX9JfYppUeoUURG1
IBTIOTEbCmJcaVky+iz+Yi4GJ8LHZALxrDZl7011B0xjD8jzS+1zgDEIZmjOiL/tfv5BIn73cLtS
WUpHq+/LQyVxM3a13qX2mHkHAjgXfntm6lUS+t5KHyb6Jm5ndBNui67cWZoPOAkq70pWUFtT3uit
MjpCZen9vE/ZTn+OPxDiqy4b87kavnTAQQj/ECeDP/K8+yf54iw7fDTNYFJ/bZcBzX9t3CgfMjG3
bwHjMGwe7UW7q1xoy5G1jvUqirQRbJ5VKySHh1QV5pmJBnJaLoqKZ/KD7bMh2b1Udvu8sYNTtv05
/+NOXRRpPBZ+5AzbsN2kB/eY/vmd5sTphJQ7zopyynVMBVaAwRs9tTBfw/aS4gguGGImLTcjUTpo
CYjVlQhl7cnjjRRSVrDZPc8GIdFcJ2pT1azwGEXjC9jBMx4UMMjkSsDNfNQ9UpmXKdeaBAABFmwD
7b2eXXR6LQcQMb5Z57wKg/6oWvp9trZb7NX3JKXaafM9vabTpJNClSHD3KUC/lCZPH8F0VTBkSL2
w7ndTG70wt35evr+7i/iBd9rwFnph6foGQZMMzlXWVC4wz+aPd+BG36Tw2HnlWYvueJnAkwUFxTR
VbWB535jwGtma4rnYrohefLoD+zb29dxnIbwR9oOeZXJKhWCPMtZaIA9hfMe9feJCF/7wbjb4jgb
N+6GuR20j5b7+HkEXHQ1dv4f5ifcMBDlyXcNHFwJCSfNT0Yo4v9QPQk1hmvXMDeDJLESpAmlPlHv
vnGliX7aO1HTwNFhHJkFCHXCU5Wt70xWSKZqefZ8o3siWJNN8O73pHqFaRSSGXCd7nZK29s0FbHQ
BC5FNm8NfCKANOIH0ylBEsOe2kL3ouEcne+Sdi3gnbaEEjY8EL13GL0X311gGrNwTVb29PqJqC8o
ExBRz546tR+wDZHCvA7z71XICtsyIC2vVIicrFs4DPwmeP5g+NURmkIfQ/lqRk2z2PmywXWajCd0
t8RtoQ2jYZYM1xyKWL2nD4i+owvatmJDXandvgzTfozWmUyq2BqpVP2RixcgDAGd53d9RMGDqmmY
ZoxlOIPo4+jCCulvC2BOvUdZNNKc5joUx94H180dyC9kCemvvy510724XGVYQzsS0VWi37RJ/RN9
gZY2DrNEdE6DJjwO+fTpsu/Jg24ZlCFEpgwKMgF3OP3/jlsBaIejEbyJNQsBHjoKSfb9fIgz37KJ
l5K3Ge+vPubK9hkYqy1jlekQoScbMeoVf2t4dotY2FZhZ/r6CXT0S+dlNcqVkFzoYyQU5RAjg4O5
LeseTuMUFjXAzNJEeydPGthoQL2DXYdYe9YqArnsXuX2CM2A+ilcCc5KZ2rP/VkW8AN3wBJ4WFB2
kNX0I++VE3b+vXMLIYE3oXzMG+pdl0/DTM9al1Oc3bxA0kS4eTL2PrWYKhx1mgjX7eV5ManNy6Uk
Bz871qlWcJDgj7M9OIJbxk8tuz42kjqrAz1pVv9vf6cpSgNBiCS7tIgQ2B14Lc7Chlo2y3ckEzP8
D7tiVjrOL2gx7JdMmhIMc+JbUgikaXt2cu4qm9ALpIfq5dLumCwHc0EujO9mo/dG+XirgvXFsTe8
krKmhB8cqIYSDQhj4jEbK+TFFwMiJRmgvISjy7dxzWwb2AhJUmEuKe06c1neS8DZ/p3OZiKvnvej
xLzgTrHGr3eWwWDHtG70m7Ocy4c6HET/UqzpjF9eR117SSRl8ClXNU7ZWdKqZvzaJV/JCKSylaub
nC2P+kdGQ86+45BNneGt+EQMook4VjT/6e9EurZzu/S8YYowg2uYcdNz09ygEs56WdTSO0PYrPL+
EQnX2ZhtQuc1id17S5GXfjapvWsaUZJ4xg7V6L395jXFRwhiD2s/rn6Ud2AKOKMqziMeLwxYgGjJ
ChFhRHWJfoD9BpStGMVwUHE5TtGB3vaGRpbScbyfF3r61n6JIeE4RUqTZ6/ggR9vS/3ct2O1x8BO
x2nkiKRr7aSTGUvBDp0ZqF9EzfViswMRfv9b9WJoNqwJioCcPlWR8hCbaUWIvY7FtjER5JQbL8do
wuSiJz+2qYgwwygeIyFIF1RuhL/slL4O+2KF51cG2KxRc1FbR0LbWvJ15ASjIybHIFvkoETS6I+O
UIEWa6XKOrnFuKZcaVwThasxQfYOZ/qyYt2mK8+hiXV5IoK8Sgk2oGBXyVv8d1hMYNJHbgXOzX4s
cjkYTKbCTbhEAuAlGQmW7u2KMja4R4eHKcIG0R3T7EixiE7IJEJE2+kVJjB3wDz5fV9jGHcoK0xc
r165kCwJXWdYSICdfcNhRK8BKSdE/WQ41MFhWv83D9OfC5piN9Rk7Dcmitx4TO2N9QYVr0MzeTSr
PXJrAMLzGV+2R4W6ALRyZkXQ9Drs2iDEH1pM0K0xLofQcma03Q5kbWsY8p5vGrEQ47evHd44Tat1
CkdLSp2X/OMkYofGs1lLGMbNSGunKxRPRgSHXmjmbrjq0i/aS/+iik7YXjQEzeQRFIxsyAsWqesd
NGR/TGXESXYhtg43oUeJXqG8v5nORf/Qn12QCKMx5yPhv9mORfqiTod8m2qgHRAcpLo8AGdc6fRq
DlFO4tWumr/BW6eHekqUk2b5XfYGQbNFcSgJnqaWrL6orKBbf95mU5yzrv1jb4u/VCivVUScZwhn
WjetJDUIsTevvDvvNooQGJFNJ0Ixao/+tznb7R3iaZLeHdnPYQ2ODxRNjIbWGb3JNtOA7oBD3nTR
h9Y5zI+bzymQjmD9Q4p4l3OPRKJ73PwCSaCH4euj4lnLrai+vujC/wff+Xru6r/YIcJy6V2TbH6u
DuGTQpg0CQbHH85Ar7exUU2sRZGQkuUvflhYliQp43iJfW9V3ZghZSW+ZneghhT/GiKlHpSOJw+l
TbAV358xPvLij6E2e4GlaN82eGhXgdLU0eOwl/ffbyQmqk5c2yQ1KqEYTXIQ5Do8caErnnYEpL/m
x3GRybIiAiCS5lyDUWvCS/eHX2kSmW9Jcfuj+prAifJdr4vrTdAbeXzv+qwbFQoR4+PkLy12YuV/
8o2foZ4gTJWb9t/bpQViovJKt2B7/4ZoELbTGOtnDMS/sn5ZsjFi2eYfX0jIotY/xRaJM+jZpuOj
IY2D6ErXWh4ljL0vZXublt2jXT3FxronmcoCFXpT8SJC3uNUuR5cg2RUOkFMqG33ol9PzkrYRZD3
tfhNWTuYJ898GPHjm/RluS2aVpGcCGIgiDZXIhN0Z4v3LOnFuCyVKurvp7YlGmLG5q9rB0Vz2Z9K
3t/K9/DD6P92RRnntwwbrQbVIPY93OAyADK4s5+PeohIRv5D8B0N+AR8jKIk26TlT2hnY2DL2n/6
mkwK4K2Q8JwI6M6u3sNqBaQZ77if54q8Jv4wGam9laIuLNifjX9nBWBXR2UE15HJm9RnjvSKLHGB
EaQ42/kTVZEI9eXVjUTAdGAooz0yWUEk+FnnLf7EZHGidUsfPzLoD4rRKDX9GWAAdXh8CmlhXqPH
cSx+gpep/J894dhOmLLK+DPRSPcYOtoK7YySBIu6ztSP31dhF3WGAkDrHsc0VwzpTS4Pa4c+Dh+s
0ZM0Yk/NqsCSbijFijHGNcgYibkegQjL1NxEKLMnhnz85XycRJeFZ8YfBxh1WQIZfRrqP/Ht9YRT
pT/0F8vPr9NhGLKZ0kMfOxU7fe1Zra+S8IJMYvSObL4Jrl6goZHpL0/8q7P9UoQ8FQfZo1iLeqlB
iYoRLAkEbOtlPLPqfA6ffeoZTv3dFplf9jqfV5nvUcRcUQagVRcYgAR8CDbqay+4CABG4a9mEBsE
lKTwpgdJW31P8j0zV5owxHn6hsV/a0QsC1kbr7AEgYYOghTUnrcPyUvRuHRh7GuzPftSay1F6zus
Y8R5BlekOqtLkZrxmM7GCCrQ9nEUhudcPt2Z9R6+f8zPOcg08+cB0r0NrLLwwbzsgLh53Sn+cjg3
p6czq7PmJeKnoPID2YNr27KaSdkHgRXUItn07bprEJrOlHv6FQ+FSlui0kbdg2B09N2qA+lR2WeV
fbw8WeeV2GlW5SiH6GOTchyTzDLynHPwfLg3zPT0eBbLwAAmNfWJZfjOzgYFCwopA4W6iWLMY7gh
KV6akep0UJWYzNOgjkJ+J1AnkHN5qtuhZDsT0oOVBo9008b3AsSzF2en3F3hrYyC6lDihIShJV2H
gngvhQL7v+l7itniCxx9eiQ9weasceweIoyMgZpInkZ6ES3BfFPNDpbG2yY9H0ZVfg05Dd+0Dy2x
Og7a92QXqG7VEEO8AkQb1PmGYYSGSB3DeU/otaxX4OhRMii5I+CPTrtvUMzb/H0jmHWuyB25F223
NRuyFZbgmrcu46id/xk9RLY17zsBlPUObSM248zxY4sWYirzMMWlkt71d5idPGlKAfVcGna3iXIk
ZZz18wBXP1tEVFmTJlpFyupUoguHG2nEWNZgVl9OWEZKRIGgE+NFs4wzF4N3+vzXGl+3wAFehWLH
WJdzbvy8hl3AtPKg9J1i6KCovYKSxHbkul0Ibge9r1o9y9KUC2NZpMBAzKn50VAleG6rD1gDcXId
KZSvYQCLi1vdfgKCyaq385oks0NUpAlTDwgxAAJ2ieoKygnV4X1DiWEy/52dTnuvbLl2JI423xq6
EHxZ5rJkbiJWCFG5XK1qAEKtfSoYOEtbB1oPOqOtD5Cn3Xali4/Ll8XxKZriySnF9t70pIQkxZy+
/7kdrhBOtPo94heGVsk60dTGWP/Z8Olw/mUHG5lXs3cz8hPKtfxxlfFou65tdM3+kcT7p5KaD+xf
9Jv5AqQOSHcG8//IScAuvavbGj4auZSves/Tgoxz0IHL2eRqaqBfq/1R1DfHbYE1aocU4XsN450e
m4dP8pqPC0EV5SWl36HlW20DyNX1Xy8RzGVU6wg4JUYhBoYx8pyVkgyv+EuErncjhxJLFiLP0Vga
z8Mox3LLbDs+gfbVS/BsPXAT4vCgpPfYyrglDMQWEmxMqV9EqG5LnlqBfAIr78m3Y2i794/OKHHv
H85j95ff+sLLPtXMSzG5FsV5xweufJ6M7WLje6gCmknYSWa052++SI3ikjF1P1idNDXWKBy9dY/5
VNrWs1ZnKYnoDQP6AzZMg8UF3u7mvykZaSDFuvU4UwMnE5/ZgP5VQqsCNLGE5k2N2+H/ENL0yrZV
/A3cPbxEJWH5NjQweoSYQGqYWZTHQVznTKYsySKpLC3C192T9A7oNLPTy0GWuV95PZnz1Roh6hmd
MW645yLS1vouvj4USjZogWyQ+heB0pNcvM1RMlyTdtq2bynSJS4AQSg4lNuJpVVFghiXhGOByBYg
qV4Y8TwB3ofavG7G9N4jChvNnvZE9yysqPF7YoLq49bKaboE4RHM/U2xonqBuGgXjiRjbj5mccIe
lr3/2vt4JfPRIWsM7HrarPaxy9UvibeYZFsOU6o6HgSnZa8NieVGr85Rt6udI9/jv1JxmGxznoBy
r51YU7Gah3CVlVJ4m+YJQNvEy9l6JX7I6PBmgFLbSmtc5/JNmDE/0X6EnPbzBMoL2l0lfL+7EExy
5xDwIJmT+7qfIutTECI5FIkBtWaIhTkXlaSIxBSDwTDIC+AlRNcLkp7wSkVXFWo1scCZGB5Az0Md
6QrUGGqe8UmPJWyc5sB2FFUK0ZjPupT8G/s4PruNT4ifx1hlyZrilZt1V9I1KPgTjpSlr0F0F+IV
ljroaL3+hw5BXFDgmvoTS+/PJQpVZqX7cG1tywlm3ghVpBquTuR/Uuy92wpvtYntC6AHycbBu0jA
i5soO6tDhwBD2Sdo3H8GS70zxwfxlJaSTheK8ZFwTmG9gqaMvDWsTE8SzR9cLvr45LD2MG63qH81
mBJWROWiWX+NXpyTPhHRz0H7KiFxDlBynqD4Kdohi9vFgBjSIYyiscoPte9ePBaJx3HAxh8G+DTO
lhssagDqN9CGHaL4j2kB47XJ69SkhBUt2TMxs7x0TaQafWKM5SCgccrB4DllFMr4RCwvGrZfkqUc
deux1U0A79/1y1bQkMmzinrMDgxvmFq5UfY5oPNWl9sI3CuAFohLTwg34wyjZ7Ko1/yfMUr5Qzzb
ltE648gjzrjrrODqHvPqpjb2kiFtbUmqpxJherT5nzlK4rbYou6ALckHPBW6M7rQ2IGPLyVNhEbU
Vp6U9fYwaCPbNOtjOhXCXZy0oUuYdO2H6nnY4l38hcID2TkIQ/QxYBIIc1fB03LG+SdbNH6rB4d7
8Ueb+Ljl6p/i2ZjcSyD1jILa/clW2cZs6zdM85GRumDKZ20CYhm11r4JHCpcFDP60l4o4qrMLtZx
xeFiG2c5HQaCg0u8PUGKrjKpkv7luf/tQjkI7uaWMAI5d2h1VhAadypKPjlsrAGFJeLVHMO1mI2D
Sq2vAr9x0ooa4pk4EbfR0jdwFrDN2m1SEhFMsH0mon2X3LhSFyA646RyBJcz9P0lNdCoCiRy49X0
3Kb2dDK/L/cGDH2u3eoCvRj1mmFGPgk390ON9hZF3cBNlpkxQHj40tEYyYaMet3xiFwdkjuQZ50c
OfZJnnXmvqxeKqmDqfAildYBnOK42y6aM+7I/93+DSvpEz0hqtPc1tsvUN95r/0oWgNvASpGlBnM
9LOKkly54PCYfTiV14jlPbm0cC5XCNxblds0GC/dLo51lc/DXPIZ3uCZcAtN++liNm1JzJGFLJaD
DX80HlMWKYxMPXua7ah8YQGH3DgEEwbqxHg0rj5ZER25balJKKMIfnPhGAjGfWzHOorsotVscSgl
LTxh7UmaaPyN2hECeZD89ouoE9zNWagYlG+zHL1jP8hBs3Heky7Oqna43kIekut+Jv1LSijpYpg0
eFgTgcB6yO2I0KlssGxgcSkUqEfOs8o5CqSBIMAkuTLJwQxoJ6a9ZWSZbudHFee8f8/YD5eLe81o
8EACw5ttqpep6EaFUbj5wk/4p3EvcyCdqMWH33rpL+b8fVAUOBhzqNu574eoIiqeL4uPNiF7Taqc
/Wz9XJ+HJmYXpdU2BpgVpnLKfkZeNU6zKlHhy2AqmjQkVOMW7kQ2zo8z0siNBZlOvCeS13TiCOTt
3c9Q3RpjX0uaJlbLWuwa1N3hmxiBnY34fIiKSIxXxrxV+Q5JR6MfNSFkZVCcVAb4TaAcWjMOJ3cI
vgLRfc5nj4DnfMkQfhbjA27T7BsCZO5l3TM+8IbWur0pLQeYNLRdNLP6TglL6Z7cKOv4/iXzLda+
wbNlzjiW5fKSm/bjuTpZWgaa4eG+eM9RoMpNxkqLxyWEBMjpk5CdgXW+QmS56EMszjAFckshwGWM
dThV5VyxBGRAMVyKresPgqYW1ftq5yGjiufQBkeg8Rh8/sRvZZX+QS9XC3awh1yfwikeF1ZGjf1D
zocjCDEo8D+hBYfPA4KyCGRtO2nLi7zhEmlJIIqDrra7G2kwS+NAIQfnMJaR0MbgHPqbdrYQXjDY
oYEr+Enk5vm8glXM3oC2SMRCguqLpGAJnukJBjLVm5piWJpL5Lly3pNMAonkoIefBiCL3fPu1coR
qKPVhu++rcncdbFLOoBcLTglFeBkn/3Gt7V6aH0hO/bPeckmIl80nuHQui5XPl/DJPMy9Re/wEd4
D99Gc3iiMcTBbgsDE4glm9haTN5QcAbxrcVPyuQCSE0y9arjS8imvZUv/4WnmUu7lN3aN7Apukyv
ic3R2tfHdWQostX1lmaBQamzlkRor6DX8B3xdAT/tf4E/RO3SqBSYtA8tc2siP0gfgCybklVk8zd
3bmt8iQ8BthAkXc5YdhPplT9oYnkdIGVQ0+DQ2/vY0GGF99PNBybxqz/GFkbS38DhKml3+xHsVBK
yULFMvzKdD4I0V53dTOzW9OHvd+x9CXdf3Ud6tQTtKvgulUKJmpqrqEc0QxNusMLWyXRmTEDysYB
8PXq9KWT8TWpFggeZx2tDe5M3fgts6zfuSAtDkUAq7Lz4egz4IqzslsRal1ORXzr01YKp8wqVM8s
yGvi+/Rf6CPesuGKeT+z2NqkgVD7bm3Pcysu5ZyCdEs599YowsHqB1iOQDrOrasapDGV0zbSzKnX
slWlSW8U/JgRAbqLRTctvMcyPuMqG68MPUKSUjMJC/DTCzckfnjsMh+WgRNp+RPlhX2aFC3z3/Y9
GTMPZVyrLmy+4CN8xToSrXxdzlRw8S7t8ws9GN1yKEXdpjwdUxPwpbsixTPBj103WzEKteam+kVN
8F+4tp6rSnb969u9KS5I7GtUqgUXkorO5qvVMYcvEJPidlnt/K2r8BFH1yP6NkLSjC/LxAMoYL9J
ZrHEOZRLnRQgE5klvHoHbp5zKg4H9+nRyqmatzyEaxr0fyekDQvHdRnlWEN87+UDngX3S2FCrbXs
4Gt3RQ7CMLB5aJVWCoQKhH+iIa72uvJ61VP6OLTdPs0CP6xlWJEi69yBCFYkcwUtEaxhsbP7/fEU
ZuK+gXDzzSqrm3mrVszSVjUXR/bha9/H1QA328sEsJ591HasAbulJN/02xhFconhAvXGCW7X/aF+
IYl35Ac7L4+vWAMbGORqZvTDC48jCYjIYaxwGqb4giALSVjsGEg53Ta3/wrPZJE2pCNmcxsXRwjb
+xYBoLFflgpRot5gn2quOE1wwHvn+RhGV8kI3Dhbtdq114iA1wg0IF+pFcwxvK0QkQMCbKRZNKvA
fcb9uisTyxczke0kZG0KW6mwMOzPj0XB9Q6EYA5sERBcLF9K/7wXVISESmkE73i2DfLVDSBhqTPs
arV+PGFtiUbeR8CpZxAUZqUps1wvnlNub2EDSfJIcpQ1mHJIbp6y16368VisxVZ8xc/cHfLr0yF/
dvLUNGNnSvPX5xdbQ+rMrg5PEHPt9cOAkpraTRQqnA9V5qGNdxhqyod5juvcVQBJY/6owPJmpZXS
moqXaWhWTYkLgY31M060oLfsvaYtEH28EXdJhPQGQ2P2VA78ij1aeKzwcKmbA5Z+l5A8KvEQN2iR
g/7OFIiMKD2WBsMR8AAsLWhZR0s51PYGXNEd/puqvpyyvbzbfY7IzcrfGNUnSzzEbApNAvR2K6tC
9AIWgJifSX00Pf7HlEcsgQ/KGG1OtdShMZXTCl9fy0WhucO9YpNAFB7BbLkqn73TgzesfAkXoYDq
8refGr+50Tf1YCKeOpuyVHeJ95ZQiC7mGRJyt1oZnWhATi37xCsJttECbjUr4C3nqwHe/QqS3B9m
kVp4Zsjnvm1cBi55xyovizg1HtP8bTHyoF/bL8uI2pWPdAR+t4mbPqyvnifooQE7Kp2Aj+M5wR/F
h4Nx9WQH+80K8rk7kG1NVqd10q3oPKuk5C8liOrzfoKEZ4auUBgk+Dmi/+LejJJQ/moY5WoNbSt1
fK8EjaB3cq2mHQ3fm3zCqXD1Qbbdztvc2crPCzTOX6x3/uA5ysr37iSXqbJMHAxGe58pEgA+raQZ
Dz5GyFqLYirXNZcJD6o4hUhO/lJ+nqThSyI3w0fqqrxN93MQ+SaRnR/BhyqxJ/8ot3a/yqaCi7xA
6ka94sROmnZOQMXmqE7xqdMG/uLBJOdhlQmgT7uKJK3h+ztanXJ4ZOfYskcoVM9IgYnvngllC+Vp
69OUE8lDB21jdvRWdPP/Oq9wKyIC7gY+UF2CtybtSTO0H58M3Qe1ZGacCs+5wK2S9O9s8Fb4tFxY
9AF51yMLa7VmRFl2WEf9Iz4onZtp/O167SKfO2uLqEmpSnzBGHMoa83fS3lRTYyZF9NHpeS+rt1p
6S1FXHMldUuNFRYqLbgz0tlF35dP2kAH4EQALMBLVzSgM2VAOpUVrig3V78bI0x8r51Zf2kTOP7S
k/CiVCkqZweVVSjW4oqk0n1dVhp6l1cdRDKe+COe/xwwR/jgXhSo1WBmPhEgwFf+tjVhV3n1UFat
Xw+cnvU73LDcZVFbEU10N8f+QsW9iVv2o9+3S0LON7gwOT/KCrsWAVj5w9RbGXEnmWQHSrMZ5AWV
BiKHb5wWvmqYdacjeeyRjfut90NOrRF7wr3+DSN4Yn0rANDzaob6Q0/ilHoGBqoL4gN74yth+sQm
MCcRi6Hc+4JvBJG5L4srgBynKKyk5aOYIYHulNEYghP2rQSi5d9mQ1L/RsXXjbxnNdNMyG2K+ngU
7l5AVXXdpmMUEyDwUxbfBJu3RcJuHdhoahsMN5I4tBHK40dlZBupSElxgsmjKy0iyytc3uwqGv3d
zG7CXLnllpddWem9glJ5+O0p/Om1qowj1B2WXPgMUWDc1jA1XbFLOeBTf2cJDDYF4Wi8+sUJsV3E
sLgKF9U62oSyc0+xuYxJRUwgXApz4X0ijNJ4QR0XSDMe8Ck0J+ig6ez4hAhUEYWiNa7Bm/hkNl+7
Gvi8HXJqB0/db1ASv2jVBfaFPCrWVYwZ+cudNpDRkZxg9XQzcdC0vzULw6wWuWMgU3TTxarxJ6Kd
SMwns4CJJWB7aoivaqu7tqgYO7GayqCjUl1ZtCFYa8vLUWVb/ubr868SKw+MiTvHT8aFOUfxHcAS
584HIRtCfqK+rfFMVSLCEf2XPhKeJTZSXClj63YN0Fk42Sm0k7I4nBUK5cxAVyNnR1T+rsWeGS0r
YENuejpnrRut79iFHffMwBc5hhmT4pgs52a6LW+d0FEfkY/PgGzzWvV70sA8jA4shfo8v5SWq/XG
S+W4tOt41QBK9fT4JWvvimdW3d5F8f64OieFDnMfCCt+qNZ/bkFH5pJ7P0fYxTpLBtpy18ps48UH
/yTSaK3i4Y3VaN8ADYIcfzyryvlbgPXODDcOjr131R1PDA1IOJujUgO0YbkznS9IPcl9kzruhpHK
Bj0OsP/5kJJnLFo/vr5E0E3FA1AI5jhgJDYVbvTvvrQiIixUG0khvleIvQQC2hZL/l5mBqYLyeSS
/qIqbroxgrM6z5fegG7tY9fO5asPwL6x8eof8AhUpe6keprYxSG3Urpk7hEcQJ1JQUlybEm2fQxL
/2lJatSzNk4GngNe3ew2psmag3WbzasDhVV2JI34z9+eln1TtMtACMiKrvZcP0Vbe3oqRH9aY4ca
1oLOJZYENKyeki3mOYgyw91IABl5nqBWDdGPhR+6I8R1h/FHN7O75r1PWGxzppRw5JzOE8ADdbQ+
ETPA6YOFSfuFlOIlPXGklIIk2RlW753MsKzIkVX/LHD3Z4Cy5TW5r+matWlThK+MmrtrQJ4D5gxg
DrrVzdRxbGLwTABhfw9j01ufy8Gb89XILUPavMDsmmLtI99fXADT2b/uWPKtIcL/1tsz9/l5Qz4/
LNaE3Z7gbanu0k3PiAEisfi8lIrqxFxQRmBQ2dWQQY2OrvlorhfCzEhnj1PKB4rfKOpX5x8b6+PG
h69/y8Oqm6z26hhGIpfH4/AX9QB01oVPHtY+lzeWuvTaOQ3bKJpHX8iHxHtjAeP/YE9oQBYGEV8G
RbI1VzmNwiVjjekCZ1L1yQ7dZOfprY/3mUejFinhNmNvbNTp3VVMxlMC6AvAw12aUJWsy/cty2eG
enoktfNk6ley0ekM42RnyQHVoDTh6tt5r74Uwymf1pPt/Wsqux5G5PORsIQXeOPt0xrtAKNPvyMa
CeIgbpYOVVxyNwfkwKKfM0eud6NZWE6rsfuwbktAsOCNnCnxurMaSAb+twQ/I3Cld6n/vxXzN5Kx
6weqnvom6VljWy3GywC1TT0vgRnZFh0mK+/tEbdTAJu9ul7ZGrG8E36e4emuT85KiiSn455o9y8N
16OGyLOguTEFxhRFQYRvmjOTJET0THYa84cjNGJz4SIRiQVb8Cra/y99JZBPHdobUDsiG1Pp1gKy
XYHdWsWKUFEc9GSFO3i1GrLnzEJPuMOGWiAgWS0NLtV9sB5aIcg7uw4SthmvOqQUCewM0rccUMx/
HUNgL0cRbta2rpDBD5jyE6Pl3l4TmuOxWKydg3jXVH1QyclTrmuzNbe5CkP8s6kWeboHL3EJwhPv
ekjeCBQmHj7wQp91chkrSEz1yvXcP/wCNigSlR6+qnp/YYppjbq0RKN60rVXGIxohrMOJfBuBJET
6nhAhHBqjTpjdl161haYhFXxyophUZE4+cGZiGllZLixC7FAfV+etnUTekZqPZuY7psau0rtzjB2
XtscdLtQNmn4JRTlVHrzR2yrmQAhTFBTuZPiH6QJx0U7KoYyEfubX+56984AY5tsCiHGWE0bW2cx
uNCbKRKj/PiyEVKCNTTd5ThcNdmSdtvwcsl9spuRT95hFkQns64u1RS1gMGFBpiXl7cViJxb2fW5
GV6IpF8pNFTXya44Etbv35047SwCihmCq7/Cdvt6QMwMmLA1LRhgFWg+aYhE8CvJix27bOFccmBz
WplhPFJRwgm02TkmHhrAzIHARIJuE6lJV9S/7evbtgUWeMsVhUdRk5c9gSsR0njhaoepzIvP8ZP5
qEXFIllQkdtcd3+u2TGTbuDIDd+H3IckJ/L/ldpp+ETiQPbBrv8zVZk0eL54X10tvIaByz69nm6c
6ok//NXENPKsc/QrIuO9UMhuJ6JxV+jv3GdOpLWQswkH30Sr1Pp6PZNEl0B8LfQxfRAvkKce11nR
txS/+S5j2f2d2BAal68tnRFXC8mtG2vGxRj/McxE87hdn8XchcaRPWXL/iLNpuTemNil1abeE+56
NIsQzW/A1Bd697F7cQGHPAb+iXDhl3Fvndm+u8uuXt6U3RfbjSCUNY2JsAQK4RasRzNmw5B7J6Ui
UHq9VjPOmOravI6lGg2hZZoEHG2gCT/b1y31TEsFJ1NCaBeFltATfc+dm5kOWvVgbEzouQnevuOx
wO3Xl9MxzQJyB+gkn8NXuM2mqlZJcd7sofhFHiJK9iE+gqOgyIRPFJjoKwAUkTSCPE3kUT7PWdT5
jFjjlLw3wEO97tuwlGqhZ9xo6SqmHppHwX8gGK6thhA0J8txMV2IcasOo3n/wEAMDXQs+ukTcLNp
dqf9AWvGO0p0hcop7azrWjM3D1RS/fclp7Z9sSxGocLPXZ0etKz6O8FHZrg/wdujY2rd+uj3W8A1
LZF2JKSf8587ISdfrq9iR1VlQR+SpH3PddMUIwVOA/Sc21d2mFrpB62CvKrMcg7l3U9x7/XwOQXH
Z+dlSCRcZnI9SVEoDWhJorr5LYoWiXBE3j+44+hwJuhNIhXhVcAiXTdOlJZWqJUcf8VLUbszPFxL
ZWHK2M9w87cfqiRP2we7FUiCqVsgayjS9SOwRB7ppoTIV7h7/GYKtd5GdrMFHYrFarat6X7Ecg9j
j9DRuPrWQ+aW0TleDZNhRN5kFNPA/iXSQBYl9sL7VrVQO+u9EVvjgSW/aHysr4IBMlHaUgihiN9m
GVNF34jEa24m9MjeSizudjDSH+Z9fIOGGrepUVsoe/0UmoD67IWIJ86BT3jCnn4Sl3fKg2UCImhd
Aw3nk/e+jDemaI2HI0NGvML3RRosu08Zj+NBWdjnba9zmko8K4TyfhC3vhImibuMmvoRjg7r8/jZ
3OCV/V+FhhSrWcpWeg7S2P33LAcif9s05EHfDLONRjWkwh8/bR54SGgF4leYyIIdrcpLZap+56iJ
xlhZzN2+c+fmm+ZVJIMpCWXPTzeNQTQ49HGWbs1FYnTulaq3mNy10QI2OhjPN/EM6o62YnimS11M
1G9Za1DgkXO5mMYYAI4Tfc+JuyjYArLlZV7AxvB+xGo+znuUghHuDE1K/aDslyC3BTwoiVeGAsqJ
ikBuJH5OVeDUXGgBUxL+buRGbcmvr+52mRUaK/gCIZDeserpi/GRc90TzrDfES38M4z/v7QwNsBc
sw5N8VNr/H8DtNkAoDvrQHk3VpPqMboTt2Q2zdplhDENzar4C460QMMQI4RSfeOlWhLbpQPovs7S
5i+kS7n2cl2SjdjyDYJFc6Y2GIAByUcEjcyVrPGfaWJsA3EkgEKyXrdF9GZMOzy6BFgoOJwMiLjn
B6qtiki7ge5AKyS4rRYqattpUtq4GHLDbYIsbYTpmR4u4ooEUX1dNDxhs8WHi3nfLXVzQ7bn/2lP
L47O+Ja4548KPFeH4Si0SMyU9LX1vd03WL/t03z072SqbGaPNLYFNJRpu5znpjSJktNwVMxJyCjB
rm4I8wvlZtBmknzjuGI5mHcor+g0BiY2US/+J/pufNCjZCfmH/mARq1+QIQyGb8P4zHvtaRTMXwU
dRM9qVz0OGRujp98i9abe0vdms1PeHTRLwVOC9EXjDrz+L6Pil8svra8SBhbRSjdVjKMPy35QFFz
kyM6uu05c90UucENOiP5ymIJ8cDKz9nroz8UVgJYycfFq1RokbYS3U1iwzMTL6cPcX869L/MxXSd
V0Nkjh5d79Z22daShEQSRBHd0zruwo7tkAopaM60EDI4anxtBx5WiLwb/9QWJKFGPHoGKsLQECSA
gO5ucEtKPMWKedZo2CkLg3ZOaettDrSPLUAZc4pP22PknRTlJFJNGC4XAXdGuwEGpcn/1mDW+EfG
873/Lf3mXqujVoOPGomWDd9gyqVx7uXwnV25lFCGhAUbnNLwJHXA6//EzFNsp/K8NQX4xiHliyWh
iSRggsliGnhY8kXlSktNtLmOuF7TKUYUpvVlTOt3lLw0fP5tzl+LbXeEEUQToW29v29jHYB/8ZMA
JbZnty97llpeuqAGVDD0YtZ0Ad8H7P2zvC+Vpwh9IznG3+WJKuqn9gTmuUiTHhp6OuL5Z7sjk+n/
mxy6fzmHz6eZUCdc9KGuVCOsLq3dMkvfhhWCMCjPImUuu8UImHbuOINz8+2QimIeCHi/KBJFxhoD
1SE132v9MhcZBIfvUvZ0tnNGjC4VrN37TbQz3ezMcCi0l0y0EvzN9CgeoE7IwqsHWuHHnTc0pRk2
UuefJidK8dm/VpzUh99c4CCgI32zvXX+9dFp8ulgO/N4vfvQgW9sh2skExWu9DJ2e3Iq17YlisAJ
AZnghuxiHeiW1xiiNkW2qLbaTg7OAkZ/c61ywQ9xMpDqX1Iui9T0XAXO4AkHJptuDo+6LCeXfQM7
/p7PDpFzdxANxeLXxrCdy29X5ILIBa0mS2es2tArxg+4WjyAR0d5lRyGTGTkpI7i0E8BkxCEy3M9
HmwSfwC0RroUzEyeccyDG6M6j030vNbuSuLd36wb2woc2Y+++ieS1PSjJjq8LDvY7vRsoTR+0Fj8
wjNy36UbRVO9BM6rYh5nhELIXjPK57f2R+eAcLpy0cPQ99sszb7Tq4odeL0yxXd7mOW5ZlHwOEUC
NMkD1y9qPBDcJxg7JP5d8eEcYwzLEoSh80f4BfDxIAIt+TWtqe6/v2VlhsX/woUR2l/3cjgXiipr
fd+AD2i5h60waxGX7j7dqj4z4ELtT6wIc6RBNn1SdBgGLJ0+Uj0JGnKDy6BvYqZlVUftVJ7zvZqs
2puQeUdZhyBd6MbXmIPZXMCJ3L7frSj06ZXmNcAlEw7BElXGukpy9Rn7oCdmtLDQnOx9jHohjNzF
UGNlT1ISgNFy8YwIn1EnLpSk5abciLsF0qetx/AksxPqZzFIUI/orNRHZzmh30TMsw0GDHc5vo/B
sde8KzIwadQVF9+vbi8q9+xlCdRKLznLJ/CIk3KxBceSy7pVaxFdtfyZdnikfbbdCcDxVM/NVbVO
/XNPIKPeK0uhMWRJpoVgwBKq85VXxk94oXj3BjDk0P6mn9l05Y7ip/imfMFTBLQ9ja2k7AVb5Vwt
d1LNrtvhZTzfZZn2fo7np2B5hW5eXc3OVmJ1zjT/STxkCcZWrlJaEl7EF+PIA5172QvAEFCRYvfU
KPV8LNodboA/8G3LZRDLvpUVclWtuhsUETFrlf+IGcfemSxRNx07jfmlW1grejVlQP/pWBmDW276
kQuTZPRKo4zPeXpOic0KARg8F82ilTAYjf5jSkCSBLdI691/K7lG19ppVfDy36w7hrkJoLCf4hpy
MTymqRwf3NvYzGJjUw39oM98eqpV2QQ+qRfLyG5KvxGbfliHm7E0YI0ymAaKT8ACJ5jVAg3289sD
9Aa4JoA4hR4YiF1b5MItZENB60+1+2hctJ809HJdmV6M4/8EsVgmNMnUIlJP7Crg74HRju+wmDpD
lAtRn9LdgrJYskBHQia+VJhjCARH7v9r5o4pDW+JYyp/ZM0ljI6T0Q7/aIKYKlc0J/QlGqsOlMrf
GBqoUxPMAL8zPqv2QkGaI4wos+0kzOGWjKgSC8CIZl6seE/CLRJSJ/1oobjoHcq+xHUgXiYQEi1v
o9SZFDnwQcJhHNNBtcoaY6pt9jYKlJuquhlVqGjHrGhOn7mzF14U1R16vTfWeJ34M6ayu6YtWPwO
9ootL5d8YGZgI9W11nButbi0Hghx+nNwaR0oyG1q5jGDkLlnVdWWDklbS+h9DGquMMo3xmNBZooB
kDXVp5EDUktFrl0oPi2RYgsK1I4McHEs6VXEVGk6fJJAesGc5cQ9X+S6L9AnJQHHqlGTYASxFbkH
3C+Ou8ehwaaUQiaA1xei/Iz0Wr8wsSSbnoLVscuOT3tMUKmAJyCPHiVNghI5j7J7N1yOgabJ9u5i
SaXuJMB0cRIFOwriF+y+GlGjp9Y57+3zaNBNIVeRC/tbAqaqRVp92T84OTxQaoALoI9QJBroPknm
KlUjJpvkj2eA3pxWNzExMNMqTGtdUKWYHV9DE555B6uxWYqS2NW/uDBO6k4FE3ch8orGW3Pjn8vY
sK6vPbzg2uEcWgMpruMWe/Z5d2QOVlY+kMKA5Wj/ZV4l7PogrjKKHmP710YmU8BUn2/iDm3NksTn
b/TT2frzM5j5ezU0xYwu2QZZh3dhuiYI7rpZ/gfrp7+rGFGIwHUF6wjn/ZtgozyWR97Xna4UejER
Wj+oh6rjH2Cshyem96o5qnFtoz83VZ0jsLCPGKg7gmGlvrSwUuL8Bl5zWBuTKYPojmeVFTCdaZJ9
XxxO2Byximnu9DfyfNNDkU0Tj4H4yK+9beRhHImrm1kWdVlminMNNpqQ3CQ/axNI7sdk+4OGq/LQ
Me0djCGuds3wcpq8Z0+8cNv2SJATMFG9F/AeFP6VPjBnu6Zp3HeYyvUEpQ0+sVWVqKkyM03dafjg
ooaETiJ29cfNUH8s7/nXne3L642Dh2moIVzSNM2GYvfaTREPaHQ4x97bQeOrLuQEeovH447dlI9P
ule4GW616fmJFU4Tj7RgZnyqqEFPliC0SovRN1PsRGZwo+8ac78Gm0raw9scUWqttvJYndeOMARF
GH47Q0UaNO1kddDtCvZ1U3G1MqarBHN0+Hq2FT8rDwVqnIikTKRp9vvP5s8hkFrZzj5MVJ83hI5l
ye8w8iVVcsENhnoX++PdCltEsJxvsHDE4UDq6LEXxQqKpB/HKK17ocq+bHsiNu2EGfTlteFNz6Dg
RCJUTeVkuapfi5ZYCFvEbTXPHeKPQ/B5lwjWDRO2KdpInRU8bV/rlDz29eVShl1QzgeSJoCGW/ha
+Ny1qsmg/Q7KDhKh5oudMhiQU8UftWK9lXKw1/qz4EuJGeVjmprjcOCmGEZFpi89AkP7J1iX+Ch9
CowpG3M104h651iYBu05+fqz43NRCaYacOecaxKfoKsWYGyfJkbW0qbkatKxpR3m0nTEZq/52kld
yNPLUtR/WQ3YFmVb1bEWpfTZVFsPJip5bjnESsJVW8wUoo3iDyhwXytbESE1szBgfqQj76IWnRpj
1PGERETeYd+9g6OHRkovIDZjBR0CZhiBuRL/C2osMRfR73Ztmbw+wHfE3zvI/qYlqg05mq4nCqIe
bzji3R4EvEeuLYtP40TZtp8WoxfTq55BCNYMS635RpXrP5jpipshB06JHjpUyuEW+77cOkKJsIie
pfS1RWY9LQJ73QX2i03nX1Lc2VZXP39/jhdwMyU/wa5xoWnrSrXweETEFjy49ji6v6zflWISut6+
gItC1o7rmi1tF+Qo47x98y4315DDWhJcVB3xjE1yRJlytCzYbbqv7g4ppaz8jUUuCdymeqQIX4AQ
lF4XrGGi+XppPS77DsQIifYyZrd3ks5yyVaxFsNmLzXW1vqaXFsxRWLyaDIcFPdZ/5kS9snXzBGf
2n1ekUJn6Ds9L/XdCShFWaEdV25ScLRitjaRMqHSkJMwQyyL4N2m+RIlS9qNasdQ/5K4kn2UFhb9
uQOytwUKyepCV0P6S5wrZWDIT8D7Erc+wJY6tiMFYOkZ+z/FGLvkBmWnTClioyRo2agq2vl7wnZj
9HLPu0/YYkak4K42+ev+j+dlGMNEw6ZVq7e1FdRO+QL+DRX1l27nwAjr12N9vD6hamSTnvjJB5ZM
z1Tk+1DeTx2uEVG8XqH8fFEMhTSonAXPbD7iNFsJyYV4CDPUat9TpX8/wzuesNwOQ/ajfKcruby7
z+9QZcl7g7C35+e341eSdLySM7I5mpcL/d53vp75mM5bXZ7guySB1P0nHFwxHXma5wf3NppDklug
NWNSKpSYgcqHcSbxyLyDeqlUxSgQ7Ec/MquStZK5MyxObl3qzjlHJcW0MG7LrYlb36dKB7PQM1lw
8fsVhcgbOINfi0JSG6e7Ds/6IS/5ERSmrw/dgNvjSZRZbrJu/VhfITEiNMRXrbs3q2eSHItApaul
Zr6v3sjcOJCGrVTIX9GnoIvOMjZRmJ3utvXCA+hf2MKlLVYhxiTox53qFmjAsP6kP0xqxu0y+D0E
VlbhXs4UF4FfQcZCY9giJ+cV5p0bFk32JySI0+pT2W0TcNQWiTMAmClWuUgRFswB/DdJrFwLQQsX
uyBob9gXL1FVTSNk9+JhJcnw5lgq8nyhVxXHQw6ojDgE6BS8e3cTcVkLHPF04LuF7NzAB4fPLSMT
DzLySZjhknSu1QH0gOxZlZHWysse3DL890zv9q7MYkV2XhgyRBcfPiggbtofJ7UOU2VgeOovYgyX
cwXAOMaL8RHz+f5xYH4dff6ekh8qbwgunNq3LkYDzGT9va3XZWRVmm7qfCzp0/ogvMtAa6O2XmhR
9QHmEseXWAT3OWws1qdUlHu1TPWyQVrmKrg6SY4UujWblANd9Z/Q+DeyNg5J2gPVlzn6tMtabfkk
JXPSQA5jJCfs2oFLedvXJ0dKhpBPHyuCr0ettzZD1K16chVZBBreCCK5f8a7jxurrq2P631VWg80
nsWDphB3pOcElewYHOOELXOS/6sh5wpYuRV0UgmR1RNThRXOSB3Ndjb2Z1eklh04SWELTBoECp/H
5KtFu2JFcqcEFYbgwzekIwCAZvjVhQdg0tozMgEtyamBuhwcYS4Q4i+fq6Rn/SGSlLsoDrw0TgzV
CJbrwwYCUcVZdemyabbIJF48mRfcgEHkHngIvP2l7hKUjXmlMkMq5uXiX3Yrzy9i9c2u5PoWNRzu
4zy3uRk2i8oqf8HiFDnQrrIfxRkgdFVlyjiH78toW6hZ/oP8UKd88k80RSX99DMUmXBl+ldE/gbg
Ku+/wqmIhNqaFgot1PxN/nYR/N4/30F0mZov8/TT9DNUQvcAvO1PV4jRLMIybHA68Khn0HEOjN71
VLcFYVs6FV/hZ9N+NvzkadDSfIExzHzzVDimH32uz1MFFMWkit8AcNAXZ6Fprwd5VBuC74Q+B2eO
Hk4VzP4k7eavR0LiF1zpYa0Xtu6od8WH37ChdI9tE0SD3n2HglxDTa96ka5T1eGpbe/ZGcNDfWZm
wzP9KToLPGBekcA+zy+M2iW1z8FwbM7Vuz+ZmKByFSuMxxRTLnaOKgvVWPFMBzOZ0UwzoNauZIQ9
kOQzEdnOJrHy3S19O3rDPojgary76+zJhLCndPb7MKre2Ev6ndar+wrCJIIvi+FsBZCaPhL/b72l
4z6l19KIHCHpuQPG7HytLFNkYJoHfrluyk/NWu7x6A67EXqu2p+1RVJ0WI3kuB5Gs0mBYv6AYDVx
OIFKIJ/NdchgKct83dMo8Kdng129uucm1RmYfuY9/IFzcdLdk8ArMvPhjH1lWyT00m/U6/FdtIO1
k3qQ4P2SfJUhuxjxzejia5Bk4+I11KAuutbfQ8Ynxr3mfWTTP3TRYqcwoeq945yOP58RH+C313/I
roehQLd5SSInr79sipTUb/vvwV2YJ3G4uQ/4xdxzs7B3G9swgn45SsCsi3K96vG3f3bf3JZcVr36
UcHPvDepBwdz4OetEZuN7FHOxdLhZQAIUhcozbCDXBO0LCtP71LXiFWCIdx7M25ue50L32/HDkF3
NztNRL8YnKoizZ6iizOQ2CyfhXKCsKVQ/Dovl6CXCpv6HC194P1zHK7r+Vmv+2K8tAI8WarjjjKs
A/HQjnWx5SiPA+LG4UXB+YwwNAabTtpnYv+ahTU38u0iHyuwanQFedl2KDvk6g4tK2Dr495HsHK9
QaBl9YQPBtT0t8NuaWh2GwL3QfN34NgbhaBmORVBmxI8CBrGxm/D/dIpQJfZ0K03dBCBsyMwtOL8
x/pUUx2jxsQGfxeEXvF/HDNDgDXSIkI77GEYVcppSeBpLBaezy/y4CrZHTcs3Jdd8mFFuG47k3Kz
GPByqaFNaHDzW5dEQKPkEXNSQUm2rlhxrYyuVCRYRXSH1Olp9eUi7Uvt/CaW3uJH7epMvb6EZ5DQ
/707T0INfskTrnKfNpN1cOH9oVgy6875zgVVMlS+7iUWDMW6Qvng44e1VazdkQ6141VSqpRnMYlJ
BA/9G4WN4CAONkaV7vAmE/9VYi0W+KHFY/klXJWOBh4d8Ahgl+K5X/puiQ59DdjphXfKiJJZAdNi
Rmr6wsRQ9rxCXdzc/oNiAoAF+qQE1wR0sx1C8Sn11GqBgADeFoDiMmoQF3UdAasr/LoTC3O1oU9H
1xZZw37A1+ELgiIH0pR4JEcvdV6wgCx2cCJ0llF1gh9aHfOIG05eFiU48zTkn0QX3p5EHC+CXRiZ
3a7juNTXDsxN8YR6x4mhTzGR8VKbHVhqQgVHj2hE0E+mFsHkw6bHlmYIWbK5X4DsGVlFsHhzwkJl
sLrN3oxq3WDmLuufIw9yyb7GQFbEjolcBgpQMu3YU8X/O+xbvvTJeIirNGS2QKElhnmRssPMzs3u
+F6p7L3l/2tGxb5953BxZf51ni9sGmGkLrAlElc7gjCynyZa9uBvX6FvCNlYR5bcJ4iXDRZIsxnF
BnPQgjYVWAyf1phHcBAm51iGImoo4mMiLvuddR9SO2UMnn0Qrqa55vztU4Tp4sBWtfE7npuECjRN
LnTDC9rKhlE9rebMBD/wBF1yQNnEN+Tfebb9F60CkXjnYAu5u4/L3ngt9egq1QQ+hP5Yw311Sqev
Qro5QC86iOcNmlySmpB4WSdwbvrInql8JLcda801towp99jqXGrdG9NEJUqRx7XOis+aji+E6KxR
SRbKLns0/YGe8zS8p0s3SRIriXYbd/6DXK9ft0zIcAGS0iBNTdf98tz2zQ6c8v84Kp9c/DixyQFN
e3EBtIicdf5BxMQ/B+PfhBRodiV1Ag9x4A2c3iGtVoWRcj67tleNUg2M/aUroqh+iZXJh1wDJU0D
iL832AZ2DILdOcOaZQW6FV8nte/RablsnxXdwwdXvY5JSDcSZ4weHZEOGhT+ynEZ3jhryoq+/cHJ
cdfR4zEm3JXFSQeZfAfnIpOxcodpERPh199ZMM44PGzh5zUPQp3bqQ57hcDwIZzKQWHeRoP1aatU
XGpv2BIhN+KLGgMcOiuxsFF+Ev1qf/UnB+BN86+Z1scFDGk6PuWf63/kk3OfNPBHsuCjcI9pZj6k
K4RLv+wKGB3af+jRBGY3yVFsscNWSAVr6fBwdoQKSsMNZAZ54RrLAhPrTHdmCM2s2+oIf4x/OVFC
ykmcpTQ7BfzuLoikHYvGE6tQCgWcsdZ6q2YMnOu/UsuHxMh6ZHrxdmhm7stVbvrnM7r5S8Mb2lf2
0h9mgIiL/vBJxqZ1e/GG9Dbh+krR2cwQKSFNV8dZiwKFSlijNICRrre2+HHJIN0WnkSO4iFt2jJS
m8sfH9TzVJWOfDqCJRmZpO23/O2N9/Mo9k3+wIvsdZmYmCuKvBGhlZT2srNnWHR5Tdt2rhcIwyhn
6+96JooUc6T9LuGRQEqRF2pT7Y9eNsFbM68PVeZHP2oKu6/eeWDckevGkS9A8i7B3yvzLsvXHwll
3W2m8E5SQDXZp0zrWEC+acTJXKuDXlJQC+tNHvAbaI3r1ZUoIYYsE+SOsqr5xlFXh11Nd7J17/Vh
M0jriLv43uqea23UXcZlCvZVHzuxcdBJQ39y8lM0HNFj9bcJVxu64sIOmICEE4ud2Cwbbw8UrgUv
LqmmqUtAkqa4ac43lllPr0zwhajys0UMQJqWuq4UfIlGWNAwPkb/x9P/L5tKzntZsgcjLUquimox
tRpYPA4wjLnsZ/H/mZHFCaTTNX32T27PCx8ZVg5Hu+pCMaccwGfC4Wnesf2RQtRAopd9fZh1ry0R
IYilCKx4kSfTip/C7u8YZbda8BEKJtiM0bq5HMoIFmCb1Wtvz3QVO8Cjk07skZt9+UZgQVNy4rWr
SE9ODlesK+3dUCvZbbxWHkc6pPgxAQEifgHfaTRwG+8Z42asGMS6kTrielcexe3N4m16hxU/j0QR
uQfNP/Ca6DQ+Md92isTfLm3n3XZvqj2PiQbn6rwmki58Ke+/uemQvnbfiTva/D1BbcLvqogbclrW
iKs8XiUFMtJm9+Azp80UQz1/DPAbyf0Ef6k6CJqoUOnO1pLPmckkhA99YiOKn/VxLI6xi1/eIL4H
w7ugiatG8FfxOIJzIdd61bc2GJixsG5D0Eq0XbrJ1b0hrzIgxbKI1dPF9PGfkvoFrMNSYbz5a4fB
10l3oymui8AovdWk9u/shwdL7dXaI2hHXni20IZLyiav9ZJfjMdOy/6XyM/u6sBIXiP+Y5Qop8pI
s9Kd8WKUH21cFV07JW5QRTGJeQzQo6vdsjeEsiU9ftnQOdtSby5RXdNIMTG/ZaRuvKg0NdSrwLuF
yqyf2xUkAEKNsWjBhmCt28Qwn/wbpS+7hLiNNanSbDK8Oe9j6w3+m1GtEFTV7MY5Ox2LCL6Mkbnp
1HONTmfkuOOFC9bfta+iK23o/EhclVSPnsRh7H8cz0dUcj+KAxLzawldFKjZMediCiN9vIDrJqX/
H8zQQhVwZOictPFfAiKCuhAiWD0tzHDmC4mRM+WZgZn+1Qg/5fdaU9470xjSvWpeiCvJU7ILO/z+
yqzF2et46Sp3Ed2e1QEqr3PjtP/u1LO3UpfJ/NMTz4EA02EHxawqNidqacQb6TPR4X6Lp1NeGMEZ
R8zI5WvZ8Ur4xsEoUVXh6tL8xYVae/cc/Dw+cjaad5t57DIMPqDgPrxREElCPHK5zyONmhjzDcAI
bRBZ9cywjaVCSqjAaLPzN4eAAiT/T5S6WVDUCtmguibcqQjBl8X64s0c33Q0ZpzRJo+44vNXxJ6G
bTWnnWK4vEHEqzk1zWnJ9X7V5HwiyTF5HV6MSAgHYgioC9KRsh5LKq/wsYKpPmCijxEy+jXOJJr0
VnvkwKRk4d74rmHyWrdDKgahdC08KCmGkxEwuYUQ4U4JLvTlDuO9JvIv4IE6ANW2z+EGaN3iE2AQ
KsE3aamJXTlD90oTS5sAIgMwqSpYE+rufBnfj9Y2Nx3UgcNzrJ8sXWxa/bC0/nPkAaYvFX1POKTy
KUxfhxObqnmXEUny8QIJFmjnjvrI/6sdchqaNhOgMHjQih7rGBLGXHGyLZltpgUYyz7G/xaDPPQd
rnYcYM+ps5pCEZjMasNyA46gGGrpNYZDHBc0oiylTHTAa89xbpPqp5LDOGYpEZlorsSA8rKqs6j1
uHBhvYx4ZDRUU+hhMfGB5Lv96hnxGH/8+asGtOg4f1WiPeOVoKhAyqSzNWri2haaO60Ys/p0h70s
Xv6gWowYKaomTlo5esyAZhZkc6ZtnJ2PemsVPo8jjnX4J9njZHdDNbyCgSzpbmwIjuJvdjApx3gG
ZzSI/Z2T93jh4XusvquP/O+phyAt8Ot/5LUtfSCRh6IRFivFEZ7z18EDRwBP9yZm53xWdXo6QDxe
NVpKTqKU+MIYprdexlgjA7dntXPe/PPuQkAkk+UjKIxPskgu31ScEK+vKNankdOkdhk3aMIZsAmm
hHOjYlJcwishGI1VwLs5omfipNMrvqMY6HDw7UxedyGX3jVqlJfCZ5zUqdUfADRwfaGTwt6ZQT6D
t10o9c56Qb2I9c8Qb0rOzGllI0OtJUY+aj6ecO5YQZ8bLD/J5GvsJKd44p/kL/0AibUWtxsjSvcu
s4TCweA4E1o33p8KcR29VI4r5KbxNnP/yuhg1eNZV3uvWy09/Ut2tRbezwNtssdOF/0BvWm4fHqK
PtoVaepNaR8clS6jsnJFFVW7VI+jtHvumWofHLOEjpTILcurDGmKHLBc0xxGXWa9sFsTZ62XsNta
PJkIy+yi4Rp2GksoHbllhq3LgCJPk9oZyAz1cuWuXsGB0tiwmHVHg1WAw84h5NUfFZZSKqezpSql
OL9PH4IkQV4rrJ8/uQGzaMaW8I3Q/Q1N4x/DBmZhYEFftDsWddRZglfE/eDX0QEDjoEHUGsEl+1f
1jxnfXeODuBM4JUxF1vUerQsaVZglTXobxfb4hPz+qjeg6bNFNOr6O/yCZidfZpOvPl8iusNFo35
lmfzMq7LrHr5ZNAc3S2R8u77wadf138Y1KKULiiZBA9Ca8zli7WNeSK/BSKxrHp+lZV44Hskg7sy
mKQp5K2/MfCRrEcWjZQDcW9K5lTpqj5Snxp3J6BFAqRILTgUAc/pcoT7odQv7KzXrY1VVfbc67/x
y36wApDCYFn6ZVAnVxFzoLVHUvpy/+PKAwDcdlTXFuxgLVG2wVcAG3pO3nUCJWd5N/+QETPg1BCI
t56eifZrcNhQ+GVtt8WuUw9cuO9lxcSiHywCBhJQBsof/vF0e3OqBdjkFDzShQEXH7uY0r+ZuMeD
iuWjloyxBCuQKp9rcxs2zGrJdo5kwFc3QUC6Bj2RbCmMvDRAUQ/A4SfU9Odrp3I6dhdzEjXdKPXU
d41lfSTfxBC+T9UnCdMsvUglz2/zilMHnLIVipvbqKjrpB8uRhivXrWkjowCTedjAva3iZMQ7TaJ
vWHeEY6xmmrQwMHa4ErwaUBeSoi9qC8TiqdhEJ5JITitgCSXJ3KtkrqJ+XQqlM+jByNJgqDboQLa
2wImasxOcW6q+1FqZsxkN2fKpyXFtfADdV7pE994UniZd1lzL1kXleM6z+rBN5lb++L3QWEsA0g2
j/2GV8TdhQi2G4qShqQ1nw5Rw3yQJssckDtY5L3D41aGJ72rUUOnypUAPDAYDzbPZxtAyE+7qBCg
ROgxuCj9y27gWD/2lb7UeLRvP+6vpQSx987Q6JsyQbWCn3S8xaKgqfHbSMl1ogAy8rA4L3+AUxOc
9q3ipiwPARlI/0uQjm6YejZnkFjNclETbYhpuO9KdA0VNoUPd7RmYXNNldM0t8cOMWA3rskepUZ+
WjE7NcoJKKAGSQ20O9r3PNpqlioytQyc6lQC68e4HCDBmLqITmTu7QDWoqvRvrX1AuNwbMDxyag2
4r4O3sE1ykDzODGkNpK3BUR1aAaIyBYWzWaEFANoMLmb7e2wrOeJSPt02oKFYv+iKWrCw3/oZSEY
nbNK9JE3SfsjnyyRso+D46pI0zpOgEm/XzEsdJnNP3xGLEheDk21DeVWQkmdtSj5YKj2xSDNeM9K
uWmdzETMGmUhOlFAKnNTc1F701VTbiGG2q2UZYlTPWprG/9VQnRzoweBMhnANKQiee5Dexh7yH7d
hz141lP4BZFvy6O5TGWsRiL3HVYRLpgSpRZFP8Kq/sn/rqDuiQkMs/kRHocHjNRWC1wFcXmtK4bD
6Wb4r+KvcQuf2mf9TTPtn+JSmWKU4Mw41VhSZkHP2dUXuHp10SiMrvtwTqX6Vl0RtPUb/OBAY37X
8w9PIWlz7wHH6u/yc2SdA8Ro/cbhYQyry5zpyf1K0esuWrUOadKd41h8JkrmOdzgL2C5ETZbjnJ0
6Ktd1EDOM2X6WZXyZHk3/jatbP2x9VhpEHT4NhKIiKiFh5krHYn67a5XeVsv9th9iagxurxVd/DO
PztvYlbtaTegCUEA11HklbxRpyeieJYnybQpVintPefa8e89E56RuFzMCti8irwwcbflek7alG4e
yR+/6wfGgPuVj/2J6DNyraCuokKbdLg/p8GvdH88D4VrUDzgrT/2GMYNcuzTmKqW4Mu4H1M5/5F9
U8F7mjTzXNVTEKR9udAOHmzcA4dTMsY70zk3n8O32wqxYW71a7KO7AJ5FCfZKGgNFM4bwGZcXLos
kx046Q6luqsUFVykr4khZMla643uZ4wXqe1B0c4i9oBFcMru3v3ORBF6iGX39o2PjLFinmRnkJ5r
AlPDkKf5uu5FoaJ7+jpqwq91nYdGgastECeLgts0asdQMLVczfELjh6NW4Jf2vIihdUf2Tqq20/t
66/uwRY8sdCcT5a2UkbjGt0upguj37K7GrF0XCkzVYDaIXQCTKlc3AFdyzlzsKenL8VjEqKJNxnr
cLCs5zI4Pf8PHT11HDH5612BxZniCzwNqEaOyWditXLfS57vEGX96QxfAoAMPhbDpfO/icwoPcIG
Ssgb9+LIQEZ22iJyZdATgR/lpj9b+KGNuEARK5soqGax/pDR/nr2tNNj/eLZL3hzN7TrJHbxgeLu
5tU87EP99QuppzZ6zcdTr1SA+s4zDVgD1uFkd5whTlztg2fWfBaQDXq0nepaZgtISMG2rQdJnSn4
egMKif2TRM0Fe6gKQ0VtDayxeLZTs38p3CxpI5k+BsOtqZUMSFGTbK3IS3lL16LEbiUZpgeW6mQl
smrZUQbkaWCyRDCXAEHRVVVs7kHc9cjQWuZ3vwZNcnMCbVF928mBOdrI+9nAOR39Se2YVxFm5wl5
U0Y+xmWGALGLfmoDbCNyG0sja1/gNS7E/9kIKhB8IFJqrVr8etV9F0/nXyZKibZ8vchKacA3JxfF
OX/GE/ifxjjZIuv6vf1OGQ4XUuWgn543qK7gOUruEaIjoAd/18icPQMp+eqviSIBexuf0a+bSix9
N3IS/tLqVWUn/NAE5piMVsAvR+kbV3bSXzbNWFLLhwlyKBvSoaGXTlcpDxEyZOBvzRPVQjhsIaIh
xbsilm2QDcaSENvitk+DDPDrjB1kG5c1H+ugIZItvLr+sRkyv+SX6f9JJL/w6bh4MbjKg22BXI+Y
CXcY/oYni0jhGMF3v29Cs/Segu5BjFGWHCfpIxD4kjw5TiqKQqVmJl3+sLY58u5MDHVIXK/UR5At
F78DsMCHu30K9WMYUj8Ez7Ot5etedX1jBCOswKR0lEnEyGoCHQ2Htcr4jA27eQk42qQ4RVkPdNEj
vzCCvqyLgnswql5B0A4GJP9KAw3MOGjLi1ABSks6259dvjP980+ZFhp8qGeAG9XMMcEQj65fsbmL
HYiosekKsxIRcOzomvx7crrjzd7doFwGMey+S2zcUI+RUp2nOK7yyXz/0eN+Uj0nhJCf90nxFODD
KL6rneS1bAnoxMWYBbM4SOcZ6jLPhsX0bEX7PK+nERb1kMUdNMAhyYuyUkt83cQ2wDaQsP7Y2FM2
HadMSYdAYePHpr+uvzANn3IYjnDpVv6MPAbFfHkEWV6kPQv/IkvYnCDb4Z1Q68tBNZyiVLeI5VBE
B9HE6ttUmN/mjtfvK9bm9tB5/ib6PMmkMjtfrWAnApy0Akiv+iceYL6xrnTGyxPceVHUQcx6DaQu
B06oc5O02FGRjZmV5DcGOHxLJX0YT/ZBWzIWeGqU1PbIHJ1OOMsfzp4HOY8bnqHDe+DwSoO5gjBe
Q4oLkfVHWgtgY1ios4CQxWQzaEt4GEdB83t5aoJunfF1Cp+CJQVxBzrH/DsKlD3ZvB5tSF3uFJYC
Wn5Lex6zBUK8Wo5KyJFq/xbt1ogOI12Ht07Q5nODshszCRwhv1yBKX2zFvlrh1spx4e2ItAxi5Mr
bzqG8DqI7D3r1xiRLXtXV6vppqTwwtAWJNOSXkzyx95pc+fOUvWtC/cCV/zk/rKKmPYLBLa+0Epb
k1NdA9jVYxhCbXPn4w4p5JOK53p4xfTz3g+kutevZ6Vo+/GLpxNbQswAJXQrHy3abjoqO/odz3cJ
RKGHJ4kT5Ac6Sq4kzHYqoc1bi8VWmt4K5sJdwqw4ydzqV1DwSNqtSaO0nJk4QTk6hennPW6KcVyl
ffHKte2ixS6bl8ZtTCOmu3ha3etSZ1QvfEtYcwcKCxJV6Q6GeUPy3lO4jsOSZcDHO2hARCtpfECD
2k2Us1ab+DWdG5GSl8jxPOLoIwUt33zS1WYRDPPqmoJ0OgbJ3tuJQYxNFiFLsSbd0DubuFD0V9iX
GT7s8YZ65JzmeGJRaCL5Gd+mcXOiXzKmJz3zg5JGP2V2GlioobB4wV/Q05M+SOSObS1wgYOq/JT7
Vqw73zNumFTgre2EHO9AFXEwY7N4IQEEnhhSec641waFCu28aoB9Xx8rcWMeH5FqFPIYb8iJTDbM
y0JTZZG9MyqxloNXx/qBapYhcbXg5NaC8IR0D+//xAuUkvvy+vz6wtz0AFodeXygpH3LbJULd2pv
NjAE01xxgX+gXgvwEeGJ1K98XsMHHWHCU6TVsiJ6VRK9LgJNAG+6zn8+rk29TOoS+mza6luXjrKv
s+pnJme3hepmEPiOm1wNlvcN0Rmn6Mt0+yK59AarAtdJg54F/tWgTxeIyiRw+83zZohdwH8ltbTY
tNwG2oyZ2CVOCsATUoBfOuGhwW1ZyZ3w0owDJ/a76yaF4WWlVpf83AvCKCwuAQGnCdG2S+KRJjTz
22zgwhaFd9+uvSTqIPcUgsyFUnASJWPf3+OxPd66HuSUlf8/2a5LLZ1qfWZxApEM3ep9OxNFjAvx
ymBnUwc0irYoFpXEqPJbFxQCpIV739bXGoKDCq2S/JLk/fG73LMnzs8F8XYWm8YU8WZjboH8GqVu
OuZ/4o/dXqLsRsS4Hn0JZ+3zlL32bESeXApWrDG83imBPLeRFmfce0iSdCvnzICgW/ffEGY+3u0O
s+tyYjp3NtrX72A36Q0ndj2FnX0U9oPxasjig/MF6QFDsCNQ6KHPUL7dcQF/qwzDACM5N1SDB00u
J4jj9GYxrE28cOUKy7YkSwxcsCNQX80zJbTIxgbV4eSRfD2xO4RdZ3CCIvwJSnQX9khS+YKhsrob
xyNX37kSSfpHYuMVf0sE+sT8duD5HyI66fwAe3wVfYHwzTdLRf13u3zDMdPQ8xTCX+f0VsnbtU2i
Bsos+6D/e+JfbDXSgfS7+bNkSEsXvraURoAT64N56AShlwyZl1emQC/NZnicdDoydNHYnhOGU1eB
f7jMll6LyvXTIPb5PpRd/uTDXwloAKeL3gur/VxDhsiffMPyV1VM/CfuBo4XBze33BEHbk8MJ+mz
aJIiHDD2cP7HhPCxnVcwSCDWPLnE62zV0Q6yxDFNx5Dv5CV+TejJbS/b87Seev5wzY0Dv6kBc+5q
qeqxvudvcKvhfmiuViWb1bJMlDiMfMWryiFLUYicig7msTeY0yHC0udwyqzNipz8zIEOSwSOEtxf
94Z1OtJFphd2QeAWLIsgVuX5S8BnZ6bln/CvHsvEiV4FPHUtVKhYL4USj2EN2Uys5zx3YYAOKP27
ynfyktHB7OLsai0bCAqHT5mZTO2HEdS6xY1cn2L+CScQhPDuDG6MQaILRtptXbIKhojnNJNxJCvI
vICQuOo0XQok5GoRRixEWOaZBzDp7JqlsrV1LvcKQZQdXI9qGtCBaT3AK3uUUy73AQ5Ty5lDfyeU
OZx1W/c2AYS7BcJweVTmLJOAZaC65Fyq313xiMoe1BD0NhNpI1/fRZlgyUVQs3NxkHoZPp6jGxD7
gVI43q4fsB0ijjrFCfxe2g1N74xWlC2rj18qH98c+vBsHIz0KWn1i9VGqfgskQqul68ktjwakbvY
qstNlWLOJemlvSZ7jn5K3GDYMnJO2ZHPmr7uNBJ+9F5sQgd5BCrnZQZv6Oh3ZgLaaFLNr1CwTjiN
e8UYUJVav2RiZYAW0giTai3hAnlAhDywMl1STJVN4CVtsXsoYkAiDeQidO4Mh4U0cRAeSpQGUygE
M8InLfLbcHxpNc/Xdbi0PTWqPda8nMFoRySZ3jnBlTLePHpMvjxrUSEv4MJYq8ZcenXyQ40xKK+N
UegoJGXy2lPTAFGnwZ5BaxQMLAtgnRRLg1VRk118D2s0Q9ZY8QT8NwTB3i9kgQEQ1OHb1VU3IEdK
lyyyhM32g33LXM9a4JC/3PL5ctIkIhTCNLv8kyXl8Bgt3USRJ6WEScv1/xZ9QzAxDxqDTT+VrYwe
827ubC+1UB5vRX/7yqSw0owWq6Ak2E9Er06nkOt8dABlw0O8xRHgEpuN0I8Uyjd9uy3XnTm4j1BT
3dv7M0DdZjGZ1GkL/6VhZ896R4FOooan2aW4oyMaqm8OinaENCL+rcpwmXKd0RGXT/9vA/OZmMNP
IlCy67vRnnXztd7AK4h1FbGiKF2ROJlERt9lSQ8XgLAJglvJUOORgedIaDL+hSVvcx7HCWZ+J4vY
Jl85owolMqcuTSiSnzFo/BlBCvPC8nOKZ9Zo4TxjSiQ+0D3lkXIfUlIcKiJHQfY94mHXirn96/0T
B++fYAy8CLFqIZbDwd4MUKvQ1ea7QXZ8mN/4iTtpdszYOOEZQ49jT+1IGcgvResbkxokKfqF5Y0R
/58TSfRECNlR2H1Jhz/Xyykb3/Boqaq28fJGZJxPMds+NBBdI5Hy6a7CMJCLcKtLkOWwTMLUlXoa
upotlAyCmBtNnEvLR8d0jw3jXySetQZ0PfQjg1cLYXFWbWMCw1VwkjP3Kp+zE5fTvuu/BvtR8PBU
ZvS/KMMuf3hBsU/tfOBj0fkyUMnpISVXmUEy30koLYln9P2GbNiQa9Ww47INIsz40CWVvm9lucxG
J1A76d9YZAoL4GUoJef/1amLZUZyl/fGGMYRZdTwFQP2ocHc6U/OgjYtA3YYqaBc6pU/NUYruS5K
q9CX4HOrtnyVzuVRAolY/KqPfG2dJIwVNEtShNJvkYCiQAJTcUhqHXANyWr7MTze9pwaR5AQws9L
VfKP/pXdK6SvEEHrKUu6Ce0GUm0oCnrN31vre0IilrFTbU7bcNUC1UwRgogVYk4P7SlEJCINfhNS
y4uWbizz5q4p3wRLhPcpzhcKx6qlPnCNzDCfHIKW6dsyz6sXAsCzLXMtSyKbMW0ZZkcBGpjCghkG
M0rMKHQdMYXYZ25MfO8fxtrGEC9mBLb799O/rQRQOopi0NqR//GswZn56YwBrYlvODgYjKdBAIRY
KyNM9Ul7ZW5q04AQVPidCWWBPYUjIQhqaoO4YCRShaXtxhtN2k3FUE5T8qmWIQc5zWh6mAXK8q88
TO8RkFWdelFDUsdosCNzRJG/IPXAI3aEjjw6QV8Gt4rL/g7fWSYp5VHrjOu2BIh1qonutSpjbRWI
HmkdXutDpNsVB10uaPNsRbKIorbqSUrO3K5V4yKERVF8OK1GNKcZD1r9PrtuQ6dz7jNG7XgL0HpY
snW5OHPtgENhf0EC/wcDqC5Okhx5dIqdsEzCEXE5VwBILLBeu5aF2kNn9F6Atr6pC/BC1qdws7R8
/UzvzTWw9VAqIXpkDVNfqdkRkK4kyAPEKePJ+uPSdHXzSWj8JbMUcZz6jeFwiFwSePNtUugjuhka
5Nm5xg7y2P8yvmT0locVBHk8ARSEVPUyR0k1kCvjOGPY8rbt/1zPCmrr+oHA393ukERpYOmnKsAr
jFripebjAv5bBbse9S1g1pFybAydA0T9LhSxT1hiziN+arQ/JeiqRjPfp2gWEG+TzbtKdJaJY5zp
CfBXkOTdqa83mupttVJKMtd+I5jxuX/9tpiyk9iYWmCDIk3H4xTwi8lkUttPe93CRnedqBbYtSVl
Fx7p+YUq8iDbMgy4s2xbzjKl8hR+9QzISXmhLz3J+sbz8yJMb7r/LQRIK7K7LLe9qwuKGG2jKw2o
Q8EWzLeTtzgTtVv3Az9NJ36Dsfd++DJ73W392WwwdT/QSCwILopDAqP3gaPCOYkNQZcV+x2+LioT
gKSSE07Anq3yPV37RkivyXhfIZGUParc/HUTl3jI13FQNMTqlIFAGuxm9CSBO5SZ9/CETWxqNa0W
xlqH9Y2IA7NjU5L+/O/jcRHPr6vZvXmVK10fFbLzDsOfhDtb+Ra/oRxn2JqpeOOPVEexnppaWfkx
kftoUBVHC++ODF5PWDlEPKi8/Z1XTPHG0wApEfNHqhXN10jbe0m4VDua5DF9/giIY/2bFRwkWYR/
ZUMnmB7tF+EUoeKHstcFo93uPoCoYCIsPeg/UpXSg8KGn9dKR3obDbacflS/Rzd5XTgMfN1R8dKr
9fJ49KDAceaVj70m0nt2TsClB2uw55Jrabq1wggi13hkviQ+rDlHthGQKfBWQDqCxcBahBqggFrE
X4y0TNPakWtVVXxyytonq4yUzSB8rXkTY8nsSmFXil/QtWkEqUchxQBifGo3z0M8xsDN8TfUlYkH
lVGDKrKAnXbh7Oxy9vuVI1/86KVRXwDbm+eaN2UB6a1xHihhDuL5CLlgIVwmNgrTMctW61U2EuE/
DRC1Cg9puoxg5EXBwwuQn7N2/N8ZyzS1913T+TQDujtbB2GUHiiBIJB6T6MG1FOE/eznrWRSiyQH
VW/o9FqSSsKhqd2sPEWDtft/A1e+FJdfqIagtm9mAblK/w9hCr12GBbY63+kTuywI7lZVrqUWL7/
DZAI6AXXSjPr7vEW1oN1DVOdr7r3nKJhOXmT/bMHuAC8xHYMVWzAJLawALq2A4aEJV3hvrZXHIYj
lkgV1CAtDrFX47D2yB1GeKjnlidlZ/MtT4NAnLV8ThT9wNOXRUPMLAfsTQXHagOVnFRBgx8RoW8a
XVXpLIMKAPeCn8vWpwE0jD5HrdUJimdpqUQ8E0mx5oIabVnWAN99qtySTQsZiYoU8Ymn71IDXI/G
vjGNNYXpq0CEGodnwda9C59vLqCnvDQpvuvzajk7iMoiEQ1V6Z/YMWDBd3dzFBzjlsuZP//wEk6C
u7rDO9iS874/9JK8vG8egbijkf88MQc6FtHX+Ci9GqZ9IHxgxfRD/eWzF64vQTViCrhrYYdnnqcQ
pjy4ifQZ5AADo+WcDOXcE6nhzMdTc9aVi+9vjdaTniZNCPcOGQgVCqw6RLc+BW/vxhPSGL5n/OmO
961qsWe0b6q6nUIxXngsDX8OVSL7RrIMmVG+U+HELJQxReIIbX4BxiXmhZPy09FcgdC8M6UH+kR/
mIFhVezMJiRSfUR+utUAWWarQ9frOsgVyprxE1EEbSeRgOwFdEpJaSZ705agWPhdMepdMNHY04b5
RoNS97Om9ulce3v1JrFtBuGH0JeO8Sa8DC5R21n+RvpaUbbEx5mmxUSB+JU8qt4HeC5pDwKkoJoo
GXcMVIRkV6YE0Xyw4v/TnpyKFuJhfRxQME4aB0UdzC9Uc6rSNjD8IGKr3mP75c6TVPFmYM7PhR4k
iwYrvaNw+rYQcWSIpZpyIV6vUGMt/KLMm12N2Td2Z31q2jFyWvP9J9ExioG7464qLgaF5bhtzGp2
JPH/m3/+IwEQ6FjUeYk7ilmEKyqOLQgYZzTtmqvnyN6zYkQKvf0yJiI8TbPDRFtlWnk62JNQ9gL3
JmZWZm3qOyRiCdZ0elp7dTbuNRdZzL5bEGZH27ANXKZOZiwjHd0kC3No0Ny6HZ4xi23WD2IuJuHL
MrhEPuV8SE7mCl+iUz6flEU+rhRWQO5SpTw2qUXFs+gFw8XiCHyE4ORHwGUSjqMnPNuuTMUqVxWj
m8BMD59be6Vaiu1YO+wVHNs3KAnG7kAj9OxyyRC3O9mvOqD8XoRc8l/AvgtKU0dxJaQ4sXh7GdsV
oI4Kr66YswsPbEPYXab7J2noxs4KDoTJiw2xyZrvkvISKHp31qGpojArDxEsICIEHYp7s3vK5Nih
2HWWcJuoVrmTqfjmfffyXIioAcpujfqfWat2ND5SdFq/JQtGhLIGdLNIS6tirAKKAu7MNsqO/Oi2
2StP3aQYT3VfxJNeP7N4p7JRmE4SuhIUuY+4TmHXToP8ehRrTGH3cj56P2hlyQSLK+vqkjiGi8+f
Ba6jKi7zIK6b9dYGnA3IDqJiHJ4aV/pWNXjDFkmL7Dp2xD7Tgps4oZ4S2WKnUaS1bm/rFwRixFeT
X9uN4SfcgHbhyu6+VcFbLz8ki1ELul5kV6Up9pgNvcjehQoMpfN4wSbCvhHTKksqYcSpa1cuSwfE
D18n2mZ0vCVFpMXnH1djohnZfFTO3ws9byRBPWs1yUUAQA8F6y1TkWK7d2Cw2B2ig2GD9/Dxt8dv
CnJj6siFLrrTNSUgopzfDpvtRYMXroM32qz8TxmLTyADpUqAzFOU4liRwUz7vg3ufw/nHHtTuJWO
6XdpdhPWmfCoezMw85PX9DRPRWhInL+NGiT40DJKrDFEob+Bm7aQGn7b81dkdDT07KcQHeLdMWJQ
FlADx7zNGJ5prAjU/BK7765xtK/MmYzun2F10pAq9pG2d2lY1Oe7BbaqEi3RWsN00o+ta9LrGQxX
NIPNZxT8x3Ztcg1uQuuKkAhB3pAUPS56YF95U3QGwiWsIgptncqgD37hLC0dzMLDFqI4vQVGAivW
UqZz7X9eA6InqZx33nNK3+t4eMHv+XEiTK5peMUnZW+GaVxOz1vMFBiDUr24vCqt71C61Zqi4yNI
b5BcwR0MEwu+vNafJyAcwiiIjElYkacB7bGOGuonLYEKhwUj/+IWSdKbUmLxDPjlvAVknTlaE7kk
DZ2pzro2ATMnsbrIq92lrTLS1q9pnHYaebWAs3vxWey2pUfrzzd+4fdkhlCKuv/puXG3IIgyHj7D
Zw4cjFiUNgQUlmMoWSuoM57dMd3PczUfBfMK/GisTHO0NvbV/YjZWM3hIU6PB0qj698zA0AwY4ea
8OuCpk0m/YniMziIvi26OaOPXt9Vd3n4yrEb7yGas5UCHPDEfZjhK+ebL3Ebc0ncBt7JepSalUw+
S0Y19uVOlhGzxZb2Rl3TIi7qQYWiuUBdB8e6SOEqXky1XYOpNl43lrx95jumfIumu0Rx5rH1DA02
xH4D889ix8NhfITdeLOwHx2EhmEs7j8XJtoQN3TU/Z1lBn1Een7cqFNDqc2a4RPpAies0C99VQSc
mfJHQ1pz296ABBKROd0UItKHcmcEoQoACoH45KMuqLbDKfwN5gxMwcACIxeusmHvQWLr6aXvphGH
RiR+sS9/oWQNY9TOfvZULQbop8zURSZ6T/MYzTzByQ5oSiiawISHDvRxFKQ8x0c50XuIE/JiLPvV
PT7oMv4UY8R5aImJLbE3tfEzIMO9e8lheQc9N42Ag1KukW7sLeXtqahwR8IvM8+SzBNvAS0yZR6i
lmzxWxgxRqe0C0BEt+kcNuJUHcj2EYEzfabbXzDxgdZd2iMIAyV5rjjnDnIxjTCqb6wwTTGbOt+b
WHtf16VTX7jtVgxCpJQYrflsN1igDHVGCZhlQUsJahCWfVIIWeWbDjDOzUt4UpH8z0O7mig1pz9O
nO/HcCjvcvesDyug0UXwKCcXXWPIbRepZ/3lkmDBO5ycAe8cwI/5CFoal99BL9GRRWSvaCgoX1ip
iyPT6lKFJ/80GQHlrvksyGn2+dSPbPasUB97r9fvPU8MMlksIC9p7sD0tnkT23WxlPFfmBlGrDcZ
BlDt/3qm5ZXuDNQUBW4VPRckPhqH5/OgVuYKPrS9NN/Y7bwAXnMGwsF3rBs0rKErcrpEzvK2h2BQ
0AkcicJvpmLyVFosYgIQk7JokEtzJZNMXETqNzGJZhzyRj9fczGuMhS9uxoFnKE9qzIu/w6a2mgC
14+k3eKfzQiY/sfUngDkvnoY9E1PguHuAgOuN9lk8txiA0m1xmMbuq4Aj+wfMJsOuiHr/fuPBAEk
ghpJoj/LhGp/DfZJI0XrDie81mLVeLSreKgQxcC5AtblEco09YW9S4/mJff765W/wnRaHPjdvqyH
j1Tn6lgmmUmGhffZFqt8lQ5FshCZib+LPa+wcfVsGGY6IGSQLRCEumWme7LrRuKfRsvec56JI0Za
NUkx+f1/rDKMnBabxa3i/1A0UKsP1uYPf27MUp3bM9V60rkpqB7BZLV22ed8quckuYG+9V33QXXE
5Lh20atx+X/VE2OCNm7JUWu3EqWP6L6WIhnfaTo9ADRPZay+HLwwO2ogEqgQxTr1XhazxkKLyxTk
C+/SlTijNZzwhzDFzl1rIKyMVjTgxfm2piLjemH+jsTGBvxn+1FxlDj3TNci+FARZUgayVXtLv7g
OU4OGoCYCxV92WHQGBWPjZhqDJRSq671n/mZvnnX2E+myJTH/Dh3Cdpsgk86ssR5IpljDBDq2yA6
9c7JsD7jQPFDyZNE2MGxkgfWFiOg8+A3e0x/CLeT4o8QWtg2mhpQb8VEJrU39I+fKqdDr0JdM1d9
MVUVnOTxsti99F+q2CSaYz42hEENeGo6q70X8jmCv2K4PdMvmX3rBxJL6p9zSo129Iy2s3QrpWTJ
JTuoSzmUgG+nZLnhxKyYJQE9mzME+QMq0aFbZuAAzv+cumeWYfZJQIvxdiGJmkaOSPjGmYtRUrtX
epcs2cVl+E/GvOILzKnX40a2ZbfyRO8t8gdVtlejj94Ftoc0xUV5qPRHC5FHHTWCUKvK3nOqmw1w
BvkA4Skc0CCnvzOOU5wde/Af5n/rs2SPhq4STR7h92ba8q27MZsHXRbuBAAvVR1ta7Vl4sQDT9ZC
LORzDPFCP3LzOymLz9DrGYVQIsIkHMZelp5wA96U3dH7lB3jPZ433lU5fdAoWD5MSuOrDwC1pSDh
565YxbSp6A8l3NykJLMjyrX9rBbG67J0Tk/2dnKchYFRHIWDkXNbUrYWRTg6JwJp1tRVo/Vk5onE
60EV1WkCHGbH3/UO8z62pJCKlgbsT0iMydrwIO4bWmBuzrUvalr6M0TYFIChfN7LDKuwXmImDgx6
PB9/SeWsPAjiwy77op7sNLPkq+O+JNL3d3vciBm7uxdAL/B0DIaqPT701q2Lfl/+nrI1TlVBsHb8
+0u5sT2pRd+545pmhreWU58qf24vFkIFMk9PKk6TSA3cSP3pBFSFC1TarnfCe9ND6xGPLzLcobZe
GwOkfJFcwTdMqp+6uX2bOTUsAJn8ce1reUYj6ho92uvfhrldvSqOr9wuXUS+Y4UCuxLMEI4ex1cv
Dl6+K87VPCkKfBSrCXF+7Zb7tHSudtruZ13tZOHsgJG0bpPji76go2Zdcy248g8RHD/vjLBzmyMM
DzsSzUt8OfSc5t8IsKK1LNtZ1d22DAlm+DqtL8FnWFSC5g1LgH21atjTkXV/tRZSs+ZUQ3VpsJAe
2hYcRfZQcMC99Zh8tvLZozB6q/L7eWSgJb1Y5SosV5q5yp0D1K9/jTMrwTfdMzahq1jhu5nRNSjy
TgMqmAgn+q3wIqnVScZXYllZF0bvUFcAqNPoPSVDlJbP5vNv0gDkavfy3Y1eEKG/3QibtMO11LcK
mIRhCdjDDP9gBvkYzUJ9uX7FsC1Is0phIVONslg9egfms78DGX2hWRGB0CR+GRyLMUNBtCuWpoht
1b81JSv0LEh4p0y/qoxjYH8VrPOr4G/WDu2K6bD7svN7lLrewmCFhYUO1ULPWbr5o1Uu+6sBVWNa
TKEdwExWK1YGVuBkKvjlpOsuz2bxj7Rqy/YP+S+upK3YhtDZ4SuaszcqvtcsE1bc+4onlaffhNDv
S9mu3Yz2FWqlg4trftyBvUPG6YhVcXXU2QCRjzyxOoPuQUHk5zqEeqpSfE7d+ZobI51baKmurc3e
dPrDtxMZPOZJE8Sr8V2Wu4jc/bNBe8b0SBEpp8gyHAnSqegQWH/qAnyCl64SZ9TswlvbxpMUVbXl
T47r7Sknt5xiG/DfagYN11IGFbBPdI4cyLYClrw4c5P1hgqGmEfbL8AgMGa21BNa42/JohDRk2Cs
ZbKjhfsoonKBFUUFgulUyLJpoSkqa6nNxQGttgRxUeN9KhS1sr/l9Z4DTnWIJnOelKCGK1XUunGP
A0enLaG8M6aiXc8ZVL+JHhY+allGI0N8IP+vcYLLTfhq2XPxtRDQrq0f/4w9WAqLXRzals3Tywba
GQZw5mTwsCcmu9oxLvW/vPwoDnrli+s7qnL9o98l4MqBnC2kvkh6HU0i4lqA12Isb0w14GK1tG+L
/cbhxQBHINTqfyHFZjMOvt+AusQjRKe+spabYzL0DLaZLdA0KB8M7qriMnFyNoT9DjVnZ6rmSgF9
UJDGqs85XvnqtkOI/tPcI8BXzo0dG4q3v/2jaUv8lXsuNfkNUZdLIDEuAwQMaHa8ScKwFRSz+h0V
7bFqsYj+4jowXCBg6PWM46T0Z0eJmSNbksQfA3h0EC43GRbj3/rGBz3W6f8pjZexTBnpB6/D8EQm
WcbVr7u4QV+Od80ZZ+oKWWZwXQBKJ2PdgKP1adHYj3C1o8HcxSXZEkSFIQ1Pmh6Dbi/4eAvtzByu
86tY5K22gBCVi/lKzNgWlUxcthGvXFrvcwca49MqrDcr08+FCEsuZ37UTkYKW6RpjZRm1M8i5NX7
mNMTTNWNOlvcQKayQCA2NTC34WnUmG6Ybq+UGwJLLJ/lUDZfOylhwU5psyhNVBtMteQ3N7tBGM1S
fWDPdI/ESttSzTHMkIFgeRT5Ni+kNl3Q0ODN16QRMgzDqXzFdFfulIZ6wPBVwQnQsta3DEpWgSv8
O4cPOX5976dSAWelo15WlPKAWntofHWGmpeEaLaMgKIV/uJ4fhjjrshZ3Ua3rOwId/2JJ+trrXMk
E1IW6MT0aTA+R5Qr23LAIQXcCSZGU4WY9tpGuRVpvqnnwwX/b5rfL6peDqrRkyArr0woK8AY7nhQ
4PEognfMjg6YvXrNAGHeycc7xUXn7ow/i7VWILfcqc1D6Z5+0sPmU2Vcc8mEkHE3lfo6B5orAb0b
aO0VTjCQxGp35x74497ezp4XnBvg4OgzEhpKLRCULkNk17NpDgCDTI5yTs+VTyiSqSoQfua2srTm
AtfDzazMMRbpH5QopHjuF4Qt2jlfoDtdzW34Kt1ep/2GUziVTTXqIi843DE9k/uFJ+RQSlpVLdKo
Yy/jfd6VLvqM+p3ItGYCxgWevdNdMNNgw9dFrWq+Sv49UQyMmSTBYoosCo78VsN6GFqNtNFpKB42
c8nyTARHzCuYj456XcxqqKm/5ChtSDs1CdyuPziJBv/oeg1MtxZhPM0KpIJXpbMxr9+IHbhLKIoo
nIeLkkTv78Wr3CdSDILsZoMtuFFWFTqoEYyaw1g/sdatrOMma9BAF83kYaqCrtaYrUeLJfRoy4VU
2XTFzS/NjjtKrMCm6Mp7pB3jVIEXXL4guyEL2mLxiKp6P62MSzF8ijeeZwlHpY5BuPaRsz6s9YpO
j9w06hUQUhozpWxHoM8Uyc9JoBREiL9Lt9/FukayUFR4EfsDztt8bilYUf3VYiFAiTqLgmBPv8ia
X+JViC8cYg8qJD4xt/c1yL1q/p9yVVu5i3Gkh4nEn3e2Kjogssl4q+pdNzv+dQ6rHKED22W7Cxds
uZI3AStR6dyfyNfxQ9H8PDXna+Bapbuh1A1uplLkWssaF75bcmZCSujAkWsPBXIec7loOuytY2XT
z022Cs7rAwHw2vsUGd3vKU57mb2KU+uagB62+SloeI5HA/qvICAwi9w8YRn1Qp/feWJAbhUk9NXb
P/6Q7nG0rD5pJANQ5kH7ke6UQZe9WyYPxBw+53lFaN+FgPkbGsFB4wzKyHt6+hrzuvy/LbGXvloW
O0UedDysssdOntDfLZAraWILG7XDtuETAYEa4KXZcCzhjq23EDEAAaxa6Fq7YJ7h+flDTzNY7FMb
D8U12Mse8uGKmdkKN2G2zxlwFGNwoB9x6CETuaYCLMv88HD59phnRyBtHRdAz6wLSU+679ym3jw0
GtsNun7o46LU1giJorR0CnID/Z15Zz2hnWYUsIhjWKg7tSvvAnuYpRg6vTwRBpbSakD8Hk1bC5Ex
yzbNdQ97/pO7NYDbdB26cF9Ls5qwPZQMuJqLL6jMt8epb8JYQq4b6jJIrSpWXGGEkntqy6H4RSpl
kYY66lqW7mb0f7yXP6IhC+flplxtfIT0tPMMrIKyLxnABcrb0ioKo94KYLo0M3rrorlhGnktPhkr
lKdv3DVIs6gSD561n2OoSEzd4WeCCtoc8ERhZkV2L4TeEBa1hKbBgC412syWZHrJonxKCVwBs+zj
Tk6hYS1rZimyenXZMuLFs1dyIJFPnUmncBsQtKF0sKscSGfgxyrxZNAxVtWvAnp1fgqDSl0O606i
Un9p6H+S0oV+h8BP2HUC0yAQEtSd+F4NurRlT17xdSEAkpPEcC0HbYDJesnBSsgrsrlcbAZfjp9q
Ymffh+dJiuas7vDB0vHW0IlMlc64HtPEFdrOnOVDI78N8FiKFxlGxnJyno6ge0SaSCznsWhpSuRT
fWnbNAsYI44nBkcVdXUoFxZvIc0jJf8+CNv3OLMG7VHWZ64JYbEjG1SXSbpbxlYBPZWgAkhGW3TS
g5KH9/Vpr2UETLOz20Q0tIFedZTcdMwTMWOgwY6EE5i5V0Fwz+cVejXtveh5lWlsT3qMroTnzib8
gQPV4XeegkqmGSiaQdUqxKkdw6q2HW8Ri8PgJR6KsMqDUt/8UP6JqlToLEd3yx9rS7EdrW5hKwxg
H6M2MufPs6L4w+w7SnMkXiytP6GKlwgG4BqTfdS0FnihyMs2WNywt0UEd5Rpok+S3Lj6yQ+2kAXH
0yWKYypELdh35dMyNfcVbisW5yKPIXPPhSXP6KR1voxxMlEJcI6CGkNrQx0RssQhAXPF3KdxGF2J
96a12EHp+2VbHEIwH9atdY93uEv4IOUQ5BNB3EzBQfvyhppOFrNNsLCA1vcUgzllAC+czdza9WnH
9OCJm2NdEk1KxQGZe9KZZ7Q4+pdCJZ8Q4Mf6x9p/i9wUPq5uhQ+BxWO/rUkpV3WsiH7J3pRkK3HE
Hev/06+Tj3Kd4o6QLt+3814uD3TymexakX4kvxjBl7j1TabWRN1S0fuqpHXiR1bfP8CQ2V6H6B7q
vswl93Uo+W9asfgSJ0nr+abOZqStImh7RMxnqnjAGcyFm/wTXg84vikSdw5NURMTUm5nogmiG9Hh
dOWJF8G8Q6LUj83PIHBUWyp+TJSWDFb7763dhJ6qrJnfoSuz60oTaawXBZGoclQHzwQZUHXHaS+G
EJI8E6IW87nNTVkmXPKwGB8JuZrLb4WSaU9wHXXi4BNbQs02E1SWT7udY/9WMVjkhccIo9vj/xzl
5o0At2e8ElqIBgheNFpMBQphlPGwkyYKfDjAUBrmbRfFVlX+d3UNAeKwBnuOaIBrG40mfNUfM6o5
dh+tUZNPa+GvWxefjoOB4tf6ax2RWdSU2BUWdb9jKt6Fyc2RqcykdR2imM2i740iDEEI8jIuhuhQ
nKiEhN+P431QCJ/+Jka5W7ximyo0ZrkLGCeph9le2wMpXaTikFN0ujCvqdunD2oD2bcqCSKn/Hu1
5E1YmRvW2hVElK7yUD5ZoSSWVEDI9VTM44wGnQvtJ3S+O4SEgFT6iuRmiLee+4tuXbDpFm3lnQNT
w5BtvWyKVFo36pjwOkTAsYGpZlZgTC2x3X4IwtBoKnP5JUYTmNisokym0z/QdVAORJ+SRAKjh443
qGVEbzBK0olpiHdE1GA1fSlYx3v3EHQpHe7/cVx4/RLatx1g1YhOWrnUZ6eeGrfOHV71fr93GKa8
+7gbB3DQxVv8K1HNx/vUfvc4udC97DsfvZTgMBL6WV3FaeJlB4LFmrr4PvFkl4tt/2HD0G3utPQy
udeZuy2QdyOyGwuCVOg8fSNpu157+sEgY54YywyNBUmtKnxT/SOAyhgVdceWYj9sDECTfC2rDSYb
s55d4RprO/ylGDsrI4j8IduY4EOmaIUB8HzXiR/Nbjy796A/oJ1YCVcBIJm9N8N+li+CtU4sMu7X
7BM8PRMdXpCEIN/O0ACPMrOzv6OA2S2OXmHJTmtLGah2rhs8Ilzu9ZlQS1vBSldE5s2gMsVzs5ST
vzeomgwLDmlqtE3MOuNh4wx7zsOAE28dcfkMFzGmEjDcz/AVr5IpoTNWEq9cfzLI5CjId7nhxTlh
Z5EfxJ0mIJXxS52VitRfWbcxbYQG75DZW1LMphKJ9qOy0TT6FItiAFyKXM6HhXWwYRXIer3xBahX
jEQ/hdmBXc+YIRC4f/5P+MKcmXwNyYA85no8NJwkkA9MefVDNuFrTfLaeUr9baZgZXD8fvo7iqEo
28nWCnIzVMMOy8wb2NkUcTqmzoR9ZqktBAudKWp8gHX7aM5ShrD15brUEs/BoEhL/RV2i03FUnF4
uMipbSU7IVYIF5FuK+hRmaItdw6L8qouqRYpqqjOfit79rRM0HJgtU7chAyzF+bhTjYNBrXTV1VN
tAWgES1csDsbVPWX8nw8v8PPbMniFLk9CaQ3YCJb6X/72PT/5AhQwY18l4NmisDeMDL80GomQT4Y
zMhQsfTbpowp0OQsZIqza5NHt4mycaBWFBAHVV/4q6yxhkzASbcc8S9X65wp9w9o+1YtjJVd7rlS
mv2zDTrxF3hdxVWrqFnxI3RJ995LVe/xO5oax3wvSF4qpMyfYZ6x/XPGi6c3K4qyqn7ZARDX5nb9
VSgjnbi2kERRYnTDBLAt5Hn4wCxeCwkr/Aw5AwnLfzu+NcgPZIpG/8X6Xx01JVp8NHEmgZw5g3Fi
cHVSQOR62Dn8FfLJnwWnuX9ETlCh9JPtYlz+I/1pQbzgAicBLgBqtSuerWAW2K6XlE5Xq4mIXexP
4HLjHBvjrVB3ENDHLNvVT00Vp8Z/54MJ2Yd4G2k/oJDZUBW2ZbvgG/CaVQYYfG1dd80osSRjE7HJ
wUtOCmysmzqixvJpe5I6fXThglKnyhVwoMxwULyHiQtkg0QO3HiAG8Maw05Eil5b0geu7QgHJKNm
NJdkF4uQL5bOjy/M29ZLwyZv4uNoGUcH6qa0L5wBsUaWVd/nX5Sw5txDvAplPcPY/NRhtHwxer2g
QIVn7qu5y2u1QBaG8yVBNa54PhT7js3RKSVlGI+yA025XdJfm3nyO3gAOM0ehaUn2phzLNhdNHw6
MICZ4X4miao/Mg+iRTQQT1grwZOOUjUchC86XvotXX7KCFqrgAd08wzBPx5Rf/4XQVaX+M0ImGwS
doFIvHo3D64f+kgmcsi9LpfIilBKRLtnKn0W1YPWr23b7CCgVc9K0ZZMB2HlGzw+tclO/lrAbt3m
DmkwUrZMWCq84rWV0n++RS/JtpuEgnU2Stof/i3NEsCxo9zHiY0NqxHE8azntfeoywVivu/smAjE
joinkZsk7GQvHlolTLXoWk34rCrt8qOVhxtWrK+DxwYtISZwux7IZtJdP5z0hh7AGlxH2h8t3pOX
bvUpIE8WZc0pZfUIB+0gdvP27eRv1bNq59O6Am2bEbFDmEwZmPeoU2PXBFZ0NniBQaXpCAUiineU
k8nns34nMDXf8Jqf5HicCoZeUSQ1p5N5/V1bPK2hMv1z2iRkb+zTIumiYJ+oMEapzaORJTDCANHZ
jCwuI/9i26IodT/jnVWwgVLvCoclINvKZUxlqa5PYnEshVRYTtMKkzyQrLosMt2dIqHvSg1EILvv
GZ/OWwJ3/vQ3p/Cyh6zG9+oUNfmHR17iR5Rg62ZcM53fRJUTptTnmv9I4X0/MTKLXMLVNLIX9j7m
aIa57/CHAj2ooMEsRd6+V/YroHfPre0sovKE+E7nbd6WKcO38d/gRjMNwm8QcvqmmfoAAofNdZCL
9ipYTY2njUW5nKzEWBP9AzsMf7KikMn+ivpA6RjpV8ocFS2hNIjvCgymXl+VDjyl6ZcNqmt7B0NS
tBc9aVIHATKk/zzlUDhbNeSAQe9fKGt+uiskPBZbNjAVNwc8QGHd4GrunIV8G1JmlILG8nd1BlVj
LQkOJdQZnWgQm04cDP2lAE1DlvwDuBBxcFfoLwCyQYAvHmj7hY3e35WhxEjiKOb5xQjipiWMkLIQ
NNolyBASi0dTio32oPCvG40J4dSQB9kakkT/Vu9QN+zys0zeBjOtARY+OOrPxcGwkVpHAUviQGpm
ZT9mUd38YPBXnL4P6yn9yu83NSKXf/UijANh7eASTWDs7mK0m8SvGzs2SHRuXaNLop85WgDOsY1a
XrHybCz//U57sT6SVnKy6MKSRYpJcc63TCktjg8QH5LJDakQl3EVvIT2ph85NajgpbplD8psWOT1
EcO1IntPtJgjhJe6KbuU0L+VxsNgk2oMB+VnRIaJCWiMr2cRRv76zcBJxXgl+xhdhuShAKpgRuUP
OwLebYGkXXbDzMmL3HDCwf3Zdx8CaE8GbYlqb6ygZA2RYEaIHiWU3SBgqYjeCLZhlMupvaJvlOUY
xRgiwd8QUWVs5KORDjj93CcxGy+ZUP0mrfdzjT1ySfPrZP45AJoMOTNiEZJ8IHsab5UnvbNCNyqg
LQEVzni/M0s5Lg9FU2+zHcIeTSsRHbdWgdlhEtbPJxd0dL6TfHie+Yk50L5KSRaLx6+OFAMBbOGR
+5bWLofkl2+uK+PDJu2MlAm8E8q99557o6vdabSIKgWtH7maGjpOD+Cnq28Krzh2Wh4Euk42z6b/
gj2zs5VrrtWX5JlZs8P1cU3Q3VHrEoz8zxDIq34bfdp0FRRpfjWTSv/7TRUdfAzbMskXOtDkRwlH
oTjxfaL3rV3GxBKMZSPCo2NkPZjb8rxQvRc2cNGyrq9fP/9qZphbmJ8GFE/FG/MyCidHu78j5HFg
NLYKgGcIXGOrh3i4bUsph8+pQ9yBgKkDfgw9zAr10uKCsLmyKoz6hrBxiQRcdZ4WrE8KzNU5ePZh
1+uVddGbOmqhLcMh7WzKLim3ZO4YPezHk0YAgjkiuaiFDzybt7GVblVe1/tVpIGvvLZUVl7e+qVQ
QQQC/+Yi9zwsVEKDXmJdUI3V99BIVvIjE+PD6zAFdKx+8zJ111qamU22BwVLIHV9eIo0m/mmy4gl
RnyzkQmWwFkn2tQMpr/mvKoBUNdS1hMzjzAejsE817n55mfLhoHtJ0etiL3wQGxmQtzZmt45FXPd
oKRgI1XtjRs6qpFSeQZuNod2O0YyrdKvw7Q2cE49d5Sx9wlu5233ezjnDkXS5qh+BdliG2XbQFkg
ZfSiOfLDxsBg4VZVeyDys3G7jqhL/U8wcsyOfw/QkSNqitg33pKCPJZSswPo/EkVTlOkFe2M+UMZ
0TzbWTYPgRfIELu4TfV3qXZxWoMFHPweXXY+1+KUKZqC4BjiYqqTKoa9oJNqOuNjejJKCGQZctVm
SOmzceYt75pF5EAJBuuTkQMtFQ6/gq7ihLhZU3BlaGqQGfQA4EOZaAQvZKSYpBsEPUm4esDKbU0j
fwhnOjI8XXLcE4zU11nO1B/BANd/bRxl27uHWa5nlXO5xN06SPQyNDlTZslWLPH/YjydeZnTzP6a
Zzb+0xG9ZvgRVv/tMjg65kyX8HqLVltbuH751QWDqxN+UBVOuzexVN2duYxVyOau+zKZYPTiPrK8
E0K5oW3/HHk/svdgMB5gtrL1X1hPHfaUmf6HlaFs9lH2aEmOszwqh+Pisy6aQwo1Rru5Y5z3XrWv
NxPgNUVTWbXSWWd30f6rpG7MeAGmLV1YyihvrcQQ6/Sku0bV3FD5V8KLtHwYmrWdcHN9yIdzUWa6
KwKbdG/IS76q/eDtZE0UO/clVmBjj+ATtE8ThImFDa54pbqGS1t9ZAGhfCrC7uvOY+4/zqwiOPjh
SOXH7RYz5C6622JgKMSStc7wzqX7VXBQez3eOxCZ1rcjpb0fwuHgDxIA/b5gkKps6kG1t2XpqEgl
GD4jybZPe6a1TBwGRBUMJeDl9YFX822GVsz1jXfuL9jez0Fz4wsZ+6hu9YI5wUiH7KORfUMEQ3Iy
btsqCZbPEyAphX/iTUcDO1zb3SOTXJwtTjLlBQrj1cxSO+jhXdmDmwotyctKwcwjtLDPmj/qDVN1
SJNkG1bA1WnS6mZWaO4kjEQpCc5NXgr7SMiNdrLVM2OYZSL20qYz+3HWVRNHI87tvHX+VYxibshd
PrhQizjVnzf5ls0NcycZvTi7vsqHQqWRxXlddVxY79HBLbGSf+b82MZVC9EQZsN2RTWoFl4Dt+6P
d4Pf/BJiJZjC/ClccheQ+N7OJJZ5FmqqobvwpqOqoUE/zVkwf4pE4YgFeSSQ4wyFerZP6rfS/Z9S
JgNX6zBhqWNw/NULdbyytFkOdFYFrrebkDVeIiJqDPbmSUbPDpGyh8dHsSVm1vs1brVF8Ohxay12
YdhMCUafHiYoXxjf7eedhy3RSGLAie/+7XmGfkZENHFk5cbk0V0YuhzJtkxTXuxzYT1oSFFr/+Xt
en9qJINYiEmD3DUttbCx+eZ7wkSYH+sKyD+v704T3wPLgitL/av8s/wFPFoHPjGIPr3/ec0SH/L4
0AcHDJyhayDk6MdzSxtg7XiVehIq1Tz+DaR0DgK/WpBgIP4P9IhyiFVWzHM4HzkAsk7n6VgwNFy/
XWgQJt+0SE3Hs9l4IuCnLNq7FY7VB8Bi/UOOF4k9qdPH3s6ym0TvrNVT7D/KxTFKIei8/FHdELoR
HNJcmPPhfwM3RCejbLjV1TVwk7kvmKtkp5+cyVSHlSfqtSJnYNqKV+w3piiX6PFe+JMjDO244QpU
7Oh+jcIq0hFw9mI2mvOnwWhhSiXvcelooiDGzb31VenEb9kzg2ONdZJhH6WDsFUwSUmXvmMQEdAy
3H7VQOrYPh5/9KxaAYMyWwMzT5lKGTbE5U+0zgMwsMRt4DvO5J1Ds/qJGzprOXvtnaNmblUTSYx+
7LGwjXdsdo2CbPddxsLdxRC727xjfgYFI/IApDoS0DJMphY6OvjSife/xXCGRYQlIypPL7+gxNMt
N0GTrucz3StFbsg8EpWfZckbH+Is9rrfW1ZNdxmWiNAQugxHCBsxM/uCbpOOXo+0ysxQkn3H9Uf8
Ub3VxUCGU4ZL5BIcoNB1jSIwthlYOv6RT5QBzzzi17rokbEGEJy+7iqXjwkO2rUI8skCb2vCf6PG
Zo537kICBjrdLqlRPDXtEgyAcINM+0ZFrsHv63PKN9zE+qxOPowIETFHI7DY6jSGc+/fXQtBpH0z
zi77V/pPLJB0J+wjYzg1yYqtJsKAMMMi8E4OJzGlxf0ARUjyVtAS6CIXba8WLPCzqyYiu+/KXz6O
9p2rXt1Gaq+/pE5I3vKWrvr+qb12kcxLc5u5OhrE3D1wzfO8+r7uEnDzHTGyINPDiry/e0ErSQWa
gU80gG0Icdsei1hCeg61Vqo6Kej+YxS8Oc/cj0ohorlP1YH6WkBIp9Ta+u2u3H/J+B/PtTdhnv2s
gNWYwb8sq+H1arqfM5mpcAVG611wgJh71M6l0TMlEcK8S0GG56Q7Q6j6mlGqR27ls4cDwneLOD4f
lDWG5/5uBF34E1oclA3EnpoBct5kmIMNBmvfaIY44cLJ5+toYS1WnJyayI7cIxUQcZKuCeaf4DZT
FNkg90QfnKlOQFs5Me8QiY/hWIX1S81ic3IVR8JqZgJYt253Dj0db4UJtZ+7IGX7q3YdhMQeQ0p7
22EBu9yHBdhtC7zX8cjbSqnGR2G8EyPjqWwzw+boQ6DymvUCIzuFm9MgWi30LglbgQIqA98vbygB
W3hfSCPYbKYIFvmAhtnMLaInl2D4D22i9CQrVFQ/xPZPXvmqKVLr3xeUmycYuVI/8Z/7Do9NMkWO
cOMLS2z8nvNlarjhqWEgQBhXQJ/FcKNECso59xXUEZendKeGfdmbDgD/DGNAM5IrLDZmQu0L91vJ
ikW4bCpMyha4lUvZaiIE2A915AkRL7Us1d4ZoDLVe+Vwi7Z/+Fi8AHgNmXaKNx0tFDv5rWYkI8cU
G+LLkDZd75YoGcgw46lgtyYyei0syZWviybzLnOT85fKXAWZBIl3vvPnApgB5Mx/xmf9rDQbWf7L
B/Cd5fIxTE/GoVu+uSE0GVmXjzZ+OO1ZRCtX4uNelGWB1D8bOxXOTO4zGiT2zWNKViE+syutiNJA
LQw/3oluJ7ojQ4GhXSoghbS1ilBGowYgldxEP/lk9MSA3PR7SXQOEH5wXlXPNz8OjyazLhdczhvb
AudOVeQTe4gvxmB20JrLSI9bE9RNh9qAQVMm53Ese9do5uDaWF+WCNTrD4PWXoeokPWU6MR91Y7b
hc3Jlm5X4qyksswnh+jujyVqwrtg81D2AcTLQlVf5ttRdGljruNN0bkFg7oBgzslHcVIIbMP50fP
FBh/EWemxiL3HynXHCJHQycIl6QyDTR/dFi8jQoVQT0ZpioyULf2z2+0sUDQRkiDq8Q0MWBPD5dX
sc9wbnIl8Ibmhg3+tQzLY5fPQ49m7sHh9uKPFMbqZqlPWWeKoVAR/D70LhCLp7hMCJshhO+f7y+Z
KQg0J35PzgtS++FZ5Eta9nmmSYgtZlsek/S9e9Yd8wwWKBxwD7cq5oeQGm3Th17fM3ON+V3PgRnU
pOMDqQzk1UYDHKlqdjcX76v7BcSD4miq4Ob8EWn2JFwI4oFVGGf70l9XVqNZckpou8wYiV/ACj7W
TCE5r3UVdVFYpS0Rp3xdLxqt10HeRPYQKNRUfmBNNZpr1KWxEaUSzOJEyGzuFNi7FL8DzawmUxbr
siWFSpKf55l370h5D/7xV63x2mKUatkyeA7NVWUEXyKz6Ge4HSH1NveKwEcyC8o/DGy8gfpVBvHN
qRsjvSEc62rZJc2DNBpn28J2M1U5UNLpqm7vKrTvAtCLgbzwOF9r4Ww0sCuiEHUl1fHW81PpMeWZ
yVjDqJp93lomeiHNA6Ye/eeveJOtdtHTtr7vIJUgAcDl64ilBhTLr7BjM05m6jS0HGrmRUJ154TU
KleLwVBLV959wyko52ILxAmIuqGQdiQAkdjbxNrDB9lXsZ6XLNxRjzwIt7FvsD94in7lzBu5cJi8
M6j0l0MH2YZM/yam6l7lz9Jzx8HN1YZD4AyTm++1o5jbzwGQs3aPTO/6hvObC8sCHyIdAda5O0pJ
EgQJXYYpdnG/0UoeR0fiA5CLLMTOxWWSlVaKX2k2rC+I4K6815h9ftSJeZDK2o05oR4tIsAzRgP4
ycBg4z4CpOF7vJ4FXjCE+wAX1YuRmOoq9RoBbBKuMD/bd3Ae/cA0ckf9tz5LIros9Zzp7NRXmJKm
+KSayWu+HSGkX7YhT/u5b/DduWXRXf/Addf/Gj2wwOTrSregTy5tYLDpV0gfRfBuK73VZYfESCYB
GiKJO28/1dXEkk7bnC0G6/t1WNXBgaNuvYEzJ3j+fA6EmQPS8LrfTEG77CfjFKQnPZ+Gi6lfVQuJ
zSqOdmFU9P2nqd+8F1WkfgQYXkACjwp5AE0PHw+EOu6OEURmmayqZe8zAOuBFPB6wkXXJ5GxWBqa
zopMnrWzMOQefQ6qdU8EEFmD18llddJH/ERwza9DQPRBU0gX5Ysn9varfc5aWKPLrOSOgubsj37d
pDmjkVSm74BnsB25xQr/PoDVfMPHyyodmZBEO9SmULb3B7m+pQFCyNYXESWR9qSeK0bJ3/oqRnRl
4CJg/LYstG40/g6qBIClzcagGDRrcfMkMwX5c3BdAuKimsG1n+GNkJdHR8JCjhDYH8YJR5+oY6sB
1Hpi07tiweMK1Fr3N2RjKXxJSrraxMBQcpyjhWegobVz0nqSweVobJ5P13oGuYtXGUCz0XJK96PD
iAQuwmzB+ICMs4SZ2jF2x3X5XXUTqBbSy/CFYKBYwXLb3Y3Xau1Yn2jR8g/HNBstXJfkcSYNirol
+E5tECO+MIyaC9Tn6serUpsvhmS5WL9w1hl6cbjMK+J/N6Juaiza4/+XLrvD4Sb0Wl1gA/fYRvyB
WxWTkZp9wJlcyGFjXxktB6w2k6WlZaNLcS2SgEv9S4knaBHknon5dtweM7B4JgTDfGU1khWBJV95
1bpaDUNET/Taz73WNN5pdvltdOnUi3qRgjn6hVCEOn2jK0X0ObYPPeBnB6o23SJM9bNXl0CiBFJA
Tb6GjTGYsPtVnFnNIa0QuPVKG3tLkVCbVLnBS1Zy/c2XPBrQVXGqZ2FqtC8RLLKT8VkTZCestaTr
waJ0WhBuJjvPSnGc3F6oBXb7QRmsoFOA69iz2n1Vrzl49j+VOBq5Ux9J9FzIbsr4p9JPMrUCHKiR
YyxUXhhRjnVqOSBxganvpPkBRUHDGTXRdLC3GmwjFvCi4VM6gzFKuZ2IC9i2RzcxvVM+2pzsm7xM
AxVMOhbnP2fHUFLbygawutHOR3VolEYfhlYKHgnEerh+h9tkgYbncDcM4e9quBVa7lyb4zhl2Vs7
KtbT+fJLEwaW+0IiOrqtg50PRSTeKr57bulDau6S+QacLVNYC0ixZilYhPforDea0t/PmSqd9vM4
4WcuLxQVKR9cSzSphxsy35IKw3fmojbRmsq+9VXvHezn1CwQGMqJSfnMXyVFkOYFtIsER/LXX+eo
pJjWBphiwLLtwFbTSwP6lXzyDmz0G+2kaxf+rsXXaEjMaeLWKdvBflFEaIXKnRM/TIYdZnpWpn6f
nGbw2IELHdgvGd0sbhB4cSx6wE448yLhz2YSX0ytxk+nRUW4uTRziTf0wqAypCVBlcfepbFe8bBZ
iHG8sLM3blYJdQOQzNjfLDWSH7KQjVyOfr8O9b94tjvBlnrCBTpK4qbAD4hPTFu95wPVpdqq+612
L2/qNJqJeOhZ0ROso3dpQoTjPi9W5gMUXh3Jco+72uVen63/7a7/sNztlpfiIecjbfcAkoS8kJAp
XRmmeswB3aQDfwYT1HCK6pE8fLFiZde3qLQIalxaZTGUv7R8bfWW144YsjEu1Y8h08Z5er9xFpWs
+t6twh0h0csX+d+wkfH+OpAH357+XQIaxDIca4kgbfwFWjJKjnq7T5MUsj6xXQv7Pgkiil/NvbO8
45Y9UIl1vlFtoYgoBtCGOlEJDELNndfhZrZGnmtQ7Bin7lP1JkPNAYkX8n6c0LS18Oz0XnqMO+Ou
/XRjd104IoI4S1gFQQ+0i1sjh3GJ4V6q23U0tWa9XAkuiChUfXKWAtNuNNO35bYsnTSmS9utPqjP
FJa1iXij5t1rv4MOxIKU6UuSS3IWsozVkb7HG5yytEfhUxbk+CioTMLN9U8zRKniTMqWf/Lo/mcV
EfwTrGEu+6xR13ZaV2Pi017Vv2j3wZ/b1WAL24r7z+zuBonprVMClK/wlPIwvIQ5ew/CepHWXSna
DfvxdE8VAQf3LVr007GAmCwpHMh5gHdbkOvMuxvb4XKAuvUYpR/K3hgy3vT+KfqGO8wHRWg0mLKg
Z7qnalbcYHoJL0J3xu/JKDuZ0BhitwZ7z//QxaAGPX6kSRfu/GtCJM/YwBujEAdascqSsDao6ts1
VR7ELempo2rMmSCkFFp69+ZZ2qm73VnHFPRc0BxI1QnaMRhuCDnNGJdQ8qkzvpEu5MTE4yIgwwMF
5TRCIwK0ZHObmIh+SE44qIo8bMZKLunASuM/KSJpx1ZCS7yQ7lbjudmwCzTIX6g4AYJnZIF/J2yq
QkpXQk9BTV0tkbieoUroBOfLGR3oWlh74NkS6Dctt2oOlXzdnGEXvwNDnNvNQ63Y2QnNF4caixeV
ukiDWgfnAWx7eP+fku/UNrmLaH3o5YA6+B7O2NAhWn1CImYvMxP9ZT14g0cbrl5N6SDJ5qlMAwLE
HifnmWPaixM086lPqDYid4Zg9b2wX4at4oxXUXLWD5obKJPlEVz+8GRwZvInQXsmDsr2BXMF3oPR
gfsqzBCGUHhRtR5RwDgL8MTGcA5HQ0bSSmxqssKVaX5YHZhvLoQsA0HqBvxDk+R8sAQDAXqhHDoA
53/7ZhX2+amGJ6FzPB9yjNHO85hcMjbhRwG/1Az/c61S3FMxt9u6xmSYvIwlRRdXyt0xOix4QUo8
cJlGUn9DrHY+E6tL9Fj5l6RqZ7A9jzEYtUG7KWSItxVXYaM6zfGA2Fut3k6MfXxZJ4KGWKdRfCQt
dbuENhpOvKCMps70d/HBxlr+bQWrzP1u7C8mh5Z05FK4a95ASOIemLQTZYqZ2hykmqwBa9O5uIqd
DJHy/uWCZp96bG7PxwB+U97V1fIga6T/vBspMGOiwQ3kDDzilwQq9qRjd8BjNA5/Bl6Am1ElZV2+
bGsx9NPF7MneolempPmyXTf7c2v8GJsbuD0S7YwG95cD7PP1tf8m1cf76R6VSbrj6fm+xws7rm2H
0p3GZPxLuhJAiR+10qn7yCOL12HfhMuFr8vsOYvgBJ5lHIJQ8D+yP3jO58TT/S4LxzxWtOst/rGM
/Hdsx5ZltlBQPqoD18Gs32EzbDZHeFDIx2Umn8lmfehj1PCb6H4MIIIGDfJSrxb1LBF4Ox6CdGhz
qX8uHiBpzKfDjkXZkgfyunxpYklgVV+90XK0QJGxjfmH7d8A3oiosOEKPj17Lt+gmwtXwXRR7Q5d
8ANRX6Pem03ZICiac0wqiKCbcQmxsFYBo/jlylAU7bYu8hUL0A1onE7kkWfmaEtmBG0L4ocdgNOx
dqSyVOxihGt7ULfZh+opaFrQQtyGAVzNBJ71WdbIx694AC+LTa41n9V7TDR8ENa5vA76NBkmKpL6
wf+ZXHmwBl6htQpwx51fRo9at5zXn4hQdgoLCwuTSsnNQDMNHjgBvxTriuC9d26mzuXiYLw7hZZs
TZNsuGMDiDahXz0DpxakbHsl79Tb+E+mzeoibxF9z78gR69z6kvp1f92ZtVb4kWi4qp2ajaRlfLz
+MULMSKmmmeT/jj8+lEWmWVFQafjzVl77sptDCsytdcfsTTVfJru/4ceVltL9cMMXpmnd6PaontD
yC7HaABsSMbg6sOTIxCp3PGpr1Rt8rSvQSyVFEgmy28M1RzJMaL/tjEGpoaDghujliX0wT1zBPhS
/HZS8xWl1LdqCy9sLFE9gDbXM9fQLBcMD1XauJm9veyEKTEhbyVUZMS747VPanavqiz72LLl873s
qprPumr7zHFytZAF1YGvj1q67Z4BnE7FtPWFOIqBj9EwgunumWi7vhB9OjTQmlKKyshCaJSS7sPT
NcRNX4GBgknoMFWpVGNgtfy8uCTp1oiBt5E5dzWpTuvG+ixilg2XBPmWpp72YvmHoQkzWvOSziLU
2l7ly93+S3AQXRlJ11AWJt1DOEx/d6UNkR/F5wgXUIlyeMm+ihmOB6rd3io43Mtph6KclAAzsfGF
vmMXIOGxx8zGAZsMH3bYsvp7A+I8FRb5PZccPCMWLIazlecdfCSVicQzoJTuxB06dL2HkZb3oi7E
STLM4EKpXhj9AzcySnsu5A9SoPKHly4bRsJlj+YByUP2Nm4O4R9YOSaoh/BR5V+RH52BC3Hs0iAJ
SCeOfSV2YRRmtJjlPQoaq+qE0WyKaV4jOblKJQYbuiufk/d0btELnApw18zm2JLRLQHt1gDl4e4U
jVRuBfd6SB7ITEJyf04rUmMajkZGq6GK7vwQ/xkT63Sg2nuP56NBGVTqxeP3yHhOwwmWwSi187XQ
f0F85lXzZvPye2utfenLW85xTk8w1ul1vNeI72JmU3+e8tV8QuXj9xrDuuAx3KzObW6ayInNSJcH
K4NL5gUGTIlYxvZ2cY9mZmOTf4fKOUXfsYy4p+ja9cG2Q/yWWfaIa06x3FCil50py9jQMni8V1bR
vD5UWz+bxCc7SCIF2u1gqm/sbSxnDhvKqpreAPNqzsWOF1zMr5v90+PNm3mxGaFAyKltyouJrMXO
lcSeN4DtMyS7S9Yd9U3t7W1eV5CXp9M7WTtOK7b53qjo1L3vp4YUKatzTghdSdrw6Va/rZ/xvmrQ
vRebwJs2LuunU/O8ntgbr6ptkavfb23GJW+OO99qDJSLQhpDlDH2NTyl8qDrb0cmzDwtWBTZUUkn
xyb3i1mDaOa5JrEWPQggigPuMewcfKEREQR9k9epvTfek85Gy/RwTSTeaOIiF2AMQGh2oCu7uJpn
1YGCZeKOG5nldrcjo6dhUmNNfSqtwDQr9CJFYw7zgU5H1ctsYbf1juA/Eh3xsFHqrYkLeEOBnFL1
v/l2Am+TgpU0sZ3J6TN+EtaoAm/E0IrEx7owLoliVOWfMZiuzAu9dw3roWZb9rxmNPMkOh/CwxkF
EbkBEkgWZIEn35DSx9E6nMbFF00toRKmAu0kRj9eWb0Sn5IZ1UbBykb3NFBfIv7g4GrfCNKbQB0W
gWGIFjHbHjxPtguURJ8S6kRm+k8klvv/1dSpgkHov9hSSxZpfyNwHuUn64DdMSJx1/I2G+WRil/h
6f/ar1HjZSjAGFvtastfF6JGEMhdR+TgpjjM0gdvd2PqQVKuazB2jrw7W7sANwgg+mpvVzt++n8y
CZpGO8Js0eN/kCxyRmPT3WLMStgc1eH5gKDMJWPSJHm06IedWnVWHbLo6RRoZMnpSUyooisVb7BJ
ETQO1q/dtjPMoYYMK2HpaE8JBfvAJqSssQzMH54Pz0XFPY/5xfTns8qnKI+5oaHxYgUlV2Hqe4oP
E8O/pm4uuV0CHIBmia0TG/kX96MZS4VY7YrIP/vC35ihMsRN1dk+IEnpWIloq0Fbt0h0B5X/O37q
B225xIuTJIl5mTLNv+AdDmaOT8yNkKl78I0+PlPWIRLvjrbHIduOYUDcKtfkRhU5v97ZJQJ7lQod
35lp/+mbX+LLX22rjBuMrL50iYIOoYNWt8wBQ1aTyekvzMt7hiuLaIohWpqFdudBdMYzcD3vyqi2
qweMVKLtaMh0HUOwdiSqs1dvoZRBWiTPtvqheQftLUKM7ERRkUfYKBxw+322E2Val/frDB6eNun/
XRwq/7pXY2vatC6ujliKnnT2EYRyduu8dKYz4Hv/HmIUkavPiEcgLMTAH9QNHeHDqqI3Av3IGDyY
D0Sh7EVyLlhFvAT7728pcZLGKdkluCxQNBuXX+fAyM1XfFOWUmLB6VoIbmm3ZjFjC+qgq1PVjeOj
3XasdPdVOPmKYxCq5z9Fkrcm5MGNNsspWpbEtrJfmrWGJZj9tcvoFrvBZVbaG5DImIHvH2JgI/YP
FEf28CH0Wlf0FMeeqR8rQTNbURJe8YCbxSbfJOrW/Q4WWUt20wS8XJyFh28HfbX7K+YXOH5atdAp
g7vvpPIpcwEjDeozSIl1CeFzFlNQpsDkPDHmg6H5G2vpCBd4DADayMnJCdxaEkUXAi2h2atKy7o3
KvIJ252SDAcsGcLfF/JK2dC/fH20lStRhTtdZgzE1nPg0jttksC3jPyhCgcaNEfjjPa9AvSTTh96
6u4GSfImg2G6jpErNj81cP2Ue35E0kigHsUCPHz43nDgWz/qONNBtAy6FV5kLYzRW9hkSsGksUEb
x7A2fVU93zwKt5H7Ca7iCAukdr2YgtCMEo1U7zTHkHAYO+BZkhoHko7g0fYqRH/pJd2to7DOHjZy
bbH0yyMrRDbKKPnUo3+KBXuLo6WL3qbhZZ1jcS+O9emlunxKGduPAQICLIazqXokLnS9NLGuVdA3
A//dS3Wp00B9qzkkXnaPIZJxFjeLDW4PxmlzgERHkzDZN3oYA2enZcJPHhFWoAWNBi1+lA/Rm6nP
Mz8GWPVH7eMsZYRnq5EcLw3cx1bWfDUxMTaeibWlrtju/XZz5VAy/voQFUqaReFqbqwiUTFXRoLx
KE0hry0rVjLu1AA3+++VcAOjL67vcrU8jaeBmjtakskHNqiBugPxqGPtmqumErHe3yA11cIrHqyL
9302cqbhtXpqbVpjfDLqfm2eTTsCQ12Wh8uppDbaPkImbpaNy+VUlZ7guHO1/1gnENSeZnN+pAT3
2HH8YvqB/8+fwSTgehIUpOlb61QKFazK4jq/uJX6sI0XyNJWBYseAKHsvodKXssGf1f9GHWt9x0c
ner0rj1ES8jkLECYpz6LleBXjAIMBgKXa9tgNPjQKLN92NlGHPy4VlWfSLKIV+TnBpltGyJnJ8Cp
Dspi9u3KYwKbaL3FxPcN73WyWSL0v9VrmWzPHOwXjrCqZ+fydnde6rvVPdSwrFe3JbINGTP2W+1z
i5rX1vgT7REm8ttVsZ/aRMwePAKSVYMg+gTzX9KpmtecGodIvdi/5bkRPnaOZbi2sTNkBksXO1ko
QRwnZGT3OASeh6PKHUez1o6j3LzpRl5a774GSffasm/T25O1b26OdxSRqFnDk58pt0V1apjXP1H8
YgPWdvhb/CeI7Jp0jnTACIyksW94yfIEU6hjTKF7mLHQI3V4/AqThSYlFwA8ls0yAhKwNtcTaA4i
S3bZ02JekKMqRk8jtuXqqSeQOmy+Nv73436gw3JuU369tgN81oGAHXcBgGiQ3NmgVUSH/wK/Kh4K
MGBFJ1YbJJz64VkgVSg5PpJyPsT7qtvualUF5QaffxG3kYnAb+nSx97Mum/qoB+JsvbAb3YDNYjY
8GTaXD81JPQ9ZhJzC0qp9cTA8Qy2J7qmY32hGTB2BlJM/sCQ/CoVihGpqHe0EylRFSaLF7TzwqO5
jdC2Gx+/cwwZzjocRqZLEBOu8M1gFdQ0OsCZ5i+lVfQOMF6lH0pBNnpzUOKD05xf2ICIYZmUl15Q
vaCW9tmNOJQ09V99INjI9Zmw8PHJpdf23pVHz/1jfc2mJTmgNh5F1WZlMIUQIewqYczj1cIMU9fg
nQMPQ1XZGYtFZGad1L9GsfKVerqDw4u3g2HV5uWIGf4ShT6cqj71DFbG9ljfiSLGlQpCu11FGL9h
kr57o4O7PG/PCdiz5d4OnlZ9rqNq+gYMOAwcxK/OQ6zg+0/SIacj83MhsMg0j1oAyrCFJvDz/LzI
OmuQFYVVnHjVVLYZ/rNg4ByTuJlxML5IhEj05fKseLmLZBsjEV0Uja+qIiQ/Az4Bs4CVUnfFgl6B
7iK3X+NqYga+DPzUBj+LZf/NcJgwWQ5UytDvy3x0f5htjSpCRvwmdwWOIdO0SuEl0O62a65loy6v
MJSC1xi+w/7kiLfjJnQSx7a1vz7AxgnDmN3oniY+Omx2Q7fLFVTT5D6bLNmfQ0IWUtuctNmqunhe
ZSbPFT3tzXK+7rOixn+p4VSjCCWwNqCSDJtg4oQpuMIcx7ZAYO2Llgr5Kn+9w94WgWNuWqsqJS0B
a2KIkINltma2Fg8srkxJuOFKOtEIC/vO//47bc7dZe+PCB2RT71teSwCvyrwmmvlpl1Dc+kcp4dv
lRFMVoxgrjJ57LVfGuxG+q0UaajAIeRL9rUJo1WRaSg32DLzgpuGgqwgFznZP7DtruUBxoLmnRJO
jhYVjBZ28sMQaEu/Q6AQGK2ueu4Vs7H6Ip2fScrRIGo+/nRorn3Hcc/LEVtYSH7vPSxYYYsWcdab
ebsw9FLNQLSkkmwg2Tt6JEarc5lLqIoXIKzseAd5VuQztZYIyUIzG8bc+XNm5ekfLzakYgoPs5tU
4T5KN3yxczLtaaIKr54gI+/Quoh7yxjf4pSIM0V4hYocMSOGoCKTMlaPc+/r/kelwAbO7XgvwuMC
iEoBWCp87+EEjyw2HL+cSl/pN3zW5nyU2zee+g7IP962/4Vra/rRVWW4QS6wzgJLfkBS+nRpzqXW
0oTkmS5LzBijetkWwRr0NKCd08/n8iF5JQqKq7blMoKtttcBZgJL2YsJRcyU/6zol7IEy8G/oA/K
Hc4mQ3OxFMIw12oo/Z+TossIAuefynFZkWQWc1tJz6GqES6v5A5WkFC1QL+wfZww58/QvdnXPPlu
x32UhGFX6iEniQEyd6ypMgar6qV1ApAvmW7iZfvEsZ108DkkpwtAXOIFI9btKzQegxAsKRoIae4K
b2QSbqdfWL0ZMWBxL3zmlSjLpFBsV8HamfpwiLRJKyn6rsvEHtNS0Iq3YN70/LvqUhs6w1+j9oNd
pZZTWv6M515LaA6PnX3nTGB4Bqm6nDdLt4So+6s90w/wu9C+5WDit2L0Cu2gkHcKt627/fFL1h/k
ntoURKkmx1shIWyzYOr2XjHG0R5NZKUIabA2K1DStnqU8OsDRCWj7GwRUv1hL8MJaIbu37TLhONY
376mXFJGfGi3VXGW5IoTJSMLWTaGM7ZoM33+GIcOkGO8DayPGJRueFlSAjqwNXeCT0cuA9fQGyQc
9ep8tieaFi73uNXAIbGPyxRciv4WJpibk/MPdCFCTpcrtFVGMtZt3kEfcDmNPGlbpluiwthuSKBZ
xLJoFoscnQacIiSqXnXE9q7H37wR/I8+znQfr1JfP6Gv6KEwYGRFksrh0LyyHgDlGwSEUb52g9PX
HF60GJ1pstBcjRwLJ4ofx+GVDaoONYYDRwduZjS88DcRXtCoCjyOi6MCrBUbHKyzU9KwyV++jSz2
pGHberQl1K0vyQd2bHTCsj/VPT7m5HoTeSH3gB8ao/0xXPS0yLptAOEV2XtEqhZhvW/I3Z+tdMX8
o7C09hyv9T5lEjuuXsmms+VNyx14lUpRt7If9rgX7zRN59ywMXcUdT5kr2pybVeEPoOQT1yc0Xb+
ojEGOjN+RxIPbVkTiLdLR/CrG0Lhj0jGmmvgnPG4+r9mjLMZ8oAu0TL1o90JBHZ1ojq/yu0CCgRg
PYnpzU4es9RIFsVnrm25n73ltJURLlfyO8Ez9+tZWIOZmE8NYFtKrQ5VzTgMzR7DTht9eK/KYDGZ
iWyCKnG4Ky8IfY/xQvtcuNWlDC99Y7HwO487rBnQhPHn1hGDBFwweEAGgKSv+OhzHYrw57IAhjxM
MSRTiaTtHfn8Iq+A2Kx3B0ffwmxaHcFU9WZW7GulFNB5F49u5THiBT78tpARv35nx0hqG7cyuLQg
J92sc7I99TYHo5r4ADk3n7G8PUvvwDcyLBpn1PbYmC3WYTCQKEJdGzcCcFz3UTsZRSUZpFXKZ5vg
J+HIEpM5s3/6Cc/1QueufSEB1A0FHv1F41DWeuy+s+EsF9qUNUQ1O57G1f+AMCNxM+VwjyiuXtby
XOGwsJpIQPzVOdhudF2bxoSpYGLvhJ+7tfW/GHs460p1uV6mv0BSdGK3PJMhTlpe17Kp3ZH+EjFN
QYCS5Cp4DGJxSg5FlUzlNIVfSXwpvKxAExnctlx3eEXIN+mPZ1BEwCGFO5D1eID4T8uX9z34kbvC
rTINzi+gwGgvrI1tGMuf/svXlh8MGJAnEvcSL6CzS+S8EdMMccjeF260Zx9NCPmtrsU/pyCM2+El
9SsnAByfLLlhpCLycDBBMRP0i3t7x27EI+YPNU5zJYspKGkfKfIoays6/cOajfZ9bIk7EPX59cl4
AhKzDmIpSNYZVdc9ZabbVZkWXFnECiDmaGjaM2o4O8UsEHFcwzsvOsLs2l32bfZOCXWtvox4189R
fSdxveeZz8qZcKzJFPT6Mf7YtAZnmPwEV+y9Btmdg84HmLG1mHiNzL3CD5bwpC/GWkW5Z6e9IVXv
dwfuWmfcKxR5NRVlTQ6hmt2tIXwjF4W/AlWv1xwom2eZOKNuouj80cOmxpBr5pRBUt2bRqPsioq9
GJOYgaASFmzXfNjHPegKlmA+vq9tTcBD2YuHnL3kKZjBJGEZX6V2wHxq3gW2uY+U54MG9JCtqztx
mQ26I8HE6QNmpwLKvuJrIGq7O+PVjINaVtRKLl8SXFj/oXqd8KxDtxxLWKJCIyOrXCjXajO13uQq
HM+Qhs8U3G7GA8w31+AeWWkdhqFNzO3MIpB4+0fJQzIAzSMvKmQ5mh26kK93lSlOMhslOromFsPg
TMakq3KU3bYrb5GUw7cCwUntDaWT2Riksa+qb2bSC1JF45lgibFPHT/+HumXmPl60VA6Vc77C0hq
k3mJJNuUDwQvTOzuqNrmN6XpWlzBqLknXlsFgtEtmu7sB3OmZwlerliylFsdtIXjbc1xQ7Fa3W2u
Mw7snfCRkI627Kfvsg0f9kmpXRT8xgenGxsgTBfr7jEfLObq8njmImdV0DXFf6e+C2UFB03+3CLb
nY5/DGn404ckodaz5pSRFXitsIiceQvCHG2255GimuRHxuCbpBTj0fkXMWXdYuiZZ9BnR1hjEHh5
agJCFu+ZIwaMb+TaUFcXYenc9FKHMuGYgIskAOuZzxT5irQOxObRFjf2hkIWjAmwGkeAAEcqI42g
MckWJio743n9j5tcr92OaB6BqSgBhRlHvFn8tT85LpgQqUKHOen2HgzJmAqejl6yDz9GX/t79QQ/
CFOw07sBC9v5N/c22m/pNAaQk/U8Pbc1J6/kWZ5Uh9i1PjxhbELFJYUGReHbm6HQhozWhSjMCm5I
ezdlq+fYvkPPwme6TcNDoLtMzjZmSvaWb+isqZJ0DsSlVxuwPVDdC1Ssh+aaYh3ITmo4vM6F+1z3
c2efeDU9KsoyItKfLgzjse2DXIY1FVe7ju/HijXxDXy1iY4KZRpdl1qYzrFUpNfdsha1jyRVcnLP
mK7Z8gF++67aFhjSfkJGj/UPasbqphPatvt2LDWrXD0KDladEAanEFGapAFFp9n5gN/iUDq9qzIo
gTwol58fruGs00tx1pkPr/5ou+D5H0QRFjM+GOMnZwlOHmtA7TrRQBMRIvk0JU7hfRtoEjVEgMI4
uJhNHAsyqeIRnlQ/JUqkvfafnQ8+wOHLgElxYD3bU5+HF2yw5DjL0CpwTlQoY3gIsKEqYVvDLL3x
xC7OJVp5D02M4YN7cTjFcCJR8uE7jUGHDqIwAFeCdXB7PLqyDJREUMDIpVUCuYmXAhuIhl0R8MsM
7aEu8LPcn7r5/jJPQGQlWQ2u0x6CVgZpKdszVHhMWvaWkCGGaH1aknw3qw3aVzrRK3jUsh7MOy8f
BsrbIREETkr2JEBJeGbUWmu8bIAWQPGSookH0clUw4FAw38omb8A3ZEBcW2S3QfL7GVbMhB9ofoR
EKvpAHEt1lkkSruG/BXhMsbmKU5dsxY6uTfZkzmwBamXLvkV5HWffM+Qz/950mj12Z4fLgZWj3xU
SjXpWOVxLQB6ahKIhWK6xYAHUpNMLOP08r0m0IQloT+uCmDZ7aunf1GYBF8tRkO7Asx5nBTVfFqH
uEejEpJln1YfChc7u7OfIzSgXZMLzdNoWVacIOu6AhV3skfSDDsP6Sd1Bza0Royb91h0SRFYVZNE
PyLFHZw8fwk1T72KpELd/3K4xXXUmLpX8vI6YQutiRovTwQYblhlNoaOmVFjdj5JpFQEwffj3BP3
umAWjsS1Jss0Ea6lLIkLzeear52jvXYvLya9leMNIxShFuB8vl13qqxtnxJH5ODj0Y8AQxQPUz0J
zdAbw+OyjnkZMNrarJuye1NWBfQaqAlAL8+5WM7DxCvdm0hQPW6OwfsvBB6phWi4OsD0peHfSb+x
Fv+B3ua0WgRd58HvwYTCTUQPknb5w0e91fREDO7p0sYcFyf9AFeGSjynMJiXxL8xxONYDPBGN3rk
CIiDnes14bNspVJjemf84hgUw8QWQ39JRu5ce7DTDfWeNF7R25kzcEcWFSXK8Fbcya5UPLqE0iHu
XG8aaFQaPph4t4Au5IUbquhyU1HD+5FksO/bVla8oZ/xB5iU8e8LKFJ8PCcNxnvzfR1UcJIoOnnb
jfmMhERaD/YDNNPrWKaB2d6aCODFenFg7W9AGqYcZV8eO2GAELKRWNdvMB4XsHnxgtDTyMTnEN4F
WCHeIgLTWauk/bjs1ExY2ZnhZsdxT7FIm2biY66KmNw4pZ3QYmd7wKZ67/D77HMd1REFpbDNjYbW
7oxwdJtYs79Mzybm/bpDor9AFTKxpAHjGj8kiuHfqogIFbPuDPguwPZZt8m7kTT3olmvcATOP4m9
8aaZ5R4LOCJL0ssxfuvJKE5U/hoPB5n2SGmcdIjlHiFHs/Lg91DWMr8/ooBJ+AoPBIzKd3ZTc7VL
rO+anDoDQdQlAknEI2otTLR+UaE7Ejg9WforlnuRhY34J1swjbqcwsXPD4rgMEP/zoBUK1tN9yzM
pgFbWJbIede+tzceCaf8kakOeNqDEh2WgSKzQVJxIIu75gJkANEpn0PiCH5QSnNnxZxRqtVHA/Nk
1g6c9IJ8AVXS7oTSzLXya9YZAbHD3cVekXT6KFbC12WLg6mbstVW8Euw/aT/P6jqfRgAz71PG0hR
4l39TEjtCs/x94hsKymxhHnyeHoMnKWhNueDfC2uiLH1jH2fihp2QrTlwncdBIN5aJaTtKfxc/Bi
0DKkcv0O0BtIXpxvhCVVFoBsZgvHSSYfVzY3KXYN1ROnVtB307VtN2cZtf+/NH6kbbH/X1besjNM
JmYEVd1Ztpf7OGI9rxJYukMNxwVhgf1RXENPRlY/edlUAlBm482mhTu08fL/BAdhBj2Xsqw3LVGN
a5H7Na8cPLZbG8450w46W2FaG8sU6I8YZ6LZkfiqW4Zs23d5RK+QmFpUz12lUCQvPKQ5+O6dujGw
La6SHUKyCb0Qm3rDc7vWjvMVpZzumwXhwt0kZbhu0J/djI9VDq4soMt+mO6c62/gTSzM2hpA1szj
CijzuoKaLE/TtfCVU1sGkrjN+EYD/16nsWw2aW9aKpsX2EwvYx2JaVzNCboX0xJit4/H9iL0NvWf
1dRtIWm73xML2v0ASAe5UopOnDzu79KAEoq7mM5teKRI5xr8U7oA8s69UNclDtpZ6hlqsFs7QaNW
HuZte7n3vtmckgiiqh0N+x5SK0G0GOl4aJC9BA/qP/m0Nh8rH5QiJ5aXiVB/yLHF1evbRJ70pI/X
9oGMKGTKv6qE6KhejtQhzF6rJCfW+sE6v3BNKc1f6KQD9eVKI/prR68Gk9ZujjUzweheQxPYD7J5
M1bJ+sGygMyLvgbls7PG+PvdsWknlXWR0rfr91vJ9kDQ37QF+ezKDaxh3Rq7DwZhUYe360dEOMUp
QCoiqKqIcrkT5J4d+2lX9wrZLccrKgmci+nCH2jIZyAZTW/k/UxaHjaMujd2/+4msyGvRwT1rrD/
q+zCvyhi0J00e1I5qZVgHNqMDlSZm329xGKHUavjw4UeBrM42rqvuj3VMr8HjuxRq/0rL2Ykyt34
vXfQ/48moD6G2pQl/uXQTirvWdYUHV9K+HyYtAuSNQTGVEN1WlH8Oi1l63fgfmTjwsAlTNuVLJew
mZyiPXM+HkQj+I4135ui21THZDiaAigiWBL6WMcSGDLs/cSY3MM6AkeZ4fQeTO/TAaqQoXN02au+
KMKQqThnpmxZUPrj2/tDxCCdUU3ZKLCp5HKDQP6nBlya4cJOf1uzjtxLzw7/tR9MkdvZ+p0NByBg
oYlm7Xgm8csx4cbdUuofk7haLxSzjNWLUMsuteERC8kkfit43OYHyt43zB1P+PHpmp6yLzfCB3ia
uubeRmeMK/um69oLd6uAFPlC5s5/acNyt0JabDREKMU3TfwdCdZ8Mav/WGDH1b4LHw9nDS4+nxK0
9kwBa4ZpY6TeqK/WDUhG0Qo97Y0d/KdhPo/OIvrR5wveQLQwd67PgzCmGWJQo2cT0KFAFy4QusWh
yeCjD0KEkBXMJF3KzQUEGllVzGVJiFw0zFI0KTbm9u5bpOrSt5VGXi0K+mvX32RwfsiLH6sm26+3
PekpOFGxOfbLX1yYYUfArLz87Mj1R2yq++sWEKrGLl4vC9mYP9VEi5ig6LDta2uN3/mktNcrNN3A
p6plV4PzBhvKbhkTcKaqrQW3LbUevNJX7sAAO8olzwRm9yZ1Hmyt0YHwzesgFzbGMh2YY3X8Yqx6
o4Dk+phNR1jfULDgskBg/ytiYsaKOrDfCxkglbMJb4ck9egqRB0Co8HXkR0wY+qmJUCjKW/u5pto
/i6tJJ/SDJALXtTBGqz/RujbK2VDU9RCcrpYnV66q75ugD7aCXT0zKiq3v4JwCF/gLd7tasQVaVP
BqKLWfzeQThgo7qw8TJF6R2zMxBGY2OiyXuwMOdd0Wx+7Qjfn9xdQYHjOHk+ovNh3DqvaBasJzSi
n9N4NkoQLvr4Fqi422fnLiJj8kgBdBHpqaK5qcnRHbDLMaPfnxp5ydmmMo6inc4mM8B4DQYwKr51
YaxzTiBLsaiyS0GPHxPquscSl+h6KVNfdywDLoI3p0Jy9thunRPlHDC4I9hSp9KwvnR2+HGLmtbP
IikC85sES7HIvyvS430WkgojEh1+qF/LzbCNrTo89oR8lqsUpQcJYwGkbpnmhTGmJ5DP95ia+QMx
LgL5ctx1V2OSXW+TWURQP0ODaCC0fr9FBT6OBKzrDSt0tU84enPnKZ3ir4NfGrAvtVR/0toqaCB9
Enf7LQLXAHTh0kOv4Q26cgBI6CRGk23KWML0te/179b1a4belQafGjj8zBKxxCFmcb2l0HqRWMZT
M4yelPqZwhG//XYcfWGixmEUeAIZiUBcWLe9YvV8X+EpLYcr7vb4EHT1FqU+HbKvKZjB8ollCxT+
OvVvnHKwIhxEVS4udAmCb/7eK1CHsUV0dv7cDYhT4y3rSJqPK54dEKuy9rd0FKPRBhrRr4mxTErr
bqD5UYW3Qfl30yT15ozHpydU2bKEhxTCuX5C/D+4P6+1b9E+7AJYrZOUgMUz0CndeKBqMrpNMEhM
uZyoVJ9lZutE+hteU5gUN0x7QObST8nsmHi1lKPo166xtDHyUloHa1OxUZGIwayhMjov4+69Is4W
itzrxb0crD3xH5Ptr2T7o4o/xX+vQzYod3M0C1eTzwZyv1RAsmqgE3KY0Mc5dI6q5hQEePvPya/Z
k8GATv5DabIrPgg5Bali80rupuqyeuy4Xaaz/fpCLnDiIn0fBw6IP/NBJCuZKacedKrPJlb2bgbc
CtCGf+PUN+wJ5LxlnKvvDGhgAWZHRYE+5twFhLb9HoCDJH2pTjqFz9VHrDiqTfkwbX2F6BmAmGxt
ul++kWuRzhmBxXARq3p3kV/625PZaOgy9kdgkZO3bzBpmcojXCUEtM2S5qd9llCJl2oQz2tui8SW
/b26QZz0ptse6sPhXMbDxs8OiAyH/x0/Vhz9xZnYoofR6Ko8WCIOPKqI6QyHZbTdtUR4MBguAGox
yfvQRGKPqeCaxvyP/H21PK236Qr9mlZpc06IJjabQAX13NWrEhtpuOtSdxe0ThALctRy8Vpe6X9N
NCUtRPKZ2SfiDes69ZuPl8/gN5y+qYCk0zIDtO61PalV2BXp9FnjJsryo2Ij3i69wniVixaEKAHF
r+t3zIRE8ynO+KP/c6Y45YZQZh3CU9HKAdpLNs+sg6n9TURPh2/MX9oPYfzMj9co0flN7j8+Dfp/
onix+cCvAr9rXiVYeWMAYXAnUyxcDGo/XzT6mc9/ZHxKxDJa/XR1CO7vfxTy9FE+kNNQj0OtIp43
ed2ZtbFX937bcCGLu/kzhWj1jRM1lYbOqx6mHsoP647/G+4YJ/Tm16J2VymXDyXHHQEVdgBzHxw6
+MfqLEtNLJVBCkDiJdYCSQwjGtdZ/6fnM0iqOjJytHAXXo9PckyVWRUDPxL+y6ZtuIdiN5IIIjMw
dJm8eKkTCpx1y9m0suYJn3gHX8MhU8Uos7fCc2fFdietb1b8UsvX1n6RosrPN5QGTAjI6QRDM1eV
7cwEpUvgvWEVpaA8kNR7UmN5bLbls3vHZN9/hIR6B2KD7fNnqhBmRGXt7ENDj/lPJNksotaazpRZ
6tquFIiTM2AcKmKsVCQhE+bF8i9+s6DT6C6qKpzA6OxGwgw+je/8V1kozaLu657DpnL1R2NPYOpk
NS31W1rf40i/WrUstc4tO2QLqH67Q7CpAldlG9BzoBF1t6DrHNN65EGdKFZNnMWEGeHYbcRdEmrY
BKeDvLZM5mudQW45tXRgsmnzZyI+4EPygvv8lDenkI2mZZAyfrJjnlegSKNxgvvMiBv1ihEdHWkq
91vlpJkFoStLdlhm/R3a0USYlu+dlv3BDOxz1V0fpCz57eXOHlGznlIQxtr2NLP7gPSoIfutKoPP
Q/h3goEuITHZoEnlH9XZYpt92W5NFvPBt7wZIWTIACJQspGDsFTMneHpOKHg3ytBVJRO7z488BlJ
CBgDG4wH4W2v1jGuSDujY5vuZNtFdbl3T+cZsJM3hsxISgQa/8Ev2ZDI1ho2UKfexMNfAi288jUH
Ev3+qLDRMXdIAAAcAMQrg/819wucKf2QV1Gme7/J4zz7RlCgB+bfE2HlDL//OtMtXjl38AXKaWuV
cSvGHDahTZEOLe2Lg0JP2q6Px2aGUKUCxw0euVfahCOyqnvsLObn9etl15iqtwC0HTiNDXjJLQuP
Zijqzr2PGYiOTOaBStAWUY9914cr0uBTmHWkt855ZPYPlKXW5GjH0/d5FnU91HqKrxIhhIwAL9wU
kCAApcnAJO2Wpa2+nsP3hxq2BxgtPwe5urKQskGTD5SVaz1epqI3F5HDFWBPioYZtmt1P/kz/3ER
CBHbKVhhDaJvhP8lt0gEubX+bDvFHu0H8bzoYR5Rm0y4WNZakqaMpObD/n9l4pMrnSHnGnufCBhf
exPV1L+q8mFd7cmzborC2mmbgMf7bcptlC0HrSWYGhQ4Jnhh8nKT419zBnYdFHqqXEbCgp0XGaMy
gNy5C8GaynXhBhqil1afeU+3wrFQTTKkCnaJr/XyPApQOFHhk9HTmfwxUC8xifBfo60xoZfNV0DK
GvGVagAdG2/VG77aVsT6hMIJ4IJQGDtJxJeBg9KRolxyQGIxUh0/IOt+FYoWhbPlwt3MyNUmPspS
SEHkmDAM1wbt4CQz0jlUemzPypAM8OFJELJZAaI7CPW3kv3C0RktdAdWbY89qiYNHG/5x4TE9AlH
VZxMtSjywNjw23WFxBybiVaKiQjwkylE3TZqmLyDu7PwvrpP7HtoY/BiORUGqsbUJS5WkJORbtFF
a84bhc3mfEFG+qMeiR4iE3byoWb+PWGJlPCsyWCS3X+aXHoP//G9Qbsg2TZJ9t62YjBMfl0EgHy5
lReK4k9qWpMD70gKnF2Jcux/wHqddaY8Vczu0EYtM2uVlTx9dkTlvWo4LIHBYxnuBiInm39hEVcu
O43YGPHKczT62CJfhEYixWCKyrSHGtwMAxNiVE+F9/u8HWVd2SxYqvkLkxjCiuUJArLjDGzDWeta
YBSlsuQ9NcrX1wFOZYiJcq/ZobN03pIBD5+ZD1ioAc/ekQXj+YIwzCzLNtTkus5wVRr8zZxP66D5
9u9u/JDn88IvYXX4H0LAhNgCDuwFymSHbliH5UJl/Uo3WjFBshdBo5cRRsIwZSndHWGZUNRL6CnF
reVNo5CD3uorNIZT/47gBLYtNXQC0K7Zez4q1+n/8EiU3Ek6iRr1UyMNYueFFEqJ6ZkZqTTRX0Nl
S99CYjPLF0HkUi7RKmWRnGGp1FfmD+lN6abnI+91aSNGK016P3t7yjpJDntBSU75IMLvIY4EyFU6
s1ZyIJz2moIx0p+S4oLOPc1Dvoi4PicKLZAwjfv4meiLK7g8sBLAXSJMgXfZ2eRTZAq5muhF5SiD
1K4cuBVbBgPfC5jzxrz9A/OMOq8IzwDWM2VQWv2vJKOanR8P0VV9WszE+AaydAinOcG2H6su7eVt
vu/dQBuFyIenrMU/jSnI57ivXnjeTrD9Gp5+khbbvJ00XZkmNt1LO5KA+rrVeK/USPG1paXgxVRf
255NRsB28Hu4IH/EfGT44rgYshfNWWO7ntNhB+HtlRg9hgHw5h4x1YeySy3nQPzsZ9A3zGeJ4ggA
5Dz8b58dNsqPPpt0+DXJclbYUHFsm4EmjGU+UYEQTIFwUdw0DqOZHHdhFhQeBPYPI7/gNcJL3BM8
QS/J2kSqLRy+c07BXr42GjD4pZ0GgR6xSjb1sLEKv96T/O7U41AQyBAj8NpY/uk0vqnUCoZ/EbOf
mI3a5bU1XiZsXh2M2up0hYcXFwSoS9A97LOl4OgcLMr0eSHHxZXCg+FKlIZ1lqZ6dLB+SZfcG+xT
IUHsO5ngL5540aGvk8IX99nIhdB/tukbg8Jjjl50fq8pxUVfUayg3thMEFLeCaGokXBOlNBHDoQ4
73Ie+kktiHHcTdFd4Fs8miWi0sq6QJQqHsZiZnfPevCj1Xo2lbI75xt9e+Jp4l7PfSewEijZrnLP
n1ikXNoGv61H08GXgx8+F+vcQjqi2VaZxc2fUezz0B3Scm94HHrhzX4xODCT5BtGfkG9SeZ0+iDL
sxV00ma+oS7R22Y4AlhMC1Z6S/AiIQd/jw+BOCObW0orPfUjWCV5AZqiM/mMXen2TIBaEj43Gkfx
h2RqttwlGxLqx4ipwnwqql9rDiRROkfQB6SBOvmNRgjuJjdeSiZSSlnN/PmHobU19SV0FDO2y8Va
yfc5jhG0BZtNr6fCiPe1wVvkgoE2YAGmHIq0dZ8X8DwI+l4xE8l+L197DwXCI0HOGe2JKw8wNgLm
s6S4v4B4HLVZnxYwOC3GWYoIan4Fd2ncj094WJBAN0rAB7H/xaVD3n8VZRwbCYDpySXvyaVTKpK1
nB1EsGc+FZ9uyk3AY2Qeqd0uUMqdL1VyfsNDoiHTtSX6gGsGZ5ONyDjjewDoqXpbQRtSzluqyhZa
1eK6Fq5gIAoSUzgvFgK4m2GUwbILkGkaunlhbZIk8BG/2bl6oxMJYLC7iVtt1lYs4gV1j72sO8e1
j4JONxfSBhn69rsY9BSHBD0oZcI2H3WCTpI9HQXLo8D0wjg0Myi8uaOGNxlV21IWXr1MbWXlIw2E
sZ6T7AMb5zmaDRXJ2+OOTky35fFD0Urr+snHfrDi85fD7WMxJqyVGw+5qZNdNV9tpl8AZnzaOx9A
XHnXdQMbzn6wpnzpIggZyTyXe5S1WRuZ56bPiC5DyFeiSrLyXDXS6IFK2ZrDLtMrdQr3gdHy7aCp
Zg5Zv3TbIbXQss5BKy8hX+RwLVPH0FsuWCfFj66nZ4+mQtIj1dRmlV4HwjFjYHcGlo8c9vYdTxoA
XSdymRGzSYA3vovOG2PrptHeFWwM92J0oYoa7VyhnnITepLxAGOD94VDAIlfTdqdGd4cVS6i+JKV
uqu/9ffv4L88Jt0gDiORFA6MRE9WipQTxXWwtAGizXZThePjsu76tfCq6guKBskCk9AZV7oSB7gE
7rQQegTt2rahOj2zpHXQ0WZACR3qP0C2EAIvypopuQj0Alokj2xQyKW74+1L6pWrxvrTNTBe2adR
Cmjwjrp1UBAvhgt3lx9hojV9gE6ce74DlFJ305z9R1I0o33tr2aKNRHnXjOZp0gYSy219tk0NTZN
LoVGfCZL6KG1ofMjo8gad57ECtmuCeOaxOruqx2/zaRRik2AMFpszUQGMPxdYffEYWxVFs4uDU83
JCibqaS7M3oPC+SQkKV+3YQ9tlz86w+DTCJZnkZ+4e1gXdQood4tdrAWT25TvQ6Tkxgbp7ol5knZ
z2VSWH7lpuFnvPqMMfu7Vx7g/xJpRw4v+GcwMCzIAjP4YQdEQB6QCETekNBtUHhDwSqgyyc4kfqH
0BmeYTcmU8dPrGYOFwVzcjRbYweVD992lIUree4oP00Se0UUhU+lmnC1KQAuzDB+loChY09zJcLz
AKHI7KQxLknHBTnCb+RmeLR0hBxtu1Mmz7eBCukWDuX6pmsrEEiekqMJMWFh5F2fIkspzrptwdiU
RPkETWkDDjVjPXypvCl2hqe4SEHVg7IdGn0ZFLA7BzBbG/fVS5IrwP4NgYZWVTj3sHGSZ0Mut3LG
C5M7HaMZWyfxhlXz1G+oW8dSXJFF6RbdUDNv4EIZFD5uhX7+cJCuSqH7GlhoEAIiypqVaXEaHTPL
VuwTq4ktLkmdbIBU55dYGoVHRkSQ90qI5qrKx3Wdf+ddk6pg7fV31C597mV9704ljfIjSj3z3Nff
/CdvmxuzpmY9qLxSiLrDxJHMYTBSwYrMevlqUYtp1tMA/25G5JGWOMVPPHdQLQqF4/o4uTikiGrK
1/uqM2ntWDb6Q2s3sZwKHig0Mz9P4LGilFwIxrWPARAy+hcpcUGmnvSafTmm6n6B6Aq5H6xOrBrA
sC9beUcGS1W7yBggrsJpIetnOuHy+RdioQOtGTaCz2q1FbpXJzfjk0jHQnl0s1Smne7Gf2Bpjeoh
GiXZpFopwnDLWkB4bck/UDpl/SWOogDr2Fml1GVBmEdRe9zXq8f1rzw0w5c6H4KqmisxN6jIjNDL
dVtpSF26VxJ3z8wIJwrw7cmeG+RuMBGUBP9HiWcLttFC/6LuZhyXhOKlP1nK6p2iuCuilXAZeZhe
ISWbHKfGbuT7kaHelZaiSp9GJkcvEmD4vOyfDnDbgN4ziRiw6RQ65n1A2rNKmW7wNlmWWlKCk5Pl
0gpkndeXYBizW/BvKBCzZjlZJ29KMYLi4zQh2wfrcBDx58OhTUV3jvhj4g3mrgoHla6rQ/8ZpYG6
DnQ5rP2/yELfLq7rgOpJg6LNbaWm0gtqxNppfiykUpiOutiBN5bAkoLbmY14XJn0EISkP3+CQHuL
uHHNXAaMVuhFpxw+txQ3q42KGohbOjWiZqPOkr5OtfeVptOqXohQeGDATzb2GsBFz4BuG9C4ZdbY
dSiXAY9+n8RdCyYZ9d6h+wGXGOeqepgbfrA/SArSemSgLliroCwjgNbsFb9r+D8FkvNGks5MYItK
He35gcljLZBkP52s3878a3ELGme2ez4aoz16tkt9u/9H8nucvHUB+PTENKD6ECN0YyWugwIzkv1p
uEjRra5RaSZJMWJz1aSssyCfiAko+ZqALGGX9PwQo6DhPWk+9JG0OzO3t/qclSuiYl1rZe48mX9Z
xb87uoB3SfLcg3tPfNsuwWnnR+Z/MgiG+P+6y9cAwIG4Leqkk9zCZFplDELg18uXpUb04aBRCRXs
Qj5hB1L7DbSreqJZvZ4jzeLVUkK1mMT8yCG6LfBbbUSNrfizvfymDuA7W7BCGKuGjeBMvFwdmdSw
0z5DGXBFHSjXeK9xBOsgUzOSnWPCE7VIRPnX/z5pYKrgMmefhKOmYhYBAjxALSDDYfrn2oWiqOjn
MQz0kYkcatlqf1HNTlp1IHWsJnJ/7uSwudQzwXB4x8EkIX5ek56Lsc7UPxOkyzRb6fxCk+aNeuvW
fbc20S1YuP9v/tZ+axcFznRenisfmtgoK+Mvs2lEbUHqrcSd74DeC+hlKfbO1yMxaHmYA52FTxP3
Rn08nvyGz5O9DOGDShFZQO8tsOuADzIhZZoi43eQd/CgRsX512ar72C4dWX4UK7Bdp7yRSMEAO0O
HneeXiihIvPKkNSpoO87P3iW+uTceEOPUZNSvAsosPR9Wtih//jGPXGaFDZWr1tK9AWWT5DoYq0/
FRQFai6h2Xzeg2nGeUW8FVyD7P44hQyQ0hWn1UMuXQvztcxekmsoiNpGofKx30wmNo4aGl7EcgEr
U2guo0qeDaMd34b2iXNZpbBJRIqboxhJ+brooGftomcvCIcC7HShbvGYAE9L+3GcDc9Wp0lU/qTX
ZT8VWpv4RmlgD5GMqaEBttaaI/qbDf/65m5atPbFNFvbQB7lDWNhkxZ8l7zh2F6C4kCjw1/zgyFi
Ej1IqOo+Ki1g1VFk1btk5TX1sjyH9L1oXP+LmBZ61DFGlePk7j5BKlXYV5NGBBMKpoANY8RFgywP
WPvMhwomk2qJGEULWwoVOXF+zhhlFMN8z2DV+KXXZZOkE6OIjwYTozYV5mzCApRYyfrqaM9SyII6
iSQh4kHDN1ytkKRlQmAfjKfWVFWw3hmsNB+Vk2131onpYFhRlyD8EkdE8xAxGCVxVvNccCSCdq5u
nHpKCGqxfeFBtduXyTawd3VNvi5a3D1xgP/ebC/8ZNVDaW7zK7Y7snqRa+WMN7Jre1mxl2aO9SHu
wazZBYtceBMqw56ofwTsYg+Q5DTCHai/YDBkiX9TUL9dlZ/0AJeG2dqYd/Ap5u70TqfcGRVF20YO
dKkCcl+UXm29JzhPmN42g1n0O3C21DYQLOdiBWoftsgthI0ohA8RomvKDl1wypmVx7gGpILFYUwe
ZCjoJgwHO5rrk83blIbIWsNwCxNrk8wC7M/wn6Ot421IammXx3QWBeNmxgpSz61jI06IxHaa3C+A
/197+I5WWJoHtwnqSB1PsZcTmma9iVI52oRgUVofvG8cm+Cv/hDi7CG1VCebKI0kuBXfylsk7CMX
e+FUwKOwhTfJtfZBi/YCpT3u542Z1Y3iJeQ3xYCjGnlWlxhdbvE+0B5bEhY2dJsyiPJyM7FdC/qf
Li9+YwpBjEfsS3mkldR3sdUG6BLSfk+KOAOb7GQ2UFoooQVSjxJ+MIqfGoEuEtPTNS6l4NWxCqZp
x++z9Zqb1mWHRweLdjkulNDVwGmWmiBlA2ANar8sdoxFda2gGiC/C6tc5ZtAPu3hBn+TiTeaY8cv
n0it/WCGueU//7lNOHa5KNde9VlSFKfc4MP0MCRWkxuBKTAOaNSvX1vp6A3M//76r0G7ZErNOdxD
2Nbbs6nYCzCu6BYBaCxfbhbePEWQXz3+v/o9UQFDJ3UjQVaqPZ/4y2jB5QpNaToC4rHZsqEFOWDb
KESVQomlg2u7OmRAa5T1j88FiYVsRuo34BuHiBi4bXjBWo/Azoq7OymnH4G8OiYwJ41XRq8+kxgY
XI10kCK3vCqf5trhBUem5Qmg+DgSKwxLf10k1O5nH2MFLOSNLVmzEqQcLzdmxoH3sthuJ+JJyUiw
W+8sI7P2besdalopajMhh6vh69cl+9UHra5ksxHgKntruvrrwqPX/NnG233aJRo7klWkmcK0lQeF
bj6M4fY6c1bfE5w3NZRBMK57kWgRqHAieq1fr+whBn7n/jPiOfN8fdz9lpGGjARWPN2fuz91e4Jn
4I3Kx07Ot901qymC6r5j14dB41PufcOWiOBNITqOOD8dkmYjzqoWnch0U8b7WlpJeKP7VEYtHbCp
fK3R7iAkoCUOIXNf8iVRD6J7q4nkoWX18l3XLLulfj5NwlTYxxmW7078vcU8mSQASL9ecttCHkaW
OOnUB/NznP6s6SLaSrmWd48Y4Kn3yIRxfDg/dVom0J7VWz/VSQtv4b6aB3O+bt1XYq47QgUH1mZ1
332gmOvOMs0ihQU7sVhrKPICeoLXPdOMoV2xY3O9X1+iZntBWy0s9pVFsIYd0+dE3goc8Ns61dtw
IKeEm/Ck7krJW9mLdFIqNRWZJvG9WhQw4+1MFAio5ErVXX1AOUZW4KKakNoh+9zvhcUst2+jgY+p
uhXEXxCETzHvCrPaoVj+zHB9mWL26SDh4pFD0olHeP2K6k9vr0HIzRP8JCvxS/jIt9SOF8LwQqqq
gE6axfHFlMN6hmT9yPObavbqWdZA66puG22IfbWJ+Omfz+9+oVaNpSVAZewUSUzpHJc0Brobajb3
wg1ElFYYTppBFVWh1Q7K7PIpZdH+TNH7ZdklSuJiLJ8xFv8FSmwesUPbCy2u32nhjTKkSlNId3Nx
SKOTW1jTamVC3dXFpzBhis6bsNl6dt0jwq2/u5p3w6EtNRdC784D5FChueMpVdo0FKWIHkbxgzR3
KpIatLFTaW+vZ6K7A4wN2GSpBiDkIkhr+hCXNjmz+mGiGQKAbHprn0/Of2Qy+ODL54JT7kIN8qzh
1i68yThR+SCDAtH01VnPjT48Q+X++f7n2rPfYTZNaYo7hiuj5aBVviOw5R9XR4TpQ5BqnSJWmU36
JjGLMnmnl4kwDTCivqbtplc6O9jlzSrlw9Vj9HJuodJFnedG4G4C/Uu712Q2aafAd531n4XKmRs3
PoUK7Le+O4a9SiSD+iTeqP1KwuS3pBEO+TD6fFdzmaHdNOohbhlyopMdrBdaRQTISswcBMLWr74O
nOmduqJeigUhV15TkApyY26OaBvQjh+bRJB9CVwcEL+E+qRUX02fHqSiqrWWsC2mPrr43eRSipww
trHQUXAT00IBy42MHjqxfX8wfHg0LWyH/Q39EXfQMEs1voje39X9JWSxnCTaIW4ZNmV00NY8GAn1
n/pbXYNAvsHOMoeX0myjsamLHjN6gvdSYYyWfxKR/8S7eyYy0swcF2tssBHLTiJh6AkRM+4lj+r5
pU/gcDT0Ye4icfTaEbcS9xwTWOVDCS9BVhXwvX9c56xLoLdKEVngtcWhcSoaP6R4YFuh76rfML2f
BYvz92MeQF8iCHDeyRSnDxQNTTyNzBIjnRONIvt/toZbGhZGuFWahrQ61yTA+O0arve8VS43NYzv
kjP6FhmfHkoj8WoQinhCiY3qyQ0O14RSxFIfJEu/hH30M3nDpClIbVbyGn2Hty3UCKWQ5TgF7obi
rB6VdbyLyK/pAT2Pet3FVEgFaeFzHHbUM44+NhisxNV6pEKgmEJ76x08uXz7Y5eEwhYpMq6lSVdM
I1PgE9VmQi8r2jsbakm0dnrWM7MzPkEW5GpxAueuBuLp4NMdlYhOTvmyE1FJ5zYe/xm0Q04FKLCa
fq6AFLpo75can8DlEpUTGx8HabnPj8Hb1+T/0eXU+p/ZpG9AbqysExB4cuqbyjsUizMzU3816seb
i9gmSH3p7jC21WYj4cp1UiH5m4b8afJQdNxZUX1gwP/t/xmc6VDzvGO/iqDr9VYyOL13TLHBEo3z
v7UDLOx3qQZNV4P5f4v/5YbCrmXua9uC2xKaOKsnpw/N5tmpB7akRAJu038lQ50iq3wFd45fSB12
lBsGOS6hwr+mTFwExYwfC90CE8ySX6dAT06h3YbBwgqyCKyNuWnTb4w20NMZky4XdtR6NOks76sc
js/2OTwQz0bY2yiS3Ugu5dF4Pwq2umYNOjxhpXigipmz53UOo+aOn8oe2KI/Atx7DaWJagIG+soW
/cwoKqQCMLHKxNP+6vN/8R240URqOhHtgb/HT2FlPkWBiEcVN7QFi9gS+QpLdpvRTv63w+PYSLCE
xrmlK4rJmIRYbmMI0i1OwhfCMSZhrhtbmejtGr8fk6Ey3+7/bOr/qpzOZVS6MmgmCYKvde8s4uoA
u63/0a2TJEkwWqO8Pl7iAOU8/kI5V4zAx1qJjx1KaIV+7IfvKZ+JkACYMX0THgShbqulQCKPz87v
7EFe0TczsZXK+qsHvSU8ghnVm9vsvTqvGxNWieGWfqLc0QFhso3GvuMIp2vvdn87TFlbn58aRjv4
KDZ6fFIys1SqKCUOpLp+myvQOs58OTC6mHKD0GzaLsvCJxQBkpxWDtTwFVxX++SUCPw8IwP9Lc7w
m95J4BlshVdAOWN4fpxwZ/jcmomCpyinp+F4XQtzkBK3mg+20S9XsKpWzKHeT+GMXP3CdxRONZHl
Qt7IGrK6MC+jQ+5z2Nrvx5PLKq7qMo7bBSfd6c1Y2nnpnvxPuQhidokOmTGcM9d8izZ7P2ExmPYB
wGBs6BI/fRNN0mc8mUH473jt6/SXttPItontM/M1/VuNZTx5EXvIQE83jpy7dEBUmlhhXAnVvnsU
AEvid1L0f6BikSTEZXubUxgku2fD/2OiGekqhHsR/FzFzIqnpm1Gc4S+rVqVLxiQ/9UKyMydqBTW
mKEEUebhp4K4bk0CwWybAIYiegBLX8yf1D5RwH6OM3siNAbrqPX1apv4sAjOr6+zkugR65cYWTw/
zPOi3LslGwIpr8yShAX4mSwnBT9/Dwyvn6/8sYTtcS88tEz5FjCflobgjhSyP1mk6EgwJ+C4gm5b
gJHO2ia5M+7xht8jGdVzV1xVRTQixxacYRkQ+M3slernVxVWOqw5gtOSkOUQfxHgyln0Oizvq2ae
C2wS13ARcWYlK3tp04xMypevP/K3JBVu7U7U4M6vuUGn0xfxCn6WyZVIEWMjnsx8IbKZWBY4/r0/
xxyNgsyEyaewNQ6hRdjxDccf4YtibTiOy+sQWvsfGW7O+zH5OLI+jXm8dtKkyElBTXRL2RY4a5LY
SOZZepj8DaIP3iMI3+8zM/qzYN/MU7BwneVHjUzmeG0/FpgARPR0TDRsyVvXOeUtWhaVpKGvyzUU
vd08d1lp6P8qmAJfdXblTDouWX8mOU9KttHh7Ji8qkCUSC2YL4U0c1JqVqGfh/nJ0wkGheNPhXjc
iyDWKgzDm+9nFbyxFH49LIoV2frJ3UcrEd0w9ZNcFrA05ZXTVgj3jZ/5qxImkqVjvhDT15DGhRVM
r8IfK13DXnz5Cssman0Pjwfio+zYEGLvnAtnfjF/pEZ/8mZJp4GumQSDl0iIYkm1qWpxODEJAkyM
rsSqhlf8uIEvFJlOtNd7vjSp/SMQY1Io7Gr0dswafasvvIJJRkBua6/xWVWOp2uLjirv1oNYiO57
t9oXhSAIM0EYfDRmxNhjChZ/3VroTT1TFeVvWLm4xszlMNYDodyn6KNALyALBfEjRlAcJOccdltO
TIvRYJcGm6z0lOMBWtuCjVVJHuBixsmaHjI/AICGnRApoUUuw6oiL5MApjrusQIIKRCsBgRQ6mYD
OU/KnJJDGVvd/mxmK8zRuGx6qY3UHxMhOrJ1uLk3kFSU7q0UtTjdvYIq4+HDVMX3gzOSPbErJSBo
nwb2zm5TR6ecUVsWsQZUEK/g9aZR4OPY9tYQyQlaeFI5ihtr2pNaWE64YypnaA9l0xR2LV2jKLAu
5iz9267FRWM6simGO9EZW+QHsb2ntg1NTQh8M5aHwjRCMDW8J1zhYR69FERanoZtDlskG3Vp+R+L
6I40REkCUDdIsjQIcx6tEO7uvbH7C5TteEKmaJ4TYlFavG8Xjuf9M8N1zllSZu/ncy88SOQYbgXk
R1cS3qFzWtsdmBe0lnTjEWbWjPcq5CM6pkFvbp8HpqAx7oO+gjcD1jwpZR6szfZB8BUBRsuhUp0Q
5oQjHiT8nlQKG/I+t4ExYkJg6EjOPxgh30ffmDgEhSHNmGa3h5MR3D0JyD4k1zT+ZcMyyq48U0lc
8ZGenGsGd3CLU3ecaKitgX1A+PnbfWap5UHH47hBm/vY+dbP+yq+IMT22WVkwvSYZqommdfKkfVJ
X9oD2jm/E0K95renxmQMCS1YYA07L8x+ZlD+gh7KOogrR1/o0v1VeeXb8GDBIPro7Fi4AgF8cerm
l+d37a7NfgkcHbFVTBUD1vF5RT5BEhYHW1PnKRwCYd0S3J5N+SJclkoFYEPl0Wqlr93m0rji/GJv
3gReVyvdzaVxxw0PnSOGWBPS2HGWm7+ug++mMud0DUN7jW6TCIkHGoMaMlP4JqrEhwyFlYjUNPij
NDh4R5PZA0wHTMhlleVkyi3VAPLBWeZWhOHlStnqzY/33Z/xHxUnDs12Mqz1lo8vlZgTt1LBMxt5
qdT77NDAh13JnzX0uhDIi2jtYvqjza9gS66VEai2+L5wVl9lMxKd48VuG1YrezLwbVkFV8px1ycs
qzeSYkoPeboW7ioP9iZq8QQw9E4R/oV7PH+Rgdh9O60bU6saoydd0EwESni41MH1TfQ6C4IxgIJr
Ba1O44oldbo9iDpS79KZ8YQU14qzWnEONdCCloAinP1addkj5p/jImRTf56VvyzlfTYud5/8Fheo
qUNDzXZktAhpz1K6VhHenRs/zgui8Q0WZYGOQFgb4BGXazmZebFTHBI1e7gFEKlw0/atJqUPRauO
NKI0a21yOvbvJ8wDvsFBZUstdBry+pKC6/tgotzAtkk3F6Pmpvc579zHXEYV6g5t8/WqF7PN/fBx
EoiTXFU4jNPoXSaUSxqmuLNvXw78Mli7uVRLJh1KxiuWXfw2+JKnVtYZpejMbaoIWflELTiWP+w1
APK1UQN3bQ6FvJG5Q/XYEIEYZ/n7X/ihwYCGq+v3PZiZoNdJq5yA0Xe6ynkI85vfblNT4dQ/PAx+
68TPyYOYwv9lAqWT5dAdl0D7Ig8A1SoqQMM5hr668uZwFD6j22zBJuUW2FofEntWwaBZ8auIt1IQ
YNpkRfocoMrkeHD5k/8Nh7ixwDI4v8JHhKI1F1ByJYlmMOgtmMH+HdAfgm3TIYHWjt9Ize4TgKDp
735HQbRS7zdYfBKrGeaSXVr+UIb7lvYz9CW+6/sqOB6JmmW7bWx/URaikfH35sxRRlBjmfN9/qLO
G4kg6pCB/v8jjXgp9QioxBm6aif8mIskfgDklUiUFmx7wZg/fiTdS2Ixy9wBnnjgDZTuLgrVBiTP
+4oT38OWzVj0/9WqCZVbJ4eJKkp9l9zil5X/pv5TVh0NH+aImJkKLAVKPb4S0X1eeoGieAigDbFC
FhZurnnwuUROvmpMAbp4uvu4MnW5EEndtO92J7VBu6yACgIZnL2bjMLyKYdQ1nGGeN91XJl7AeuH
a5ZSn5XeI3X6dy8UTMW50bGpXL51SgpbS0H0sBkd3Y2XIjlgTTngklQSu+ueqs4lC5RsQvrZQSs5
Ydv4XSIbP6uTlbuY1NwGZd/RXY+ySsBpR47uK3AEWWdiLPshAiADEyi42R99z/YlpFmLO6p17gQi
FREOIkuPbddkQpu8KF18mCCoGmONemCRJlklC6AXDBh8E6D0Zzt98BBhaiIRkahhmu8EzEx1E1Ma
apZEIbY6u2xjPklFhXM+LZvbk5e+lLLeAgdMx4iMl6lVspBl7VifdAKV1Cxug6ZdQLvTBHMqwh14
RccstKWiR4RVgC7CjXjCZ/vdxcqG7FGGcskCJszHjKDNpyKqD0F4UTDohf681QkCtTxBDY7QPKef
wHvw8KyJqibk2yGNsJM1zzScCTVnbegB99m/hMVs4ygA044iuPW7zSeV7oDd/6qMsB2ZDN1wv2jx
s39ECEQ00Id2MHMJF3p2D40iqdPxz7bRg3mzIfeU8dP530DnsnuvKrKt9j6TL18C3uETj1m9hf8a
wuBZJigsJsgQ4/xS3CH/nmx+CtCWJLVvBTUZ7c86M6ZE4qAFL30rz07c7DPuDSJM0C/t5HtA7Bdc
5zFWHiQxLkfaGKmsR6nOqPv7ObsfgJ+iDfbr4zFR/fQ8VG1l8NY9NKFrsT3e6nviDHwSE0juy/ht
c2dVubgwLHpkdEZ5V0PJC7vWNwVSfUys0VrhF7CKHVIN6BcMbJFcIfo9A8VCFbgWMB2plPNv5zcR
iBT9RSBDLuCiDD+rSSddZrIWsEo/AzIZDcD5PmTKxHlb7+ag3h0LH1hZhZimOoTRk6fV/jpOU1Pn
hYiBicamVs6UocJfxcZb5IjDhXGTOlltWnxGjWtZwbSma4Dd6E5H3p1cjjZprNvmQQO3SMobj8Jt
yATjSjfrboq3PQGzsSsw7icovxJjWhe1XAJCccJ8egafrma2GMWKM9vgHv+W46ersWOPsZYVdlfo
fBn1X7RFbSvzYCZlHi9XmJQWI0+U8q/YeLumeAeRXgNdDXhIeUuh86xgrgr82q1yGFlTNU+6ukFy
LwkGsixf2Nu5GzKroZBOwLoJ9mg8BOt0vWMmqZQvBBISem9Sm8mbwcrwYt9szwQi3SfOsaEpLUUx
fVUklXeEd7kFg8DlcC6EVCvvvjiplpmfTc6qAsjNjUS79Knxitf6LnF5M6IYoBWHX8dJAm9SwhVe
aQsQgk44Gy/CsiTuC7l7WNR/sDanliXnBT5XL87SpiqQHBZ/P5wPO1fTb8IZ3ZrRACKDAaLjPiEw
RxHYaab6P5PK45PaKp8g6XlLODGUaBBVKg1A0C3maoFNknmDwKAD3H75LqaByQo1UzXRGiOmFN5m
C2BT+wWMsnMhYrWJxrebr5vDqcD14NhEeiVtOU2X7lL6TEk/RoemGKOJgNqbrTLqCNV86R4OEWVn
TXsiQT+oogzBJ+GptyN7bDiMqIebmzrSSl3j16/jfE5hHYVQaYSjzCTUFM5wFoDDRU639PpZe8P5
k6MX+XuTHVTTzDq6UTxENk3B6cz71ETEMTEv37XmWpEFxV411FBD9G5r4Z0hOz+RjnOQD4QJLh2G
8qNEWazDnuAmYLNvlDgELPffVydA1xqa8PJvaeswNekRdjRSH7/ohHrpveJGtgjUeLg0qHhR3ROG
JSf4U3dVeyAjXXvJt7IelKhirvVKy2Nf+ET8+gQKlqKzXvVDN4Tncm0JZml/AsNikOnMZK/w8xBD
s3J0ddqihwUYA0++IdXIqbXdRLd65YglaJv+USgOa8BXmFvNIvfsEhzcHveP6mQdrI7Lt0u+67fe
uJ81Oy1IKVpEtigdLDR8NKKhj6VONSrYgymLGS/Ir3k9QZWxXbXpTKLbHfTOHWS4dbzp2Us/QqXW
4krkuxwwI+zG0kugWprZLA8NrHw0EjLvcPiBptZsEr3hynHG2MQIVxWMLAsgz5A30pKRuU9TCZYN
MKyi8q/l59Vs852jiVYCGkJrDkvxgzmYKMujuujVcgj6EypC9UMs7W7jKEw5MU8BrEWzoULAclbx
oiX9vWaeuplcDIqTj+YNdFMdGWOKfvyv5Z9r0Bk9YH9OYAsd7pUEIgxqZ2qUZPPbnEIZUZZX8ykK
2JctbWN2l07NHLAsbDHyhpUlE8IIpEuCkKake4LUlLFEdXZdKUPANdvGGM86j0WQRuYN+95QdphD
hoQ4Xt6GbOfxKHocOBnfLPuLbveqfyaE8bq05NjZ5D97J6fE3tfBGxBH1JChJfu/I7np8/uGBjyX
pULg49r3LakArkTsi2tOIPspltvSITcFWWUQKEpcEU1JV1C4K4Fahy3dogyKdknqDlQBk7GgMbJa
cIkD62NB0UXHeq72239CxSOYedRNAexK51/AgRr/IocsLG2y+45uDKsNB6jxu22U2Jxb0+YtWUmt
On9hTxkoafB3z6X7SAtLZTx4oibw5dig/F+p5Z6c2KPNJVx+72QTmwJYjp4lsCU9Jqr7ZXYIDrOB
zRqkBBL+K9R94z2WbhODgmFwwqqVQB6ewx+12JlC4fyovE9tW5n7CDnUgw46G9uMrAr8GEPQ2usi
MTGXhWN1WnaTutpi7i9Waijn4DdNAqW1SWVGokd9jRlQX6PqQVNP5Eal/akbCySokikMj+zvz+l8
ZlxpSOagMGSjzCwIaa7OLJNEsmyGNgZVlu2yIYc4xN1Cs922RpPx2KFH8oliIXVNTXqheVzmO9g1
NLACThubfCD/OP+elSLT6crfb+mhxSIkW0DXksNVUgqGwQspr1a72VVsFFz/gQt3yR0lvrLloogG
0eL6YH6l3RMC50UpuHsZrQWKL8e0+c3RwWKvG9JOAFxXGXSB3y+lfPqSBMJIycjDVR5okDRCGLW+
yD5j47t8sv3CnO9PO2q3jq+qD8HnSxlC1ufMlVZr43d947+LSGWssQIpHQ/G3lamBQjqLwNuflo7
SY6rj+1WY4PMdI+YTs+pYXKCJWwDBHSQ3Od8fTa3XJijtLyX09f3/oLUl5SobiG58ohi7CeNfvsr
eUsWezYyTELLccAukgyyaeKmgOTbKBab8UNnwL/U4UR+VX4jFUrxwZu8Vp3G3uQb7K7gwMsPrlQn
9jUCa2+SiZKY0nSL40ZhM8dDyTW2fEJkbO5PmXaIqeOlq8a/AEgbgiXStyVjvZzp8r8UmFxm3nfh
cnf52ZVsQeoAeFxswAxpHZz1gGf7ukHeb6R1o6lEHq4Nrh3X80R6nIG87iwve/JPNgPxM7KtMtN+
stDVPvx+Z025Q8dDDMKhcU+uW0sZpCZ3i5Vl22j/x5Z/E1Mr+zyN0LayG/9s/C55dPBV4bWByXLQ
rQnO4uB2Rigzr4ZFsSEb6mVvXV7CkBirVDMRY89Gzy0vkgnc/a3NafGpf48/boeXZaF4APplt7jm
8nLsdNHl1zF3gscXhh7zT1WvtwSV4GOeiUkB+xXoWIJjJnUSGxaZNIVU28+TG7jB5044c9rOIM+J
oLqor2NTmYPLJhL7wQd4xNwC9n1TxYljlGmex2bKIOz/Q4aARDD/sZK05+bTJa8WuoT4z/2IbOFE
e6bw37nqPWAJfs/yYbHmbHNE8QXwuz4wFqZpsGtxWL6dNoFEjyCwYLEPcSoQNKNW1wryycfPQYQr
TDhKcWKI1zbT1C9div2OwxhT8imQXfZHZ3aeycresa3raLQfZWkM8HdIU21LQ8cv3MxpU5EF+nqn
Yf2QAgLl8XM0vkM9bTCfthA98oeVppijUEalVF7XRFGNnNGO/liCVjY6pHUJMi3cWZmRW0L+yZKH
wG3gNmfGlme8CdyfArra4cjIDLWt0VOMOvl8QvY+7f+UBIAw+8O1nsudFPiQLhYfiBT+IskTCtBE
dBDpY0nj9HQIhZNRQ96jqMcQGbeN1tezvdGUd/evmcwNPju3tQSfO/qza4MKFqcxbS4sFHiK22WC
PNyNUvuFXjDx8GB3pOSxQjHsTC0MHUseKqxh9kd/Pz4ogiesNyZk4aV5+RxJD4Ej95J+yiOyygFW
YzfNj8VXSi7XSmVL7mw9afIflxLfCaokKafjJvb770kVT8y6fzluPrjMpxJFarnr8+0AA9rSRVB4
7DiQsXt/7Tp0+IxKHJKoQH+s1aHXmsT3p3UroKBIJELiUUFALjwBFPDg/uK+kWfYH92Bt/ok7qgC
6N0GstiMpfyY0Oqu1+0DEdm64p/IRhOR1EBIl+NuknK8mJddf7l8lRtSKC0eanx2bS207LuGhrok
1WXaGZudU8HcgQmq/gxZ4QjGsgj33gBh11sMi6MLzDdeR6aERZv7g2cabl0iP7llHEBrODz8L/FX
0HUuJuPvkV5l2md+lJ1Hzz9bn+4N/tR2RoPtfqotW1Bh5+bsAGrf1BgiwIt2tYxZINn33N0N+jbf
TaQWenwDhB9ZSyQ2qAPMl+LIpU0Q8whttpg5bXi7m1oN3vzTH6HXZXrqMZEbc0ryu5b0XoX7+N8C
lTj6mEtK4ZYCkgE/qfM8D2GNWGQKAsNzLOaJ49TrHTFqTArEuF0wIseoa+Tz3gNwMqo9h/5D+/gU
Pgh+JNdzgIAh5Y4JfHhUav5EOv4DatqycTsSTT0d84sFWmU/zi6aMJAes87l0VWfRftmF8kNgt7i
wgOhF1fmdSO8xxF81+0CW3tJgoPj+aBpVvfRygJ+k66Y3XECKUTdflrIwR68pSY0D8OE0L4AAxzu
8pQw39u2CLfm3sVs0NTht89bXdMJnTs/VS2QC6YumRxb5UxiNKrTAlLhtHhz05tVRWVBwCZZyvKJ
FAOK66+G3TiyBXLCTOaUkjtPC8FP6C1xwzkqYVNaICIhJJWSfe3ovXkGKNvPOpo36hNnNR3o9sAO
oVIgbzVCGe/vvU0YbQy/ytkl+5OBW8PhOqKGCjMBlGxi4zQ8Yxuz4/ZhttggewWofK7qT+YHvFcJ
G7ZEKxo+xgdZm1u6vTpWn/Q1PmNSGWxGZUFdQhe+CxUBLqdKn0sdNzPHpx5jjQIIjbm5QHbvtCsy
1nYRfWD6qapWuMoJt1Ptf0IAWf0rt0qOt4ren7MMo3tSd8dRwkmfTXfOO+q8y8vXjqYnhRu0nSm6
pgBWrbC6mdyTNuO7fWp2YftrrZSuk2VaW6V8gnYpoUjs1XDe0Y26KvVrTFQpVeAG+WmzBzLINb05
HzBdzcXGBMfUcndZTgOck+042sZPankcj4SpXrIq9tILHhl9ymT53vIh7eM51U9swHzMLp3AsDXr
KxJM7RdW3v5vntH6XO/kkO220mB7jSQjYsyNji9+MJUxMZmw5U6E6Xpc7XkDm6S6C7qx4Zrhxew9
qqeezHArDDeMMAzFwTBUQtmhZ+6Wrm3Ipk8HPHggP/jwk/2hK91BraNTDemXLj5xV/NVAdqJ/Dbu
uXSx2yi8EApoNxA9SKlG/3eaLi/l1mlj2z3pKz9YZOCCzQ2Ji/f6yJ3v3RnEmnG8sMKZ3Azvtqvg
VOcNfsFk4qpCbPrBeR/lu+DwOsKKWgaZ9xRgE6z9iyyLs/r0LYe/ZCiPsvRXKkDZBLqLASbid/04
oj4j1zofMuWqURyP3LsPMQeASEK9ZccMPNx/t/+X7edp+LSKsIp6OqU8pWrmvb0o/I1SvsdCKBWz
jJOyXMilg6aUejfSHAotEwts/vRH68zZuZehacivGcGVTU0krdniJyyhsF3BcVtrgxnmmJrjLIZS
J+Acabis2UicdyzVjlQYiiOZvozK+qWUR2ybbkbwItggUME6s1yFyHUWjQ48IzcQJXpUBXihFUnX
kiUS7uuLL/add4fp8BVhzSisJlOxhHqCvhcHMGTk2Nq1lzlaumyrZWOgmIaJekfKGvDL4M3DVaro
yNMt1x5jGfYOfDKv+wWm1R1wmWuxMaFcfOHZvabO/Iam2G+7nwcsgwwHsvd3ehK9//BfgL+Ryob0
74Q7k0wSVjJoEe20V0uc0YGZ4QYxwLCWHJM+uObWrA0YUDzvexfYJOchLTFr8N95icysEhDNeL5Q
tXJu2bWyLMgaY/VyKQUNBzQO/hnwC8IB+lhxBIDGRIRQCCY2YqWwFlqkApcYbLR+1/jRViTBdB/C
SprfKjRHdGCDBKnPBMM7TNQOY69IxC/YPfUJHnlWMTUo0zIBG0bBo01P64FePj59cAdmk7vTK8uE
rn0v64uU6tOa+SGSjRzsZ1oxnWMkzOMcNMZYOoQrCZsN+nGWRUkmTnVb0f1ke1M7WZXptqK2RoZF
3s073g8dKkV3eNytU2Bs3Q8SdEc3pU6qZ6DLGWKyOQvqzHA+LG6Yfy+CErjPqbig2CcBO3LZ8F1H
UVmJtklwN+8APUFVl30slTV6jNJZkwE1Vx6RqWL01lN42rm3FVU+sIjnAMZ6yjt74f6C5qXQG6Xy
g3k/LOGYzqcw3vwwztB+SY7TiXEpPcd8gRPPDFkIH46iiu7xemQ5tVQTyEY6707RpGKPi+n4c+js
+z/1aEe4/I/VGdTvB8+2+AD/7hsUBN9CiYW8qGxuGakp5Ho0onrhHghzgnjEePV2egTrwMCOKajG
qddcvb7fcXHfgRvEVCvuLpug5R/PebXkTIwBSmrh1Tl0MZnSo13SjwEVOkRwSWfejHsvLWFt5C8Z
FLFT983s46eLAnHZl4SY+w+J5/zXoLS3QBb1ezo/B45IzdePI6wQ2H1gi2VcAQjwlGk2mQ30qs1F
ZIzWP15LgYnknW932eYtdOnIVG6k0UtsEATpTo6anxU3Zp5H1zNH4zqZTE/nYR2DrnvULXoSRPck
MHwabr8Lk4NmuIgAbt5Siz0GJuHDs/emKfpE8POmIuB1pwaMfHknqyoZ0FLucuRrsBCLT63htCgJ
n93ePW3zkW5dHwn07qQ9a5LEAMrI9Fz5dSC1X1p+hEEVBSUgZ12QWaDPbzMK47RBo8skRFTVrZ6c
9GHvhGS2m8LdWcAorO3p7J8+pM1l0tYOk3yORS/U0IYbwEgmrhD8vkesuuoBR4L1HCKdhJauDSE0
onGrB+qDHxVVfenSVQeIGXt8kW/9OmGqjBv/22x8KRV+PPARoRelyW7IdKd8/BO46bNgL9G2a8DN
JxvEta17H9n/hRgoa1bik57KZTdZI0rUNlOcmfqz6rW1h08Ze50HperFL9pt4tTYRtg9MN2p7zVv
ZxnCAmbZrEc7ofqCY7EJdlwANfb6uRj7R1EYbCFRrj2sSQB6DskgMhdDvA0XabS6Vy6+vjhVCI2D
04uHCDm0Q2N1Cd2uXg/XpEek7z5561PBZ13R1xuK56dk++hTWhhCkhknZ6uCL/iCFMnE0eQhGrI7
h/ot1JNpdOG+UtY9cSng6rsj6dx5qZxphN1xuQC9wfCxotbtGSRntzazb8yQvp/B0tFOYKsNJfPp
xiaxdVcBqAN9xMviwjnNgzgYQ1mvNaq4pFnVxdIr8mTPYrL70bnfITWGpTQWOPFwlB2HSd60IMLa
pKNCprU6GUkFELEicGU3gPRJ3liX0OazES/ZsI78HgN6XUqi6vNp+Wvwp21e4P0DoVPup1UB2xwh
p8ysUxJOsFvHTco897XNln8sa6aiT+n7DDCMW6WIHAtAYYD8Fi1oVSEBXvvJgxxnrywZTIHyp1dK
Jhj02so0D8ns+mvDB3AWmfe/R78DFkaPyjSs0Mi+cTNx8wlKdpQ1Xd+OQLY3LZKHJ1jcCd+lQA1L
9f78GI2HFI12tmwLsGWYEnqiPv5EGtcJIhE7B4C05JIVTnfCau0kNlukhAzT/hDRx0KZPRBC4DDa
VaejIz61unKPnd2bYKQfwNH/rdaUt+qcqQxphMrP4ocL/O8eze3/j+ApfwlhRTwd5ULYk4wkWcmC
lY8DNvnmPAPxzV+VnooQkaiuwZi0zMEJSrjm8gOt+wmJwurrr6Rbd3bFfvY5BdQoI7t/It0WGrh6
o51a8WbfOm61fBoKwPDmyHlnF3Ou7TCv7X8kliY6XKrFgzjsUaw1/FDBpHnXR7EpSz+6PMCiaTbg
Z56/zFPZiLSpH6+q5qPvNYAZjmy0CV8xxUy2nSYoeBR+idycHWcC23jPeI3WBrngn7eVeevNqBCc
bahnsxztBPTDB02pFUn3V8QNUW5GD7vxtOZOKTR7JkmGqndRACReqH9m2rNzYP+3OQJg7ChPfyZs
ez4TmG6uqP0hjeLH/NVyDPdHXioi6TYpEGKLQD/2mufclkFeRZhXXBjga7+C2O7A9lGzMocCrCN/
+t2h8deyzEVhoChDmjE3JlUGdUZig6saa9N4PzXAVZ9D7MeYKZ8IsiHc9w2UVJpTIf6m3Blgjnzk
VuEGw9acxazcvm932j2fOlcVc0wiynLCGkJVv7TahbYD9mbhCOKUDAgjXHSQ8QxrkjYYe+pNw3AU
HWh/ejhU9cHU7BdFBRIdrKpyDJgfpkIAD6b7EtnAtmCCdaDgAORQWolei4qQsRws4IprtmAtfJSe
16qQL/wpQaEau08Fiev+jPvp/XGW8o9h535PxgcClcLcL9r0Psol5IjsWuEjqbiY6FMBpA+V/NBA
tAbjLsGNKRAh12YZnm5fViAVGJwUqi9v4tHnjSYJXKzri/4TIwIzX68uwMM0sN/I+OFnoLxZWUPy
ZwlFCbrvN2J9/YxNBVr3flAwZ9clrR4bGslHxyxQ+PBGd/5gj5xdxAeI3YL18mcMErjxAwx119aO
5MpJ7oLksuOovXqSmgompnq6O5fRrHBNXTZAClmbUtSTGfzUbHuOXzT9QacoFmZBa7rqcpEOVzV0
sWo5HqO7/ZoBs6HbbXqOs5yVfywngi2Lj1Unk/+bmICY69uQAuB1wCEp9k4bjUWXCp7h2Usva0gD
IdR1C+FDiHC8VOuGxMlTj5pA/6sxxATzQu+SKXO1G2xP1W83K/MA31ZPoSI1X/eJtPUhtcoJRvyF
BoxHzaYjePRJV8zx42XEBCTMaBVrpNKIUs82oIhIGsHOYHETwVcH7/mmqagIM4XwXubzq1rA/Tlr
CDUIRY+OYjayb/mnct3PSvHquI16WNdYfcypGkO1PhKtgH4h/RNYkl2l4i0rDbHa1hbLu+oMg8Pg
+n9je49VzZOuZutrCIla3xOtJtYQ2jYVwF2swf7zp4L3vJd2qcbrDeVirdd0SCdh+NNXB+25UMyI
z0qYIYH0br/6uQ/JTLeA/eIPHCtpwzeOLxtfNy/sZ8DxQJxzJr1vfxtRkBvQUV7tXP0qBGjZpLO/
1cluaWjQRPYRG4Zii/ZpJwCQyOJvGBnyUK2kXexvyOqDAmRmQc+D9IXSqDUYXki2iNEJ2e33kHDI
YMFzeY7L//eUR01CDlWCjVBkSNab1l+Mw6RmavowGU2q/NeQIoaYJLt/0bGE1SA83AgzvrxZDGQA
xFoGSC81CH5cvKihQScXplvbNGYBrajyM56CR5Dpv5NicBy4wait8Ewo9fH/0IiL2iGNKRly/9hb
5hnQZA4f1tShFYFQDFqKrXf29JPSL1RBODrsniYpNdU+Ovh/3A5U+9e+5mCBLGKNQH203oky6EMO
wDMTb/kFN5+HG675FmtNkWHu2Wr3WHcHr8VD+sKQFMWrKtVKE6vYhX/HnaH91X8fHYDB5vV2xoky
Rty+lOaBp4FH9qICMLpy1VGr28FrnJdC36P/DBgx8lgeVs9G0tmXQdJvr2YL3s89b2drRpfmubJx
uR+Iz/371Nggn37+c6sctPtHvbmzXPurX7ebvXr6igOSEystmomw5cdbcoaOFIQ4P7Sp/raM6NrY
XR/6dUNyXh3/CCq1L88bgA/1Kyq7bPpjA70AsYLiv8wKF0lXgIdBLlmrjVdKXq5AAQiPQQXmJnGj
pbOIMmLWsYODz7hISD2TCnLbiUE23/NUIvPviNzDyTkF8+3iunxUFYo1XvNql+G3vzB7iN/tE8HH
qg95WjALuJEODniP4Ei/ol3JDXL+7ztfhdMbOS6el/n8WdTTHVC9D/WlgPj09uIxE1FYlnTr3Cx9
+PbiXZXpxt2dRFQ7ds/HydBzefIqTqqtGK49Kf8NIf6pa74gUurLNMGg+Cd9d9kVkFZOzlivKXGD
pLq9602MHTduh6qxsbJy9puH2b1wppseZ03+SbygjhcA3uwZ7LGIKXOz25fM8wW9i8uJdazrcPlv
K8wt2hsQHsrVFnIA4E/JNcWyl3QsC3SjFQeOi/PQgH2Yj1ddyUJvFcQctpcK2WlIQGbwsfElk/u3
QtRh1KJEMoC9aduxej9jxMKOGW8oflKF4ItbrAXR/E+DZhS8NQi6BORdCmIj3hNlld1W2oF4I7h6
l00vzLCAtURddQivB3irYB6Trfu65xP4NG3ON0ZHZLIfSsV6myOrh735xN7RmVVW7ZzQwJ47DR0V
c7OFrTefXggf+YB58cfXC1+T7qKlHC7A5gPPCS5MF+nqKxYpeSQcOLDrTF3gOSLtyhuPJDuT8DGQ
iqEtwqOwCk1vbA7WQVXriE8Rfj5d+tCIIPGI2j9+fapd+zQ6wg3k8iLkJ9of6hRugN/LmP6clLfy
fwnOEEnynw309Nf1zY3eVkBpG2YizJIUdFE8r9KWorKVDgAWqGgC0V6/WLnUoP4aSP9VqZb5FBdH
iRawZTTTXa+pWKk1FCbs0Lix+oqIIlpDe1hcA9cK1yNgT2ikPK0PaUlSFuiR56xu7xJ7hRO1/jxJ
FecsD85dnEIls/5mtFmYXbsTHjIGKw8PRQJXOUcivfdLv4UYhbp3QYHyHhtLovjz2nOQthV5p+tK
7FXmEOtWeOa1fa2JUEfo6NPUAkNRs2RsyJvjvSvGY4ET8JC8xGYGkerW/baEe/R6RTwP9tOd4mNk
mpSwIcbPHEPiLcwivJYXTypXlu7B+AxZwAXLY6jcNv1pbInoYpyKfn8EiARhHp5dki05N3DRPxEN
q0kOlevquv/aPNe0gAxXmKDELT4xTPXo8Ob1lFaEBofFNxyCzVMP9Ukbed46VaYramM8NoaIvOOU
oyv9xbY/TAHJYARaTlCbzCbCOr4C+T8teLg6XM8fJk8lRwE5n/Db0aNaVpzXsFrZH1PWhBPCWvwh
bwWYnWI0w8ugPjWsfglmsIc3iVaXdh9BEoREtcLIT3u7rfUOV0XH9oY1DCAxsIjue/3ADLmE90DM
dwne7IOzuMbWwJA3PSOLLiKW7GvI5kMwCYzN6rz6A2qwOB+ZOU7mNfGgBvrHqKkqJoHGf6PY5+3t
l006m93CBEE6jknsv6IInGvnlsVpYrb3ar5l0S8kgwNf0d7B3qozE3Gqh259MMPoCV7fcGq2pQQE
a5ce6eDl1BXKPBV7BhQL4ZgJOkdi689LePA6wxPlUN8lR9neOT611RbGJKn0b7Hx8rw5OMROw2v3
qL4gCzbb16Sal7ZJNUHY/9wLuLwnIl4bHrwgcIhET+myrXppeOIC2uDTz7PHRqStv5xDbHbJd+H0
KveSuDMcbDvK4ONdkicf3XFCvUwWobelK2R6a+vI+KYiFJmtaJ9+O5hspMMby3Vu9quUJnnHivPI
ap+5sBVDnz0bFpwmDBgqRuquEeGJwSpNPpvoAcV/Ct/sicErchB5T8tlG5HH89CxeVBlazEeFKig
4Rg3UZKsjqJFPTu7ix3+Oor7iLDsK5yY4eNBbpeX37AkeAokFqrUCAUR1SlICDar1m7Nl0j4jrUe
69kVW9MLAtUKDmSyduK4dxhPIAOA+wbPWp2vYRhibhg++kcna/sfUFzMgVDekqqqPyCuUwGgx28z
Oyw32tpxgFifyVHOffeOi0odjDy4N3jm0bldXW5woLy9J8T0FXvTe4aitdtvU17ap4rh19wA9GIw
NaY1XhyGQgjn+OBqtbjE7IxsBnw6awA/ij44yIp4lnnQFOxTBoBEQljZN9MKvNAMdVmpdgNoBQe3
w8Ku53kP4R/uev+QOnh7jnbq2y9vS3xfAdEVs/HnQAg6/eWeqxObj3DjLVSoejJYwbeQD51uRznb
AqHPb8qDRSReWW95sFESUmzatODgJbJdcjSMoKzIP3W0do52Ycl7keiYy4aRghi9PK9rhFWI5wh7
UNeoMnIT4/Kzk4hYZHNoyiwSu0bzvUl26f95wFTEa5zIjYUGXQ6BGAvBkt4crE90R1xrJMNCPIpj
3BdIEaSqHAlcbnWW+exsb7LCjqKDpG7+JiYEmTdpFvVgiBmGfWj0gwA4xqne8vP/Ll9rHY+LCfbB
l6+tDpz5tI1Aw+0vhNW1BYqmmpEA+YMnX86BJS7mUAG8ESOTH4K6S5xFf8KxHjTyCtYLogVOnSPJ
HS1xntFjdg/FPzUuBlQIn0fIyQadlwKwjMTOvMq1l6bRZ9/ugeEOLC/46Ksr0IM3NzZ5UXC8con2
flb+XT7csgM5ZlAr4sAJ1M8oJz91tcFaqu+M46qOcOroR/Rri7p9EFBvG/Gq7BL2ZJAa9JtyiXfV
9mWpS6puwgyKzma2MWareFf/NTJamtv2lgpKxBOx24bufk+hi0qOq3H+4yO9jchhdjFaI+n1Tnbb
UctWxJtWA9KuTLWR8vUlICi1hIl4h45COIJS58xulKQS0D960O4Uy/LMPysNhQd8CnQgjc9iJlCg
XW0UjX/NltRQxtOkmHMN4+FFu+vDLuJwJHDTOFkqw6gkLZcESdroUMgBG749zMdQPTIac2DaxBPC
lJ3Mw8Jqp9DHF7Zm7lm0XY8zhJD2NJk/XpyOR7tgJrtxBr66IkiuMuVRrJAPDk1ClTaQtXzFGneL
bZtr/ZDJ2XstvzbkMCW/2uqExCFrxnydn8JriLZgmIk8e6cpiZtslq3AWU7ciBFe0BUTVH0+aQR+
KxahL7Hlu8OuYas9TdK4+82g/tG/rmwYyTqDKKE0NBX5A/P9gqJt94vdKfGBjt7lPSgDthcUZfCs
7E9dXTet6xuxlqXLknXhQGISwVbNEM+mKHPJFaUmGE1p1/AekBcQGw17lPMFgVwXaLtGCbbfvYpQ
seXiQPJL43iCV/jFTGup8CW8bWUAwcOb8GC9joK/Biyhwg1Uqb2yjXOx7PZefjGrVP7BfPkzhUr9
588EidRpoQDqcIJ5EABPuvO8hUpAu0KKc9x2QxPGTuaUACITy5vhCzGPpkZ5GI/AlrVzBucfO9Lm
3ykbEfzggQLA/lRyaA648nIkvCsH5h+82GwzMDwK98K2XSneX/BJzYyCutKTaoadq9ySLTrRNN4i
wfoJdv9aTu+TvgEHMkLwD+RoGmkLm8EDghtVG27zhjZvxObSNSrQMJE2Nro+WXwnhHbG/pm0YqIk
LRlSSo29n9dqLE7TfuonFlQ1eJEr9TAZF9fGZmV/pHyIZaHW1nUps64b5o+btysDnGG3bq9x40W4
CNhucteDLEhZq9XWhemgiNZX4NhMMOBplT/EsWkgmpcIYRoQB6o2xGRY8rNjrx6FhW25ExBElNF3
gmHAeiWfXPVwAklq4rhVzrhCSv9WRkw5Slqs71n/9DwC5p4f/iuEMh0+o8Fh+eIpMO+ybwOWnQiw
3/rd0HsfnFnIrC9zJiixtswtiyVNIa9WygWYs+hXAd/81jEdMnt7JCzHXxp4d60vLMmGDjKQQd7f
DYmxK5tcP0YeZd/P1NJtHbGC+CukPb97eFWA/H+h+Kfmn23W0xeQQ6OMT5H0uLl4tbghyiA0HB8A
U/n66hOcomsAVAKbTeU1Th7ySB/5PKQjv9Ci5YIUkHIQCv3w5JZktS7R1RhgBshB11WcTnaArwaZ
w/vgNTu7e5guY/Jt3dULUzt4rhh0reGSESXgg0t27xNuNAHGQR2HZrH91Fe3oDuHn6DYhuz6YqVw
8xbXT6O27CFOy5O0tsGCOdeA7/FHhiPLN4KKJ5fFvSr5GvS0AwsIP9XQaAWe6m4jmOGncqRQgVgk
5keOAFgAFtBCwys4eYWLxGRxy7U4ousYHvX/l4yilxZlP2JH6BoV30pvTfWq9EjmTkmD8jWE92BW
OjMBVMdGumR5Kp39AMb0FlxO4/l3g5BKJrM2fU7naTGN+k5r9syqm30bXzH7ZAeJ9ScHstO6uljy
hsK4qgFt6euutKykivpxsmcpCjVBZsXidRuEfvWb3llFMPq9deUn0RShYBY2T1zns5cmKaTOhF+T
Lc+LbjjCSz+47CODRu82A9MB4T27XZ31Ev/QJrLCNoKn33MBKv8o6gcpoHzEWOjMOSWYRbSwFsPv
glSSe3YW/7biCB6ax7v1ZUAOe0T+fos+B+FInN9mq1qh+aoOr7LRBdxlRoiDfusjkqp+vowrtYPc
B+UGNnouJubjLOUC+2g+dul38LGPxIlF+Ka5KmSvI9vNcZ7VJbGtiLcvJRenJrsnYhv8IfhHnwqU
XVNRs92Sd3gsOr+yGUqy9naEtTSVMBCnyuSSsz/c71osuMzSWIerzUZP44ufBgrFhzMVNfEV5zU0
7HEN4WMC3ohe4+93qtXzcgmMQuQRey8YJJjTTfefQ+JJm8oEQTpNpidHbm6hcJaT1+303DB4fJS9
VY2jCgZ0ZpAxGRiCvOR9CIpTnGoDSGJnNm2UTDlK6wdHRZcXBPZiHJA0mu7bZRiNjOMj/EynZR+W
rCiYLXzm2OAS6DwA2Z6NCFXFW91FUlSU6z8p3ufGcBT1C8b6PP+LxWce2jwuAEGQa4L3pQCkM2nI
wgKjS6iaPz45/e05TOwbUyhwAoH+w53uEFtZew+nARhpO1CZ/TFDpYzhCkJoBaQfs7vQWG/NMSAB
7fJ731kCjVmT4xAWxS899qzxUioW/SHNp2B6DXVzZ196D5Pc8deS73RioIoHbwI2uoTRPsyOGBLM
a/G9eeMbTweGbAu0DyZmWMDLioYKuBeyZrJeArtCwP56PV3U6KO8WMzW6DjzuQmh5cmsqwgjMqdj
B5yMZuwuM71lNYDezxJaXmQgo1jEXnFTaqvVc8sdChfIUCnIdJ7O+Yi3wYEKgzXsjvWIaM1Ar5ls
VAQNYJfo+OHDLMMzfye1IZjvM+2y6nbETnYA+0rY/0SVitPLctlvXmimnumqZE+JVyGtPZ6s/ocO
U2OS2jj/qMUUt14xzU06z65/NILYsd3ewYC8NrQYEEHEzzGmStoF9E6rEI1NFeRQAcxuYbSzCF2H
tRMuCObs76Vive2ah/rqWa1fHVsis9M2sKH7UvjQ4/G3gMnk8eoZWMVk0QbC5b8IkJZnRufkCPIf
KRqsOCFRnkVZ18147+Mobz/iuzXHZQg0MbpU42OBIEzLV1xic0aUIZD2f3Ja9efpTJfIHV88xDhD
Fa5Po6RxETcApsdBesGtYfebPpLZ2+6c/frJWsvkS6b+uj/lhTT5dH8wYXiplYLR1eJvH/rzWUbc
0cw5C5NOl1l1K5kR6t2f64aP5vfC0UrSsARNSQsJb25HDR0sXItPzG6LxGdcwIRF32MqVzpiVcZz
v4qlWrVmX2bPM49ZtVdHBQW9eQoxsPE4ukJ5hpNJ9ZfNUjAps+063xjjBBSANwm7LkEZzQedfQ5L
5Sl0jX67XVlwDLAoeOYMGcJOSNpU7Mj9tMtASi5RIdafPni2vSOinPK+uZE22dx4+8YnsPd+qhkX
wtYcE2EbAe7l/FzmiTtrDXQNvQ6mp5MHvmR+MV2YcwoSMDBR5YW8P8wP0/PNMsNw0iDalalmsv73
wt+UdKP2SX1ghkYJhfg4KK9UnNHvg0dKplf0SVP+6pST1+ovXVbrFumleHsuqLOOJvsn3ARqsKP/
pSm6JyjHo1tAXduaemoABzXOhYEXtwSiwsvoRZ91+v4bg7j2P9LUqoyRigtzpT9RJCMRLBd2W5tX
Jbj8UrX9iKrHBcWFtmXuHxiCpc7fOcvBKSTF3EOt7O/CpOdFgAFR0gdStCV8IaSy75fQxxayq2+4
wRwzjDc/CTCn+rzIlZiKvluaxCdK1BTbYBGlvu/UPbD30UHqQXbsxZBTbYwoSf3XWWeM5EwCCXbN
9QG+5YrXYU6B9AF+XIqJzf96VTYsh5SicE7/gN6UXQmxKMwZIXu0HzKT2RAmt+vE4E9/eK7c5fq0
08sEhLi+01YTD6hcg16PTmfZBMMChzEStAClbJ+ooI0BnB0h839WkPLin+dPEG/Xj8Sv2Q6vJv+c
dwBbGtvCmCVGWuSxHE9towMIQQlz+qdNvILm1esL40xYam2E/UkEofeeEWB6Z/Qxk9iqqKVYYVNq
7i44Sk7IaXgQ+MsgGnirFV+yinyFKxu87XiWUHU7yttHrkSNUcgJbl5do7KyDcFvtTHZQgxn+N8J
2KyV4KD6sMkg+MKvlVFJzsySGQLKFiYYAVoKRR3CW3buU25LEsIQlbumNDEf8wQHwx0xXaFQGW0E
StR5BtjI3Vxb5QtWhhzHaw0L/DSuzDm9xTM2gz0SgomXmWiYSLfs4ntz0iSNCxpo0xksJAX/6AJ2
sSDjlUpRyk0INEjo6Ai5vhwli3KCKQq8VLKCezTQqAjfJNOSUGvK3CUgWudMUPjOTD6P2Tmhp4FJ
qPBfv2EdSTBz/dNck1DeyvZh8qmhrJDPn2pur+6IClhwNNeAiSAzHuRof5WGYKKEvxbXXZm7IzE/
45YqyB0uKcbmDjlrXtkSrjlx5wMX0ULK7hbbxYE0XSsVU3mojPxI5tT7XR9ClnP3IVF6CpdBoVrR
71sUfeEECyuxAhm5o6Mqq8aWd4/mvehChcJRC9d/6bhECduO7norZiMZ1XPnbg+oppoVW1wnAqff
DHB504D2w22ue4DI3oRh8K0epdcv0+yXaXqcYUKKka6daWq2OROZNs7u0dFJIBTrGPa32HDPEQNQ
qz3Oe4YESA9Gd1dGnF1AYQXOTai4ZhiCzyigaawgYJvxbCDXSv0O4AS0b9DjTONBY23SPfEaOE69
5V5QInQ8VYxVcOODtq7Ik0/tqr4bgKHW1jR79Xe8VNlmi7MsnBeInnz4+n+P1cubY8JuDbvjfLuN
FYt87yI65/zudXvP9QTP2jDCynWqSsfb0IvXu3Ulot+/vq8tlkelKxWAdLqbnH1SlZcvbSu4RcY7
TRPU2G0duRS9IXRVqKGoi538rpG0kniewJiq+Xu5xmin1lK1C9vaH0DTZfYxqq/tsnX1eRUIRf9k
2vZ9LWRQsMxhLd3z4KcE3mexel9OOBBRKTr7q1RwILSm/9cgfEyUk2UITf+NrhLv1jK/CihAkk4y
dfsfC2DU4vJpRq2EGsw/Jc/M+IKH9TOzBtaZe1YxU6a9FHqM61w7YCBrhgMiJ3rj9BZY/YGBj/VW
VqvYLxOFypAr4XJPsIUQwa8slmJkj925wQe0K4rDHRqSE1ypDZsfbpvgeaKvESA+XXqwNmKuGvpZ
QL9VRQwc06yJjULbgqDX5SCLH1gnQHPlqUvoE9lPHSwqy5UCW0vlrS6LetSSs8kZpFSSsn0r5cvI
rikiDrBsGhoKpKjqB4AyEpHOVkBbdrkw4Ac5PWJZV8dy5SEM04AYjTAH4Rf9Bd0cr1cxkOa/BFbQ
lIx7IXaPHYMUmS40m5QEz9u1J/SADlPfqyWcdGPt1clAKOS0AQANbrvqX8Ztw/hfuvrWYFsRYo78
1aa+vPV1807uoXbqOCx0uxNWZTh0Ci7IUce3zrR4rhNNGlXsVVNVI8WTOOOtLaxQLwKSm/cPnnqQ
iIPu+TxyHipF1WrXBGmPEqd6dapUkw2OqlErguqxz2jWrcoAyHIrGJg2dC2dN5Ppbl5lrzHHCkrX
IpV1EFVfEz1r1iIhF41qokIvnOl8xmKdNy+i4nD1F5UZ5qlSyp0LlHn1vS11Z9yOaCkVF7ES3L4V
v2LizX4+6QEWXJjSfGLb8Tvk9XfsPkjQBFHJoP7nfEjIAZM9ajVvhOGWCJcANaiR2GH7krag6QAg
hrJp1oFXrm/Gja8JKhZECNz+gk0OAqiiUnU71XWS7N5jNy5UkHMrS0xKSCoum4DG7mMJJu4HPhTA
gSm7tYXXKq4uhU6Ja7eV4iU/v84qUPv4lj3PBe6R0votzQSoRnX9FuKGiZW0XYugO0pewtxAr1Bi
DQ0wcCfuH0pM6FCV+ieBo9x5FJOv5HM2NG65eaJZOntTpDC7pN0ezsQqHAQONDf/3LK1cskg4W2f
JiI7aa/8b7tIdPDe+jX9+vTkyBsJutWiBWt+ktK6ecK6f8fZvSgUvKATmuhL1PbVtninAgunmUxn
SIg04/SzCloG//asNxHLuc+tbNWn0OHJC92MJlyqGbhqf1n5e5CdNklF6K5hCUC+YBJHmFx2CkIQ
Vi9nhVX2Ga2eJLipEQLoENvp/6axGAvCbyp5Pqe3ahOBKMtfPt8N7CnMEwCHCKyjIzhmBN1x8CXT
3kxE13XmOMU+9huuDEVwJuSTPY7w5BWz12r3AA6kmCKO8lJ2IwjGIPD/3Sw193T54oABovjScdYp
O1Y5rnGCvcjooF/OOWh9i7jV9cB3XfkHkhZtvz2sry0ffsE8oiFyvm1yKdfQpZrlCZWdK5r0VyJ/
Zgn4mTSJCGDB3wVodvBYR1LhxMsgP4Q6WujIofEbn6Ga9OKFecAEctmnrXlQTcUgf/0GuY3tnmot
VKI3ZDYWIGqhS2bjGE60lv6hB+FEw1SHWYgbF6eQoWDeqWAXx6mToHoTccRBajrRMVBipqmn7KvJ
gfzk9ldFsCeSo+cDbvCboWW6O/vvMXZyQzwV8tNd9A4FzoDEghn6UiWdGKSPwck/9nHtAQjw0Upn
xJVqk3T/JMDu8XsB/YznfFVhl8DENagTggdxI363hvqMFGPX4hlbauOCNZ/X44UWykkDpzae5YZK
LWzwU+UYaE2DHB+U2yTBJkZ1pyBWMoegcIYxUTSfeCir1nGo5ByH5uPD+mGBKaIECBnaq3No6Ua7
2gbDdj0qSfIlVuM/i2QEI7aJ8jI7ndp4E3MTuOolABhpiU24V3QRkd1HytVBhSOaWZcBPOHOwfAP
LoUcJ1flacW3YnwWxGQh2oucxdtZg4VwjvyUkF3/VhHEl77XkCOrq/CzYok6vD6+0x4T31vgurZq
PvBsQDU3rP2g9M+s4YBRwP8upURWOvyE2qG0dOQUPnS28bSli172BpgOvL51u3WIfrfcb8BYpLX1
398gNUNz+0w742asbExIj8vkPTtu/cvawcDAZw7/NT5LKX701KKktNxjhuG9hnHeXmrI+H85GbmK
XiJ1KoYwGHgd9UJQobRUqhyKop2drSSL6JTtFwh9NxwiiWXxyNwsbODcP6L13HY2NoqeTq/J0dBl
xI0uP6cMZ8siMCZEhw0hIaHaGdBOIprPynV03BchB7O+PoHtvgqh4eHsfZgCQuxnFzOv5JWYTLQg
PeQ/T4lLxBQnGhigLfPrzcr49SmCknkNXYAT7IdU9u5jRTQxlYvIXZtmD25S9+Dy9HtryNweTOa4
194AxkqZCXjB0xYGMhs4YXNNCDH73zd0m0NVdaX8lzA370GF0v4ZE7YduE1hyRjuW5zgjRdEcjCq
apFxebxCucKQWg8cD+KOmH1RO5yTLMwI5/GYpsZdagYquypuK+7VAvwDbAqKe7bXTh4DNbzHZHR/
9dXz+XG84cdWtk0Gpl6yAMD4J93rJCNI+hKTqVat3k1l0ZWEaFbsoRTG+0NMz17Xqvc/SdAN/VPS
rAk5uzLNPZ9jwlkfWke9Af4HHvGdzQlO1cP+R+3dDBJQ3VZ/zEWqqs3nqcPaVw8PSSErmJKyjYjI
XO9jU28G6jnygyQq84v4GwRO6+zFFDyjLXZjGZUVVh2VZOfVCKCFHe6nPB3OQC/2rQM60tur0pBb
HfTMajohBuJmyMnSitikDC+2AnV6/EPaOmhBVMMSfVfdP7Gj6/FiVfy2sw10TwVbRLrUVR1PtAEv
XXdWYZoafczNs0xupfMOJtTaVm7E57gIDEqdb4aAvr2rGyTVOTeQGfS+fbFzK5hTUVRA44cFllal
a1EyZxDp2aIhRWMfdMHjnxPPzbBtsWaIQPfRRUO0wPl48Ln+iTV0HAUMYT/AEl5oydBetc1EvxmK
Bv9dKRlilWO1Aa+DQ/83D7odlnn5wbBsJKsXGpfIffd/yOOp9z+v8m4JaRqqt3INc9uZAYtfmgT+
gdEc9wglXBrU1evjzkAAl61BqlUXc88SrHJIdCM3N6Ug2te5ZzfKGayk2zHRkZLc7WiWFiy8gOkZ
Rz+NLY+FsYmpGHHr7C/HcuTtNtH/AzmjtXa9qkq9g+FxZ5rLLlLxEYeERsYHtDjqhknpPk7wcCi9
vdCfbjQrYpx7eO5Clv19QvbfCcyMAGjtNSxU2J55sgH5G1FvJES/oBsaRl3zqUEjkX/A5oPR/9dt
tRuZiXBLcKWsx2IsE7RNG5iCUrXDlxGEoO2Ntd1LUs1g+wxz8CO2KzrgIUVe26PX/zzP38lAXJls
DLe9P8AQxcRIl6A8EtEXQkOXg2Lq0L5eK5wubMmfJ3lQh+3b+Jm082UqoSsvyQ511Pz2KLmnQB2Z
Uj+BRuk0UoPK3z5Pii1FqMASTpPJCOWx1bcdAWD/NHzZVPp5zDl1+ZgEGTOUsxGctReKyV697X+4
KFmSmsPpm8RzeZdVihnO7Xh03AO1yfQAXCF/XtG1Pry7pB6tnPEQYN/3niarlwTJCNIohQJMIOXb
fzmzjBI1WBMm648Iu6v+OzmQlfR911+AWPDCRrI6m6vbBx7/PaIHWAt0iHKxpRwPd1D0w9R5/CsI
z6cG8Z15Uk10ToH8xr1fnMzFg0n3FsMz/Y1j4PWA56RcmtOT2DLRWmt1HO7MhfYqhHasGGBeJbLK
eIr1zlq9qoc9qD/aIKpgp1MVvoxi2aWTNcf2wOyPcxIUgi8LBILaQShb8MjN1Cc/U0YqvaLCQwrg
OCdT2aazb7K8iMUdkb9IBXeroY1/cjanL59h09rzn7Z+NF6t2T+rgej2amxvocyNZ95wOKZsXz1f
PGQdpRZrxdDpd/lvHn3mvAp6Fc5H834NcNCe3N2duaMqSBrT4g/e4xafXNyKs/o5du60BNBnfksp
NOKVjaaPgjNjtJJ89Me8tVO0T2SIE11cnHxfs8BuqkE1P2ln8RF/c1wJv0R/Gk9/yITfOrBxlPrh
kuuznPm6dyGwzX1JdLbanqKOEQqsg5ZU/vajkMLDN6N/okhotr7jo+quo2emWCBDI9zYB8G6hSZq
pK84S5KUAkt4GwQFWTUpNbI9dWi0bpRQCckIO4PixZXnggMUUGr0bmnYp9CduERLS8M+KeQpY4XS
g6PigmuYNU/DbdCf8kn8swImxPgFan2rq0c8bO4Ln6/xGEPGJrEj19kJ7sRwJh8Xz3n2tJbYry/o
nBhqbKn9U5eluKlTgKLtAirbwLyEAATzB5s51qi+tRoy8c1XbwkiMk+VITvC1ohaB3Ju9bFU+0az
NwabSLUYplhIk0M7eLrpLPObGkvmA8zkPozSsN6HUxhD6TpcIm7tsCxrNTXrvT7Kn2YeRrCAdyDj
C10NnBq29uj7/EJBYYG2Y+KOhW0EyWSU9Vqlknukq8sEBD7jIjE5wOjxdJHf4s826zWQ9ydp6O67
ew4p9RjznhqQrbY3YKt87zTm+44q/cps+/swfSh/sigLKvjl6STUSBEWPleAwl1Tq0f3VBVAxCO3
Zc6gr7jsSUHuyi0XsF6P2jaw55J+1omoHDaPb3BpI0btcQohlSftfhgUHqDzKohcwmpz0BHBGJvF
g47H7jur/yCQI4MNlKNy4/uTU8wSiCN+CWxmQ0bO5Gv7gIsv1Pfnx9QGDo9JsInC6XEqN80aJFfS
BZ3lYV0UhCvdfHJyBhHSU2KUMOCEqpEVbCw/KZrSrQwImY0Z0ZChetR2C9/AtF883tOA8KrxfNDN
9o6t/yGU+POKeLcMcdWbPd+WUaPrOIU3rUJoeJNvXqBV6ns5Eoi0b63yDwQwBvySo4sAnFTwCJPG
cUjoEMtBZTg36ay8hxPbURfWbf2ZTxAbo8qGCggafQFPwBYxMPCGgrslm/3UArFp7sWdY4PE3DH6
uZ85EhmyO8PaUlpDm5llV/n7ANewK1fB/g6iLFIH4pECr8Eyl9RE3b7v3YxHRZyEvty5cW1zBgre
IhLDAwO6QlDhL3VNlQbrosyPCv/Ptpvkj4qbJMC7d9++PN9DmI2nnuUvLNeeJq4ZpO6zInwmVVDF
Vo8nr8wdP/bv/OjqOB8B7PDOmE/9YEx6yc0KWiSfIgs+XJ68Aj3GP7lw7bP7JmydcjflcA0OVd43
H5TTRAE7xyFGc9dG5CTHApOzOy+OPo0PrAyrb1t/qvLVWvKoON+KiGJ2mpN12NZL8IdfSRQYe9FQ
us7qF8g5wGKYR9XU0o8XVNkZ7fmK4KV9E5aXiUUb21xqQCNeiwjgUhguXPp5LR2f0rxs7jpeBD58
KEqlUyXbiKEisX8+wBbatrIMvLGegmb9JmJpY/1JvoMbaCCMJ0buXPJw2eg0RFBXvHCHUtwqdsyb
63Dvpe3Lo8z2rCM2CCWYU9VQW24UDcxjhOsBiIrAFZAvtlM4tkNS6gN7XrqRuqvEDERTrGKEV6mz
iJhkL8+c2vDMS4cVDXF1+5DGrhmwjKPnyEYrxKfT+HiYzcWHz16/VXenTjtMN6e6yh0KsDC0fHP8
19fSibwCNH+Gw6E3yHV4tgGCxuMs2feCfh8eg9ntfzdZwXgngnJlnc6o1plRIEoFixJlpKOQcsww
Nmn0G8s4B+JBYeGfWMhtapQU5fmCjLiw60hyBQmWdH14Zcq7uemOw5TKy6Jwde4fbzVd1SBczz6b
Z56h33eUgzg5JamU1vrog7QXSuoz/hV6WC5N1wA0lpsSKy+duJZtpwDXysU1sSrVhSvrp3p2yp8d
wC/8lxcKr8DSwH3IRqgNTwstnqRAVMVfB7wyLNwATRB4TNIdQie7lotSs/ZgeVhmDZVxRatuMJ8J
DDSo4g4nZgwOuzAIY9piIh724YPbQbd7umBYPePGIHjvmmPKPAAqaNcbYEf9rAJtJdJDRE2awgle
ZqJ9Ex31tiYSif8ydNQI713ouNc5W/LtQgxNo4IKQj50dA46C/aQy0w+pNMVhtgiinJF4JfQrI5s
FkKIqffa70aer2h1oMnC4ZqCCOzwLs2qkL3I6vhxON1+4umkkR1uVIpBqS0Leq0VaxazuzbgBpK2
D5lMnFDIV6EYzYp1CgO6gAdabN6f95Sk0tcGDolsn4qoMyUFJLu1miAPPUuo0b2QSkJ6x2+CRSkQ
l5DALJkPjY0flyXBq2AwDQmZtdH7/RxoSpH4ZFchY6+z5PhqRdoFF1/QKmvM3fm5PS4rIU2GCg9C
783hzLzgsiCMExgzaHjODeGkLauNdgLY39W3Fcf67oEwDzoforn90GUrzFyK0L0G71WkVXh4Pc/B
r74Bu7nqoKanmSRYOxGGm5UyiRvn3PD9J3zbMxvpW91ri9PF1k5PxjB74nLDZi6PGCH2Wpq/HZfl
X7uCXX5aiRhe6q2EE8Y50wUZxOb53qFE6ttMK1DV9BhEH5Gq3qqrkizjeP71+Rsbrn6Gd89VVLgH
aeIq3H3uc/hygsci6nd8rAk19DHs5CAVmG8dYMTp8qJjl5C3BatNoSSLmem09YinfRYydOfKNPiU
SaIUi9Yn//TCyMiT4FPNiJ6NeE7FwusU5Tq6/XKWks26y1kbA0Hm8EqDD+veyV6w+3iuNRr7b9GM
+L83DUwJI0z4PdpyUAPAeW4RrvIZ/6s9J7DOIRB5TnQV3OxQN+OaYugmM+Ylw2uxafs5LqEGjyf0
OHJ8KjbFAHWBN4BsM3qXlUNsX/KWNs9EO+qUpNzn6oDFUG0Ro+iVLJNKXfLxpR3sYxAVl23Ve8a2
YAHkdDOGXgXfvSHCsI4y0xxrudk6MU3StfVDmtuEkCgll+0kGt+KqXZBkSYnxOfMPTjaxHlWKzS7
F0o1Mc3T22+UCwBmH+ywvtuQgM83hxMoQFx3O++k7ll/BtlMJITRX28zk4N5b1JYFxMPjfVDMKTA
/3rHUQ6LflX+gBPMbQuQStB/OdRnZkBg1vC3ac2IgktHPG5Pfzeh6w2rv7Sr++gB0Y9QxWaDi3Es
K4uGgTO1KbOeHP2xJcEr+/RrFE9HXQjoIB/nw/R+Xus5c8pgMmbvleRE5et7hCkULj2wWuPoK2Au
3Fe8CaZLHNjLvaAPMYwos3niJJDPV6IcyXIvv/ufrZHIUfdfBjhaoxoSnjmqsNcJPCsfOmd0Njic
xJBKrun8ktliOqEfdTNu+D/eLcwBTuuyFmFfeMQmHh/Mcx3rB+z1mJoDm555jqlpYLtmAJrTUL9M
OtN6i/Xndh9c8bReenq/Am1uA4FOmB13aWo1OME9Ad7VmMQbG0eOsyArERjVjTDrQGXan7wqdikX
kFYndZpuaNwqJqyYiO6r7A7toY/MFjhDFwq3dRUHODZy+5WwI1jIx4zvyJ9kPhZAi3HHbbDp+pkX
yvoKG4tXZGH2RXF2oOQ4YgysxLH1a3Unv/TWRXc7sUXQs7KS/yolNhOzPDLGuC2lmijY1FBV18lg
R6m9TdLeYYbhfIcdlPJNkU09WPN+Pr6XZoitGlFCHZgvMuXOCep9q5gMxZu6seqW5YyDIgMYfWGK
Kfh5YsRxFe8rSQHe3UKki7y0Ebzn3zlE/N5lx/wbPZ6l9iAvQudQvtHi5jeF4AfVD+s070WSDBl/
TXmALzziug60tF4reK1H1jjwle23Yqimohcliqa3/vUX6NOZgVFRR3LsS9zgW58joZNyeX3oUToQ
9bazc31dArXCml8gjNnHTFiBxu3V5FWY93T4p8ct2rNr3864IzlhZcxAyi9ZFDM/G+lMv8Lijyke
/Z3Lcplyik4n6GFOCSmv+z9igr7Xt86LIEAEgiPp6fMDddXPwHfvS79vyJgVDdnVpyDMzKJpP0gk
xUU+SiUYxmu09bbLOlhRDeyHxpE9VkhKT0Vz1hUCXcPzeIp4gqtwhxqiMVX3xzGJcNk+nuiMb0Tn
t65JPze5n4M5G0zdyyZhTQmOT87MqHlQ/jDXPd/tAX+IgwgnugIFxsREwoqSABeMHv42WyU+4M6/
A/5auOnghSQw38PUsJvMo5f8tu7GdQ1exvQqgFFXuyG/dkEf+sfLVbJJH88T7lpCGOdT0rutlCUG
MSOMcPXRTyn0jkWEfBMs50IfdshZmIeSoRtHTBa0FtHlcM6kBTHJ2yj+4OVMhMuwDdMcA257GIrf
Y6CjQlOUyfR6NbXIouiljgMqSK4wsv6w/fkQeKXm9V7FEVPKibg3hP/ehaLjnzicHniM39azEHVf
vHQXZNFOduH4MR2di4nJB1kA+TKiW7IAL+JKga8NW2McmNL1GmYzaoc/tlMg19G51d/TzvjiyYtD
xekZvFZwiTJpxz/Rzn3n3i/ogGUuAMuNQmLWlBLhcC9OcEFoXNwcedDBS/6maaW2Pnqo7uqHo6tV
FbFDB/yVa3Kcr9GEFFw8PO+OpcHpXGgUqZQx36lghraR8oB56eKuyhxjvKuVICTwqcmRTSs+FXNB
gJYloktbeHvrmQTPRjQVJb0iQxgK3do9xyRXH4HNvVL5C1UJwV31U79oxT3eI1Rit6ChAJUj5xLz
4IsgbrkNgob271yc7nQCI7CEzt45uy5nLanI05mKwLr2AmbC6Vmdh2eZXtR56epKa8M8bLr0ef/K
00q++gBKboDdy2ycEYub1PwBgLiMRawGW3TUFxqPfIGElT+iWC/QPBEAHp33eYrhlioF0Mnfy+r+
epTKgX1WDcZVe6vxbcDf7+qm+E11tBI907iuj0tGPrTMbsjPJwwnaK1Veq2YPVrmpDgF2qYeOOWy
Y29v/5qkE0fymSLYUnldsnDDCMGR0r2W1rzo6CPLzRNEcMK8SydL7oN63t8+Xq2BV+cviEy6nMS/
fA2Au0TeIZNBPsgt83cBCIH+MxxmZLOLhJu9tapfZMpuFL9UJXmInwod1l+Wkhe33sorTtCqfiYZ
gmAdImdPpSp7IbYvC7MetZHJ1zxCMOfvUGOIsF0cL+fHANfFIOJYjaByrohWfXgZ0JVMstFOQGYi
xwMUoEWTzU1DbKnoNsC3J+NPP6tggnxVa79RojpcD03K1nGFjqqZiEjOHh99iAa16XYFebk5FLW9
bEtdIDJFapZWAxURGc/PTM2bY4Ikaa68KOHnWZ6yKo+/ll+/jl2NlQfczg6UxQrjzmO9zeMYvIVa
kq7QFQ+jyeSagYGUUFpvXivRrZ4tAH0mDYQQtHDNIwKECBkvGbneCY+JoHAm63zjnRKwqgKZzPED
Ni1A55G8HUTLOGb2n+fWr1JxsxpkXN4ySE/brrxDkUb2DZv0r599pB5F/6/MDP2NxZ8TKzz9tj57
RyPnYxIhnq+dhh3Yl3YJ4XrTO49JC5Lz1gkyJDuR5YHcgXW+Gs/JArPPVLo7FQgqhTQmuDbRNMI+
6kUtUbgl85T9lIJHMHpwWQw5qk9rq0bhGzw20pa/Ey+z/HIW6UgbwQRVHNaBzL3nJ1NXUwGGbKz8
UMRNKBS5Gxm8qGiNNSH+unwJ1Hj+9KtN0I6mz/GNxmbDP4tmX27+zM9v7nVqQa95I5UM73e4uYgJ
utCM8Cmq9Nejf70CTV9SzDh9IRzXHusPc+tJKbsrKfE9waZlkK18xT+bQFpj1D59i5EgupSK4CAL
OC7tGpGd2V6jVIM8GyQzN+8xQUxWMu0dIIVtLtUz9EPQn5EBFZ3YhCQhHVXP4smHCZDaVVg2deDm
1tjX5RANFlUoFuGH2LXjQW7VtQ6BUfhn+o/rI6Rf4eRFlB48fp7lCxZ+g4vLSjcozskhAr94sEk6
ycg4dxOBiKPXrR/j2sog2w48HCYSz6O+vJuHfhrWFiqlOWoPR2RZdYRCWH+u+vo/fNFoTet+yLTS
QDgcO6n0P1+Lv1GhO5TTvKnM0iz61totQ3ZHsnHixFjGdmz2vDSNU1t3Gq6U5HUi44186OfVasmm
MU+EdmtJ/++EjKetH45qvGHpFiCwBpt7Cao+7zrGCa5cA1tCA7taUEJBItZ8UCCvqMhWxgYJ4PFA
aCo02AmnO9lEAUdQaP+ykZ3EyvMS3UyB+z69EvE7zxNJnUNyymBbb8j+DOUiMxVm8z/EE3uZlrbL
6MseyFT+vjBsIQ706YJrvnISqpC+apWchBCTu+331qtTgbr5gDOdPGRpzCjdcrzoHQezVYF/QNJ5
iERHHKPDor9FOdZ/hiloHwBKFUnNvlBXT5QiltTSuaBdHb7ak6bKTr54lWJobvwjwy7SnNA3VaCX
taHYY7NmdLrsgjWEDcDyWS5lMoiCKmTTjZuavVF2UY1qqtzY1IxYdzG4gEAmR7zBFoI29EIiOVou
v9nqjP1NLo/6FBH/IT4vxcDGXjv2MielbOtvAAMQ6DC1hwyY3JlwBsayWGT6FD+r7xST5hWzHh1a
jZCp9OjyHtyMdgN/Ca2sF8ECWPJF/IsY2wjs28L9pDjhNRSPyhfDkTq8NQgDC8yyDEXM8NGJfMED
p8JZA1PqY5tJbL2sAX+aT0uNVt4ZpMDQSqNCWQqJhmjAThzEqD+Fx9Pcww/6EELXvguK6a6rFHdN
UZxq6u90U/OaWIobNzfyqAwTTmDC9n81QSx1+tRrPl+IbSxpGgQtzvXUn6CcYU6ufuCPNd4/Xn6P
8LqiCMLb2DW1mhCFJ0OsvULem5MdvVOy1WjpuOzfbivrDb81KwUy9h6En1qc/U8vyLXwSf3adO+c
TNs/mHjmyTIQlD6V2aa5ABRxcbdZHxSH7z350i0sTKz2stJmLOGFfln3rSNmRHW73k0Mpwx1T26M
y6ZFwm1V1FQ4Y+EEWULa/aq/eeG96U4gPwWPaR4ZVjgvdtd57BKXFDJXhUXwwocRsG0fFCN+ezms
DY+vnUtXPmzZA3AX0DtN8F2SkoAqg47MwEmWZ62uSujd3/2hycUJOM9cyx4gqzOBZJXVoVcxXdBF
+NNYf5HgItZ6Hft+CZvEXU1B1CtCnEuDpunvACUgtQdZCvuUoinyNilvOCAQKbJhLTEcgJ5oUaot
cZLpgbG8AEdmoMMBURrUeuR3pVTKV3kofZAJPUeB4IrL5+N7BJbUAwRO3Fe0zb6eccKLNOd7h6HR
E+pLgk5bcSPUvx98kaFbQmr06NqBohiiZrysJrjkRImA4r6NlE8Npk22V4WP1Jv4SHdGWWhwlBrp
hLHaU1bLsiPLp9kY7i0bWsKMNaXdM2VYh0uWpgbBgMGPC5yDaQeoZKzPjjOzHNpdwpJXYq7z8UaO
27OLpF3fF9RIoewIr4XCvwIeQKQhzlT0ZPyp+A5gdxBiw3hFGRgoaRI2qiXFA6YTyBzO8JojzHk6
ASDQSR+W+iIyRvpDGWIMEVBbY39bJdv8xYTUbGtTxtpimskp+402K96NgWORxAhQDMve1jAoG7Jy
0j+3CfkdB5cUKtHKNxfBnlmJv1XE5sGzJR1WVmB78i/yecONLI78Lpme+FsfNQb4aSPDu1DYTcSS
qmUfnntgjJdGMF9KQPm5fAlkmzdLRUfIJDuleNzlxaPAiQQaLdClthY3lqVZ8wlL/iYjuCXrbCwo
0gQZzHFcIs4jVvJFD75vuqz9Hk2ilia+wovtHNOVoCEyti0dwQK1H9wvIwINwjTqTqZvAonqBwgx
tnPgzT72YVBMgkknaxsJPnyogpvoJpfU830Orw5OiL9LOOGpANNvsqa0Sscue+Y1TL/IRhDEGp99
X+nSrwLyB9ZW6BVmX1eUZpLXXP/NWZLvJbu1j9ZlePROxNDym+g4LwMeBkPL7yDuo1znsU84A7Qs
UkQ2rKAds02qjK/VzNxZGdFNTdOQJHtG5XcVr6pM0rLT/WsFIps16F7hKJnJggu7NlvZri78N2k4
0kxEJoemPB5gb2RNbdBmo6XZ3COlAhtvsnbl/dx5p8JoZsqdu0rd2aqJGPVQhZirSxL4ZwPEB9jU
tWR06nYxA/+SaVcJ0UhIOfRSA35cYPgw1GrXQBWesOC5t2nJ1RTg6Eu4Up15J9kW5hCpNpZTrNiU
vjycgFfY7N19HLu1APcWn8kM9bTnsos0xOOb1VYGNCqW2AMms05UEZvBJ7Z56Ihr1pAkVOSU4NqB
0UEvpbrIdVK4nZlv/+EQaA3z1rVSNNx4anoCPjXSIUgiG3Mzi3amK9MMKYg30rMdKEzu34d4s7CX
geGhhUDPlQvByQoEQgByTpg7g8Mm5x+nsUqHrvPGf+/DfiM9wcVc5iSWQkvkA9tewh4uXsou5xpv
eyNvW8vpcZTQYDn+JLXmBpjXfCceiEz7mHT9uI2pOwK8mcUXilcj/GluNyoen42JoM7qxSCv9jl9
0BNmOD6VVX4JhiF+G6vPYrkW3id63BZSBfPwroyb2SMest6M8kD2+5/+5gi2aZLXY/aflKFZZLvG
wP8Zk5fyaH2xhRFjUZHEhqoDJ0D80xnQTjLIEGnpyY912t1S1Nzv1PHLYjmkv7YL0zytUJyvcact
1rAFy6/FY6+IDJ6AtrwUU6bs1XQfl0vN0eYZ138AtS816smSzTPIgXf6KEsWMawaA3Wst1ip+0D7
C0PPcGZIdAK3AsOd1auAvtQVKMppusU2h+iRuszSugW9OX+Osb8quh6p+04eSRHNnZMDcw4kDid/
XBaj/H4rLRN4ReAWwJeWo6Zqzi9FnSTg/+mbZPFQxhRSABiZibFzsILWw8LKENcZyM4y1/fJl0Vw
rdQovjID7cotkk6ADaS3UvzLoxVwu1qPiwnojIe0OEMPUDg7SZ5F//HKPw+b+3OffxqzqNGpeEOe
iH3lK+Ux8Xz4OWDO4lZoSM8TJZuN8eXiA4PBoMtvjfcWf1MYnZXXD5ORo/ybU1UYmft5uNswxQPA
ClW+Plzmf7eClpTyzO706/vdNUrwcbLawmOpeKnrkitDpKs97hMXH7q77sw48YA/K68jyikhnkhE
NjgDnKVTvmHkPX/YXIDdDWX+2DwZbhnc9ltJKuds12kw8gHAO0jEO38Q9RkE4/OlrB52yNwmJZ4w
lhCbvLLCZUWs/MzwdwqpyrUkCrZE9a/wZusYvLUB8aBfjaeu75598lxy0Ua86/VNXekJA30TcQ2p
mmPteG3H4YoqC/v68/hsEIR3VVvOuv/fwyOu0X/F9GJlhwvFmkkubyhevUm1ag6+5qI3Zm6yLsTl
xNvRJNBUdcCWcyz9m/zG57heVjIV+hyR5S9rBbYzvjjvsfYExR0SEwiFn2wSZNUK7AW/t55UnGL8
UVT+7kGRDd2eekZmJ1rjRD3FV29iB9BKfPJwekTVtd+DrXvh9VzNrm4BZGT1CjnbOjrW0tyB1qDJ
A0szGyCVLE8yFb1xMWvjAYxuNcU5XDlmK/k9GZDYy5L3tp9guBuRRvfsiCQVV5KwzH12hKuy1gML
D7XdTFLil51QPO8NQV3dltU1m0aJyBDYvuHWvtorNFK4tUPQQnrMbpRBShvbBiNlbYRCphqkiv1Y
ORek3R0OQFDZe0FjvfhplMynMGEL7BrbvDyajW2+dErzlWKsecvsTYO40cISESWZMkWegbVzFBlf
IjnlRtuenisZ40cMGFb9J6WTbzmOVbnPiyI47H4oaSGX2rVlxNyw0THiaT3O1gun7YOuHJWl1Mor
Swztkmj2tNj1tEHEALdv7FqQLcvc5UIVQV1oEkw7LIZlPPJYyfHwET3Zh2K+P99hJ1ZXYhv/Q2O5
yObSTgB7J2r+Roz+B3iruzgk2fXn9RDapUKfvWbxcQTHhbkWEKwUKMk2zir9BajztKV8qoVP6S/M
rVVCfKdJs+SWWGN/7fq9jJdHvnspnzl+V+JD1ZzaZuynNfWjzv6EkAQ2oJ5Me3C659ChvcMPb1mz
yD3iNQk4aRLicXo2oc5VmuhYXPaFgiE1LMgaWCE6PomwOPXMlgvDJZYvYAFVvOv+1NF5n2GxGf3a
unJy7sbx065Ejv76RkJidadOSL/1ywAgPNICrArpT80HtKtHMuvdB6OYvo0H6f6YTMDQFE/KoNk2
UgvAK+sWzVdOGU5zfyNNEDxI5TjOGbkHeEy873S2kJEy4q6CE2QST00OpZw7afztpTh4QDYvDuiG
MyKlBTFZogvm2s/WlHGgl2Am07sJBqnFhi9i4sZZwul0ZK+1irkX9QIggOYIvy8qo5C48TzjBQ36
h6GelfRVtH2qpZxrR/4I7mx0DLCFFZRiLQHxgb9x934ABS6cbF5hAPt3VL/TgEI8DD+zPOzw/MI9
2TMOcYvsyX4Qjvtg5/JnPTA7O2asTIh+hP/qdwUooyBw4BWTLqflC7CkYBapTTgQCP32x174EhxF
1VgJ8KOdK6vJMmjko70hCwPmSSqNh/GrcpV5YMeLsSXpiEcDCxWx9675+FJbZ5SGeD4Z7S5jgJmF
8HPBj+qU5+3vKQR+QMEii2X7HyIRx8iashg3nnH482vIUgAsSB8nHrT2kC9Ag8L7HjytTRDu6dH/
K2N8vPGFS3i5UYK/N2iWrVg7KK0uTn2XKqWCksNjDj51yNER62oCRQOqyzqqM9V9SfKS0w8hqTYZ
a96H/LQhModghAxSNKmk0b6mAqZBogUdNj/W9FLdRBVaD4EAa3glC1OW1mJ9NoeeyacNalSq7zqz
gmt3nOSudV7K1zQMi9b6CVpx3bKIG7CMv3HiD/FNeRlrUW9yvlWwrAw913gHSi+5uq2Ed01iH/Bb
XRAz9bFv1rnogqYysKBoxDhf7zlcVkQXcTCzSHaO26eP5aI0gReosxjspo2ynGAG7RG5sVuVWqN5
D+751jDWPLZzp50seOIsnkRDP4yetuhOyPjQfq5qMo67JGyTNP3v2qMVbA6KBo2yTtXJzyZdpE7K
p2jbzx0tPBMYQuHUSwWiKQ1qEjtVQFk0nlSiVCMAWtQ+ColiIq54w1hJaVt25yqyy+OsBoDTYS5P
C3AxgzUqRoeZbakYlNIEmYj3EfkIbF5iIDvk+c7/4QPUAO/wYnBwIGYVwWEfNrGhCuiD+ajNJiow
+GkZmNKGBiw2z6FEnhVRIslhaeYhQFYt047sxxQ7b+hAyAOdI4oRJEecMYNr/iGiLRs1+L8fVheK
qPaq/HbZanKDwwuPxQA1xqZw7Xb8/0di/s0zYVzvWAy/ITVipJoZSwM5HV5N1xMAPylDJ7o8eqse
AuTRBVWImNThJ/EBhKidvUMJeF+kwIP2aksGXsHtFXFtKlUbfHMmwaJaebI1jrocmOGdX9J4a6hX
zDBrOXIPZBHFW/IPFiDh2m9WKgDPnnSvnFOFkIDes+fpLm1R+rf2Ta3mIZR75jZ9+WZowkOUbDLc
s9CLDsL7mNKregflc2PInEiW4G9ElUKTF3PqaB/6PrxUdZhMkykT4BcG8MqRzExkemD8wItOrh8j
0wUIqac6A/77HODwRDxni9JjVfVjTY6Q/Le7ZSqD2F91Cks6yVDk70zozhgSWaMcVY/2f6vjnu08
KYv45F/zJTp98ZXpzgefa0cLNv0OCoqAqxkYggiAoz0EoDY9RryDUUpNmwbZpQ4t+7zFEqaZpBpw
AkYwyeVWkg1Mcb04GQnRdAFp/fc2J2AWJPdGr3p4WN0MdC+cPUMkhGetz29efXjvjNfdok6IPl0f
vifvBSkcKLKKZPHilu/+rQvFhVCUNs3uhJvAgUSgjae4O2SV93YZVVrZg2s2OFDyrxCdXsTsdNnt
7malh3Q5JxT1fb/2A0yjSPXcjmvyWMyGIF7xU0+An4PwhtB1Bp0wJjHfbXSyFH8e+52Kd/EphAaz
Lb3BZ0BHxaMtJRz4j+qz0wI7IU7atDHj0+2X/6WynE9PgMrm0ammFyOgRa0v6ipY+D6us44L2owc
kUYuGb22yf+GfF3hVxGGBSw0qwbdq4B7gQ9a3vs17coRriK5gAM/0Qy6UgkdNKPBEeH44D+8B1PI
Ebo8GqhB9YvaIlLjrf+p1BXMn5K0Fc/tceYg/+Wcnn4syX0GdF5QCVs68zvR9b5dkIC/TJuJJiyQ
qN/nu+CFZGwrglzYQd2do50Zb3I8VbR8gw+LG91V+m2S0GmXT4MMcqHNd0nN3MS5bmoDYjnCRAHc
Dpwb/eB7c88vqhW0PlFLfBc177bpkTqcGVzstwmDu+6UbJZYLjHuJveD1WjoId5/lJi2zN+QSnK8
tOVjldT+3Dy5/oEc3CVDD/n9UIXjW8CmqNniRzh/dpDvA9ZwYDihH6cL4XlauJj0rN2yTluW411O
hc5bVH1VJBFJZzjHbT36L2AZs00q8j5yxj3OpT4YMnBU72hNeE/ENY59dqnePcPppTNkdtHBivz8
6wsiZ9LYsU8CyIF7VpETPKbbRyUwLJk2QX1ftFWFT2YHss329WmP50qcJBga7In+hsm9PIhYZrJU
sunQ9505klvw2WeIz9vGGhSzM8yMxgyU4LFJX9VeOaS2zjElGXfusinLlRAIS7HKBRwFJVchYdVd
E8v3R3iQ8hXOtr0Rh8IkFpN6fmgSledfRdR++eGwNnjqGnx0Fzmnt5VYMi294SAjdVhEX3mHJJXQ
nZ1Txef0kQeXrfSuY2Y2Z5gBhV3i3ss6KIwTBK7xLzaPc44OiXp0Ery5tadrVHJUdlwwdPtNqXUs
1j2Rl0Au9nmoS7yDg765JaEkApjgHTJIeI1DXxdokqCsEo5BLG8/dyCUUXHeejiv/hBzORqqbKTG
C6TXGt7uP1lvIuvUQa6hXwOcqalkHS2ictrgIxebX902WX9BpJsVjV68kwSUYxACYej8YM84MhTH
7Cn9qr2wHSo0sE80WFyXcUPX7vSP1TjGSfEEBW2m7C1wSZbzrCgj9fhRAKONT4gypGssEGrUkjGm
n++1pTsYwi5mEv0b/5jGab83zFvd9bhAWUUVbUF5PPIKa3F13lh8eUVip039hT63R5NoiqV6Rm69
3PxpAWSZPxZdDLuL6enYepGddjQfdvTkcIcd+J/uIp2PjZdQZSJ3hNTEyJ79b80Xw/U3z69zyoFA
/qOobAeC8CFErXci5pQCZ5+Ug5XrpNmDS24Rk7WKncZmaqg+2FhYNksCKd9Y7LQtyTs8l+d9wARJ
4/KHXt2YRHHZqiK5AebsDJhedhPDA9CA8Xsqw3/byT1oXc8x51wMKXkpI9LjrWrylCvkPpIzcALV
UsLbEZX+G1EoylSv1x83IlsJKNx0FPYeAol837bOj/HAfx6WC/P32G+PaaFxSWHMwx+qyrIIMs1b
UE20Zx0G6Ure108E7wvGHlKmhO/Lw9zARLgUuOeJ+ZJ65tVYDVHKksXUMyxuiOYtnsNqKMlkau2W
ZRwpudh6L5LKRB1+Ke8V0K+ugZE3pNSoQnQlYL86ZYAv7SDXMe9gG31jM2VZIL1MYHiQnFW5EjCc
U6+TR/VT8nDN4ynANyzwkBFbIlE2Z0OzhmvhrfnEEv86Vmz5tgpbp4FoHO75+UaqXHo1YMeq/6dA
Rb5L9c/zLe7NwmzMO25qLcn3qLN1wKLAb7wNxI4akp2RDfFPezCa28P8lrzvslVNTlJF3mHZ6pAc
6lmRbkN2lrN5BHe83KRpTAADMwaWVFovVx3kb892BHvpuy6LiVoW4/SQC1XZ0hRxZdXfW7WHSqz3
TNnX1Fx0Gm2v4pFW9Z1eRHdu1XGzp5IGIX7OL7kyLJpVUzlujOJmd6YE9q9/YlsJdiWtA6JfKa+w
krAJJHFaqE/zj72fVP9zbvmE3cXoOGu92GcgobFBGK/9R7Pb4vLwNO59KColyrOL17J9OirqAETd
rjUDCybs5L0SjQruNiMOEGrn/jYHi8bycKGIUctdPdviDPHGuaFrFSLfFnh6JyU9Xv8y1i8ZHFXo
N9kdlK6mKQdy8xiWk22d35bgWpK00ouhANfJrcAIHUZoTw9AJGHxoLvfOmOSwYaLtEPKLB1NtUuW
7aksoakJiAjNp3huRvwMI0W+fjXDyuBfSmuZuliPgWuyhAI3bmTzP8uCKWKJ+NtYVCcOk9hiDGz5
VsWdatCvj0HKj7BFAmfj/fbM9+QGywWEfZrXMra8bwBpnEACJWAtVVkk2WMcXP3GXOIqXA9766ML
6L6KDErtxiXgg60cv5QRczRc8svX0Xj9kcH5MQL8eE0k4ER2LqNcIC9BuCXhIdCNvK2ltM7P6nTx
SOL2xeXisVW8ZBHIRV3Ww2uIJ/T0IpV90IudluTrNqpSinnOfha0B6iID6RyHU0LHijlNrICcCG3
yMmkgK6Q9HKf0g9AZyWh5CtHwjV9bC76KqeWOlgihqOdzq4kZ8B4L6UjFFmMhm9vVK7xzvl/quDW
H11AnPKcMIJz8sAiGF2ugIpqd8LGgnifiILmqxtN/LspdT5YjLDj9bPSldHCBqjS/RKhrxxGbSbC
fO6jnLspRikGuubrjPV5tGOlvt78mpaQCwoUBFWdBb5FnuThZLVvMBcntXeVS3LtMf8cRWBaNH6r
74JELbfASlHQ2TzFOROctih1bG02cql9vJ1aVItYhXeZdpozuZZzDxzp0W479pMqwe4Gbt1jFW6r
jkg/FX0gZgXpVdci7Ea0UvRtFitSuB+pepr+sAndQDpCRNO71MzK6GW67t21TS1eHCo9h7GiJOkE
EcNUIjCcN+4xlyoUZDKwzX+9xbPQ0ZgSiqyxcI6x2wf3NVu1kNzvwzjb1+MKqUimhV5pD3gkQs+R
3OscMA+rVz0y4UukE/iDuslqQJ/8Tr0byTlIOPuTHDz9+0ur9HLMcAXoZDEs/bypHfu7MZIZQv/F
XLSop9gXv4S9K1IMzCaf9pP20pWSv+tVoUTxj7fHnj7ZRu5kzg9zrnIltOwwPEQYn8TuA3w4/1WY
km6f5psaXI9YSWEUN38hAYaWaBZLRrCrO/sOCHJIkngf/qx4ipQ1S8gFhSuMmSBi2HFPkMgt7R6w
pdn0vcnAbmFJ2jImtDuHkcyggdcJAW8UYOPmBu8UndhAc/jVNo5p8AjKrKp2tYAz1BN1NDtGWQDU
+1Qu5MmrFlAs2vzsC/amayXO0h52UdLyvJQDL1JHKjQVsV9KP0pRjju1qcLMXgsAJnQy2iKdCls3
ub44qQOuUB3JnufkblLKxQaPNFR9A6R5GSgZv4qkeZ4KH4AAuQfQO1xw5wtO5/PxTkkLC8iAr0G/
SOvbW357gEAd+in5/+wIZvcuvJ0DecWvVC/+u1XASvoQI3Y4sTKkzV+LMEaxaoQ5yCUx7vj24Z3U
8SADuG0ds6zm5FCH3ZJU55ZYvebAMUff88QUi8zdH0naU5mORQcBLR4IM/ERwj3WVwVjW6GW00Ey
TqaISSbFxeyS+0ZzRtz8JKbB3JgScoei9+5iWVfQDW0mhxHjfLbSr81ZCI5m/6GqdzVCyqogYabf
22aqNnjbCuv3o/kNTRcQiOtF4SiSIcFy/UnKjGScWuweN6SRsZbzZAHgPwDNVyMHfwZIpApLGR6p
8DZroG/Yl/vYH7kdL0ykg1kVmVcUycDVD5iO2+IzOie0O5JSKiMI1C3I8T2UAUqbEmZytQ1Sb7kA
eBx56lNxnXRsF7pTiDmumQPJjmkqjA1HXi0G1TAV+KBFZqqr7CvEn9qPuLQqU8lpul287qkbwugE
88nCQWxjtkqaPaGGONQ9jzRgUx6/0okdwpJ0TX6Vo4IOj4a1Bjs3d6+L1ASrANq8ERzcmma4ifNF
3Tzjo3COwIT0y4MsIGTYS/2R859bGHThr739nWhVbJFzrnWlpAjUlZ+68ZklGdYyZhXlBhabrhha
mUGfpIGD9iDHFmBrRxwBg9SDTuoMDnMuu7WDmcWYDRLtxNqq0aWxTdousk9H/dqIasn5hE7pMu79
vIjOo+JmqJFYod+kBRek5LeahnlzJMKDAzfY/qoUIOc97t6WRsdXxbXSLj5w6CKgjPGqBkSII1S3
LOQ1yGN/2m4I0/oGeV/bE7BNp+YcnkzlE/ChInRsqmyxS9Ry0OABLAD1X2yFyZz8lyRRySThI4uh
b3S6FvWz9/Gt09QW8PbrC/ZmFe+YPJwlnUtEqyvum9rXfkZfQsdclwL8A9LbCMntpopIThO87hbG
ViusEJUexHWPbsj5lAfq9X9ZS8PPQnpDu9nDeZQ+WLHoKaR6mrDg+dqsLu+bKHXhcCE3lkrAFyzJ
H9aBbMWGhKLDRNAHkvl6uW5RMVL932HXpN2GsG6Pzf1Yh3vd7c4V7eIxDzya+c54ibAXk352Wg6a
9vEDEcf1+8JThe5I7UpdFEFJBv543yBgdCGcL874eywWeAIswS9T1yAXRKGbPVwkpFyGiw7JYnT7
Ae0Awp5Dk0R+DNtimc+u8OmqvtKeHiRcTn7A1Zwr/YArvmlANt86o7dephFbQTIffJzqSigDVMp0
1hQ6vWEO0WBkwguL1gyREGwQM4Vb33q/djjzOTtFAmPP0biAPc2uoSia0P5QqiL+9VBJExCypOzX
3PKSaakxIsXpB14OD+e+IpIfehfTNLouEifqAPzA/yXihw4o/rTy7JI6ZfuZEXKYIUO8oFm7Dlm2
jly6gUDSGl9nAQr8Ui+i+ANxBhV+GX54qOv+J5TtkTzXvv2tZE7UNmN6lq3yZKGLybOs9m/bp2G6
/9eo87tMu1swkaf25atq97y4POoCxfwvnSBo9haAg3Ks9SE8O0iJ6wS/Yy1zoYODFbyqXorESnl7
XKPQc8mnuDtogrSsSfRRytx/FsK8hkwX4JRK4+qUNxNcO3+9cDSQYpwOwMbd+qTVQR9DM9eGcp/g
FwhkSADgAESzduKs2CUTkfzG0hMTj1Y43rhkzPiOhrab3gkadsUUcdetaetK0DCVWPYgLXidu6+8
vVS2ER+2Px6Y44DHp3OCUCz9M47aNZW9gZekVBFzg5iL69rkdmTj3c7TYMQ9A6WPaVYG7GdHmln7
c1CP40WpTPB+QIbTbml9QG4uDFwI/3AIWEgKKhaIxbpQvfJH1EnjWP9bYY9HKH5zgSDKMwHdX4Oi
wD6UE33gvGSdYwBs+Ut1q8zTp11NrRyJ78xiGpau5wI4l4QZKVp3mDO19cQT4kLss6ytjlkVoL1I
jkYsot82362ShuNhAMlA3uBU3WUJRKZgwMQQNaQsAwSgw0a4jOCqzdH6TWe3MQZBETzQPqLIdMBA
jLPSsE6Ldjvmn59nOFj7SkSkMsoS2Gy8f7XHSNN61JX72X4o0IIWLnmmz0MmQ20i1JlBEv5I5TXu
2K+hgsk8aPdrij5YMCITb87OwYjxSYjPKqcpc2N+2GHcptyNu4swq19GtbHHQt8vBljxLlfoSG0t
CatIEyygPaBSpBbouNYyi/NnLKhRyNSD6xi6v9W1Na9/XS+hI1CcY+qMv0PruAe0rY3mSnIHCTiN
/Qbq8MKxO6/eem5cyNPPbZ2NBxyU7ahQTK0kWZ7syG17eDXX6vzZkPsePH8/PnFpEKGaLJAA+EAT
bVYVSrjKHikk0MhEL5Jlu85Xxb1JmIqPtmw1Nq18xVyuoe7fVnb0YXP/GXpwBHTXNgFn4fqZHUCo
1ci2MVW+LZmAVxjtpHXho8jFe1csPGDnj8ookmasGokmXpWZOLEJOpVAaScrYPCn0DLfTf7ZdbsN
ceyAdvjKD3A0vzjjCH50oPA7qF1b+3ERrGxBp3X/ODuYtUb7lTW7zmWuiaEV7i/HRUmOyyWniGuU
o19EosfCRrNnC4yOH6onpugWIXuhvD8LyEDLXimbAhtWTLrbM/drig6vw0/u/guGsKJuZrNfXlKK
qTzoH+jkVI/6CB0DMtgkYEbirT8vjIMM0TvcTwlpwLFbHaHAZH13B6P8MHabkKZc9kIyi6P+elL/
oteHd3MV1/1GiVdIwd4Jqma8VJspwSfqtzQ3ZhsyCrY47CQhGPDAiKXdZKBxMuKPhQTz2m/Tc6Af
oXK4h8zMhULbqKa0ovMdDXVDiEREMQOmV1xX9/qhjcp1YGaBxCMh2hpGhU4CGu6qEGbZpYqhLKQF
9Yo1R+8N2D8UAzMKIvgSmL5XuGOQQTQKufNGxNmQzD20iU50qRWxzlSZ7nV2cixxcybn9OYuaiS+
oTqoCQ7wSjVh9H25+5J7IsgiqcFOJEVNLe3ikARYPlZDqZV8kFd2nfEk6GqKl/e4xSRuAoVo/HqN
Wpp/RSwgopeSkOb3ybnhRvaVcNIry9XuZPcJaYori3d+/S0+nd/y6r0jI8icxRJrG3Kmmyhxst3o
wYJ8WWqK1ErU1Z1WPvEAeb/ZVc4VvS1QWwlxPe8yZj3pNdCyeY7dgXcCN0H+/9ck5N9p7Y0EtmSj
/0S+9eN9rXDDQvbraF0lkOw4jz39cumlmyOrVuEf1S/sZYE86XPVyvo4RZVu3lm2Q8Vr5gRd1nON
wwS135FJnHQO0wlBPEY+SMtG7bqLFqeN9IRZgTiQWif3pLPD0FTBzHGjy9sV6Hst6OR4Q8wR3urv
KLeQlTbBI8Yvf3KteHW2iI7n5046ay/v75gGQorl0Nt1+Ycc+qwWYJgddxxUTH9qPjx6B+XVs0Jy
bBjQiaFrmq2sAFlOSP2g3d4PGgX54UsmAOgKepzDWvirQBPkazqziFRbH8ZtNR3rmE4YUMq1LnT6
JgAyeZBvlioA13J7Cmp1GmlrrlUCXvcwWjb/YXDu/c+DTJzA09QmGOrETta3ZW+6KsVjf0Q8IcVw
r2YUup4TsF3zP6k/+Ha0eTGHqbDR+dy5OG195JqD4Gr0BrN5g4O+veQvs7ybPfGrx+cZREas1Rj+
9L9FmI07ji/iDrJOdMimX2kj2SBqwzC1Om46Bu2dKsg9uIPxWqbE+j3Gp+FoIqqn+fonvhfQbmUF
7VK5CGj/K7WW2RWAuo0CDSgRuKyy7UVXZFcynsirkPZbm/+gJVAQCTgLoKwz8GgzUqcZnaPvvnjz
HX9YMpXAKMoMr/gZgGnXcM0K4hcdeJGb1QORf7fpG6D+Tcr1sCkdsRAyUfay7TcXCN8rvSUfZk4X
qeZEgK6ft0FW8GUZ/UPHT3Rhr15os1UKmuxw699VYQL2LaxhnOPLIC4kfE6NNvF3IDnMwgCcbMJB
wfCVG7k20GR+xj3pipmYApo1vBTsJ3qe8PDX1LKDHVFYI8Wj3A/KO/UZvDtEPqIsRVaVCp3A7ndK
cOJxndAlzbEHZMB80GJH4mk2ztYjtNb8JLNLoCREbvD+IABPX5t68NJ+6JKmaLn8kXOEC8Y2sgJF
v45iUrMxpTFv/JM74agyQLUIavML58+NedDAHlXMtDq0VUiLrUvG8OzfdoXuU+i853xN1kw5q2UT
Atki34hJZYUyeB0CyNgfdpk5wtTJmi5JRS8DDc/a4VHraZTh1qz6YI/xYKwsroEtPjhk425sU9yD
9eEF0H1smwGiIpQFz/xeZlzoMG+GPFetS4bCFvWJrx85SmdmEd3DRqq3RtUME5nYdziqNmVE87LK
rf/67MQDt+GJANHCrNkdc7H2AS/Yv4h0+o/aQFWJJvpv9xs8HzMZZ5y05GwHxEFMqTJP/6m3Nzor
O+OMvQCQKSc2kOXLX8713hORB3j+rmOaH0ykQEUBTid7KhPJ9Hhk4m+gVdRragUy+LTE16z7emsx
Xw1H3GOv2RzLkFMozVgBt+J8Tjh5Sid2G1Y/VwjhYuv/DhRQCFSRHLCKQEA2Z9+moOtX0Lvuic4k
Tsjph2ZUMPiOi7nwZk25bbfwZkZW48ryjkDxvRlYXiOzFC36R7SLncfIivhDeucSXOkl4nUek+Pa
66YuSv7WF6SjJ/eRo6tR7NvA4LFF2sor5KmJUQuMmII7iTzKve5Nn+0wNW9vd7IxVawKZhWWkEXb
RMxWbaefxToWnXgJhLgW1r/0lvzlzzNp9Zb/LCC771NgtQjK0VS1PSu6PfXpV0hTnSMOMrbzC5Pr
Q2CX4ALxEZZYXoPfbiwqlWrRlM31bhtSszbYNjiBku5bPipfsmUFNhtF9QToTMKuVkCo4zDpCZi7
/+GnlVZn8ltplOdngRcwbUKld/4ckCMkOXxMvmNxXGHD4i5UFpWfTW2gWQpXrWCMyPlTIptLLW6L
9ZyL7Tg3N9DdO9gWspjpreaL8bUm3Lr7CcuZ95yHXP/W0Jk0Rgkn0PMnY5UWRvF3/Ju417sFHs+X
RseEeOTyMIzP5W1cDzlsDv95731fhZZqlOGtFgnTomY1pN8tkgwDBrGFrZUzXgNBOGCuH9/Z0RYE
XDSiK6063RQD84tDBqLFXD/SvqT9gK+0wwJRZ05P+N5iZNt9CetZR3nlMaLxe7BxmegggqOAK/OP
SEgXJQEZV7mI8XZ/HIHOn+5i8rm4vKDgHtnINdL/H4lioFBwxJIcHM72gsF8j5LrL8wWlrCmXqqN
jJqjQGV5nGxfdcwg8cQ2ltT2sYP1dW829AZT6cuvkaDh1dxDrK9vzXbbCKkwCcsfKQmNfyz6c+eG
ljkp6Bb3usUMPIwn8Ho/pVemG4Klvv0PZiW+2z5lTzjNErIGLRLJ/wr1f97jrSeVxERCjM79sAcp
pWh/JDqY4j1ONvdh1Fv5hwfwBHu0p4phJhB0ZsdpecI1jsRedCsT2ye0Sf2N4HmTp7IedNf0Y0Al
WigBgtY8IDP3btScFyCVGobFJeD6GeG3XKh1/uK+r2P5jZVKscNKKgNlUXuQWNcW5uYwbBjbYbIq
Zy812qCpoioXwyAg63HS1/dvbcXm1S55forDv+802Rh+MvBDhagm3muIiEG+EHut3tmF7LkghhyJ
2eL8QqhiTaUiLm2H5KckAj3fmvCDkFVBLTArTr5R8EtGvOVGZcmXMAJgGEUb7DEIJsbEyKfOK3+d
Qy/7cgo77SsUmQ5XsvCZk+Nc5kzBIccZ/Qmy0w0tPFDS8zUsfdQQFjPIiL6DviyKTxgi6nKUio7C
cCZ6sn3c/ZGcen6SYrFLxKTvRpuzZ8KcOwC7DvkDyjBiQZEl8inwNVIcXkmRmZQ9X3dwz1yiHVaB
cjUhmz/Nb+mv73VnLk/Wd40MIhFirMEPSM+kRiMBdeV+gtpHh1XumHtqdMfOBNDAMJnIRa0rfP7t
n5MMAZlPhc/Xgaod7mRjCvS8cDy7VZvpcFg0xk6xSrxD0G1HfCqWR3q2zIP7u4yoM+i1o9oQo6db
owHJEMlt3E3cwDtTQAb4h0hiqELpZQRG9ziFuMhY9gdf51OPWVbPf0oQRNUEeFR2ZAMz+ed/dGRn
72VEncwyAe5HlzEJlxfuEOo21/HhSaiXGpEKTssOPtMipO6NBOSXSDhUOLMLGcrLhLTgRzawayK3
wsc7ZrccGa9OrT6heS0a1B7hdphH0k2pMymqxfTv3Z3mY9qoA6lWKsjKeZlO2SyYIBSqv9Wx7Awr
yKFxNbgcuh0SK19s6hg6D/BSffldTBwEbGkkdkKS2c625f7mqEa936NmLskusm7LZ0HvpB1TJBC1
XTtMxnh3CWRMEQijAmvZNcBAFeZVTp1itdaDM0zXef1n+1vKNd5nb8Phm4hw7j58pQZ+4DOUoF1C
aXDJickzLeX6iK6U8VAADjDue1xM/LNsQa+A71tpojSp4gScMfsD30SywaEjpDukJ+bvICsU/oAY
iSSktT356Dgh3jj4QZULLeZXSGriDD0PyxO2zixb8uKZninYzgK5jBG85iu0C0XP5E5UHmlgtVIn
CtB54t3Ppw+kv6ytWxVemIyTTrKOpDdS+ep6j7jiz6Ek7eYi1BZexcTrp55yTkL0GNuF+iSXSOXx
k+YySeLpo89sICu/E4f/Ey8l6pxUa29nChEg1hYySiwiHEe6eBTtdrf+mucwriy7b8DyrSLhAOUM
9Dwba/xfotBkmSu4ul6VS882jtefzOpa3eKvPseYNKDRLws280F//KmcvattD/4cEow/tQvGPYq1
a5pOmKb23mT4XYIqwinB/1UtPoExZYPW5NiIiiApQUeg333j23/Nali/405UiW3QDQ42dOzlZ0uC
M3qEe/qJ/wSx+XZxwaTMQBx9MZjQ2hz0UIVLJojHaw/hkHOgu9T+rES1DA+2ZeHMcazBHa7IRPku
fE5BuNIODNk00wiw74zVC676XCV/9J20I546+CGsehnVctA6YnqwgnMU1Y3Kl885eGn8kX4/yPE7
PTW94ELakMu30pUGrrbom9jWcnMZ0WYdZME7L1FPVZu66CZ9gckUh8em5EuAKpohGJ0gFjnoOt9D
jpW+KzS0Tdj5+C5dS4a3IvIATtYFCfTlYOfM0Vxuz8DxBaraY0b9Hh0J2mbE8WqZZh8NRDy1/sfX
zoEs7UTyR+Dh+1WQaAmfaWelclnE3mdlhFbQcku66hxbfFpB5ypRT2VeC7euUUutrP7W6FK6jE0+
pQ/Va2xAeqCDi10pi4/05c4YWan3xKgwpkVUtMwQ3vtF4EJ9tIhPAdEIa9TVTCVhTWx7zMmTXtdn
d/ANBQ4wpzkJm4Cm61d6ilcPdV1PVziQVizNujjS9h+S32oAtnAAcO5BMK8zRE5RRvig+OmYer2f
5jDuAyC7Ik0EJHbkOG+CNgJjCzj9aoFvFIUe13d/vZTZI2eeOMUvA5h9eQAcQ0QWsmv2GLt3SSDB
suGkDIpcMK0gb+Dv9XMiLILqOxiKr+0iFbU5H1Rp9w1XZ3xcIS8GpOIWSPWN42MWkQajGgmh72NT
sbm+ddgd/sQquV71C7cAop0P8JL5amHkK8XDu4UeRBHqh51zHjXfaYDivQp8ckOcMBhcTwcZroLb
7xTVTl+bMcftwMTmTxPDUx8z71ZZDIcOq5roCUvQ+lxdrpEw1YLKkrWzowdNNUi9BGO/1xLjHn5n
OTCo+UgnlZ8LD5l1S3w95UFQzyZhPdS8AhwI0KV/mxB+N1PqkrIVguMOlMc3G+aqm+IexpB7PCUq
o1/WglGsXw0vnftBKH/P17IvjVj81B9BMR2Z1dtX2ekAk84A1SmTj/CTu5n2WhZprkiLUFBXO/bT
hgiuaJvZCTJUP7zcP3MqQuFXVpPP+ofywhwJvZsta438lL17VzZlD0iOEalQGcmLPjj72iSym6hs
vsNEssGsNVW+6yLtVVkPYgtaY2eG07xmEfC7WvMDDx7RX6gp6+6CnNkaFey0MNWn1htHXNU/kET1
w8BLGevK40p9KLKUIT3008A+FSOw/B2XuZJParSBpVvCNJ1EBPmrKeJf/IedMhkQ87L0z+5qtfB0
Y4f7HbqMZTfH475d/LVUaQL1oJZ05IQXPH0oFRgoYpAKJ0fbgIosBdQYuZV0bQo723eb3VtmicuD
5u3cOotuubEQoTM7l9q26Hc0DKnzlK5NUzxKRkre7742ANu2prSm5aA9kGLPJdDWIwIESOMFwg0L
0vhJvDmSf2tF4KpA94EF+EGatgVOLkZHd5EQ20f9NbcrEYEW/TkY9O0UagWFAIFjzXMTmGLer/OV
IZ1h/XoFlascypQfMEoZJVnRknHHdGBW+tDu/CUoNtuMq0nZTo/mKFOVUZ3zasD8cOPgciyOBBkE
cNjlMGuSVc6B8bjFfZHEAv7X6O4R6a53aqKGq3i5sQMl2BxjbwE2weEnDi98FlOXy2cEGyG6/yEW
QLMXDHCPgbjnooWzWt53WQEszBw4dQg/KmfXc10zFKegScl2GjQzXCXL+kA4AjhWgHVXxfD1mn5F
TciDh3CAOy4E89PthkJXFg5SnMxLRGAQCNp7BL2si0emoCTVZFQ1CZ5Pi6Ju0D0eBnLaP5hBnGeJ
RnasVrStQTkCiFWLw1wh6gMiY6xdtJ0B8NHmHz/QycJ/jkp2WQBHWxzsynR8wXMmUOS4JlFTBiPi
5DynY0CWdsmG9r5J7rLYqyNOnR3WLD2Nm1AXwyP68aza4kPHqYTmJxBPrmm07VG0y3HhF7IMNvZ1
tzNr7e0uvsv7ZsR3cOjraIRrxOxBLhHunBuoqLASmq/TXHGpPZW2ALXWLQh/W2eB/S6VKhYHedbh
GfFx1uXpz5w8v101o7MsoejHpQoTbKJk9XiEJZ0/rAmh9aBL1z14SzOscRjmKz4Pxg9K6m5DHcqV
HMDEkhv7t9drzvi11Iu1OPRXV1F84Xr6sP9omoQQt2PAeh+VoeK1rzsQEYc/mldMSYqU9ekwjxaM
1qVJAjX0dHWl28yoQg+h4gd2jNra5zDVrKGwwd1ycR5F6pisB3ZTzIZW0nSi2xXQz3Qe2dg0xgzO
7V7c8mpuC479WXfsYj9avV+JzJyWUEQj7weef2caeqLh74z89Y41nqr0Mq4vLrSb5HvwA5QZyBni
DfLtmHPKsSEJ5h0O7LDNQ5n5MWuLq7Xqxlz2ap9h5F4fPD8I9Vd+iq1GNPQBQ+oojAeVzZ9x26Nf
beg6epOIFFAZVGZ9CLi1ySpKR95qZVwVGHeNF+pKWZ7ZMvGezwPaSzKBduu/peyWTUfOnsyzLCbM
abEH6NeMUnoBaN0p2u0q0NWfG2loo2sS3OLChs7KsvcK62GON8aFgAKRwjVfVS/QuOE5EqFbM6x6
siulXd9HzSuyhUdY/F5SVJVWDuKy+1psxGEJOmGmmzOofE7iFVaSHr4iu4djSVPWPoqsLm8C2Ovw
yt0OVONO1DQ4vgl+La4PDS89o8M2wmKt7vUGj1CJyRe4ObXF9nhz4v1GkYLqp/6If2QuyUjSYNbu
thg5aKrClCYheU/haBAbi06nfRqDMoLAi1icqCMcbHK7npdfBdIKxUCeTDx6TDvcjeMaZByqYHN+
D1AAfeA6xfmbS5zH2aV5kBNQJZ+1avza4HVNm4JJ51pRskCq0kUoa9qTsJgLopoHEpJIgLoFC1V8
xdhnK+pJrN/yrzbq1PkgyMbvG/6wguUI7/ys3T+cEihKECVICj08ZXJk5pNgyzQsNG29rIXJOcRF
a8/pYqXqJwjZfyTw752SLIVlAifzzYYFBJOpLfdgQKn3UXCyoX+exdGrOaRzn3s2P2LzLIeILsiH
qSmTyKlAndAJNgD3Q+14neJkW+5UcLNicR9vL6QhVn8wWof5PyFXmpZhIGsh3T6g3xdHNQ1IvjLe
gVjTN92SzymvA38WwuuwKQvT0qvlmn79nesVm4xSaYddTT5Mcs8ZWGIzM3dbs7g3E7OAIKGqY7Kb
bPqznx4mhmaI4b11muiXrwwqBmHtfzgjaLNwPACyiX0m0zalaLxfOsM17rKSW7P0De0uGYXcK1lv
dfZvJtPhxUVzzZC2tSWyFfeKEChvG3HmrXVNoKvVuuMzsRHAcfgwkGzk5Kw1bDTK106lZiav978E
VmOoOxA6YS1cv3U0b06TPJu4fC8lM/1vt1+q9hkY8CuD34jm0PQYSV0BjgPI2tuxdT0WeKzIo2dD
aV96s3fmVLGqSNn23WhgYuDx1qQrQl/IUwkTeFnDXfjVpXLJAkEW3nPq7A2hzPz1j73obp6mR0iM
Sgt3X1t9sZ6xbpe7yCwL/wPpN/Hg9PsGJrsy8L7HZjPCAWngpOQaSvgB97rr/egejwFArkI+ykB4
3mvcb1xsjCUHDHPseGiXrk/0AiwD/nO5yLDoSuUpwdok2JhxPHc6TPBoRYnzFXXFFzQGfXGgGRnQ
agDaJRJO7LgQaJ4vmoykqXyj+VTllL3oo+BXo76JZSOjopcr/2qA6c7gFL0cjI+MEHobUtNek4Pj
mp0ZvipaeLlrOl/TrQrDsSXN5kmwtWOkAzySXHSH/PuvUv+nqTuyVh+Vr8Jp6eyaVR2tW4lhDEdM
+3LJlDHvPN52/v8/Sd4vA1xRaHl5VfNWhBxrjlUD3duLKREkJJOln4dMz/Zz/Oc1coDQIxGB+yu/
hpYiEJ4CcUP3RKuDTD6qVZWDmBxc2MZ9cDHrWJEsmjmRxJTfkYJGN+uRXg1VMFI53LfLaeESFZP5
yBT/527OIDtDdvwWEVBPh0qNgK/184QXequW32URlnfbqBmBW5uobMHNrr0c3PW3rVPdqZ3FH56i
J+k16m2rdCvtJRL95D2TLCPu4O4Y6wP8o5dj3ry0UX3EHP/qg5RDeBkZlFSf+3dNlr+sLjzQnBK6
afkaZ7MUZl7Xb4ju/Ol2xyJuImOEC4L0vSGOZSom8LxVKJpqzMNWJBFi6inP96FArClu4PsIUpGO
WaqOPXL2YsQfiqSF2SkSkCl7aewQFCipHHKRunlIcwkllA3hvopZEDR7LiS6N1yER9PbKt3g+5tf
eiZfhxum0QJtZgzItxiE0UbMoLbLHpnmREru6UxgnR1NDycDxLvrrEVv3Yr/r+9PSu9ldiJ6xJUd
rEZYH2Neob+p1FwWckzJiVZaNNqXCS1D3TAbijoV05o7abCGT8cRoUBMtGz3yxPrudgsHIFjNPmP
ebKcniLdvSUOjfrfqrEiQniGxqAL4nUU/XRlq0l55+wV8EfwmZLvI6EboaHdRbLbm5wtksy5xCH6
vnesqWeWNOBQq9sU0pp3Rf2KDfCvvd7XhnTnqk56N8EEIQBeeJ3DCaeX4+ILnz1FW2BM2LxGvrjw
1LANQi/8NeN9U/z8hKL/iRxQBCZ3PTvkRprl2uvPXp0gwR/gaNvL/hTckg/jedp4/pYsBdnvRE0h
TOp6UM3EZiWwDGMpKfVB4R3b+OZCETVkhgMGzUhdJNVq0r9FfXrDyw1c6Zhzh2xoZD2zMkU5AiFW
e/6XsurM3tjGaML4/4uLiJF9ql28GBeNif7Px265DzMXrTslIGrDRpUMvxx0+EP9SUdHgDh3GyXA
/XcrnbqzM8pYr77eYRVFHK/juqL15i48BUwjoV4FQr7Bt6vjLkjsI5qALHv/N0BoT5t5p0cK6aLu
QG7aI3uc++Rtmemyj10Sswo0gPk/Sz9dXn99Zm8F7/yZnpd5SL64PonwFa+vuMOBWumuD7YJifgA
utuQR6MUoiH+SNr0bEK7LgNjRYwEyeRThTREKwltIGETfwiB56DKzgGaIDZreAoJ2on+Z0FB7kbw
3MYil4FyJ95l5S0DmsZqqQvLfYN64K41Nln0PVZkW7zL+fAsSOEIB7qCUr2YyNcET+pOzy3JvpwY
0p0RV7aCvLqDLqa0Wz/UGELBCbWuzgfOnt9o4ki1TS66F0v0CzTbQqmrIK6FIDyTu8zTlHVGLR2e
HEbojhj5TF31x2/7mdCoev30z9ntDTK2kKnfFluWPokw6C1JuyfYWbyyXNb1SbGgZsAfEGprUMzj
v066s4noBf19mx3sN0NJtXLGMs4ohaFqYXQFXtmY1sdgBJirLO/d2udBEE85dKx+wOv/FKK9zJxX
SoZxT6Ds0f1lWn/c8BUwRuwBro7mSBk/MDFsrQbjRpdZ4w5rPZCGb3vJCvJY9m7G5Rl9pw0QGbZ+
+Kgw5NZx2hLjxjtS61fHBNO/yB2qU+UBtdndWrYBMPFEXql7deKnSKYzQqyZ7+zaNC66Q00f8iO7
qV99jN+0aT3/N81YcSBpM3uf4EDHmBpwLjZppPqMOKESopj/i7aZFCaHot0zBFpnUkg28hwkeL8g
GG7Mm6HvdcCbQ0qc2aM1bkH62UU+5QdPJ+5+KY0KzSp9lG1jWpJuAvoQpe8lqjhitAigreK1g0k1
zsrfieOzMJ+OCA9FlA02gXEki9S3SdjLL32oRpG0bzcZRJe8/KwnyP7QhwbmWZQymZVOTG9erP2k
DaYZmMALBzuLnvGQb31SDMHCbX+rQA0PT2X/a/AsoPWsFyNJMo+rTiJogMs0ssO73XUw/u2Za+lm
88GCm5sJDQ1q+cHdph5slm7G5HE+9eP8+2/kW29nABTYDV1HPbDFUoEaxTvRwRcjIdqPq+NK4P8p
SzP9GOuYkwwlFxKJ7EdQxBvIkwzhVw3QWtzggLl8z0KICm+344Izyewg+8m9Vn9/EFtADuBtq/Dx
+VN5aMilbyQbHdNUscg/q5+mT0myCTZJiB2vYCaLD79X2JLi+5QDguYoPvGYxAxh0d5a9HeG37sC
26Gm4FkJPpEFbQQmur1JYyk1zXOaDqlGfexqZJxVWs1fUTijEmTUwKRh9DLpDgbh/ComFrLLtHat
BK6hwveMQA/5vIZuMBP2NLAbWwsXtktbDeada0c63gcOFY0JmUQqDSER0ZhZvLydcIW0Py5yo7os
YgPkhP8C9zEDs1b8ES5+b7I1d5eMFEhRbYbKF1t95EzzQSCEjqOL8V25h9B5JHMVoB6P88486/8N
J5oP0v5MzJpY/BsXt01wXkUtBwIVPPB0Mk1cfoW+5IIjU4VZqnuP4ooFZvyq6R2JYiDDlEFdUo4w
Y0NPfC/x9ffrVBOml2qYZa0OUJvBl5ulTjBGZ1TtdTZih0UkQtGZXzwimmGinxUWEo2LTkBKGdgc
IT4M3r/ec3/6HwWep1/ydTdDvFlV58Bb8w0+2zOdlTl1fRViVBXtfFj1s8xLfjLlGSHWA0ydDRyd
ytPUDAons1zf9qymcwZTdur1gzOUa/iqJv5quMuOG0YWQPXY+Km7zn5MyXviEYhEcsTTbaiF4jYJ
BNQ4JMaM6UFEv1SIsi/fKwIsUmuxaapofLokxxPMqcuBIA9s7H/4S/M1YCHwzjb+u0YmQnooa26a
wfasgmj2iVyxv4vFjDh40OcpcaEMXWAmbaaDlkXjuMABnD7BY9/J5l/AhYE0gDbMw4GYw/+MGL0v
YY256SXfRud95IM9xKRipm+4Vs/qZyPOtk1pwTMMx98bYlGNd+xWFLSI1ZM9B6ZyssyFbTSe3XHD
TCaXigkRL73KLHKzltbse/jYySeeWFdGWraNQYeRmR8JD49SgYm/JbwEL+KHy7+Q82Q8R2njEtjO
rBopTVnTG4KwSJXv1FHzFKCnE1CtY/Of2STTELEtq+YPEMj2VK7O6/HLSIby7y0krhBTutvK2/Fz
XUdosOnIoOphvyPP0TgX6wTOB3Rw0Dt6JJu5EG1jeQyTwQw3ewVN+KkjakOPrbTIOnUIoekHQaz5
l0reNMwaODhmtjZ8uvOZ9puxuzOZRgd/ZncWIiaOofDgWStXVaHH0sl6aS3sbEOXOTewnYtTdE/M
LNGoXn7z+MU6v0RX/SbmpxqSn5ciJVM0mN9UDCtYyiDWo/5HgVn8aNlqDcnQ6YufkWJ2oVWFOOuK
l2lr0QS6ieZAkLL2yCV4lmBeqsSuBYu2p+wz1J5A6E1YAg9MgaamthYwY6JPPQAIqN2II4qDXlYU
12FK40q1YG4Kp9dRTaQ+Qrtb3gclIkw2b85xURhgWYyPxccRcMOr6SePy4ZCX+xiyGkN4EB9S5cV
ALlwOVnOXrwujWjGZ44YmgHtXy3fCU+B3iPZJz21/o9XIDEt+pTE1JHBZCQjWt5mTkGy07c+hY++
tBe4BqvMoxwRg3SEOOnWY2lx5hhTNP4YFDSuISnXUL6mrk0/Wszp4zKDHTXEQivdydtpl/Ot2l+1
i31W+B9gm+M7/DQlO4twHJB0UJ4ZdI/BhVhgzirUZRD5i92u2zLvcnNDIB/Pn32nxgzbHh9fcCs6
zbmWUbu412oD/woQPCXxOxcPTXysNCrP/99yenSHsFxIOFjUhnMdK+b1HcMTicH/4BJ1vnOuyTJs
NskBqMwacEBBySQjgk+SiB9fmqOjPuiKLYxPwlChQSp1UgrBe96mKb1iKO98Ce0SV9V0l3I84soz
rs8rCThzzkj4qwe/W8jVQ3xvTa8HChIpbvgtA9jUGseQpJu6mUHEzzU8AHzkEj7SxUk/WGg5HKRr
LekJNag18XzbKLh0sYrDMcjztM8lIcoZGn+cqmgsJSQTun1OJF5gqrWjjR/e26/hVy01+I3MCnOh
0rtTU4BaQH01no5rUQkvPN7wLgUGualiQbo6461CWIpFHxbdRSg2shwbTTBF4ZJHn4OWr44vvLnY
eR5N5vaJvbfHP8kuk3/KwCkFAIaqtf4JJ3EOFFUgWDZXJGTl30xwMPEnVOA+NLQEfJoiEEudSzZS
qTDQtBRj9rd9Ps9l+hb4OWRCEsz+y5BGxm6JozdpNI5RhbnRF1qf0lE7g8xmCNQ/y529lhVAl8QI
cw/j9jE1nKcCR3UVZt0uSMpfcno65YpBhxYtS1hmWEYa4MTNhI1S4nTOnCTRi1GgLvV4azKrU3HU
pXxHoFhTPgu8ycy53uj+3RvUp5Tuuu34tOH87wvYBmVwpE2hetiY9sK3ue6kCT45iWuB3X17ehin
cPofyzrcezB3WYAxxpjY6sW2lw2pYASMeUgtztU+DLVYFZACrz2r4eJBvs0US3Y5GxFGOUzqAk1I
a6eu5S6jrI6/xTRbkbYBigQFndHHv8Hu+UCs7fTr2t5C8V+al12l0UuguhPy2E3cl22JqHFJrr98
VayycRSEjPE9xrVBZoBGD6ldrcwz87FFt1k60AsGuUsM/70EJYr9Nmu7I8W1XnHz0JA5dSC+pGZe
6FqXqSE6vt2cO3tboQI8VbReIST2thtRlfI9EeGipM0gjdOylHkJ4F8W9Wk1k8QE7fBKhMLsjVEt
b9UHVxyklvTw14kqiKLQOmWwZBN36MwLQAmJy8u+5LU2rXTqnySc19QzEFzEe46nqK2f1ETXiZ9u
jUXf9ih9k2YT+Cq5wIlco/6FpWDS0HXkwTKnVkbwd9tnQc8VN5XNIEKBzsg8YzsD0KHlAF2hreCd
xKAFkX1hztx8dvvxV+/a8tjVH+rDxLiB0+sGpZCN6XD+dzvHJXdRezG9F2brkKp2v8omQhdwV5lh
oZLXvddvrq2myJh539p5HA7u5WYPfwi7W6X7zL3nnnMTJwDyetYFLSOL29zjjnpju+ijFnJqeM/N
WhFtQuPsJC8R0okrE74H8W/Q2D9gKDkCM03QITo6pz6I1UQsxigdwwmqxoCw+KRoccLRiB8VS/v/
eg94/mh+Uc85b8Y6v+g2oHo8o8Nisd+GWN2led0fUwbOS8vkfbRPhsuLqMMBNZzTYvODxNB4Uhpf
LsNVCn2PTlh14vqzpVKZ28E2QxTSuIfcYAJwP3kCB5zTaqoSdReOt5/W7pR9N8zsBl0+7h+d8zou
a24UZap/NyfMV/1/Orqlf8ZplOB1trd70muKA2ttyt2PYu3abq8DNGPO65Evq/YNYQWWe2ukGZ89
i7M/PjknJrZfyrqo1HcQ1M3NpqODpMUjRAqamh265ePvm3rulVkWkgSdhUAArdLoxwTzGaRLDKfZ
Jb5CKMOEdKwg7aw3pEha1n6cobbNp+MYWlwViNHW+TiHucIpHB658jsoH+rxbgqKG2ycf3PGQLr4
EacmeC5pZiwnvyb3cxQP24jc4GqyKBrSVCCc+CQUQvV6rJXXaM4DFnHV2r5MwMiwyNVs4I742vfg
6quvDKyDgzNtZKBj6WW1NtnWrlEwsKO2j7eIZvVbE46XgPbAVAHHgeCvLLImS9nF/FE4fSzoohVu
VxfLN04VZu4Z1reX2aQiZPPN3MwsaA/8cMyIbTPy+mCgfs3tCI91Y6rgTnCjJOKr9177INKUFDvh
47fU/zW+/Oud68FQaFEL5hLSUECmV1LfJPGOfucU+8YKCEx/+rD9X0n6Qt9VAFGk3MNyxxeZ02Ji
ZZf0Oy+5aVV+QqbWDp4VkwnDsk67YUI7lyDKk69Ew3KF9P7jq9aI9hPElB7TK7tpPoM3hU2QW0eA
MCqUzX85GqTbe8EEiWDAAVKHc7JETFW8n7B6uUUbGrRTUJpuEzMdIWlHBS0QckQbhXtrqlUQ/5jd
P/SK1vxjiNaGM/q1QGIYmaye2LDM+ZOZGbYYyt8Suu+DZpoP/FOxn8XHP/OB97dONZzBOd7vBTwc
DNdYPcI84cuSa/GW59vDglwBMJYogcFsPHFtYTisYcZjYcG1FHoeEsRB1IWqCgExldeHSXtmqOQH
5JOqhXIvkxOaZYeTPii2XsYSd/iUWGVHW7BNyUUaujLeGfWEPpAuI3PXedOsqTLvRB+iPQJK2NPv
vJatqPIn69pHh0oD+6YuRn+dyn2gK0FyXQG94vfLJ/r4LUvKZ62L0v6eD1CsiVnQovQnCTURK7B2
RUWYrbBShvf2Icyl1M5KF6/tfGaaeIKGu9HrPPAv2n5U549jveJ8lw3mczX1Q/2hPoEcinLYKA2o
jvZBgQUH1Zww+6298uqVF5X/2QlDsw8w/tMMvdatQcQ3JeNZio3HnRW/fHMFE1A5WiokhnRXfqLO
wlisb4gMSKKmekyVceBfvOKa1pyuRoWCBZWAX41xU9RN9BNegdgNX3jN6doMnBap0Ixv4z/DdCmb
muw7isKyJzzIbI7kTytKZ/OKyg+7yJLYxWeBqNMH9r/UBWu9zgmnVNQz3ATQVxPK3lUMIcu6tV45
ybHXAhMDR1bH/TInUojZo+Xkntd3X2TRfpOyRiTwY6BJa/HsIdw/uLAp2rHjJ8Zv4GJPPKzRINDe
O+3zbBT5omNh1qhnRQszKV+D6hryfXSLtay82fijFadLI2PT+DXc0DR3jykcbtdZPe4YXaVnQ6/I
krpoVF6/U0ay2Oab+WpDG5kjK/bCzOlQgYYmn60xx0pwyQwcDOVqWAdnQt9CxGgnv2Cx4SFq7P3t
losEQY5MvtXddnYAySfv4eyTky6XfRNaorRbiURuGNTUKqfEKe64ETWFvytcCzkeatobDVLLrHsI
qDG039TYIp6CsMsDAAjV2+K93aZtXQk6Yge3ddAWitpAdI6kojOq50mUNoojjFEF+/2okf0sJqdf
o9T40LOXFf4d0BSm/cij5VosxpcHEjQHxHmmS7mCkWGPmeZkkGavNrxC+S6jGUdvSwnVQH0+baU/
YSnThho3T5Amqmbj1EVdqFI7J2TOXmQ7xhPrnrqxmKPKsOpbumgHJFSLDhiK/a5X2aLKT4jA6p3G
L6y2LuLwgg1e9vVyHD2UcXwOdJ6uLQxUnWi91EZp/59oeJ4BRGosWjWrJAOxpRFGpybbXjhQpfri
AY0caslkp4RwIGMbu/lL4Ab1qrg8W7jJpmbmZcDncU6jMCk+Tq9dgbVDk9jPZC1gt4NeLfGxAXfI
9fFrUMj9xY2FZ0NBSo9sj09etrtoOvk6lzaDBLxcMoiO5EqCypalpuZDJVt1kYvE//EU1SxmdJvY
GXtgQ6km4WALHMHjyVqHptbLHP4h9Wo2kl0VNZY+Z59GdXGVFUtzcbWQ7BLvATmAf+j25Xs+zheO
px1LNWOC4Oo3H0kHMrqrYH8fgb54DfPR6WyiHfwPov3LGQJUiLO6QdrMJLheHlBOcj0qFZqPYWx9
XSL1gL40vUKV2KQnAxwAJwMZyLzTP1XQ+cnPzU/1bTgx0elcN7l+U9EViDt3KDP+1F9fKtjCB//C
rp3zUPiPv/JD/PKT8lzFs7fEXWFwKFtAAe2V+3lSjFaljB+QBkF+fhg96+jtzjoIJERkbRdrBQY7
w+7j2HQYhlMGiyuKYqbTAkMV75sMR5F1sTQyYQtYjKXO14wO6wNS4SYAnZeRZxQEqqRuz+G/p3qD
ws2CYbe54W3zNeOSe+6LVtSbmfcL9wd38vTFq3B7s4QzUUuJl8YrdLYSD8WbsfAdPg7PWpwIJNqe
YCII6oHQ1Kc3bBTyBWbruj48R/JSqW25w7AJ45m1Ee0jSu/xYXg2/twA+IYjBULVzyWLYf0kErV7
2naRVcGfsyIWxiZ4IlCR6jWmcAcWxfMHdcz59XhkjYHgMWLtpSK4ueumHE0nIv2JGyALf965/vf4
tx/u+g4U6L9VJh3BwxZFjr9dW/8rMbgcm53p+gqBb5RrdR+1KsnBUlvm79soir0QlBMaiHp2QBp8
yf+tvvqTd7eLni3bVmvOlf8QWmGSrcVPYJHO6BCsLkHT+F589ZILGP6ExwuvSMmmMsScCz69t6k8
ZVBrcJCqFkm4HZcZhKOXWXSsdAo7JWz4Tou0fQYSl9pOFCtEiyZSqHXGlQZAglT7SiOWXimuqa5i
u+d3boFpaVyf62Te8k8FBfPWS21AnzW5ZhsyC5KmZAYZ+fnnfbIo0Ja1RsESiZK8/vbC8qukIow/
FKpv+97UbLbcYjlliFsUtBW8l0AO+R+fUhSsjX0ihkMiBCS9LxvqRc5VZHqCzsgXI0Nu5VpNO+64
Kc8ANtLZglNtnecB53l/xyvLLCNxn2n2jeiZuniZTpjTM7clyHOecTGXfKyDYrC3AsZYGIsyD97Z
NokbP47GnMZP+4mOb35COjxPdtrqrIOqwdPU11MV/ahsVFF+yV2CerOUqHNCZWWsCG+SnfKxckFJ
sFXDHBstBP6BIccEnvSqrhPuL2NC5VG8Uipu5SAo/xY8xLrZstAwqaI61Qgl3UtmY0s6bEEgsl1F
VggnSZD5heRFlfhUT40bYZ9LDm5rgc7NsaS1TVx4aeky33aPYKQnfVbO4TkWj12oVx8rBTKnqeGB
3nzgVMZTAXRAoiM2l24c0jpBJF+xPZUbgWxoB0aH785EX+8VniTdf+/OFqXwGXd9a1f67dQlpP5Z
jCFztB2qKJP+NhshDY+UHnevn58hwni3JmvgQcC3+zVfONMTnZtm6FDtuXLez4ooBNliuBex68Nq
RCaJLtTVHsc6fcdb8w0NSa1bouN5aAYdgq3/iH6cbUR/6jE03nqElq9f6X0gd8XjEkTxL0PHy4NB
qOb5p9mpRxGSNvJU+J+r/mam3kSlJoTxKpPKO/YLoSnlAeyBWIGsLs8cK0DIqiELihchJCa97LE1
v7JwgUfp68ZUXLm/IwEAEe53o0ErUg2HHV4/n70S67ntDscxPhvA1oWUmIB2iyjInfDfzMWCkvcX
ltxndIZpoEqHNbSvjmemRrNB5QrOAeunuApDdcF+In/3TDyDWSarsrJLg2Sc6ljwGcdunDA2/V4/
qRiEOmzXSV/JZsyPX/YgOIHXY8Ke8kKPpZsxg0OjxNqBKHX0bHMTrReTQZCt7bs5lfSvxOp5WZx3
uyDTcCcG6W/2mL0edjl8Jy1K4tVDFmXIb5/APZELxm7e3jvS4Wb3+IYstxAMri+fOC7etPlztrVr
Pb6PexUNG8mMwN/+Sd+4LUa//8BZto6QfxpGaymcZOoV9lEuU17U7a3OkyVp3XrfHVhOCR1z63On
1UvXM2ycA+81fta1MDqQBaCyyD9ka49oM/dIYUqAeGiyA2z+dmPaB5W/24eXp58wtbnV2GCoMgDM
RclwdqCRdruYPKg0l9JhtcXQW80cEx3fCuiDbSOR7OETHC29eKJBWtywQ/bEUqLNy/3ZE57OZe2q
LEcQqxrCuNmvkzIT77VPsScXOOUR8YMqO1AUVNlku5FhcEfk6EBjez57ckJ7SmwMuWVa+/VJfgEu
Z2iaf9S5YEq1mePqNu8gzgaNH4VQFYlIAc38OOb07yQ0y2nLh+7F8X+/4NOymhsrf3LGYiI/TGv/
oV7KyMO+gfxxrFIomFygRgj7xUO5jjbpY1KEPsDUIXPThROwLPB2ZVOiP7smyABewZHXavLj+y6n
Svfs4HSHngTYmGn9YwgDD+SSauhxpHlEkjOg8+lrNpSUBtfzYuMIZmPbW7RNlfh3fzQG+XCAyoom
BcxGWRjXVck9xYCf5erw0SoIWGuC/2GacKvvWlkqzHx0f5eU+79NPf4Sha6L+UIA1wUA7dUx+J6/
Y/sffE7+94MjM77yHH+VJsSx+O3pg4RjIIzeA4rL39pl8WU+BKYa61ZysXJK2n4BRmZy0/ZtkA6J
YPPLRQherDn7hGeZpPUnFqTgR/jPGyYaMQCH7CJq6+WVtqJE2CbpXoHarQsWcjA/V8DXB0UzUFgI
Sw8hQvlyvBYaSt1eOmsamUUDmvQqz59JVY2OpxtivZW1/8FuXF/TIOdz3dNEvmTLv6NxAGHmDzdQ
/yW6miyLQzcV5DIJLZ4HtwBPgQ43xQq//Q5Ysei/QNtscaLV8Pw+hFenz3WL93ElzibmrNbQP3/G
fTpHxOupPiRh3nk6Mv7jzFnSNgTMzCXSbkNCcVHmiOav1tXpWFWRDZ5Wjsb1tOFxtTz2D6PhUj6Q
bL3j45534WnHsIliQSp7m3JBu+BshdtvjWavaoWKhJagy1Jty0Zx6qJfMWAz03/uvkejKyEjwYnM
l8FnFKuH1u7AYzwOQuOwLSH4xD6DUxyinhXeqPeyxE4CXYzLI2/xGeP0/SP8lRrBzvRyN/hgWnaJ
4hGXDZVoNtm/hxPGRahWuW2e2FkPFxfsuaIsl6pBNqhfbwQpMhxLMRy7xNezQ9MhA1t6EAK6BcQD
aBcN6V5/o4OrEvetDH1XeG75g2Zfr4niD9KufmaQahhXd+D8cGV6wGuIHYqyNia0MqM4u1lCoV6l
eAwvGUDykXkzZH3RO3QNQabrAfe2fuXEHkKj73HjtLYVWrTUbWwqubQgGpX+m2IBdVtW4o4qWmUL
qM/9p1fhsESMSXwvQQHfAMfJjbw+aYuIiYPHiTf7MrBZCu/aYDV0C9Dp17SX1w/I0oXVHZYyr8u8
JWhLsLy4XINVZS6Q3lwkvk0KdyLzTgVB8pQ5W37PzyUe/tA88BbRgyJSNxKlr17KMmXLun3RAGei
fijqE/KuY6OWr8ZryYQHv7Ikq5Xym7hfCf1nswbWIQpnF1EJLep+yTIoGcepFvSXw0UDHeUq/DLz
TmrbxdkT8K+LW2mDwt6cbAxrsScxnsXox968cDfn7/B2Sd5BIVTMLJpbRs8hhCPV/kgDtprUimcT
qpMs9RvdGGLjsC7h0Ni/90atcOlYcxBxbNyq/VFoLQyU7t2S6+DasIWAavqg+/LAK68crutVQEEk
OqZG5WFf52pZDUHn67PldlOjb8BEoQ/oNhneyEuuXk22j+2PhPtiUi3mWMgOvRYeaoRCpoCBgZW4
p4GrDAMGi9CIhHYt+U2cJqBLfYr3LhmatRYY7tFyez+o+VkJQ+CBIKeMlCWV8ifz4OcClxzIrXVr
2LGbTLWU+ktk400UvD0px8OcIZZ0tSHvovkyh21PE9WeTfc+cwKLQUsIkksRUx3mJGu83oXVHZZH
LtH76ICOIurgtck73fCfri/NAdlDm8Apj9yjMNYTtSrNnDtZ0/8+91mKBG/z0sM48NGEHKAQr7bu
fG8u4j16BWt4B1JBtieo2YZ2iPqdMMC/Y+0WPe2yc6Nubjfn0M7XUfqOkZl9z8lkyuKv2J3XGIQL
K3bO/4BmrJuujRCdfYvHeYv46kuzCUsuF/QVoS/MUSa0g/7u7XYikRIouh0hb595/Piiatlbu7nQ
X729UxMw/q8oQCfdudqu6E7tEW+QXHKOYRaC8SEeCvSrQ34sErGTpnPWZFJalhdAf8j1etGIEqEj
bJiYCqPNjTBiTL+ZG4YnG8kCCOJmZ+m9DbL0oJO4fac9k1VCRpl7dcilQcgqmJPk7Ei2/lugi64I
snSns/lOGL4wQjHJCPA+bfdNHpgxw8q6eAxNZEfS69sYwcUqy0PJUsDCikr0aKq6qCkID6z2gq0A
C6k/bG0WZkg8NvKPW7EfpnMa4DqJDASnPIgpYOupvawNotkX2QFq8QO/xS9a6mblHSNdAUVXAkC6
TUYacFioJNOK9OenQE1UbwaBc8JFbXfWj/SGq4NmYU0LtwIkUUIu/uvv5zTQcF7blYHuaz8Lt5DO
p1dcmGlaSzuR6sHIGRQ4uu0N+b3fjp2QtEr1eH4YQpdeGqC4JK0zKcgWgnN/CSqaIGXw4FtD5mmU
Yzd1qrQciGMN7u4DsPpTKVxx5aNgyayNF5FhgjwmLAzO8J1lRXXAJZZsjHXb+LLVrhL0bfELppMs
18pH4EoVJZqX9vRFq6Ox24J7w5h+jnj2bCuyjYvBibi4mScNEtbdoTwZzFHIXzAAQ2aHu3Q75hvA
7u+ayDZpp9/IQ+FfsZYWWYMb3N93ivv2dDkmBVJ5GYiwLwNJglBUPZz2OizyPIGiyWv4M1OZbeCR
YlpB36P7AA4J7NCi8r6hQSxzfYlvny5YdC+VU+T29PD8B62coYzyODKDgcZgibjo4tptore+taTi
UgpP41czDJDCbRQ6oHa1JL7JvwthCTbo2l+f9WU49IQjUEjjuDxhc1kIK1yK6pUSLW+VqeFssTBh
mx3bxYGoR4O1CIRQZU6TNsQL8Eu8m6J7s1W8A6W7fl0AIPcOb+eDEB60hm92+lA9qDyqDTCDNoWN
WtsDjNDTJKKp8bbfAViGnJvIo3ZusplCIwPMd8FOc7LFQG1z9rOv7XpMRIHeC1eUsBGkFsjAfCR6
tuZEXtb+fGa8ZLQWR/lTx7h2gsxuDNnn/KnN+THqnENxdD7i3vnLPpv8HMPE63tPBdW5CWrhJ7lB
1ZWQ3aKQK/mziDJph0K3L7VQEeacQDUlQPZX0DbkH/50Vab/V2y+yBUSK9wcyUWX7jwfZ39aNvbi
TA0S/xaUgGaRjQsW4QsiPDYtsoxbFoNg+DbelyREdYTJ5oQCspOfKlXLxkpPEbMidWqv8aOQc3vw
WVyCqjrVTmzq8Yp1V3wfd0E2y8DJc0tRyBPe0qNlFqg2L4eaUXCufcVQaJdmvLNfFNqf7XqHnxp2
hcTYnt8gJ4Huu3CMr/t5SK079xXkZ0PuhZB2t9Pk8zk7LSXRSnXQDxIWCtcGJCY3SON4akpgcOU/
97j9jmDRjmNLpAHxCgs0L5hOc+obBZs5U37QSlppARTd2lcsHGcsBSPp94Yb+pYp635L/uemMnuW
SpknQG//kF2ZtsV4JlN3+X7t2+RIOixJj0BHIRxIUDIaD/kD2GyiUuapu38nBCPEFMKB0pxhsPCX
iLKG+jQHWLb8V46bIasJx6hYxa/VnFGkpBEVaJokQxAkF1S4unmBvT0OqoTn1b+uOFFK/J5Fer9m
azpoEBeVWy6KVZ1EYrpOWtOo+/esUSumzLL2YLWDjjNiehaS8zzN7jmVjyLV1BldJsAy8BmQkuh9
hhDxVo6NkcHu0c8zq18gT9qljeMAqRrKiFR3S3p0whJJo37XZiOQKyqc14z/1KM0IyGDGLgKPKat
hkAYNAxNFgMKHwMqZVhLnwZUsHRUiDTCHeCCvka53/dSiC0B/NHuiTiOI4JwmNPXk2NJrYtJuMX5
x/A0ZvUEVw+QExrJE8Sgcj1/jwwJBZ5Pyvpf5WTgu6W1lwhwzVSvVMywTniJY/eA5JlAqpfKHk0d
tf+S1hc/eJo6tnERuAlWIBIzUvqi74EI0G0Yuv+P8ght2HoKjZ+UDkLFHydCwhPfvj+GlBVGNyNu
4xZ8+V5/E9+yjhLzr/E/fXKKM2fJuekG41x88f/mojYfrSgRA31BrbZ1gh/yxTPPNxwHHdQqySgp
rP8Y/84Yb88syyfXGqL+qaEd53A48uKs+MP+DJF42Czfx9KpAuoKKOoCIiWl1GlfgEZZvGwvP1LN
pJd1cc2xpkfKvGwapfe/x6ZPTfwc/3npsOVbGDZMWrASgZx31laOqn0yRoINTUidaa/cNKbDsM5m
1mozyhxkKofKbGnIgneRQ7DApG5iwU4qivFjoWpRCKdw5r4JE1T8v8Fx/+HFcOZvFas9N4pHyj0M
LOjOfH24iJl+jbqcf8g3V+0zA9h4dKUevzE4Wf9kkPad/TO63XO+oV/+dsWhWiaoTFke8uyya9f0
/AJIlhIYUoL1V4L/kdWs6EdLSfDWUHi1U1lVTJQ7PAXipOIioLxfZaBZBbUaq3krrc7h7iBjwSV0
idaG1cmXTcf3L+XFB+xr57rzfEJ7trKOT1JhlrU+TNLRleBMFvEeDyrfwhoO8qnq4NC0yRu5qdzu
M25PlMZmhqbaaiwfXrmg9Qo6rGPxuW/q/+gbebO15r+nRepTpBG8AWWk3iMGTBl2tiQD0gci8plB
Cm2UfEiY1vsQOIlQI3VbQpNgDd7Vs6THOgLAJ/mVnjiuPTgwrPR4srAu/E6NXO1eTUc+4v7P8Tzn
RI+qWHooZalP4MLEy2HNGTnvfgDm7URqnMG+qG9IqQmNfpBRiiynP8lM+I2LH3R5k30HD/3AcDbX
DCGMpI9P+iYw6Ey23p+MJhaANv4JcHGnC4oJuwt8xXj7C5adBoV9cQI2ZfxvWPNkEIOyq79tbbwJ
4Mz4KSjBq9L+NLBBIrqFnMUpA6Tc3u6CUL3/7+tfRfj9E4hH1mYC61KESLNi8+nTHpaGZiEgJlE0
Fvt8PMryT6iStOHRJJJZQcOB6cR+ZHFK8b46GIFbD5xthGHRS0KrHKlv118qjQSXMmeRJy73C8XB
+jy6siflGVOs4IzjCTiLYHweprsP0YakjIaJa0Nz4kB5QKJQMO9HVuXDU7mFrY7AFbVbb7OQGkfW
odOEsCb9SIF3V7OSZVg7+V5xsqDqEhC5bCYurGwmGbLwo/J7T+iwwc28ora2eBq6UTWZ8O1ixUvt
3Mx3BrU8fspyXxlrEXPZCi9r5XanrteZUnk7DE4f5ywXHnESuMlp0sNpV3KxsoMZSqoWMJRhdWC0
UuQR56ajeACRFH1Z5wq8rg5tTuPf6bZZajH0yyQj0/8SVJBPjVTfWFu/BXoQg2PN0gJ4SE5uGeoq
FvorBq1UuA1dNxoxpiba/9tqzHNq1oAdptK7jAS0IxNgpkPJs8JPKycGznsGN5ptIiUvG+fyojh8
PSP9AJslDyAbbIT7ZRWYy6u1rRWOW7JL36ziZ8cvVQQYh/VerXP1/uin7t5pKVC4LmI1V1/KrgO3
cdO+RRCggqUkTqEqLCtLnhho+1RziXwMk0Z07MXkzDK7RoDfeiyBVNVhg/bJfEXOiy8iPt9LP6wv
8MY5oKnp0o3yRQw1dggU4geOm93Kv1ObgNE9ZkpF0ZyN70TxwiIIXdi6eGvm3gEM1WZREu+2H4eo
moQ+VUHe9/+6sML4c3YnBdNwJ3C8nN0ymls63WGJ0A3OZAppug7MM+/RtigMeSj57nrIj1yV1yvC
6QnhNDpRqADv5GLhGDsGf3qfujj6ia2MCHWrbTO2cQ8CdoZoo6hQxRWK8eLHUgOK97LeGtmUbsuM
w1T2uMF4SspaBBTPJlcmDLqm1Zn/6jCHlZxkPNvRGEBzo+vVK+seYdbVjF+gjqVjm1YMPIv0mO65
u0nG07cBz8GWvZ6UQdNEIt0UlLMJfoZfPZzrMju8kc0ew7w3Tdy7Ahcwlmfwblt0gX8jZZC+cug7
Jb6KtGnKuGOiV4cCnUozDRAvUHLcwxgIs9Dq6Ra4xaOX5ZH75Ligw7rzGAXKwkwPFAqnZX9bCBXs
8DHlkHp1+3eFeSGSSFTghO4FJCtWx9j03Ot7Gsko5dQ/MIfWX8rP0rUZZ864sJX1TUGKjwoexMmQ
qZZjORrKozB09wPPrz0pnl+38AiKvP134fGdvKL/G03Fywi4/9npE2+CurfY7IvtbKs3DOHVN0oL
Hj4jowGaJGFy76JPV5UM/MulPfcf4dmqu0Zf+PlhEd/VR1i9dN00pHoh7/4qo9LiPxHhf8eqezIy
hac/Qp4CjqDA09NJ6w9/wkp6schlZz74gL3QOnM/Qr33L+Tu9BQVmD54Pj+q6BXzE+6gCKfc0H1h
oygfuyEVcP6L0t2JcWZvdbDQ/ZL43t6wWzMNfRvWth91jswoT+A0KigLU4ETxfvNNRMep/zdtvXv
0Yd5/4x+DYoFIDr3Xyd4nbkUAKAEY3gfWx733+U3SCwbwugUONzkIOazkSDE95ZeiadqT452I/2Z
WaB3zbWUOwk/d67AhwiBRh53bN2UJUkTPzCA05TRw+X87KD2hyP4J90VmR01mOq8h2GVb9ThcUrx
08mPvwlJPMvNFBveOh00IuJGTMrJMo8Z1HQA72vm/1YJmmeQBMJszJFZRWJBK9MgsUo1cyD/0tT/
eYrdJBc/C25AfHNMxIzA00BKrTDOpj7J5QJjvCm2a9wOdZ1G+f2DGwC5woWARnBFoT4ykTzStbq0
qpW43yroFzHzL8qSTYGNgj7p6ymlyXjttQr82efbbbw6YgtCifK7v9p0ePaKqLSEFEtIHHX4NZ6T
UlT631n9fcSlC+GPczu7cxAaVl1yPNR4amQ6NYJPK84WzMkr//qlsQQBunVWtGrv4pMlTF6KZgQh
tTcziKKBG2b76bq7pJqhSsvW2KpurMpFCcy+cblTLOV2IHg8yNWo9G1MDbiZcxhZJ+EXx3nMNJJg
wjdNMGC9bDcbKGqClvqCgFHVufsA2RzwxBU2GE+VxKFHYIfSL7y8xszG9HI8ZTBtgwDZq4GSW7Zj
lVrdnrtfj1FsN8zoo4tP/Tcuej/Gjganu3b4PJtpOFJzd8g1W+d9kelYJOPMIU+/ItuYCP2/KkJj
QBBOycx+oYolorOsqDfTCcc2uTnaDIk9DNV8UtVcUS/5zTd4xhu9ekrhKGg3lQ+uB9QxfH2Xx/1p
49HTkuFyIATFlWQXDv3kKaSAKNEv5cvHnyV8mhmgUkJkZPoUcdaSEIGn2hcppnmXe5X8ps8tRUgb
U+W3Qb3mnitne2r8EKObYKtXQPBWSpzaA97+vsgLB1DGsJeODPnkDNm3CNHp88PBHOXYbB8zHQXg
EgiVfd4lOy13PDdQ2h479VO2r5JIYTL3drD4857pK07me43mahu9keCY+NKG8TIZ893Hdg5z7LaU
d+SKyvNtd2nCj2p0QZqBN60iJhE4Clw54ug7Un3uVTqj6HQ4qaFToy9Skv2gxK/wKlttgCfIvhVl
kmhBeatIGev8bOETAPQypZrUOIqO3Ia2faiczn0NA6dGNh+oElHU5vZZtJShUxiVJkdrNyvzEAhn
pmRmfYzj5sqQPl1E2dPWcwOPVlYjU+1K/Zlr/6sMsQ8KtGKDPJhd6/Riz5MP4ZDP4Yxk6fXYJbtd
EhDeENXCfhfpCwhuM56niR1OMQlVgJZO8yzhoYxcVwc0QRk3LsLm6Bp+UHCoiXXaigGY2ilPLmH/
A6hYWzvyUENdW1T1clvO5aDZfVnuEZ1KfHLPaFOp6izoKc7WRttkVKqsvZ1rkRDjQakdj1FCxk5m
1IJqWougV+REiYD1lUxl/pQJ+bWu7l6QXfMpKcxHfSBI0+8EMJQ4r2IWvN4dgen7AZ1qM1yIibKy
7c+qt0TRHEQmgVeRVKnscrpcIXjVWpzSkWLTVRr8z0m0lFIFHC8sShUisTguZOYMHcUEoSZdRl0J
R8RozkHl4Z4moGF6dFv5OYb7Ul0Hr3rWXiqh40K7pjbU7FJpLuRnpvmhXf7rgcZZ7dO0dCev3GZY
CDKGIeS6rXa3oAdHDtxAUQn5yhbI0GLYDsQ6ejFb2diwJRiuZLa6dipvzn/nty388fPdonCj+pDo
7LK+5xQtZ3IkgrCUbes4CV/yMzLvdcJ1bDAZu55GfNh3Ogg8HaYy/bMWNiOTbT2snOJsYbxmr2l/
NSi2Mzi4nSJkWSCmNIeh6Rx+yv1LFwzi3z43eKtcLww4Rwaz1oAkgetlY5OU+N75sJsi3OgSwUvi
PeECZYnT117dVlW2csApt9P5WIC6VBy4KrMpKqeSB+hiIIKUp9gIwLltkNjwsiQtkQrKCI5hwBjZ
1qEdDgclmjmytbGhZMH6GTkPZ7VIR33NNEN6GABU+vkaC4N1xmUBww+JMtBvejcvRiw5HyKMpLQ1
H+YKkz43bF3xrhFPWAXMKaWMGcKIvIkx1DU6u/DwUGN3uVAd53PvBQ9QNduv4PN594IV8tt9Wv7s
65XDsyTQn4/xYpEpf7BDXu3UDfzz14Iw71XfJJLNKDcKLgdiJenWX4iLrxIG4YyIImP57Gv2ur4O
6eCURY7WEphTvBAXVSRmMedo6JwCiCfqr3Ui9P57MyWGEXMdTsBO/itdoRIhmghnSN3A2O/cbXPt
Q9oExzEyGr3tt+uQVbyAjEk4UO3BI0EjxrNmvhaSV137dEWTR+EEVZw018IvracCLzPTRm1+o8kB
8XTCPRbzytCHq0nbFGybzuKvyoDeF+XbQCtV7vhtP7+zys2ic+ALCqraYgcMkGGtGmIhPDNpoNlF
XE5pFBUT9+Bpx0T5Tbxpr+n6Y1rbBYpaJGWHwOEYeLvaXS07r+Rv5Evf+u2IPeitP5tVIl5fjjiO
MIlfTFOne4XbSaPq88wFu6utgK6BagTWD0+qAz+nIX+4Cln2AxAjgYQVFIvi7aIw6aGw62CskUhV
yAYTNrOLsQAXl9IVlTYsYfkueZpjmYBUYvhs9FZYIfhVY3QSLF/hrQceyA8XObJkJrjLkclZYGU2
y5jpnDaeU/W4LA2pW/aXAfC4Gj3+lsDPSiwyfrfYYkpDtPqOH+5OK46QMBWp9TkfQ2HZvDA2bJ6+
IzSuw1KH2m5BPiEX+shwSExMbbHGBq8yDi9JHKGovCyJXw6K0+0AJIGwPfIhhz9CrWPYdH1dknaP
kTN8Q/mMQ90kHm0sdKfdc6DBIA5SSBwGlrkWjWVffDoEKUELqcXAk8+IZD6tg+iBJw/KQh4EJ7E1
QNjEouzMT0ev8cw3Y9X1toe7JAlTbroUxKNVyDc4BExkgcWIfDbyUWZxT6h7CBaNgFK/e6tHE2sj
QV2mU6l3YTMTYcAJopJGAmdd5c49BpUT8AsiE5HlxcBvF4rAEmdNYqUyM9U4eh/THccoFo76mk0l
acvbhi07lH+e7I11Uuk9qr3jjHvSqphH+u7/Ipwc66c7h9JK5ammq1jpMCfZ4I6ZJvG3Lv5pucMi
YrgJEHkThhiWmyY8V02Qvvm5rmp7+9AACYAtvJqYBBHjvU8XPJ9u+JpzvVKEIfD9l3owDBSzHc19
vaSn8XNzki8CqZ+3Y+zEDP6VoMDSV0HzzjwXeLYmWMLfhByzikmPCFiJgaEdJ3vh44Orz5KCYtFz
JVhwMxZAulYzKWR6DCwe15YPMIEjrIFtw9grzsJGzXvbJjdhb0PzqCZoa0HjkjE+r43PImxQMtOS
zpIiGCck2DM30d/OJsYnFrF3vIAHddcwHZYt/ayM7KbomW9vYm3rqpPOLAbLhhxBaZdEJuHB1n7p
lq/003HNpBEwI58YpCFdNsbJSRxSpZQonsmhqxvh9aZONfKwB1ti9Pf8dnXXJlYCZ03rdINsCuuF
e6RjOOzAI+2+T559fhRCBnWUVFEHjFOUKSUWrzJnE6OoOXipDLH1IPCGb2SKkRlKfWCmro/5QdvH
g5v346BYXG0NOxuROieqNwkv5FjsXKDx4xTiORznWu+S1VYGp9AUSU5xmDlcrBDBQeSLPE/6usxo
Wm1ZvsPJcdFNfXFsBUKjuPR2e41rYop58XgCw+h5jlZ7N4GLWwCB/lL0npZ5+trSgp0vmUqjgRO6
vn2MwT6szNmdv1MoX1hlwfiVy24IZGXaAnBFLmAcrlRV2laqG2s6MOTs/Skoau3hsyz96hB7uADg
S8+jrH4s8zijWyMWn9vyyGPV3IY/f2m54OconzykhxAQrkyF/5POwa/kwsdxBTPfoCIfrQ9xK7kE
6l1PXh6pFqVOpJHpWSnO/1YWmLERLfgoi5tYIV3qRYPjQXftKJmcF+avL6AtCEhaJNLX9ZX4COWj
jUfJ0Jr5DZTGVKhmikS3j2gkLxBAmipo8KTdz8EWyeUNTW+O+ZNOyGFqq0yhRvA1d2MHIrMzpp/8
WR3U75tnIYhVdH5X9kxJhL3JB0j5AhThRG7kqDAAtS1qvU/Z7/QSWlUcZdvF3obfwuMkVjdbLQeK
/L1HT/EjsVTPl2ERERC7c/goSGqkYbGHZjoyC2ZBrnXyjqQ6JcD2jWtYJSN8SP3lnr/rVuZl9Rpf
vlc0ez7m6/d1OT+p5qjk/7c0+xuaoCiexOkadixMpt2l9QOb/EJI1KEto7StZDSon4IY9Z4QuHDS
bJ6XziX+I30U3CSefL25uKz1PCZnVft0mWhyplep2xTvJcBCCKYrfHC9AYQX+SWkEaXmUFR9oQFj
NjYAnvU4kIAkkzbI1RXyFMQSGt2/IfAGvrwOuc3uoNalvj/Tl48+jthqgiuHjfcmObEdiHMsgAag
lGUuiqrpY/csu952NDFEQdOrBbePKwn7wFStXKYAudqmBuXTIfhTJGaoO8wSFrNtvdNIGrl4bQkX
atyqbMCu2q8YPPUD5apFrtOtivgsPvzqHvJawKAUKEUbWC4TUkCBZQjJxZdHcayWgZb/mOxAGXdk
AU3XTWC++wRim1Fyv8JqW2bWCzX15qFPXYXoEb6bhG42fSIbMZGIcE613MnOAfBUEokdIIBnBiKc
OGco42Cm1ugBos0QxyluEtxO/jdaKiDnjDG7EOXxLttmYfwSv660uNHwGWxkP2j6fePiEjsjKMdn
ryHS8TCMk7JxgTlyZ9J2DpgXVYP375kdNG6ZIGwbeVvnASc2x8w44UYRZ7zLFDwKa9UvWg+EFwXs
LrdxpPe2Tq6acewgqDKkHtHiPb97ZlJqKyhY2CuE6OplA2qZhMMj3PNES3Bo5e4pQG2v3ZBFc3/+
hzS/x/MlKk+t3RQZ35xtsTTewmCWZgVQgFSHri8LPPr+RQobsN7Lik6AbMe0SDVXeRShrkUs1uCb
lrBiZl8vuat1bQTMCOOEA1RwWyePndnD8n0d2q3L2xOsAQJU8enWURXHofm0m4o3On41akLlhICj
0Y6//u/bGw8wiCBb5hlY35gH6aI9eVBnBhTbwc1+2od48lpAPze48SLZISuk8vJ41VuaobC/ySYx
BCSbhXY4AJrek8JYbWI+W2Uyqbbw4Bi9GXZvTEqSqcfMcm3P47EQgj5cB1ftXz9mo6KuoZr04NvQ
w95rX7NIzaus4dT4VCH/cEuxsN3J8/7Ch8dkclv76YftQeUdPgA/pJ3MlYilmjLWgy3DDdW1r+3z
L49WY4TTW0BviEa8Mp+bm8HyGyjMHhIN8sGOB+SSh/Kii7Ir3FDa+ABZuY0RNaxLECZhHdzFDdZn
Skiy6pQBpuCSvHIYOWfBmWWEMOJW7z6pWJfB2p/fNcydxFSFGMDiYgjV0OT9w03Ik/HdoDhfxfsU
BJRU+hDnvbsHXLF89GkI5nhn5FOKUqBUSu9JvY7Uphr8ghCq2o94fixrhW/n5xNVLz+IlgLXoqoY
A+Ta/JgyFJ91jJsmDiqFV/xTzGJacZPtSYlJENPdq8pN+NFC9VcGWn6Mjwsd9Sed+wb+lsogyYtU
Ks2CSDm5zaaUjdd/QeCf8eYbyqigQwPmrzYmq3Of7GnCRugtFypgrVlKGgBi9f5qwZt3xOy+9uB7
r0H24Pd65GnfIB1gohzlSZEHRZXPz4ATPszvS+uCJb+yqNYVfEuLhNZpLb15lP0qnrcn5LqiIZdD
sk527swPu54B0QHY8xawX+8UeE4fYTcZYQ4hwr/FHlwuRTwo6ftzUjQOfmub4x19cOUX754oU4jT
mCkRkeJu+JTZgi53silqM02teX77JvjEquttKCZEbbjFL/VEJ6EsNf5hJ06kTnZ21wG2quSHQE2E
JhEbM5oGwiCJUcl6So4uIp0c37dHKy1+I4e3c6bEp1bUpfWD2PfrMUeS0BhauIOVT3noQpqumlYE
r230c6JeBH74TiS5U/zQB2Qg9ZCJNlAv3Zui/SmS0yB3xaLNg3e8i3BZiwWYQ9vbjLvHvf/XCPtj
ON2w5Y0b2UUUgN0ij9/qqEMeC8wq2rzErMc8WatpderI7m+0XJWLLNZJ5Ifx/lYD92YSAwysXoS7
9Z7ZJE+5UuGb0qIWaeA/7qzVdYlVwUHcjh+7Tr45WjfdzKPEvxVXtZM4mLm60zqkT9nAzeUxBWRg
pghHfAfbLR2tr7o5Zxz1qr8GHMfDdW1rLEXIlLuJcC9Hd59VTB3HvLWVuguV5YDxN1zC+8qtdNqJ
ngtdBLpDR0E3dLeqczc/ZxQFWzCV4RxKUhfG1tRQI6I39QHu0dpZpXgIuJwOlkJRJQmcXli+bQ2o
lzXI/MQV9t+tyHs6DBF0CrUXd1J9Sj+1M/9Z/J/5kZWZ8r11qIAckFJpzqhRkQ5nUnrHCN5/bKMB
gGfYySQOXTkstjlTNc9KJVL7lPwa2VeE1j5PTRLrihIbPlX7fvwEA0YLz0GA5R7ODQG93XC9wlLr
IcO5LWChSE9g3Q4rkvGY2cj284SnmeUofN5iwHv5EDLOFdWOhbcB+CW/AHQtPBRUjSBEEBjLvjEC
ux8fCqDQlUZXZuitCIqxzSKI0UipC1uWyFn+CNaG9vF9n3Y2TTB1x2ruSuZQtpbGeIESmtGstXJR
5B9jY1A/u6AJnSgd7MuYx+EO/KHK/fyf0uR/INbgr+HNqd03z+XMKmZVsqL54qw4JrCSyNljqGna
8w8fznm8JVuyD5RVDNImTkt0v9pGA36Qm6KtvVwXfP0lBGp1eO1h77Mo1jHaZaG6TpCMnW01TKW/
jbaZ4PZRN0HpMNXOVI9/MbBUyJeclQatjXTdY+WXT+I1hgvnoSkWmuedv+aIooflHPw6fHNcoiIG
6ylelJtUuO+Ie8lW84SWtrcgjC9+jBQHUo63y8trchmvNWrXL24T228lUHocSG8E5LL4sh4fnH7U
+9Txkp9RGe10dXekL8hlG1+eYF1hHAsNeMOg3wNgcGfDAnfHKXXNyf5bZvyHBXbO0oKMkjKOFoc0
dVAMbVAXU2aMPF3Cow6t8f/eQepWYiuBo2aXj8EBJ/JWtFPh+ADbFDoUuaTe4IOSxNkqnDcQrnk8
xA6QuexfMUE//xfJhAw+tqpzzMJ2F+BneI59DxAhijsKQLAd3wJMgZ40WyKxm6+RHv7P3MLr0JDw
FFEe2suPgyKFk1INngsI8bTqR3mrEqBjae1wTi9uokuKYUIk9geV7aSrIlh1HKmfZlTn4e2oFvZ2
h5rJFdq+LB6pyPxQK82+uiuDLr60w2I/8sFwtzR2FqKzvGlxOJYCVeoToJGuuYGREQhpkksRq9Ya
SDrHdTomwzFadd9QN1SDvH/iIgulWr3XBbbNUcQpH3/hUeYsN1W0DQE9HU3J2/j4DWJ1vxDBIDvH
AfVGSeVfBiDP6Yf5meBaGp4iGIXFtKOPoNQM5vEVup5pSPjmOKQzIRITKjDf6kNO4YmQ29NqYYWS
5NWrCbjsjZljzFnbhpgnVBt6UqTpppg2lOhvr5cZiA/J6cgY9dM3m0ybn+sNUVzuKTHkHvnf0TFm
F36UTEmHN/TULnk0s9qmEsADrjm1liQgZKd/iYBmnzZfTvx7jnGd5DiLBiDW6+kgQHMOZXZSY4VQ
jpDNFDp/+s6ARrgMNI8m5jdvytYqAwKaWQC5HK2L0h0UO7RXfe3c3HKS8vS+GqW3wr83eNXk8L3M
AREhTnFD3cXMK6yZ3/9j1rUdh/DtyfEcImpLm7xEIulJ9ViCAkaB/vlkFKEQESie1wEw00O+HrUQ
FvMu4/w/nMe0+NFHOJl6gv+uokMGoWaNgWe8uvSr1Yn2VU0GSM2MtEUz+gGDIlTFym0P9PCSt7Gr
kwXNz04a1I4rm5YIcrPKl8YUEh9s95oa24cgspmwqRKYn86wj4suOmIluUnfXscst97QGCeJ5RmG
Ns+0Nias8eAy53eJkGEPm/gX4biEXtTn0E6nWN96v6OPoWwvyGWd5zlxv4jV3ebFZLfR+LVdungq
OOv1rx34h9tg5SXHHdO6DcGC+ucnKR2zfJFBM9tMpay7BCv6fRmHiwA1iezWtHGZAdqjNKKTtdLN
4UGsUlks8M/zbpyGBe6pr6SaJy/TR0FfdZY/LEAcPUGjfHZORt9ZQxN95zAL6Tt8ErYE578R/N9K
hLif7qxfSWubiJPAdqvLQZ8MzolAbnysryjde8j9zPmkoBwgHB/XkHl+BmMkk5MJglrqqtCzAyFk
Fp6sCbgZEHMRd1FPpfp2xZKzTVT9JRIPHitw/mmRLUx4Yj3eU8+XYqkpUhzC8/R/hIiA0mTOw3xQ
Znk6zOQ/2Eem6kMe3uOHxcaHcsoiFYQT19favPBaJfYvwyqtjqve1tEZb9zoeOhgks7CglJw9UVv
tD3HR9v2d+Y/E3E7q49NExHgqGuoX/AX7khdG0RlOksDw+ZNYE1eKEfJykaowrd5Oyo2F3ReXb+X
CHGl6MhpVfKWsb9+rOHUX9t5iQe/zic0Runs/GneRwMX07/m6HYwIX/rBrw4qIEcX9y/oOmBQ1zp
c629JdMGM/hXdI46ajQM95Kb/xJfi2Q5xZRHBEgu+FQlW8bs6vY/FgRivW5k/ZMOnCKJMJHRBY/s
zhMKNd/OPrOVPurlBYc/xeNIztfkP/TClRqsJQZW2wo57cWqNm+JMHoUy4fuDNbDlD84ngpFtAvH
yvVW8UJfuDE20llGfKdUWFl/ukKt7MsT5ot7g9d07suH8avfZPZW63CUrm0him34wubIahAnqDB9
i70YmrObT6VrpG4ejQxAcYuIxIjz7gn1dJBz5MFyBgT1Xl9bxyLCgPoxGg/NvxQx0sjUMewkHjiA
JR3YzxF2czUNprCNWGto4FqUVqk87H8sNz/qjmrSpWUO0JaSvelz7GqfH8JhINk/udrT0x46aR7F
c9rKrybcexwbOZP6UBAjFZt6/gQxd3tmwdjVyFwBOLvA0yEe0397ZE03POuX5jxCm4umTXUwpPly
lEiZfO7E+E1/XgEY7R4jowS1kp2A7yIi/IGXJny8ZFBprQiYsu2zpWSDwcA0+TV/peL+ul9RaHM5
608gSh63zGBjrcr+CyBIhCTAGnIKMR56feQlP1MIH5kmDQ7yzwZ1+St3hVaN/DYvWR/qDy/ZpHCM
QbonKStNSXnnk3whhA8l5vBdmpDsgQyY3DPmEbdYM7Rp4cRMlPcHk7Ewf9xxH/QfDBvRjqSt5bYc
ID4OSrD41anHlf6+bT9c1zrjloX4qlXJQ1VHVoDJB0n9/ocpkekzMO8HIINKAqDnh9Pd67ScESDZ
JTLJ4aBH2sDUBOI4XUszilTXWsKN7MzqLQzYpRfGqK/QfqlNPvBfoTIu2azRmvGPacQEP3/JBgKP
/7SofsxYTYfKv1dYWaA4BQ8dTtiXq0d5XvfiOqkf1SnjYc8cUElpJdUMxuX8XczAcX8TY8SY35eV
Dwn4uoyidZq5KPsdV+Pav4X5NoveRqhpys/b0I5LeYLmKMCYn9dWIcP9zqZL7KC77nsIrTVOMX+1
boNxq8J8FbKNZ39TYxqtIlKuyNSSX4SchVWg0vLXkflpkITEOXGoAES3nremHokWM9Rd6zdo/W0V
N9Sr2QAYFU2gHYN5ldBr9h6/lTo1UrRKg1WuKwyreRXdF52Tshpjgh8dAFHoboDfnVyhPb+IdNHq
qq3IUdKPuCI80DR9KYiHoA7jG9BBQO//LDTxcNKdqgZ5PaputXpZf7sDvdkJZkjaVaWmQNsuHQnq
d0SesI0d57sgBBGSwVha8QIfvXOPaySk9h441mhnx7V36SNjYntq6LChJ1mvJ74m6WJWWkyH9I63
BSw4QJx2UykA7QuvInrsZgIc/OW4x7DPEgvzWpng6bGivJcOoLGB9fwFeQSXpVkHF5ntVi6ZdPWq
1iWpqwlLQ5TPtUJQLL+LDCKYP60v+c4lVz19iBer2gTbhOHkxEgM0ah8/hScSMdLc8MmxvNkkQnX
LkORdr2sl6zgX68DUrAfOUpaS6+ZHezZ0eY+QeJMoYv84Ibf95TBeS2n48KQqZxoEYdbn83gtGYU
UeDhivY2D1afyeuhDWaZEmkPD1uQqMMXd5Yqwh6p9xQpiKycik6KHvCGLmJchFejXItTfsVETJ2K
MzgNxPryH043x1CSBwiWSKPuo+jBY9QT4QB2dMUJQM+JPd8DWJGN2zmVGjJjpFmoXXfZbpIdFnri
VojiUD2j+gx4knG6bu0sSjC5aHQYoa8hsd4ZdKP+/yXfRn2tTyKYqjAk4p53IERq/Ejr5Vc9qNVj
oUtrq6dlX+C2TBTaAx32gigpu9Y1VqS3fFs8AsteWo8JV6Xw5r6zO3PBq0us/mpoNs1+ne1baDC4
/JoXXAEmD6A3e7NJhmlgGG9KtVCX3fQFhHTpwl8inaBzK5aGsaQcDMM+iXq+L5uTdqPhqPP5xmjM
eWjy0ThIHhXLXRAElmeHO6ArnIE0qhZXI3CVLaEFRNqyltX1id5xZQv2knaSnXGIFudwe3p+DKnv
WLLud3KwrKcUw5GEnxUvHQNSgcBEgWiChDjjxqOxnuXPKLt8KrQIX7GJuXrwN/+VXP1paOXShU0D
E5VnUhR1zfb7gH1whnzqCxxStvnCFoSy6X7J8EmT6/bfpQDT18NePS8xsF5BU0CLwUNd6TsGJTRC
wpROZdeKXcDXhZ10hkclDe4dWP3UGwzudXlVV2vCg2cCfbkFEzw0olCPLIYOO4BIL5O/NHwg01mE
8uw6UbRpa75CWfRn1qGxy529qbwAH6ZQokjBo1LWTDmBfEieNbgZxw9ijB2sDP3VVT0pXtQn8HJp
c+lVhqbD6OFE3UojZoTnrGfJnHHRa//znzJtu1XEQO5V1gNwz0UYRX+cThxaUgsfYLq3YJqiF4kn
AL+PC8pMS94/gPtbSoAG5cdg4PBOjdUoXh6dJ8LCmeAwCL1vc8CxqP/Xpnk/zwTkK/AqYUSRbNtd
E0poIOn8YL83MlZHVcQ/dYEVAYNak6DV/wzVMoROKO1e/loW+5lqgZhUoCBECIgPbQmrtGy2mAhP
iyWFtsodFJlOksIksaQWbbH23CCsik4cwFlu4M7yU5VoN6YRgTqBbrvYaNExf0FBan40NbaT4PLh
iTsHy/UagVX6juh2oz9aAgm4UnwoX8ctFh+XRmiUXDF1WYbQ1+29ptKE4dvA/8TM9mC4d1Y1yq3M
pKNY+g1qV9qh2bwLn9if2kDmQyLOu/jbs6XbX3R50YPKIc9slRHPVD1bGDvBjr+pbDkUMs7CgNu/
M5St/7G7NSY6n1BhnxSDcdeSiNjX9aDq0Maf8f6x/8pg+zqngIQN55RPOCMJjeV8UpwAm0l/+KuN
cOLBGhObWio/yV+CoSMiypHhqLeWD2ZVzciHWGauFDcHbLtKSIbfbr1COG2UPYFgkEwHOYPS8PC+
2OVecmMfMwnUeIPHEodlzLxcvGJ+x+qnvH2IDxZ6SpU9PEh8YsNM4FzWN9sDCqka5oHHBCC5Brbq
5w32voOcnYOnCK1ciCd8DtuJU9I8Fc1eIyywsw/4LuTl1HpjNk2/rfa/j/CF574PqmNeiI4HKJ9E
7Dra9GzbtBcztZpKqFywd4L1Ji3WOK0rK50IykSYxYfMvL6M6CgPSDqBayxrmiV1/fzSgoF3fAVV
p9hOp73DRq7lAZ5HuIWdAyehme3C1KkPo3fRpPlcV+GsiUOJQY9TMo1GwvttJzhkQBv3nIgYIHM0
dWkZvt+OvHeCUr1ipXXECzVlkPJ2aMcMOI6/DBHaGeOAOSor4MdEnkbKdjd04vomnfgELaHm667V
ef4Tf8byi9Hl7Z/Sp3CGDmndgk4+H0yMB0RGAngVgai54fg7KS48gM3CLGVHam9PDnDYLKAK9Nwl
whdw1ZRwIHHr0JQFmixsfwhbzNktzfYbc411F3L2Tjcz8Ey+XmM8Jc8YTzMpXgRiMHRt7y5c81Go
EjSzcZh/I7HYlOuk0CwjusJK/mAK1blPTuYt6DGkfjIZhJL5jzjrkizOtnMWZmqGokA7seTgGCI1
ZvIhHHlULY1AuRkxKR7nF6cKz/AT+0KfPMvWVz4OHjvd4fgMnRWGYILVZOHmMIfdvMSSQvcaRVhA
rnlGIuWGni9/I/Aki0/GYm6J2zkgoSrmr0/QuBd2L5TJDUSeJenvJOUPnfKtLcjJgx3sfq0ISLEb
3kktIBxdbRgbwyirwdTtLFzYcNr7bRH7R8XyLsxEDHm3L4S4kpwAZEt7XfOqAMTETc83oPmFGi/1
p9LGz8VoIspN6AcfMRGmArWTWNkKJA51y4D5yAyNZVbjEhsLFlpLJKC1KwEHNRDJ6FTusTdcfPAu
0YsxFS7tLkiJfsK4/23YDo6vufk22vZQvSyA+t8GkEMLn7fD5cxD+xIKod1ylWq6sozVuSJ0aKFr
X/oaT3imLjvYVwVnK4ERRVU80tWzqDwNoWuosP6EsH30gL/NlKzOQe6MN8X+KgWX307s/5io9f/v
l8WoSdHCnduBobPm7dQv37BrlM1jBAAw7R87NPBX6fXyWOpIyOjJ86FCq86uqzFD/8c0rUAUoEOF
9W8a7mFyAdSbMCUqqUgU64/QU4z/U7idfyVKxEnKyP+gbHlIedqlOkUXpJMSv8OihWupnTNIxxhM
4dOg6YWVLS9wt7pM8kNN/SHVRwRHoHjU9V12NgIXG/KkGZjinnrWTfyln+Lx/0VSsiHy6Q/LP27b
iZb5d9uAF1PBpfo561a0M6crcmRHYMMVQu53HSN8n+oUI32WH44eJPoJoM5UVa1yPhdS8tjcHXcB
Ab+8Z08RUzooJuqgUukCBYTRwrOHk7s6c4wFRjOqkhkfg1NeiyGWs4lKnSb0Vi0aFrch7THyudUB
qAZAMpJJAQnWHO2PhmA2pbFAnJ4pgwMLkhVyTL+eyGjH9dDF0iir7s9bOUjDpr5Wfx8vKOBANYdG
j2L+QBwgETuEGTooxW3foNJz1aS8q7vo5bZD8wXj5QQq1+uBMQZMvVxWumRv3TD4GIHv0UXh3V/C
49N9v2MMQENEmfMIW0vUO2DPeUPot8SD8SEUpYGNTqfLAi83ZXu0EOPik9BBIgymqxO+TE5HF2PN
mxUxxu6Rvar8o3mdJjgG/3lpk9tdgOsR2EyK75igJiHfh/teDK++2YOW/rJmQiLgXVeVUTFx+7CS
kBr1dHE4H6F4rkg/7VfVj09gpeTkHRlBufzjYTkKIh0WamAV8iovwrgfxfSk8tUjvAldrHDj5C+y
UjgrCjOpG1qhTX46VSPWm/OjyemCHalk3PmRPMgbPp0jTUkIiIsho09dcYGB4DvJ+etntRQVpZU0
9/DOVqptk1lMwxuae7KRSRCc0eomFh5ENC8J2t5UJHMJWFV9cli94Eb0KxUcM/HuJb4WW4Al061H
fabMaW54RZkkZ5bdJXFirqML1l78s7Ovgc73MH7ILVAUa4HcLYTSqe+q+C8zcMnWPHHfHDGOZMPn
6unu3m/GU9b1vTiArZSKROaRo3HoEAKnNVwwVOHJRzP9gJ9xtlIystBaj4Pde2wUNGYpqCfRV95U
coeMIQ19b+4ZmDrnFqFnAKO853YL1tSENv/1anqlhakxfbDNFTmChkWkEyynW0z3nJhS3vqBYAgD
nfgHCkLQqQDfhm95hh4Wv/dhP1vslYRiF6X9E0HBmOgQSqlxZlWp8mLVq9zFaT0D566VQXyP0V9d
SGvc88VwAzhU3qU476lkYepRNheMDrdRnZdb6wN8FqTHsX+wJapwd/Sl1WTajhAN+EHUVao+OR7F
lk1+Gf1GI/Z8JEanxQbyvYH0D4QzWDWMT7j3BueTjVNICpihDu8qjv66+NQV9nSn9amIftt94yoo
Ujbgle/gMHCZDvYDm7n28USK4Dwp5J/FzNrAP4bS+Jemn93131lhc6WWNXuX3TAACDoAHf65X4ht
xGeVwPAIgj0H9SaLbmVcWaUWPYwzdW/xTPxtP4oXW62FP5O9zkJPb2+5NBUNi3lXoRirKYyrt91i
CzEAcCICc+klt2te121JiyP9gEJK4lKXUFyBsydD7H7wRpsXYSZfEZSSXhyD+Dq/aK+HxdP4u+4X
wpEezsH8zN3hNijfSK+em/g09T5WVN3u3BfNeQDd+3CiQnVQff05Vq7otTT6in3eC+HFgiuQmxB+
zs8arp5/Xc7gFLLoyrcdYXVD8Z5fqTgFPiXCc11e/ByMNMJvBTmPSzPwLMgWhZq3H6iTQdt/hrVo
0791CKwf2DmQ5IN604KHdYqlD2o0ieXp92ga2eozIPii4TrNCMGWGqEvCia36jjk6tGwlyVLLcLK
cUX1XPLbCjuMFxwS/39vID02VmW1tVfP6Rpw1TZZ7+v39AKCYI4ROz7QN8bbCQhMvxBx9boZG00D
TLrN+i65mm0pa4z1kd33kRRG23WJNwY4d4qDygR3W2HmvFu4WpYzAEGJ+hYoQbGz7wBr4arjDUBh
k1L9Cu71GWbAauagA5S0JF7bmUHzocJx+xdGh/VcfkjvPvQULLrOwgObKmd5dF7MS3rtfan9IWvF
WqRD7FZQM856nS/lW+xua0/KieeIxcN7ZK84b278bxIcrK1TGDVVSyv6RCU07ZqUFEwbHVPedPM7
xb94qeqE6bIIe6fXpLTYJdz2IlZyEanTXispOJTghc478QhhaSmMnh8wWwoOYRHfOxB0BtKQtaz3
k7CL/inrgM775eR1zHaCxgZJH5l0Yz61E0gltDthFYcsaUvRFdi9gC9feSlHx7saT4nqkWul2DOb
AApfPSpw+cb1PWr5DRk6ffPqCt+KCuo4cHjgCburQfos3XpNju5qAGrtSkiY/1bxXxCfUTLFpybH
yQ9FXuw7+k2bvNOMHyKZYmHLSQyTv3DWEZ936NikOR2dZY01N6TMeMcQbWjL1T2dOSPHIPXMpNiU
NNuGlKukzZIjEJDaEq9Wmx2TDD25vzWQ/Mk+hxuXBSawYjNgC0um9nMIaqwYo1y6q9eTQWhK1Izo
PXL4WTGI4RyH23OZQbPPKCJqtuI9eMA6q/lj6uu/hw044Chc2OCNEMmpp/mvZqzIxvTFR0F/hW+7
5QcWuIP7GF/FK2jN0m3H45ToK1vnffKx8ueHQ0lBiNXvBp8O1+2KELIEV+/jLNQMvx+AqcvQrkbJ
0gKqt9FXJcaYCqk/D/pKsSyCCfR3haN2sARR8zV6UbiU6ekI9fV2011bR0ptIXwvoC/0/D7P4Lp2
p8k9R8FNTg0HVv/i0u+cGvIX1QXgfqQdx1H7yTYRoRFTiqpbZn3b2LzcR8H3N3kX4fCGx+8a6S9u
3g6oaRCMJLeFzmueEoiu03n0ub5v7Pc65X+iDOzRppzO7ycgxbZiPzD2BdVd78FmrFatFuZgrB9B
EZdfAzbP2yzafJgmpTHognFyTh25Y2KMFroUG+L5uHvgdYUkQ1UjPg4ba3ehW36KU/ZJfwff0qVK
juBXuc8SyjoUwMLAAFyh1e1c6OnsYCnqMHBUwn+KopqExkhJzBQOWa3rBsuNIrO3u/RPTAJ77QBh
XKJbF+alMwwwUO+O+6U4AlzTAvZ8ejY6vPDP9KB60nmpLlkZQFctxHigzqB6D4q+aur6dXEzlwmw
b2tiq6hzfPd0xGUKZ5b5vbhiIyvtzmGLwWjiCpCbtvBl8VzkDWGnDP3QKgK3e4+ZjdKn2BR5bW7k
Li16rrN/BG7PMhwdLeqCFbdPTQ7+Qotp6yeTQSSAGGoo4Ns9Fa0VoCnZA4pKjAhXDhg6IAyyHxUl
P59Uz+jUV2ee8IkgJVT1KjMwY18aajej7LLHm91Q80UuduUJBgzisQpSkPWAKAeMptkrU/mmEZ/m
OgZS83Arx0Icwiv3NJCqy0fd7725t5b0sSWO9DCY8g0e7pDAcx+eXrLjjiomMlbibj1JveaCz64E
mUO3ocyZitbqYF/CW8Xzp6vTfYqI+4uEFw0u+c/z0dd9/ENs1M0vvtrjWWNcX3kz8v3BYZKepG7S
LQX99UY++Oa23SOo2xWWUtaYakmonGfR32lvVzjpVmPekaEckE6Ih0XAyF9NkRD/A7RIlLhjlzbQ
sYBJ4/dlSdO6rH/GNjsj+H4AOxJvBLLcaaQbILj3YqKe9CR9YQo2HN8hcaMNkUAwddWhXzy/ypxu
naWyq6/bThr91Rb+gFd9IRoqL8uF5M83nwADzPQwcwrt0TRwqzkh72fNvcd1IcKXJy+YYBZbTrhp
hNDNAGVIS6fHFJYuXSyXbGwiZKotSutox9TEKIp++OLKVWZOEPQRbbeYSE4V91ZNC0HunLMzll4C
Zer+hjvdzPB73YshJ2hRJQruWfttD+M5etgA9UJcOlpNX3fGM0FklY7Z/vm5jPs562A/p+3N45ns
2ghloBLYKa3mmRDya96rRVBMx//VQ6In6nyWFT2YuA1VbEmOcY+gYrMyboEdOjc37GdznRFxHwCc
akTQr07cIi1c1EXIrDTolHoEQfTDJJPpAaFPvUDLMsF6B59qiii25pfSkQY+cL4A1a88+UNGe3t8
rK0adgwatRcp5qVeih48CrPFg0wRpcjsku+F0kJEHqtAL9Jd3AsjST0p9a6fGSvhmYq8jwrgSdjR
t3abHjSZuuUi3PdK+DmlxQSNUBm7MznBQE57iK31Xt6OK/wtKo6WoA5og+oxCg7r1rIjew994H1S
9IM9eTcHHdloLopruIq92W0lBGVxPxF47Kld6rMV9yxmlbK0pqaobLNwWsIuKHAQCcmqjIJQ7kJC
NonKaiT3qKOvilgew+WhleflyXNsH4OfEtaE/z2kIrKbN1J7qRcx/rKn/Qta20k7PdcuPAHnC5eV
Eer8EkPM+Q8pMeo3+c9nPypIoJAQaSo0jvkDIaxkAoTzeNT8Ho8cpl3RY5u/ZQY03wjOhjH842kv
EJmoGOH16uzZEQ05ZKVX1rtm9jqmjjVuLwRu+U02Dc7XXgNuu3vnUBhNt05pwUpQKtKOtbtWHXw+
oYN5mK3voASNHKC/PcR8X3raAeGdxAgQp5d0P2Ert2wyaWmKsAzCQjMajFbYrKKd/CoqG2/YgNtw
RyqQIX/dKkm54ohXwvaaYqb0HE+9jCsfrvM03vq5duMpdKsngTeLflNL3PIu2y1tU7bYBgB1Z6lu
ucfWcwovKwj7vY+8PXDb/vusDlzcfOMIb6IMb2jFSnGRfXORraNRgJUV+QIjrs9J5BVWLC7whdp9
KlUV/C3Q60DVjbcY+F0sOHPhzpH1sFr7V+hETp270PT/tQaDbR3SUVYLWXN8aVo6BNDZfihO9+1C
QzyVJds5Ei+BkGQBWSKV21fDAS/u59eN0EvmFh+0BFy4LX+wmynXntBn8md/mTXM3HhyuyXu194d
lb0PQiZAgofwZnpDjmFUt7WLBvOtzCoiPhSJ7EPWALg2FZ8o7pb74XhwRvIamS6yEVximRAIaz97
QYOGqZV0I7tAuS8oTZ8SOqpbtB8Kh73YQiEjTBINSSZGHasVKJge+NthQJTTAFURnkf1+aowta0Q
cG5jH1UVHdPx1EH8D5mi84N3og1nKQc/t1dgs0XhFfU/2jjUMthV7JMJBG4C9hOxByyH657S99Pr
nKaOFUrkg01XQh1Mb7L8xW5+A/CQ28+cvVfLZ1Pk2JS7o3xcmgb7izs1ozB2ZA6hkngB4GTgZYj1
G9eSkSReaDgbHa9ESPFB/LB972NMx4V5SB/J+lFdSznORj2E5kU0me70giXIWjiRtw5+wQ92GytQ
HS1hEbnua/N41STiAtFdVthIkFjgiv6u36UzYmA/2Lrnr87XF9H4ObTebJ+qrDVtu9pQiJEaZOnK
YrFWOa4wpFH9PlgxSRyvKOt4JXdDxtbM/0u9N85EDnubQC9TlKou9ZXkgyxVTWSC3K6lVq1KboXH
pVApVy2v2pv7zCK3Cnpa344KWOst7jnU7s98NfHHsW8ttMIsY3AO4c/eZwL6/uzYhr3Zkd80Epht
tRgdptVEBqSuFg3Tvekfr4xbL2Ev4cMp9acT08bc/SX/dOVe8aiAa2UDxmO2A4/+oyVmuVB1pIT6
Y/ag6AW4tcnmeiIuW3wv653M0l+QCi87t/ot7N/xzBXnpyNAau8+1A6VHnvVj9QVbrPN8WjtYt1J
cSg3eyrF1UNOXcv2radscLxu59aleSS1sEld3InS2VW3ejIKsbM9sFcjIaSvPX9Gef45LueETKce
WppC/VDa5tUqLhj2hVL6vhK9Je6I0A57JA2TPAed819ZoYl5Zoy3vFt0nyWDoVTiwwdk0HXfxhk3
JomWDaD+KxgEZEoD1ANtEiinzgee4tExGkhwgAkcCU4gvd893Hs7E+yiytOa1Axdexl289ewD3zn
V1Q1eNcdVN3H2Isd+yp/HxrBCBO+xekofbIQCqFZX+RH2XIJEVvdaW+FYtOyqM/FJmXzZvwDXuT0
2PWhfEXeg1cLsVHwUJtoMqVQmxZRU94jAykv8/rjmFOLAMvkizP2tH8qp8OnNfoOdtIvHu7Q+gy+
/gMEWTjQvW/dw4OIHQr1LqH5VFXiBL1srWtmMdNjQZec1pFxwozsspDx5k1eFjHU9LccZwjmwQCd
dxD1vxY6yse9ZJ9N4J8Wyfc7uFprUm6Ne2UP7qf5rdAwzq025epbehYck3luIat6Z2r51Q8CguO0
uUwsPpzGPYleJWy3dYjUlmecP8b8CZ5aCh4EO96xRmYMO4/yPwjsPozIKcquYfoEn5hLEsUIqkJy
y6gs3VhvPxjIyVrXZH+Krmvsh5clPJ37eveHvXZOsC5LQ8cUoDHeqzhX/2gHZ7lAuOvCEY51GNqk
feAoWzzCiPH4M79SBBA0X0QpKHVMNP9nX4EiZt4f0mvF0J48Z1lbY9IoSKt5a6MrrWLSrY8glOXD
v0zrf02qQYriN/sA25LyMNSSLpCKJy382ejDGxSaabr8NE9QOm0orzBfEgb5zB2AGfBTw5nvVLPR
gelhnInuoFDXwd8e9nUL3KSpYsnjYLLFW+QoZPAJqr6urQ2EbsAZWRqqZgy0z+cu52WqxjNCT05j
Kxah82zWBXWpjoXexcUsIO30oUMm4KX9BmONa9OYlbhB6GPA1qCzJvmCGWY+WNjeOmckowHKV38A
zDrFBCBjIdmi1tkOudjJ70Iiw9B6ocsYVVOI+aaP+RiBxbm7Nlbj4QyE+KZUBVyF2s7eurnkGtg8
6j0ePHivz1qjhymyz1ZeQ3e0ZuK1PfNphSOF+j3KP2Zh57tgHRlwO3wLsXrlUBA6BriJU7PDL2W3
wU8dGc8pbwjBKT8WpUC430VT4XdLpmfR9MzB894I8p/fZLMJoeK0Qlj9GhROAoJPDA41VP6yevBm
rNBoLISyXJ+xLEqiqNz1aZuqGdQFgasE0pfO67mp0EsuurJmtFUIyMaAaYcOTWffL1O/spx7mMkG
zancgOD3pLoHAlZjrUrtqudyoMERNRtcjVp51o9/wwzQteZMKI95DqhuWHRHhFBs3cbQXSJ1sE3j
unNItMHgu1qIFOWjwa2UVAv22mZqH3pYpgklXRbLk9bi0NOU6TQupbi08ePr6jKggxtspq4BaKnx
GvIOsNBW4AeKzEA2eL9cqLHOhrW/RcgJdTApR5vILGqGoGrVyPfjCj/g3wplhoO9SHvlo4VjM0WH
Uz2hbupEsZU0xUrGRyN6VykAfyR+jNqPuhsftgeioMzkquHMybUYIwbzH4qpjgoE7aR6/JbUt+LQ
GNwUubXy9j8/VInutass4K5FhC0JqKvMGXhBasHtO3sojXf4LfY7Z3SyTAN85Vr442Y2STSzXkaR
yH2qSn64Sv9D4wb+RX953TvkkrEcVio+EpZiIRV7zWJSWFUjbQlBGyPgFrQblW96uKZ6QkoDoUHK
gxSMqk1rkNxmBPWZNqu62RbC/fK4bnCTgU7Og46I5EAcpywBFfBQBFacphe9hlRoIMi11+49rktn
yoCZVYNQT8Iun6D394OocuHtnHpFEonFPQA/fhNf7CvRaFRWRsDNgwzJkvdHGe/pSdFVn5r8+c4t
FbaX/QvZvsxRC4jSeWZ8LHOTTmo2GtESegd2gRwtJ1xxUmgrool14lvCfiALjn2uyOyr0ntow+CJ
s5X/kqoH4/J0Sj7o+/yCJjfJkTIWhH8xGChxCB9hCKYo7++o5ANisJG8qWhpDn+LGGJe+cWmEws6
kBIROaAqtAFvCn77FQAER8U8idsRWO6to4UqXgYu8V9Roo383T9V4aqAAMWvq1abpoAKC2w/je5y
YvyKTUa9rzZotZgbrOQ26OoeICyBxWeYU5hd+sRzU8L70ZhREQ1zXl0veMKeZ06Dtk4smWYHokf5
02waR7rN0ThKDyxNf8YE0P4jNKqMFahvuk3IjO6CRk4oKBohzGJdfT0j/3zEZQ1KTsCMlKQ49Ji/
5efq64cgZ7eV4SarmW9d87eLIlKSS8Qm/evyTDFss2MKoRHtepY+rgnWMDFYuPOjaEWZfzC2poOn
tiVepF/KWwGmqQLN+ornyQoztw2zd+OTr5I+AR4qGzxhqWW4es5G3P40BXaQi+MFw3hDmjNIuCVK
t0wkSmai91WiLOlQPu0L+jBi5JvbcOE6VxbeXslsENVuICZmtAdFwR4LoJHy04yrmNz6xByjYv9H
aWe5faxtIEb7qKM/yboEVF4rUScQKR3uFEglgygcnBMiu1w4yOp3eFWyWKBMAE0xw6Hn92rrZAuC
EQ7GdlCPTR1Eit8rl1kGdSJ+P2B0PXpi9ItF9Z3pJ4IBz7qBMlFxk8P/GL/n6+bXDKtGpCXmSHqW
3GpaFGGpu3QXZ0B0bVrKvjh3Vi/Lf24ftq0pFAQXi/gZY5w8loLFEr9bUIFy92Zb/haMXbdDx7ay
1bzrsrRulrry4qjR7GZrkzsXVcT/i17Cbfu9/6HLi2KeAQR4YlaXHvUlTXJoTpWqiM9pry2ZXRgZ
A9rnjtPn8ylrhXIVYYC7prOJBWJhpHUX6USNdpP56ULT3iPcYR0f/wHLY9tPiIZdR49jXM3pf0n9
ZdVLADnKWR1H5qvvarKKojlGffGqfSrSKpxcDDvCwSYidJ0Pg5zgh6FeTbGRQUalrt+/arVHLE+U
FJvQqDYAQJQALo6q25xPmrzzmt2+mm7pTbbyybnfQYzXhreeVWojtXi4FaWhhQNFbWKEt66DWLO8
7t14pCMkLchW9UIBudyrcBRAFaOL59d8uEk4c+CxdbbDHXr94TDcooEyBOn0SGvSkQUImpBadXKP
O8QA7hooSAINyt/trDFD/tGLAJ4zuKP+0jJMZjaGCSOMSdti3qH5UTdTP252qC9CLzScuhMJ6PAu
YyAk2GPUtUG7rndRxv8Cw+WdaLNL45qUxoD0wSSXzOCDa1WMp7dZ9yd9U/ip08UXNwRfUjr4KcK3
o29M8uQxPjdfhbPeHZsYi3CLB2WZLypyfoRxYLcjYgRCehIRQJZ/29yZ5fKYJZATzTUk83Dv2IQP
UsmKTHqmwApu5oV+KjpgpnzEXNRjJ4VoH8VENBSPFfViyhV1h8lsqw0RWnuauFf0eL8Md+dbvw6h
Y7SHv9xvQBNNn0Yad2UhLYKVnQjUFxsML0FBRHVHU64ig0cDpzVieQ2bKaENrMULDy5CMHuNXex0
oJ4GBxlBE8Lx4+Wm0XoJhQriquqLRgqcebteQplTOpSJshcO45FQML9G9ngDkRvgUtdATi7Dr/Ic
NI0vu5+DjsAiLNYNWOY3BIJUYHcscFU5vK/jbFe3B4Vq0tlmkkHBwkj7qW7e9Pj2E4IDZrrFxp7U
9wkxxNkFKNVEXeFEQytnAUSGW8UA+VZ98s3TsG498NkK1Pnl4vpeJTwQi4/8RgMZBsRpcyjv1ts3
R8hAy8oBHvz/B3L0NJcOtfN0VME1LGXz5JtTHqqGHLsJvoYwxEudvfk/ZxAViFUaeLHj9/8OmIc0
x3qTMoNj3y67lhDJnUDDQZdP1/P6E0dK++RdTY0/QtKOsG0/HsnBa+Z8XVnJhEfRKlbwnYQAaf5s
Bk/H1+ye/5gT1rFZt3EtEtnDfQGsggHFAJfMPOVkxi43g8zRKO+Aa2a1/MVxMgmbirPi8Fo7HNcJ
JM9pdSsr/t8HglmT1aJh4GKsa5AVTLw/cJy6LPvkr43W6YaL5KYQNNLp5e3d9jG2YcTPbwivZ2YS
4C82YuOHA5GNZXYejp3RQ6g9B3/mDQ5mR5j8slUqoR1ZRQ4HIG2aWeJjn5K22yBUGi2DEkCzY1RY
3dADRhBFP720eKSiP/xMjcObOV+AA9q/rHqhPXULJvbQVnCmwOhIILpShT5wXNh6IDeKcTqOgD5n
PURcYao0G2A9zK0H8H7jEYaiRfP1HSg4ZDh4lY9eOt6Q9OdEbpewPz8k6YMHT/6ktgJEQtJPOrGL
hVMbErjT1puhrWO6Q+v5uz0xzrHwTKbF86JQetUtyIH5p3QZpibhT5TZA0t9VsbNYAFQoTPxZ73p
h/CL7d4000xbE+6hFj0Bzw2FquY9pgT8RbTYEkeoV04bV9oChSaAzwngeBDdwrGI1NDWllQh4VN9
lscwz6mY4wu56/8x7ceXEdPG7cB2kUQ3vCigO5ClLGw5AWahq6yVseRRJqPlvauhZPCzdzQrU3NV
ATed5cIkzFozpFQzo+6+ENwy4otW5PGcQXr7YuPggkCJKEcWjH1tOMYPTEMTwJOuBTRbwHRxhn7X
ek8Aid5eatGRAMpO7E3IuE/iufjVXreC/JgO9J6WPqtPVyy3fcrMqH66aDZ9G92Td/bx/KwP6mXE
DqfO3JsXqR7fzG/0CJoSJ00edvrCNfULF1k2qjYOOwTiO3KdIpo7vH6h/9HNFNGQnGc18Y6630A0
ymj02+XAMbai/s2gSsyDJw5ekgMAw6OKtfAJAK180OWWU+ZJM6zvJZ2fOpuLbcQzuZoWvhroTlT0
jyZdCPlLfOpwHYXeQe4POIk+S9pOUU8ae8X96x37+JV9ENZBIp6FVGlapVGdE/Ii24NfbxLJkS6j
D2AIwoYFyE63J10l/vHdZQ8jFZYjb4F0G+3bOKYSG0Pdupgwo5K5EIXbdTT1O05jQn0/h/zAK+mH
zcy3XUeMwfyHTiCrdl6H+HA5SAAt7l7GKY7ipBhFzhhr6SU2rSQn9xaTIX9AD/cndiYdq8FJJlng
B4QZOqQQOpSo8gBZIyhgaEaRNlHQS7O//4J57Fu2usc/qWogsL5Ta9i/NrE5voZgamsa595jGps4
68k9lwFp2BEnutxx1Yc0s3F6R7lDoBNbe5TD0S4w/dlOdjJfvIHqr5/KHItfNTmcGvKPaJi/yfUb
6JhCl8tBEXLNw6rIy2DE4g891R0vITG3M8F1Ft+/rp2Hd2oQdpeSd3QTn7g350+5edAxyRmavDv5
byPHPWdUqycrz1O/9nbKu2fjSmGNv7Kk6FYTXZQ0ZkZmvgIdG0ZPXY67tr5ki0TjTWu47d20uUKj
2R5pbHx5wr9hF0HV7+eXFI9tZFmF1kXt2DNgKG5lmSJxYPLlFPAouMsazRkrFJEXGhYwiHcOUwH4
S12xfncYo2b7o8iqwdp+vGKFhC3gb2z7XHtqEnsGwiYwzkbPybAUvnJAJJ2luln/+RZ06XLe9krB
K3SxWn9frSz+a/CUa2etsqJDSTrR3ekG+luk14nTBywUPGaztSACRHPITImKPOhQaPs7ytcSzPKk
HdSCz4A3j7RyrWly406FdONJ397tNDaoS8VPagygIodNEjaoAz32rW81ZUPvY2nVtimkNdkVKp1+
N0RkCM8o3K0G6M/4hnTWYXLNspw9fzLOKP6jwsaVcCcBVG4IAfiJIkKGG5wDnHiaiIbotLvAF0qD
1YFVhtsv/xgEmWUSPp//nxH5kOcJxMgBk7ClZS+qSDUPCgh2FiGqF6XsCYqgWRXNF47GQFgxcs+G
9Q2vevVx+0GWDQs/Khs5XYdDNyQEChmTpC3uQh3YaviEvxLu2WIV3TOtAMEWRWiI4RYv/jsj26Wv
sbMVIcjFxKVu5A7gLDg5JRciD26wxUaAeqcv9rmHrGc9Xzk7Q8EEnM+ZeGXKYRRkJ1jSJ6QFdqpw
UBIFyAjDzjszL+AJ9l50x0QpddlOke6wydDNDINh/sOmRPGnupeuHGnT/h85FdbD6dDEaCVvHg54
6/LE9Hv++Vv+AbPIoatcFvmcuVJkV4QRr6b1JCrcr4yMKG28wLzF2eKcee81tUSIRQ9QPAoastM8
wLYDlSsz7NabTk57gJy8n99ZsBVlrhIYr9rOvOWYqzZQ9Uo0JOgUQD13IvTtxZH5pmbx1e5QIdqf
3F7YzoWTNAl7a4gkJ5bTcs+F5fWOicI8d92m4uBf1fWecEVW8HsxXxgXgyvbTfkTJZG1G/ENDvQ3
aASNQPdEPUJbqBHqsu2JURosu/7i36Vtz7sbRxWPdY7iVtRfjehYeclrQvpzbkTSSEtlEJ8VRV1n
SHbR9hRJM+zklFd661oq0YQ8SEIVYQvhT+Ij/DLLwNy1z1ksfN92uH1d7oijqMuxDBGiEqD/dfhX
P2xaW14nyHK7Uk4s/CQvMRQJm3jg7wITiHwxSoB6n9rdDflitFVfEtKVDIaYDbv/LAzkWImWhpOJ
oCLBF8CrvRtXk/hhLuIJ3dXmeH2ZmYYJ2IuuF92YOHGBDQkm65mYAyPjgwHB5Mqw7ks62O6wWIqL
4SQTuS/f0Rrkuxst6OQIKMQUaTRMGnebrqM6yVCS1A6fPMC/vx1KoSmkpF9K8dltZKKYC61svGWv
inFaVb0nbdi8YerWu9Xw/yuyCgEf3Uj4kI+7AtF2gi/2hXv1OazYHwXhA9YzAcK+WvuA57MitwR7
bwew11BYJzZ6fQUD6nRhIMWv9gc3p6ix6nJ1ITrkD8FyIe0ARfOJXY7t2N6ZXefxj4Joue74ww9y
a5shcuoUMPKgvAouWydi07xnbFyJqgUKcltLUWvuc6Waqmu0R4eeWp+kG9aWlxd67ErFHC6o2pld
uncN21/41XNEXEhMfZibq+vl4eIcUH6eGmHTf0NhYhKusS6PtZr4YSQsr1B7SQXummWSITWl8CcG
Sq7Qs4qWyLtSNdVZHziKiti2Kdv/EkymrtRuxVuGsg04f4Ns8soexvIc54JfU1KCVszlZ465y6J2
2+ANo98X3EBzL/so9KkL1hKUVRtSBJ2eTsqN67UZ++4wV5Jjgb8WwLuG6fmXvD0qMFwGFkbMMf3C
UyTuJmcI0sl9YNcQAw5SljvoiFZu8i3tcs3mZcZqLxGyydzQxxhWucedphYbAyG/cmgZ8u6yMJES
05NcsJZ2coUKg416gIhJVKGTYlRLFBggsJb4eNaNJCHfDK3bLpDKrJUGNl/zVBSD5hUwVOpMySqS
u8e1LrJWziRX/f8+iCidCuU/PDbsLtG4V4KT4skGO6eUX+yHmjJCxh1NdN1YHR7tLmc9c0xkBgJd
xejCBWY90gEgtL0BG5E2hemqRidSD9nwq4h8+h7fQXvoootQdra/YxaaULHda9bYN67vtlCb67+N
18zZMbFMUO334mVWYoJ2HaefbTwryQL/PYQupfSvbIyDc26h4YVzD2cowrSIuhT0q70pbB/RCBRY
k9VRUuG49KI9haclsPQrazBTfdbA7aS5Y56qkeNE8s8ei5J6m/pE2SQJK/EjTMgsjyYhc6p435VW
YVEom8+qIRIlwFeH9X+nHQxgeume3eMuS7txqD+xDcVQvVP8OnA/RsjmU+ROy/U5k1fusOjJZ6Ej
AiJKEcHJIhFDQ3dBpxdsLEfLXuti8Ih+y3iBtq5eaEkJZgJgN8E9IkIpkGlJw8grB6RA5e8AvORG
Ns4q1hwc2uDdhGAdkR0OIFBGx23pqnKYs0Ib5l1Htscyd0ZPJTqQ9Gq7QE8pjTColwVVZgVkGq4C
TObYOOxh9dfT2mKr+MPgRzK4KA3W7QO9AJ3v07UEjtcaljSQNznKBMryCgM3y0KNRTc3WyzMRn3i
B7XjbFgaDELWUtbhDtKMp9m5WX/BQxhvv76UVyH2jQulGZoNaLB88O95Es9oZ7MHL1/2JbLeN5zn
DoAYLi7q4OONdhe9NE/UzuG6odKSPQS9dt25LxV2ym5LhSiLqEb4Tyrq0iMPRw1oT/ibozx7TKT/
J6SMhmbwntjzAVtu7ICOvvBf92iZmvSyHRuKRnoehkNRRaSryAzYfLO2WrjqUHPB9tEC2soCHTGh
WOcFIbArQHsa9YJRsarMK9dZUAWFi63r51fcbf8G80aIKu5GP0DAdNc142uCK1OePHmTLSrKng3x
dW893JOd1UqInuHFI1XoZsdIDgq6k19pJiWgkN5idWehUbCrfNaN3bDmIHc8lm0lfWvTpin6AqnM
K69JWNlczVndYL22Jh4J8btjrsR7bsU4Ta8lhO9Qv7b2/KIt2+ZHyU3+tqK252ciN0Z0BO812ry4
bThYPJHlpF3ZuV/MRqxkMvocbrcrs5Ob4/6zcr+FEOqPVRLGFmzzB8C+9gJWCmdC5SN10LnIgUxL
uCpz2iRT5nYcQypGakUFOa9wavrtvcCSnuSFR63s9FaiauPmbyUXyApiXHIxGW2Ilji+7yqDJ+Tt
hTDc53PJAtl9It2w7jSXSlh7hTv0bOvidOk5ySceoUTF8KjRyeYMpytkPdFAg+h4++lnt4HSGZK+
fdQ+syNuFVnqLKh3iRCUfsSOIE7VaBPXvbjaa2ATJF4OuET28u4nx+EM5YGU7Ng1VtCoqC5PrcZx
Oi5zpD4xY4kf/lgZWCVcGv8QE+Yr/KeEz8YijK509vQ9fCJNDsn+ZrF60n5H3xygZNe5ExCcxr7u
TalRNnT+DP/z2//upJiZ6xgyGoZcvzjqKbgeQCeToSWeDOWgoDTk0EhMhh63SbylY12nEBDF00Ym
SCiotOlpuUjRdfAQ1g3UjXzzBvNtPb3cJiW3CN5zOdyL0LVjVCQgB3JBYzzxgY9uj2k0aq6nWok0
QjRLfG1k4cksIOFyQAVl0afO+B+dNZkQ2ood+pZvdAKK8fMSIRF9VfRmnv8sFE89aEiNYawPJTlq
dqR0eze2xzc3cGjRyE3q8/5NwQuzqQSJwB8ZWGjSYHQgcNNTu+8kr1EUm9d5KHzGirB67nhul4PS
RhvVQ6V8ixFtvGTfbCzDYuABmuo6DLBaiN92pU4MfXvCUxlPL/V52Aiq6xIHbEX4n58Dw+6iQEe/
gwmij3po8M2+M2J5iHe9BZuiQhl2crxokICmtF9vE04BgFJBM/nnFhrZXMcwrcGyHWlZYy3grt2/
+klCyRcOslpEM+3kNog6t+Cpp2hriELyZr4CpoZCGMvrBkuKX8RBIiNm4a7O6x2quUX3oG9IvuPz
+MyREQ7ccAw0AEiSh2F79I21OxcbWEHFh9a9jrewrFovG+5SY9v6L0xbqTjGtmn9sBiuhKZ6PD62
QFgTROGKt2I0fo47Hizqd2sW4C5g2aQSc8Hro3lnu5V5FPns3nNZT1sqo6ByyLpYG4OL1tuyWRpU
qT4a13Ofj8DxO4GEh8B2teaLKGDe3fFqgWiPyRhVBwmHMORe0UF84TV2Ohb/YvQxA8E8WNYaatJN
H+E2o0+uX2v2D9XEHBCbViyWfNdiKeSCkoMrAW6JoR6sIuTSXAlbzYgpsEz8vIMUUk0yMzPqcAC0
szWzGfiCveaGFlAdkZFkfaEI2kpS5tc8N9Gy0h/xnuePK4ek4dMBi2Egvk6uMolSj8vdrQGokUjM
H3eKU/L9ch8eXSA462BKQs1O5tEgNN/kMY69tCQNHKelzSIoF1QW363GC14v+KT8w2RCulSmnQA+
/U1w4vSZ8LPKGEzgFZyxAbHR5o2CDWLFQrFUOV6XZsYLXyYdReHri5GnEf89qnEKstkyVodxUbkx
fTo7p3gos6zfHRXNuhOVMWMctLD1nXJziVv0Ll/YDZEhthTRO3k+RVaws1ftoZmAQLF/64tMXBe3
h46OjBX+1aOPF0NFvCloL9FnTwXKWsfi4Pm2QZKYJaZ/DBkji397HwqGWlPvfuZKOlYuwlecVJHY
XCnKGZnd6SwFeLRjCAJI2rYnKbxSbDrqQnprKEH/oonWER+mGgONCd21WC2IaUycVVue7/VVSjPq
0mRvtrNVVAep7Zurd7Mh16tTTi3iE1/0Qxm960TRxxT3Yh/QB6obYsV5DbT86e7HJmAZ6WkUBBdS
b5Ub0w4Itom4FlFVnWD6CvQtzFWbbL5lfnQ4NHokAus+KL2ZNAz63cvisgoKAhWvnhtax1j41K//
UOLfc5SGMryr7f6fvCIj5YaD+caQ6JJ+KruHRbbaOidHjjt+OQa8eKinWf3GyLUV2Uos1AGD7BoC
3KVrt7M7P3K8FvoPKC3PazhqKicy1FdNPhyqDn9NEBz+sf2Jm5oVkAYHVf6JDl4wQm4tjo3jRpz5
FU67vyD8UAro4XrzjgssZca6Qfn0VuXZIBQ+nyUKVxhtt7YImk6MG9bPqK8piLY0lnyb+9IRY+Gi
OcadHbZjNsC6rjNljiDaOMq5BPz3h2mshxyUcPI8VXYoAO11YlBw01DzSy6XGH8vbYqHQgBJyj1H
M2A2xdV1lJ2mL2FHF7Wsxq7f8v3Nr70A/+Qw9UZo2pkRAJejcGl6om0EXM62rykD7puJB/T9vf32
6BF+bZ6t+hziLHnDggwquFmtdOHu6lNt0eD/Ciqieul1l513rKtWIAWQ9l3NTlSWVpqlkkF9kNAQ
/0CxeaPEq75r090UaGz47WIooqXAdR02moiTN5GAJD8gic0wtUyglUZTAgpUZVf/IZGPruoVzH1k
ChHATYj+FQ+6BIHg0VlBwCuek7KD8h1BQzYj/lE+YUKB8w7A/BKSHNZ/ejVlpd/ozZQKOUHl96KV
QDsAgv0U2xJcoWZ7I0Pc7DMZUd7Plxo27LuZrSS1L3aKgm+cMQx/4YaJQSs4axaglT0wSkbFkHdS
XMl8zFjBl2wKCoAZYz9mRqz29NxeYLAxSFJ/lp/TGZSi6AQN8cF/Ja0RLagTl76GyQsiNm+1Jy6s
XiuTgm9s5/23NUdd0V53PoSOtAIepARtKtacd6LhK9SI3dlw1J5GeOYvarvoU7Jn3p4kZvd22Nhk
+lEz9oVmm1Z+9W+Cm0tTXO5uEPl9mcFmDi35DwhEs7dT4kQ210IIYhtEWZ6ySCZVc9t88ewdaU6F
W6m2ptfAmmBNzox/HueuBxXTGN67IPZzSgDffl/LWonlFO8fJDHwhmSOO65oHN+F3Yqq2EGPc912
ena0+nr0wtHIZmOo0x7fikOqpehBHyLuyDPLSMeH90uww/OZHkXco9Np9GkTOiSTGKS4bpQZITiH
mvLbaYuRVerJ7Sk8weY1SYXZKykbbIJ4v5g8Ix/jVVmHAi3tLUUEitkakOQTotzQS3DbJX9r5w1u
Icbry/nzB20EpX2Ju5Ayb3RDx9oHC1ui/LZ6wKqid+gvY6aJB5DNOsyBYE7+rmxz+u9MTXjfEi2v
Mnz4DacWr71fIteXuzwlabFY3cYiWRjt3Zna5agM9s9+R2t+JJgrxiFBAJnYmMSf0HZdOiuANuGY
mZpHm/VVJVKVL66Ep9T7kI30gVGXSdyjDqYw3kMlnERnhkR2O+Gg492KJzqqpT+vp2zrc2UdDlx8
pVHUD5Y5CQp//1apiX9lbey3z8sfjxbaGBLIsVta60TlhyqR2TAcTegdb8uI3aptcEdYlAa/715b
QarsXxhcPQ5tXCjENzvgpJ5AJ2E09naMyT55rNQNL8oXm2igyHJuagcUepus9vozlmJAJGu+H+gz
Iego8ENCZQfr9vamXQQVtlIRHYkNkMxigoW5Y+iVwJMZWs9eeu+pGNbokkXfjzhoRp+MqGhMeb3R
GjHbhCzIzQWj2lkNEBqaZkni2rQrcpixditGnPRqqg92OFJa8nQEQEmCkxJV0yGQUsDexovJe/fX
nn66n3/hxtXblF6cky3O2F5wDBr+q6cZhQ+GDISoPcOL0YqwNFx5L5tjwXfe+p1A3NHzdtWw4bwJ
iFZIJLbpSIOw2RD1IQGnlYcNFSFi7hOPdQmslW44y+Jjzdt9QJb1ceOIuEk692cHWY0yystxstVD
5SO49oBQp2u86Lh64DaTFhP25mocGANpQvldKivMYKp2FVZDteuWWutiSpUbi6dsN8UKFqQaMiNR
s85n9WrpmAqNyaXiUX8P6LRQXzKbePXs6s3u6/l0LXQInAVXe3vDHMh/4Bx03R0DuqTLSvHIADTE
mbGdfe7yLfSIQc+9KXdzKdoD850IcQoOA2cjApZr2i6x6PWv1iADh00Imc+aYyHM7yvVDYDhle36
g3bHynsu10LQenEP3f7G+L5Ya+kSNnD0/Os0Mjaqi0tcQ/pZLelps+bEQReaf8g1AbbrFcB7Avwd
Oyh41W31T9RlKnRtFwtA+3ZpWeusETEWmCI5J8l8I6tarnW9doREFADandYWJvStB/4WjpUlDIzd
QK328HnrQ0OiJhgY5LdCHwKj2VJKCLuM4UkatohZa3w3zyMudw2XoMAwr4tBF2+t2bJ0ZabncbGR
6owrMaybr9SGaPfKleeHpuWcDiObCsZkQPGplIlY1EPOJOofISHkj6E1NSvOwqqu9ToCZrtCdmah
KTRzz4jyPxGpNLU+t/5ziC/PdEkLviQUb8004WJcsfievMSxLg9TgKUnaj1si0v73sBoKLP30d7X
1xG5UT4Wsg+UqYhxIrc4EYrxxUoColX+SnvUyVZ98OIpqGyKHdRQOxdek55Mzx5/h0+3ecn88/qV
0mMWzfuu6sPGWH2zWG1uq6t0Gu2W0qD1XkrqPavUvF6zGvyYAi1wcjdjcJQt+DCllNaYypdgr1eW
pQz1VkwZ6Nh9dJQBO4GjJb7j4jGe+LzrD617d040QhNMHF5E+wOHcgZmklC4P5FC604gA6G5BhaS
Y6yzKzpe7D0J/e8P3S4uDJ0L11AAZGWVAjFwK7abhJlVcE5vNbIG7rFPkjuYpYuItEuq7YLzGW4T
lz2JA0s2xBuLjaRBO23vl/CgSnf1LZuQaKk4EnKAoGCCZwOZRhHOF0tmYXSK35BgXtEVxPReCzQg
7mmXV7WbgofVVhmO9Fb1qUEZPxKdlAUyuNJ5FPyM7tgZbBl/+KgW9MzHiIElGdgkqhz3inkCRp3j
+C65UbIxryHs2Fv0eiXVKf85mJpZuj8S7xJeeP/Fy0WjI2I7Umh8yyaLLxZzrjqLbCGwGO2IPWhc
6n0KEHxaXQY6xulC/dWIywLlL96BgbA/EmSsot3YOZ5gKWu3Luq4dafgDJeMXXeKrErXbYg33/x7
VNDJGmArgDL8adWNakw9PzmuYIyiDC9X9zHvXnvlCs9KUCtFAA4XP4p16+a711s/uMBEQVKDFXyM
8w5YJt1BRMTEwUt58Hz1ngkks/tEcYYzgWqO3z9rypisnNjGzZfzPHLg2mZkPkZrVjQs19KnOJsb
M3G702h7pBin5XfRuMA483ZlCII2J3vHUj+CYMm5ZwWMU5+FnG3XX1KkYZeLIRHW1KwQGJMO+dCl
Xk8XbjEpbbE7XBmZBh6suE0qrMAYz0XoH5QU3FKF1tbKusNOqHBeXfhq2+qfYVu2ajucjSWuqAvd
VzuBqIhz73c1ZxuCzD1hZO7R0SZkpC+v2FK0vqtLGoALLSzWBElCTN+aRxG7dND75bAorc4i/BDF
wc139P1rKQmkbRh0RHgvuzrKiGzHzADG4voYVLW12LiwEOrUj5TjjmR6kNAxWBoxiQxuw5b+lctD
UpVan/Wu+I967vuh9K5JWM7maxyFV0GZRC/wwqtethZpTzoSZiTatc3gB7nkcxdf6d+Ti0uZ/EAh
S+VWP5OBuR4S1SqyzPUQT+DTpsVfPneo/5ktxMZ46pg8gsGeaKThqzHN5YQ5PeVa+f1GVr7LInZ8
E9YYWB5LTxH/R4qsCQI+U13FqH7ys22c2mVbe1fMpZAQ1aQsN+g38DvPTlG94b3JCBfvq4n+D7e1
YxiBQGznYgYUVQZGV7QEJQcM+7NpF/iKoxjHAj4/Q2LAjHCL1VaE+Zk5i91v8Ejhnzm4N3xmedvi
hjBJpHG97i8dG9Ymm3DiE8ycJiRudQZvn04m8eSqaPwEiQ5Z4ZgmzEtemwFY1PAHkcoMjqU6giC1
Ys1zg9x5ffAAJKsxSipLWM3r+dAAX+RbLLeHUCbDM4bqJ9UHtueEFMVyJ3MHrZHFmICJG1F6yxNC
til2/4M38GPUOrDKvaWRCVUW06SLANkP5wrES46ZAb6MSpdKTVitF15gGGWDGrfYqEI0YYwm8wuL
SF6c/OyLTMW7z1GfVZJwyKgprBz7ubAUn0aHTt6BU0Yh4lg49txXam3viRKAUaNJaJ9/frP4r/jM
lVUZKSsm/xxkidYxsTajOsOFHxSa2IgTJgnSpsEBiFL6kWStuTh6nka0yhFbMxjRSwkcxWyOtXIZ
Tkdm+mXIgj3gMEzEmMsrCKQlNuryplIAA8nbGOQYJp0OfDjTHk6ufrrzcfolrEto7sBR5f/6FsPO
o+8d00uQqRqgJrFeOli2uXGAIwgIqQsN4ZqQjja5169JYD+v1U8VWaP3cVB0gBXpNWbt1ZHY2a4u
4zZdIyDKOCs96cIrLfju5m6WdV5Cf5jPT74t6EpvqHSkykbNm3/86rt8JBoVx8Ove/Iz6Ej4xUKr
5csNfEinHVDsp93xYmMiCdrvAUPF2/AoOajEyJXb0hAZBtgW5zVpmnetPkdUQ4XCuvAGkTEDvINs
S/a29hfJ/H6chho6bmUV9Q2POLkMzXehDtjor+AKncopLQazjUthMd2GNogaHas8h4AmpSiXOpPG
V4LHM0OrqmHCgmoUL4t8xB51/mGgsN9/sd/VISYCPRCDPHq7I+POVoFtvSPQxUiG8TOzs9i8q9oh
ZMVfHwIvJ0TJsOawE6+8nwhY9PXqFgBODHRw1bpRgs7rU9Pdj8Rq07J461ySt1Rto+BgsflAsM2s
IBnm7k1cv+/BZY8xyUJAMn7OKW+64l+KZaLbijCAqx3qD2JU1B/Ye+4rJ50GwYJ1UiFNpofi0VzV
9zCS3BFOsSNvfRqq2K3OuhkHAftOyS8K6m/eMtMTxzLeJHcJKC2g9aPufZjrILroFjkax6Fw3heZ
utyi08CMcbjA0HCsiscGCuYR/cAgRGp1sw00dOrobVZhE+YyjftpYbJffA1FemOc+vBEJddDLwP7
IyrGQ+z8+47KF5EIuqarESfbHxzaAL/T/ohXVXaN7TIIiZEAHanUyWgu4ZCBdcxObaVIYTVC8Q//
SBTHZjyNsqCJHhuykTktV+S/brJ0VbmPuJet/uwafYoc4z6fFIsxz7e1vhyJDYs6XcDkKVYyZ8TP
uHVCmrb1eiI7MS4PI+m6Cp6Pmg8JGgiM4XQIk0IxOb35VL/G1JqOHW9Hr0GBAXdIXhjK7tg0HLEK
syMpaAs0GoM9sV9QW/wzzwHrG4fb8uEF6YYReXSapoLni1Z3jjfQqsrE2tnA+diVEq9RRiTd+AQQ
RFt1iyB0DPBhwM55mwm77Skp2WN9VwiPkfh5Ez5vdwi2W/SUG8VQTKOJvxq3yKra3tNntESHWuFC
F2p4W+1W06RfSoHlLFxP3OlHGPe8pOAXJ9uxMZmBMW1lNZGFnUi0AS0YBtKo6ssPsbNjiS7c5d/K
B1WMsdzJsjcx8m7uDXcHkwpcyIwelZhfiXWsegS0NKnYKq1bLHVG+WpHZDf3CdshI8R0B7FBmM5r
/UIcHhGRTyEL6Z/ibeSUkSHO6bfGv/OQnJN3lHbfpW44kKRMbY1+iYm9wtZ0p/QWVAUUfhTveDIu
rEMTgaQoDHJr/UwMEGy3qOUiGWdC4VsYlPvWi731yz5yd1Lr/urzqC3VHXQzzDypUD8BC+zDoPaJ
i/0od4zNPTowQPbsyCAQX83e9TygVlG3hMaprQghChi9Rr8zie3GpuReKrPzqtlxqXFgKqNGEk2O
MiaCicYvvBbf7QNDXbK807WFOJ9owRhQKKxtqVqPQs36shcCa1/qsTzrEBBlQDPWoLEF8bgla6zG
D0hljg2Yb1tJJIC/KZ0v4wHmvGIwro0P18H+h1TQJb/sRjqYDnK+dfYUEUM7aTaRsYNIh09t3nBh
a+aC9hg8z66BECsLUvehkIM9+yVYmO+XgdF7a8IakKAUd1l1oEbUd5ngfqIZPtHPILzP7aUD7FfM
YGnqcPEt91v30PjV3ZShyfHP/g0WibRrr0rxjcobzIWAtExaOzeF+RckakPLEpJzwll3InRHstrm
rCUB3HkDWuq7+FwwXfByr1oPcNrs+cFUTqu8ahAmR0Vm2oBbQ9uFW3lID01wP/zOD+bT3aybUuZ0
sxwcmmQXQ0cxjClHCcSQEFUsUjQSHUwn4TdKKhSfevldosu0TyTsTgbkeen4BfQw3zybRfox+/PA
HeVp5xz8QBnNpMKtfZ0o8Xayd5iBKmLSGPEoButIlX7ZjpNprAq0DEytlXO7/DkGWMjuw6ke6T4R
Ozn5zL+XVwIBhJUrF3HQEtx9iHDYtBujXe8kd2VDvdTPsnLgqKJL4raLlWqu8Yw2uy1kLID+4+hX
drhsEK4ebD80FI5GTAPzxqLi8XzqNuaGZARvu06gqNdL4lzfeavakIr9iodlKqb/UC74n+7b7fl+
I+Vrwa0Visu4NXMbYZESjFRonqlOItd+130ZuafgSvXaKLoVL/t3/owkvUE+gXixll9RVgu+PAN8
rAYFSBjYvB6fttVNFhAZyVOnrHhxaT23iR3y6x3L+ewyq2JXvOtPrSYPaqiQ+j3seLeCgxVekJpL
ka0v2Zhcuy4fisRphFptmLGXMcdI7h/TR0MQNn5MndO7CNdDuJUYzz0k2hFvjICwU2gKSWfXzC7u
c5HW/yMb/vJFHaW5rQmgriJkKux/e/Uo8ICriVqDPugkqu9sry5xLPUzsWnAtVAeuFB9b5ym+t18
pL/Cpusb8fE6LJH183yIFU1qg0iCoqYTu8qb2GEXnRKwaTgBoBV4vHHIPErsS7lhquVhJcpZutlc
yQEHLfmRqtbHRAzCTkOWpcOy1IDTxQ9HvgnGjw8dz0PTfgQlx+5qQcCsHeVjTLqoNOqH5LO1o7wG
DcsBj2B37hkkUhE9h4W+R600sxKjg8TXuH9bDO3+lkS6PmJPh6M3FaW0w1bqCxI3yZHFrA36Xsgc
UWRAspGGLKMTy7MVmZ2ABuYan4mQ93jJT32wAVod0it0oPIdD/wzbsTGXtgtOMFTsPzIzGGPXEgO
USdMnY91AhjtPsNly6tA5XWg6SMKlUST0WfTFrP8zw2xlP3f7pmSQXYUi4AkoI1WG3OowWcmkcAC
kSRnL+P3k+evNKZ3ObmWUhCZj+r+AGlsv8KtZ4hCrBMmlSarpIMcRX2V3EqHNgNUuw0AgRU4EqDV
o8Em9WM9/4MlLnOOVALf1Hl5HCWKUCtRhcuq549/hqCUPJ53lN1qvr3pWkVQtF6o6ok+9Owg9pdJ
UC+rym0p/HzvhwWliLJCPu4vlTTmhypkvsd8SKTQMGRO22CUanzlvoMKrz67dhIAw0Fflsz5ELDB
FbNha/1mN4SbIvyDf+jL8EzFOCkv5KDxShTLxASXmNoDZQ14HTMFi34JiUpeAu22JPMXcft9mM6B
PxEJqtwBC76WmV1fLrgEBHW26qDfTw74dQxPY/zHlGcGL2c4F39T/W1HA8/hEBZT/RQC9Xmu/krQ
NviYwbS0/hyscDHyS/HSWgANW/raCwX35mMFYXCcPP2m0sNi6POimKST9DUbxh5hb8FdRuB4ejsT
KCg7dBu/IxGHdf+xo+NUNDg3o2rLXM9W9Q+iYBZcvS7PjR91cfwZxXa+Na15wloxCiWuciOoza5B
nf0TRvmsEmnHU0pgQE55OUdtWj53MivurdSAVDANKNO2aOKiUpZ7TRKx0DJ5hys/WeB29h+N8nTO
EZlkE59ott+BnOCrba4LCcj/pNuKV5f2YNIu/NNXap6T2CXqH5VEYpgA027wcimGZWBHPI4iMuqd
L4jMglsMI4Sil4qmmKZ6ZgQ48T6Fp5PJ+zBHhIipLVr1LcSg4I9HaZM0NIyTh5HhS7IlWhlTqAuX
Mxpa2pFezZJo07VF2rAcK1E+7YY2gC1lRywFpaMfMkEmdK9BktKGExktlQ9V0E6fyu1O5mv3qU9V
k6z2mejVwQaGk5wthD4qVUiXpG9YflYlF+PzbjdnBNuM42iHscBaDPgH8YGwquwlOJS/7zKkQv+9
v03NzUYWouU2my1+FyRolvcllWSPtNgG5QZKHKo3AmALTQ6wyQyT5erH7tFuVtGW1bJRT7wQCoBC
mnU8YIx7v1EZ+m+967CX8++PcZiwuw1z6PUKxT6YI9QHYGBNAlmIz2Z/gnrzYdr1RXp0lMkR4sCS
uSHRE2BjmvboEeS2OVdzpLBT80HzMrnszBt+IR+jDDc9E6sVTwpiu2a+aRSogDwAEX+Qedkp4G7k
gpdWc0MiB6Aqjsh5bgynHCZ1lrA77C3EwYShvBf6gV4GPJc2WujWwUveVEfM28hBltJ+qKVbsF6W
zpVICl5W3xLE6bp7okx3pRZHEl5w0c+fJVXofl7q8b+rXp/wYAMpu3/ELCnIsxPpqmTMR68D3YPj
SkX5bpg/3aZpgngWN0rbxSim5mfKoVYDrUY97WIumirwKCnh6loGNQVkpXgAJ0HdgnXChER/oJZl
Z04mkLKlQg3IS/d7ZSW8hPy3ujTxGz0vlFeAlrvrcxzZXSEOmU7CVqbECtZJyPqGNDcZlfEMj7/x
463m6H9JlaoCe6+tl/3ONHg3Y1WrjLvWmAmfnTWlgqqbN6ZdGPUu3dKqg/By151NBJNbxcrS4/tR
lOpn/zLkMGzlljslonfq+XwX2SG3ptjoMdLK1hukrNfGgKZGWxdN/EpZopM3APmeD4kgYda4LBB1
NpaYs2PdX5jDafIEkYptxw4ogA7dGdxEs19oOjiJxLlIMarp820xNGPUgyeLwHWgGDpWvLOf8cSl
AA61smjpL2eTxn872Nm1i3C1xzTiwNxihGQpOSzgx0kl+M2BGVO9ul+2Unwqq7yhhrX4vOCxxlWG
HyJ8vTSKCTZ+A5eJKH1gtw+Ba40rr7NUbZfg0zQ489OjUGD8RH9Tzu+ErXsBZ6LKbd460HZBJUBf
w47w8sT5WoembTThYejWkspdgU8GuSgWDSSQV97gy/4Lv/LpaTUb3wxZM9IJ6X4TU2/sdBCGBnzg
zw7aj4choLrSdSqXmCOAjenyFlQqj7cRuUu7BmDwV+zkYaL8FVIw5yR+bTeSppIHpDEcNuIUP24m
1Fsq+gDdnlfY1EEXrOxGXQEFlcX87tLeo+7tq8JTF/iOUGsrEmqtG0KpoTm8sbThGURGOabD1v/A
PvGpipf/08GZ41QhathIW8HdK6lcI9xvMZ/XLdl+txuOMmit3eVgmlvT/QLXlWHDwh/z81/ZcHdS
8UWgx10Ah2RT4vE478BhxT+RH06LT4WUTBBAfwViB0/z6E0R5gdn1qEL9dQux6BONWAT6E2ctANX
oee92m020vTBiKkZMh2/v7Sb5+6Ml8tt1IG2sn4jyTUjW2d5msChuSu/5LdOHIHhIkRwcadWmc+0
VHTqEHBVGods1en5ixqzy77+Y/9VHjh3aB8eog+VLTs3l0SiBRN2tN6pN8D9gUWWJGY8WDohnrEe
pOgP2xhtUM/8skgxZReIazctllsDrTrDzUy5YdjtspgGM3FAXniIEyTvEcrGOGEN+UC6walpdA+Z
X6JO2FHkAGUkUgF0RI9PvSBbGL7rW+HvLXdr09FTD2X/PP2qDlzLLJrV6Ptg+9XIfOsgCLP3r5LJ
0sk6zxl5STb3k3o3FdbdfGvgTcrQaLSQq4WHOSruLrpYBValefKRa+g3Xb2RzT79BMvOpdhGk7bj
nzXUrv4cmgDTqUnlmRab+XkLso1YoIRtndevAz5Fpz12m0hXUfzZH6UYA1useQf4gUem64+791cY
TYemZKvUZgUGaacAZufsYaXu9m2WEmXZ91B3CRzLZJM+Owcvsb4/OJwWQozW5CYyn7srhUZFk60F
iQo3DaFmVTz6uzBRCmxso8J9h3ycDKdHsx8O9+7ZVQytJ+BiMxGJSQaYsQnComWWe5yWrUzfLLLd
u8w6/gjIqirZ8WGKiMYMN3r5paUBB1umpsWfuGH1FmGVLnOsaWHW6cgtBcA/vqxXltXxIUoDHCT4
E3+mJELRTrXVuwI+R/EloxPpR5AH/rHScBJm6hDWwhQAFOjUdlMh6RBY27mLNXvyR+fP12Crq2HP
hVVY8waOAxr3MFqx6VzR/Vk5yLO1n/9qokgeGD11SycjBZQTdlxsuYn9FtLthE7c0/COuMk8kVU5
THs+z2YbThjob/QmfTqAEj9L/EEvY8hu4COb/Ni44zu4dkzkDHthDUSfhhkQPLJpGy46s9LtEkNZ
XAkgUFcuEhUaMQnYZOHwre5dnFOuZHKnrmO6LhOBOqrXLsmhxWv0X4oONzjt+hPsFtxNAWr80iJ2
rf+DKOeBwqORkQiY2X9jCMMPCOeJIvVTyHy41Ok5DigDtV4qSON3fL4/uvYlbIrj5Zv0pMFMOeQ2
6JHeMh1shXgGa1+blFK1PddKIg4JndrnvRE5KN0gcIqkC4VNWvjFhIz5yLLx7kY0qPlSDs4RwRdq
hMC02T2Zz6B5TH8bCzHYAGPNQVFOwHPmXfMmPrQ9Ceb3ZQopuypxiLG6Zl8kjuSt4ofbllPM7U4b
QVw1VlSXSBZNGlHkGBDP6ZE4SRODd+91Tj3Hrn5dwHxDro+cJ4siG4VQu6kpy5HJZhqXvKLMr+4e
WSSgvgEnH/uZ5BXoBXrryztvCTKE8R2k3xaktnt3FiZoWiE+QJ5ttKYaWPfNof+AG2JY/XQfAT47
Ejzc1OBP1c8Ub+uciJfmGxXVnsum22yMbXgjVU9Ing9p3JTi7B6Fv9v7CWYNnWKdXSuso+e0OiV2
3s1wHvPWEJZH0HHfvvkbvW+wmenO5JUOhnSQHAcpj8ydLd9v9vVJdOGvxurQBnstCXrMMA12WtcA
jEkh2aZfk3MDQbvtp+E1VO9XJrWXWJ6I5Xr7KhCpaqKL37fBSkajpHJ1mluXqHFcSfVsDZfsN8iZ
PAhFm/NCLa4xPQ94ZEuIgnQPK7hd0Y2F2mofoGXEA8fFsxSnKu6sliel+9IyUxkG/heRFAoHTE1E
UsKUwxe99dxr0IBUiQcfBp1LP3NO8o4XB5PP+aAGpFqlM3/oqNGa+Eng9I9MBXc2MtdVvpc7azay
52HuYGaUZxfHU4ObH8Y5+gNMCeFuEVrXSjzn6ksjiQRzTYa0UzAQBdKEbKV0vVD1oDjbuARaj4EZ
0ERQGaAwaIdQuKaWixRuiygmjVbepsIpHXBrcTxomJ8N+savCm9KrliyxRJYll91mnuq5VFd4EBQ
yiDm6pljt7fZ2cx9IWWTzoa1/BSw8DKaCqQjwvgcmficsH7mcSvdIiN7pkmZsaarSBomB8Rijpe/
ynNVFqMqD9jPd0AJd5gjcrF2lhHtgvApMKy6+424F08coSC/3QWsODr9lxsBwzsj+2MzCqY/BwKP
IX8EecA1K7vaoFAFDxKOBkebUl+IY1SYZV83g3cfbYKGTQhFM++ezJ7n2Q8OGnO5RxHcO3MYuvvF
nfwxmcCk4QVm/kcfdFOZWa7SH8XfViLTCRFLwgQXoUc0g/9ud8bE7VgfVhPLeUXusBAtB0ntzXkK
AQX3lScaHvR8IvaI+QQYcQJlLZUKTVwA7bJfZzpYbnesAHiiALM/Jl06kCuebuuVBVlgRTMPf1MD
uqO3CMr/g9nPsZChsAwrlTwXB6jQ8YbxyBH/aV3if6q23eROiENS9RvV7vFbRLOaDL+hNtzBVO1z
Dt9TjYRF3PZd0R/4z1pcz5wA/GhdtgiRfHNL2qXYhj9wWUOg88x9qdL8U3vFA7hcjXLOibdUXbql
kmzTsaeawtNhOnJ8yi0j9vedUU37gDW/dB7gFyQqVq7ikJB5vu+WFDkAoq1z6cX7CBWzwcipw1Fe
E9F8icoEsSBxrI0S+xCpk/zCOEIV78d8PfqACpl36vKot64IWD8wE6DakZRi8BXJqSV8oh8limoa
+RDghOhOOCTRWwqz2y4b5ejst5CjWMtsaHaEeI8T14i23EyV55Q5u6jxqyzcCVSg5Z0nYE7IVPVo
rCxA13ZWRTln0VBPurXuBPXhSMaEjZo5HGLjoXXL8L1vQu/gv93C4Eml6JZULxFXCAHO/6dFd8xb
WWOiUEb/iGJRPIxYB8ZnF5DsAwt2sT962nm12hJ1irpE5RApXLHdi/3J9kDK92dld7nzhHC+okVx
GFsaQxRW/j4sBQ3x3YQ0Oh8XHTGUtdq0MuZZZXJHVOFK5ujgRj5FCon53hF78vBFIvimUNdpVBNF
Nf9BODeRdIgZoiTmjOpnEOYcH3oBefckwzbwA22YcmnGwFQB6FaIuAiGVFldTQ36nc95RHEF2kka
oYEcwF6FL1F2EmwgZo4+qQODzLOxubcB10GMGDusAWk58TS2nkL4K3pbMNAjAGIf/bepgjbFgS3s
i8xbAhSr0zEii9ElXbn0UeyedWxfy4TRESYHK+cgrDM81Q1+3ZW76vtCBoDJlQX6iTi6tXLmUoNj
WBxTVDZXjOrwDp1tPBlRMgNxILXV7gMmgyXNZR46aFg6bea5P+7GTc1ImmFvfe6/N5VxL7+eOHld
/gg6X7Ifs0sFMGjWE6JBbP8bAxgq2ElpZfn1a0UyWO20TfTesRcJVb5HziGcxrAuULcIdBSm6F5a
p+HcnKPoQNhSldbvclyuKwx25ZWuJ6chryHqBpBTV6xCRoopBwTrMxuT5byDgE4lM84sLFQcPGJr
jhvemSwYtSBUTe2w9v/0z4V2vlX5WMO+qtLHNnHR/MikOtpbpD2a2WPNMBC/OZmp9rUJAR6QEDGj
g7TQmgJs/nKCaTjjAc2xuKPKQQtBmbDc6WchmAwidJPMBE/xvC2flfwtbFN1nGtKm2BhA6bfMawY
qRvEsahbR0r0QhlMoExjlrrNn9crrViMlSTaJLHSyXOUPMtedC4WNb3cfJpvcc/HMWOPjN79UT6K
xvMItTOj9pG8Hjc1RRBcyo55TBCepBATXVFpu1FMFyEBUE+eMrPX+3GHqkvNTO4lsX+haROtWaxh
hsqf1Ypyu2Vgb3Zv+bdwNNNIS8FT/gMI2NMY2NoO5PN9ztukGUMpKl7ZMC223tZXzlZhPbYgtpCd
ZPrSH5l9x/sSlz1X2baCe/ebg/NrcllUrR9NCWinq1jcRYP9w56+iJMu/SUOxPZAnrkFyJmZrGGe
r+f/Xz/TPv879JfIAlfxTE3O5ekE/kUBEqH/DobUTdIC4Hx7toRmp1PIc28TvdQkt0hiI7WvL4I3
er3hQV159LTqoGnHWCBNsr6ufIjDpZMctr9ZraM83IQr6no1iNHoSS2iQ3vvsljhA4CUcUryxATO
Ec8wxLz+jKv5o9vP/wCkaNmCloWHtlN2sXH9e99SUwJsPV25j1fGMLhoiRQRDdDDUglpvGe4frha
+i6Z4d6jYsuNDOAZJWCM1saUKRYh3SsTjPnFiSHgAJE3sontMhWB0/v2KBcvIS8DjM3I8EoRWYjf
VmCv45ZUX202qZTtMSj8v3yBcAvcksxZrVXHqDpJGLzKhkqr+PQ4Yworp9N3ssopAk+8NnPmtKHW
4FONLP7ckzORd2f8azGsXDOnHDQ2WZ1gjlpx3AqQ7sqzTRrdqiK4RW6GvY040x43NJNvPquEGs9I
DL06V3BGXGWSM9YltxnQmMMHei+owvUNCuPYHh0fs8VFoX2PAi2NbdDabra7uNrb1opClxZWfJWF
LytnyHFOEIUpPLmr4qPhfIw6I0WEJpwgZe7i3RnFgi0CkRUJjEHmJiaJotVWdEU4WUY0iIK9vuTv
KfduZD8Cy07o/3pbR20pcIKjoBWDI5YGWRPG/N2z3GIExvNsQF2/mPAfKMxUDPDBH5RTk8LgfUSc
IMJpT23TNaImNpi/KCCvrOX2Gb36u/akaVaHV6ZXl1/soKHe/CIBySCUyP135fzV41Oe8esz9+vm
5VddicWSxYcl9CcXLSatc8+481Vn0ofMnK5RZXXGyU8MzyXtYhvr1njfxtVlFvRqHiNiR6i41xtw
GlQ4Ey9jlmk/3gpbZfk3LHHRC+L6nSf8ZXacXibrN6z69gMieMRt7aAZyNrNq9VTAj/3E/cjO/q7
KqMDLHoApLyjNRVwp2DOwVr3922NJdprROobqCpLOyE/fTIIx4V51jaya3ibSQUpD/2TDkUQz6gb
MR1dH9Jd4jJAirmU2JFn/vSSIGVnLzF3c4/KZXfUvpDuK2eC8XSABGEv0pwlUVvnEEPFCH08onEG
cb/krbJOCluIhrmAnTpjbZ6o7bAgDE8zzzChb0K1KkJMLS7sPdQr1K+xHdeQioVrMJ4ej1QtEfVF
qqOJozaji7zcq7ck0A87aF0mII9beReuMBO63Q+DOxtWTeyTk6Wv6DXBJ40odOr7LKuy5wnhjoDA
9QUvZ1BmgWYkc2T6QMqofHE9Fc0OmXpjuyLrCRikeWHWhxTKDd8mlN6fw5S5xmjpiCSwncJ99jxb
/8jY2QKPvlMrZ8M0VNU6bYzEDl8WerdwveDG7UeeHt/0Pd07XmtZzYNA+kwB/wRKZhy5y51sJpgc
iE+A2s52qSgB0vjZG2P1l46aLYNVve3SrDlxrUVhamjEHuOJXB6vLl7+CwLTigVAVTphm7X/4Xu3
kJAyXnIGkE8iLG4XDE/b7scIzWqjoHOTdUbzqQ+nKhGHb6+aeK8d8H/XFrs75SiRExHrNmC6a+ef
mtatp5rKBrrJA1rzwChsYyDdaxgyczh1Umrdso8v+uVmWjsh0MvjcaXF85y6RBwoK6LSVXNTp70d
slp36vt30tOcSG/cwcgF2QXHiHGvPTaEPf4SgPMJFS2XB7yqec+q7gvp6MWNTNY++lz+/KTYeAyI
PbhbzhI/aIuma9r2V95RmvfutmZ/XTeYltxXVmTKiTFWO5LEk2z/A1lTOahj5XahSuA7O+0JL4CC
/HBZOIcwWQ9/nGqwFyvMqStc4KXGuVup7d2k7E1pSGgu2+dhzgRVdBovt5ooXNAsV85zsBuds1li
EM1Gc5QqZJ+aMYyboitgwezqc7XRWqaHewycBeqYoc07gdD0Rf/sMmghhp7oFN4wB94mKwCxV4Oc
jjqMAW6lwopuZ0vJU9IJrlu78PhPY5phgLj86kpNnPtMM3gkshDp9dtr2KIveNqj4N8Mpw6rHXR9
7G24KMp0E0SczxxQUDZr/HLARpk50CbNkP15fKIvO6q9ZJEF0rmaap2OUmGa+i8SQ1fWqq15iNYT
sJszcnRGLObL8xrxOMk5xmwLwDRks2Y34S6HPHBqKOYAh1rRcuQxyBDADyoJHGw6OuDY2TgZSio8
ouNlk+LG4fYsgqh/sCiw1WuVtyYuntOlBhBXsZptSbDpyCPBxlmS26ke3tSLf7GKhvL3MM5Lbec6
zxZjQ/cpnjHmo86qXyURYihiFUsOVzvN1bhruVEhDVKVu/hC40f/5BnkP/iNOuOBFSaBQM6B4wHX
XopYY9toyoR/hSgKdvES34VfQxQAc8R9yXjD7VnKG0AZMhP3X2RP4iypckkKWaIRDGKKHPo44ix6
uG5fsdM9i5UUB/TYlgEjppvZs0FgRohpW8XwqIH73O1eCTLkPR87bC8oDivxQRAlfGOIThnARJMY
9qq8uhFnp0IZgt8Z1lm3EdNhD9EUyaFpmMr5Rq9bPTiO2jBD0tKbK20OACU8wR7FCovRcC/Z/MRF
yFKOoxt6mIi7IAoj5QpejEcMA8btzQeClpCbWIGLve5OGXM8q/q855gqVK7odsxEvzycl3zY5f7q
YnN49vPxTUA+5XbOHRABhFRgVpUO3HgMrj4GaJsyFuwcJyB9NLZx/nPbYU5bwot6eDT8qBk2O0UO
n2S+/s4lBPsXUZ/r9GGoMXutVbqKG+PUKB9J++DK35kE1FlCHnNxgoD27S5fOlE73o8eXiKDa54l
+TJGzrFdw1phzhZFuD6WTujS1nGt7BTGh40+IMAwegWZeNwaMc2nITJPQvM5fYqpzStiZCX60waa
FTaQa5vLzbX/Hq2F1MeKNjIkrLFfcT7+Awuc5pcXfMARgekRIFHQzWECX+E4KMeAbbtShwLEQqv8
cXkvE9WNeFaBUycuoiWAMeOb7AW7/Wayk/leE0FrPNG7vpWEVuOKHL8N1V8nOo1UuXfevgbgYM+Y
53VWsaj9du+x1S50cGvn3jYinaeNrXyLUHIz1Nv9cvECzyFcQckvniHLHuJMxuPu1LDL5Uf7mbHf
ooA4jNrY9GKqZwj1d3DOMly7msJQ6IvHgevNw/iBlKRjWlLzsVZnFTGkS7Ny9D5ECqfc5jDvBC4E
sEvKfnRjAV/fmy3Dn8nBd3OvvimwsWOY1TLWV4gzYym3dgOwA8QFe6ujYauN7fdPDHB3zuWOoRGo
lZ9jtUfNKZwMdyjBWznsnu2vOT9Vo0/RJwqws1oKxNRiumSSHJhV4vpx3LA2GYy8PvoQdNUYYcVj
/++bkxBMejXkGiG+/9OvW25CB07/Yu5Dv90/IO/EarmJIiQNJ6Nqxf0iBS1iD5NLHkdCO3x6Cs8K
2q29HXx3KHG+6t4saQegYQ/w8hbtT4Uxnz78KaPmPj9XyrRd9O7kGTe2/ivCqWpQa9dvQ55FgIw7
uudLY+fe+a/7xnBHw8BZ1rlR/gyzU+85GVU0Qo8F/Jddq7oLfgPQ2Q5bqJMKo/EdUxVZl5686J2i
25VyTZYpfiwKL0StkooRhxvpnFKJ4kz1OP0uGrMUJfEbOT44vKXQk9gznbazKHAD5GbXlYydRte3
aqXtoRSdEmhhevWjpQ7rRSjW/xrghfF4fiYhKMddh0e0kUMex6TMriBDsuu/G9imRSJdC0bD6mlA
GGnIYG+htgGfKrAgumprue17/TZDzcCKRD2RuApSKaL8CYzTudRos2bXqS36ddXzxxTkC6EYhA7K
rvlGlWyqlP8jvtFZQr1+44aQb46H0mFSoVxc83+1ndu5savKz5/8Txc7pULr3KclxXueQZoZ8RX6
u72ZI0AuxLjSO15uRjTT68e9lKg6iYw1Lf/nwinNcrzI3Ro+Cn0tA1myJvaIm/6z7fCGvAvdpT3p
wCasPpirWvd24Z/q7mzHiQVaYt2PzPKrjUYx268bmQe2+gcqUMIGn22tAGXo0e6OknsjnL6Yf1G5
XxX3COeIfDGkHDlKsrLXKHf3GynsmgdCOYX8SE/py3Zv1MX9N2z9E9u/WbnIstEhDx2VvZiMInWd
3QeV56q7LGi5K0p80tglGi/ORrZF8u3prhAOTeZBQGvLFU026RIhuUE7MP73uKBokWdktIv53UIo
7k5I9oWGUUjK7yOdzvUgENikwCG+VhXjucFa3a3gntOeXIG3rEKsXCDiy41vQPBINNTPutSWfDCj
/L5Uh/Uf1qioNQZYQzEmC/pnOnTl4Vyz/qiqdba/tWyftRjVAMl6jM87s5CxjbzSc9G8tXfeJ4XX
fHxVFlaKNmtE7m6N9MP9GwMG6K3FKgDLaUe2XJ43k7ADqyChYqX4klNpoOlqOcudEd+rEUTYhTDj
NmSlCKs5DZYRxs3qBR/8nV5nEUlHfJ+7kJFZNftbHMr29+n0pgzHqE6v6pvfVVfgfzxroDQla9ot
GbAJlBLSfJGP3r8eeVjccV6QksyBlPauOTDEvpi6Tfi9X7xYg+wrDyEHE0mAi9OiT6h9KNXHgU6I
N1LxOxGywPDEcvBfHAD65Sm6dF58gHSCyiWD/l44kaS2zT6dHHdkqLffZN376cBuRSdgOHXE0YcV
RxQoEa5sBhZZHJRPRCNeSCiqTY11FRyecHgu1LFXXHzP1l2UFON8HMVecTR95BMnDMulAbeSWc0Y
NCBnUcRmHc80a5wKBlXa9WP/Pk2CqWmQnL7VuX64FmQ8fCWpMggRs3cC/bVNNgK3Svo/YoE/IYJM
Cm4V/E5wITVm+9GKh8y8zqKIdcUKP50ZVsT1qSRXAjmvhaUFfKrSLzWAczwJtTFK5EN2RTVZap/1
IXI1s2/i1dSNFZlEMqEfiUu0e2ERc6ucfCviLR9W4RhWlTOUMZL/yeEDCYwHQM8+2qQCdSa61pFG
oc6VqVdPz9HTNnTdct2K3gHXOVTBNw6K8Cgb8/sNgcKVwlZ0OjgPsvhmhcmdLZ1p99fBelmqxyDi
qhO9PX2CUql0rD9wbXCRYBntQefgg4hUvAqzdauvru0J/ekKposUtoa5MMZ1J0NwPJ7+TSZklala
k5gUuOn5LvW09fbrlLIiVqeZZHVpKWb68Xd+nXpoTllQEmADhi/jSgFoGkJO92wukelrulcFVJOR
uUtH89mXVpzaAvxbxMIBYVGAeK8WkwEsH3SK1uh9n16qoD4qhCmy9AiymijyvktPEitBNs9hWeT8
U6wwD28Pooex2RKSj3qC6VpocWUJNQj2HPVUEuI01/jl8G+NSsZMXGYYWmeQbsjhafXvvu6KM++a
KsKrgGfc+mUtlWjQQE4T8IlW36KNZ5ZZTpqM1fgF9fN5W0OA4BfOrlPrIYK0We+I3XH10wlmgLnv
HVMMrqVlZdACzxXndIGhvYro16AQhRpRLKLaIA/4lj4l1d2aZqyvt4p/5B8tS+h3HzSpwlgtssTm
ybxtC6syw+/bncjirVBGP5BoE7Y0AxZ4WarzcKaJpN/C4mWAoZM28eNRL5V0z6bmTYlfquf/nqYp
secb2DKvh8eN9kiRkxrL4oCtIqNzL5fTVJb1yPrfxqexW5nfz71sTMET6FzPx05RS6lzCE0EoKIh
PYGef4usVC+Dmzgl7od9HsS0l+gnyhI6/V/mAsG7QBRfNFnGYCBbNd2s3bf/1pmLygqHDSTCQd4n
3psqD+OiE7XzWzmbRodjcjHNoL+LQTgIRw/NkrpVf7Jzwb/aAb1pIKczRopuOztFPSOXmv4ms/K0
FdqZe8IK401DLjUYc/ccVhfK2RSjL0ilSwdEdD//FgBDU5jTPNJ19zCt1m4FzrgSJ1lGk7TCmi7P
Uj2P+bsChGYwQ8XgFMsYBXkr+XSx5LeqyVLXpDzXl2Q/bA3rxHGglOpVEe6xst6KWI8kkwFgHcU+
e+b6S56liAEQIJCVtarSUI5l3uyy7BgE0lhTy+k79WWPphGQU6sVozVl936c9oYm12Z2l55oIVzd
tmCmZXDzm39deZQ6QXjlGgL4tpDP4RxpLAdb0pBuUy1TRYl2ECu9lvKX7Zz7uXv33Y9uLg/qU8np
P0s1sik4ZUlKaQpdOs+SjEMteOpUI/rMjzoeY4THIL5NOlDGHALa1j8lw3nR8MY0J76Ms/Sfkdqx
74IK/xqCujfT9TjGMAp/dUZlzndxQJvHpzlYKl5orzb6eXk7hetpZaZ4RdFNueZ9gfKUZcRZE2gx
GmW5jYO8ibPJlab6xLbvROphYr/dVR8tU2ctY5jXWl2aGzJHc68a6ftweB9pL0peE/a17FJt02tY
b7BLlqpKplL4OzXmAENlFbwHEXOIwrmOFP6K6j4ejSrxuhb0BDChvVUdZzBbbcGrqxS94EGiq31P
0qVfDc+/Lb5lAKyaDAbl7veeJDOYxzZCNza2TChWCkkwqj/6GKkv/lkCRIUk+uySl3BVs/Szh/E2
5DHcp4ZAkaMghcykd+7f5iSuZRIPs7p0zy+U4g6o9Mdk/yTJEp4tRAhnYJIuHsOX0iertqcG02lR
egB0Q8SMLJ6a9xLHBtKD1Gb7Iv5gvOL7sHTZEgzMpXtEtNMh7A1U5D95wpIe+JzahtzR/VNEM0ba
47zd0eJXtgCEoTgQUeFBagFG9qBOWcyxMkBQaYB8jRrIPpCoTWTEIO9oF3vpNKYJWJdc3i9Uruz3
CtfGPhIcn8TVrN1CTh5AUy/pi556VpDQ9twm0lU0yPPzrWvR6k+nGW+YnHSAhHmk2caPqFFtoa7d
9vDIlFewiObcAZYg6LTl9qqEk9lP8J6+beWpIsLMfMEk1PvaDiiM/+604YPqZ2yYWUljByReE9BP
DTU5c0sm0f+FMF4+ia9Cdw7GOCdcE97dG8dqW+ANIn8OtQ8MOJIbTBv4g+8BE93PKOg70A6QPLg8
dtRy+3BwBHe28621zzl7RW23BpQ1PbrGXSUYjmuCxFzkeCsXEXeSeCECC0BVn9HDSn4HjWJ3mtK4
bK1CKawDijg267hW6A5vxIYGEd/seSpkQDwAEHSjGEw77Z9JRYqqLvwJ0vpKLmL4RwWBznn/V/i1
uZmhmrQsEfzDIAZcx5mUsBsWWP2QnQUhpkjsC5h4OX0xeuZlv3/SHYPJeHV6cXq/xDBEMzuoIyaS
nkmIBdfb1ZM3TANvyVUIt0gy46E68BhORq+kYMkFYpSSMappaizCD61UpkJs/rtZycsDJzsW2GrA
rlkCGehwE3rjaP3n9ilSEIm0SxNfdkB20oJS5CpJPgUJhxa4jMyTTeCSXQH+HaHmZq2LlI0/K+T9
/INO2yZk5iMvjKD4mzgcPiRBpqM8kTMq5xuCNuifwE1DvDY+78aiOM17PCI7wf/swEJk3pIYAKDl
uaez/u0a8epiYLeOGJYiJ+0L5e4z0uMJwR/QG0UC+9BbOcz/5Vue0rBKCXyeRN1KLyNjbFNxlgue
s0rHRtGZPyeI44a7tUWRQtXVfWXnv9LB/Ipcadt2pqnyP26OrDlD9jnMg+xKJAefHyf2hm6qIcat
5Ufe/QnHaMgPYuRrmWjVBPuDvnJOoxyFovhTKzOnvQguFgZix68REdVcYb+4XEu8IYpRfPf/bTyg
7sES52QO+3Zj6KrITVbTLtlZn3k27fAkIKZ1VP4rGqYLmKurnwnmVhVZEKM/e5U3VfKstjNkjLT8
WSnb5AizGoqkbJF5HebP+H/i73+gbGWDlyHeFnSNUDq9wxO0rSEFvAYXSy2WiI+zDm5tt7yhOoQh
hdphDSJ6W2CKk8bbfDxw5KZqQwEvCzjvOf831hiHD220EAYJW5QMJq/w4NxMYj+DM76b4tN71iQZ
IZTW9QuPAsxxQIBB53Ha45bQCns09bjLrXT1Q90IVuIiH6dMANQg6vn6kIkG1IvaUsoih8ri7sMq
MvBEzfAEU8wsPBsgLXGNrci+3SGJ4+/oCTvCgCM5rWl7k70iA1WCFvsPLax1HBXIkGTnTVr1o4B+
1gsQ7K31Yh6hgxnWPOQlabofBPj7e6sATBp9Td29AWrqrMTGj2LKfC1k26fsVnsoqwNSvu+RcFva
kx3bD8i5g1By7DOdZtD2GSt4y4FHZ/7WMlyg2xFddxEWIpc4tlWE+rT/XN9TRlxVXsO1UUaN8nNl
zXYS/0k7KZ0UAwiYzYa1C6zYOZct0bmy9ewpXaTz39DTKgB6rbuxD9ii0n8oqXEA3RPIDsf5JWKD
SLLajmZJPlsG9uIXJKma/j2TtQ6P3HnVEo88jf2Pbb3KjDgzT1snWqJdGWSFUeMJXDxkXVr8o56x
UNLyqoKS6BknIL7KNQ+C71wITPHUQArKXqUruvB1hJn6u4Zno8LRzM1RVhWCfBPtVqWJDMeqmnms
Y/jJYTmBDCta90DlL0J2OnhPTvv3RAxG8FMV72Hfmqkdr0/Wt8uWtwebc72VziVGH2ULCnLI16QO
wtSk89r1oS6j/+HO89mf55TkuszQ+03Wgyen/5+N5WhT59yKCDkR94CzPfV8YQTG9QICk4bw/80Z
1abJyrwtqiuSP+w1Bnz1aMm/C5soOp27gFi/ex4u7jYOQYA9x6Wy3LstKMRgn7ti/sHcs+0z5izh
FOJfRjzdiMamBwl880NTyWfyv256pgvE28eh9V9FrsmOcvze4m4gLCjI8me826vr6MMcNNdx6phD
Sb7018Ls7/IvBrpst/WRvl7C5QRycqjDJe0BDdbWX5I37oo7AR6/FVEjweweRLZTlOMqthtLszBg
10hEDXnaMmrRSpGSEPHALmyUvpmUQponWuGjUib1yPWOtPnzvCW+vjGopd/zjsz2sFW9C9KJsjuD
yweU0OEE10mUJGx/YVvBoBu9EPJkjbzDc6biYx/mtcqQ7uMrNUaGkvRCygjBGo7PxxNzK2cO53N3
yCfUs6aIrlE+eskZ9+I6WL3rymXLCeJ51lpJybh3Tw8T162h5BT0RgNn5wIXChr8FTLg+amAlDYZ
WoVUhndiAah9Apcir44B+u0kDP99p1LDTwnA3HN96DSJdYlDSU4PMPJawC7qpDVEczlxxFo/i+Q7
9/MaC+XRo+svcsGU+ZTIMiO4YDYtZt3ht/AouvGUafK5gywQJBdWAVrUKKXjHSankfKhDd6012a5
QoudAE/B15btq119G3mAC9gA4N1eYzttnZyriIXZ2Pu5lNQoxeiKuJK89BsQ6ihnpiATpXoZbrYl
2KBoDSM4fGNUaEHMAnj5DbZTpEunZRXxAYytbzBV3UxixQOOE+QsuDBF8Em2ivDGsZdNKjj4Zhak
Qi9iQSydGg9FGZghllVOlTTZEUlNyt9IUzMdkznqosUBZi1q6oE2ogp39JPIc82TohLdaROOAsqO
TDognTZa2x6gRC8DyPncGFNCtflisey1Qfo9lcGi4iKmDjf6CtbJ34Kz/WgbY9eKydd5KEuVAbYo
bh2ZwNNdXvg6GIEYgJLZsqGeNuJ7Kln53/yNHdmplKXs7Vt8jLIXDqdYb6Jj1m7Ijj46YQQuCpX1
TvBkRjJVUNleu6KN0DvGiAPJyMDTqJSg5TvRzxiCtJ6gDxT592+mFxZkVfeBtHBQdSvL4o/u0qf4
IhPuv0FUw4knoilD8KjIGg2aVM7Uw3FnzkTKwqJef2XR6QijKEP8PiA6e69bsKWQmuI33JoT0Wcs
hxxd+fBxRUWg3JvH9vmwhVEhEmFNxAdukbsSJef02EsIMFaccqqGc1Y6b3A/C4A0tUL6YSMhUwG9
JYfmXIWyk2LIaLg6WK3PP5pXoEtu91qVjBvsIzuXyhX7wWRCuFPMaJMRfpPXRHM3gI6+09cALpMA
a40X3a+Xqk1vfwhVlVlsl06cHCfRiYpQd3zgvXMGMfysZreahpilqlofaNA3CwuN4jJr8D3nA8H7
tIzmIuEIha8XCqjkgysols8p8uzgcGr4cqwf8DzWHVRV4nl8HuqiWVcHSlWkB7qEu3Zx6xZwknV5
exOuWaehZvTOVcxb8JHJy324T+WOy187pvdGjbSocUXyDQe1i0390MEORLPkyc+YXmUb1GXZJOVN
YKsS0LcSXXkhBKVosfKsA4+umYiUAq6cyldOuhk5vZtkMAaa2r1IjbCjhMz5xe+ed42VdFZt9AVR
VpL1VD1UJbUQlgWK/MhVFFM8bjw4DUGeWUz5MmxFCXe6UPvl4DkV0z8o9njGeaq3AxU7bXBtSvnu
Ul7elF8lWNMXU5DIh4Wx+AMr0tH5UurTWSHgI4nIvAy6VYBwTEwsIQjxNfuyizylD6vIJzjhKPSt
i5VrXv1g+ivcsr04w9ROFQAbK8YHorH0QXMJyqHGGuh01s13EFzvyxZj8tk4qwat0z4Rtm2dIV8+
Lvv2dCzLFUORx03Rldj0MwumDYv8iarEj6fKSUD3eEavRDdsvMGe7rblAzpjKMPw0qZONWJ+hgcX
52ss47R3cHynBpBxWkEuDnP3mZjDWakHgVCkvq7lZsGf8PLD7ox1TK+D+iNRy4kIikhpOqKNCr0j
s6ar7nGkzWUJp3NkYiK2x9e7EiKbJOqD66ojlrAo+4kKnH2AIsTFKB9kAo1XNPCsdQqcH7NjeTqX
VTurFFb5d0EabcRDr8ByZ8m3v9oqeCGUpCWegmpo3j6551tWMO5TE5eoOinqtP79DTntqzVtn+dI
PIXhITpuJbqC/e7HqvYCj0JxbMnQ5fqUlw0k/p35A62ZX26ur2l0a2RnadBYTFeKhpamXJu288nT
AZd6lSwbKbPInsAn0k1Hz5ez+4GnbZl7gLXTp2FIIeeD2eGmAboSu3Q3Ijc6B1rAu2EFc+wajBpx
2IhFp9Ea+fi9RltyB0ZtS3+OJApEvOHk9vjR2k71uu+KBrI/RxiWcOmLLGR3u0aUB4+YxpeaKVer
dNWjO1DB/sMSWy8Qpo1fqBwHYuBn87SIGQ9KRQK5xfNFVYCarjGLiU8/SSQ6M2TmgrPCDbExAgfS
4aIDhb0H2pZM//aUhFnr5CeMwiQudEO+4yAi+z4NLkZwDpBoOtMLHU6i7nWYfExM7Pd03C5dfv+x
Km4fNasHEtWe58kgk3pe9BQQ+yChHljifkTRLYLl03or2P+gK9cX0hczzKmcT3gT/6zC7tdpSvPl
L6s32h3zIhk+NGLo4Hsv5yPz3oY9uOQpPfhmwPZ7VwII6d2YmO192RSCnBtdbvtqCfe4CvAlXPRr
+ZFq3c4tO5Vjo8SsjC00SIQcIA9gyKpSy29ZgArF+/ZaH2JQxLW6tRKuGLLKkWp/iUwzGYFq/dno
o//LKkg9k4ovkHJo7Gsj25F1Rq8hPGbN/QrVL0JHlZevMpOhUY0l8I3GIAxwCeiNs5ts2+XyHGJL
6/2S/qn6LN9oz8F2ADNRetzi/A1zFiWgf51ptxVOYTCwiCIZO7SeBS1Pwr9FBRFL0VSCGxh15+xY
rTwM8H4oA9K96tYgvBprSscuR6tmXeFabM/4os+yolYkNR8IyJZ76swpX2z4t2SVw/m0ChApKHB3
wMpajKB1qSSWvWCffetlxq4ho19b/qx9CKmTFQ4oG8DSBmQz+cYT8BLscAaD7dZ7nqtQIU2yAKc7
WjcuLiPqrXB/qz54bY7aTwJnRSYHmStkGb86qkt0zebDJtzM81YB7xex7nYOPMcpB3i93VtkEpWw
rCE8cjStdIEiqjGWJ+4AdWVATIzdBUJp1Q4HVgPV7s+KnKBptbpkSBmr3tmXtRi7thK36z2MON0b
Sa01NY37iSNG9Z79u2AxKVvVN+W2kQA0deNGfJQY5GmZ/KslTRMokVF3k5clgFuqU8lcZwHecE7R
GORdlLWPsQA/Y1bFttdiH8l/dbqkBM2sKQ23nuH7JBaSqgSucpJQcrO3hKbBll7LvgXikG+FTd2N
zhkcikVOVZP5tjPCSCsxKDQkbvXTQw+DvcpbiEmSoS3gFwIXK+FM5Qcte4cabIOcXaMhOuQhfdW0
VZ00kSppMqqUOJSanWJfBRhO8Xv/y7TyZPc02wQwej+bI5RMZ9cynL6oHdUIxuquqPZjYp5e1f4U
yNx/nQIwY/iFhXPJLdS33jjeeuhieDLPabqk5n0vEv2HWGWn884dhfYp8mXElMuc+ThZcTlNWjAU
qezA6WNZDv7vG/FX09SRbuMWV+Hr27OxJzPa3JkrQvBUtwqPpqfFS9rleUsAqr1trhWsd7McrFLG
IbgubKSwF4UjlfD8a1iegbX2ALbDI323QmILUr52Oc0E50KDQjXe6PTPWjDTLelNAltFPyXNbwP0
sdeBsShO1z9TokI95lb8nbmczORxjDHKIDItDfOk5+M351aN1KiuvPeZjrBUMwXDgi3vYh5NMaF6
ulfYYSLkt/xJTPO7373NOgBWEIze54lv3I07qW47WDtBpxcYo8aTTHkCfBnMelRXpW3JSHxCLKwH
qw495RtWLWklNhlUn4kQsztNo6AE1c38K7gCUbdxGO+6mqlXzzWYWvLeH2B0rvJMYs4Zb/44u52b
wuyM+LlwG914DK+2xkW/x+gWi/lzQR0stOZrsGP5BcddWzzqweHm4zmgelifv+8f3hgPsgnUjQWh
QPckPWJWDO7yrY4ILGCZGsmupRWgIqDQbN9sgYhJSVbNL7iqcNRckm/UFHzipRJwlsofqt3gACGD
7kjaQToaxDHPhXQ4YsWOiDAdBGuqsO3G/AvUgyc4X0WgB+pL/r3Rsr9qw/fLVkpUtV1blfOl3ija
PCk5GrzX41Af1ddvlEYYfJsW8uVY//roiEA0ug6/HYAxBVl5O3Lvk55biVdx8Mr9ZVmW3iTyTnlx
IcykY2tw8MA6oYuEfUYg6qAJFX/GwdZL4ltDPmpC71YTeeRBKT/qqopt6r3JH3feD7Y4lhXConix
I2p+jxPlQ37+U7wCgI9NRezDz2qI+AfYz2MK9D5LQkPiIjfPo/7+RLkYAT+FARpwwAlMyyMFsIbC
c0/Dbqz91io/Gs4etEkpZaH38gzTFEoBoJQviW0SNHZYDmHKIZWWyEkn8O9+M7qD6QpwX9KS8a/5
3euWwKONrK9Cp6LTt6tyHlre3HVUG2V5DloowAL6ZriVfuDXENy3SK64qfYNFYHGl8fQoFdVm4Mg
qwu9xcDjwLb5OyswAs7Yq+4zZwnf093RRHHn0lJQlcCUGhcnxJcu6nzEeKThd7N8AXPnh3yfugLa
VsMjZ4uWq8fXM5fg8f4/d5axTW7RA2+2S/DZQEKe9dv8CY7xGxS7U58blGNB3l4Pib0jxgRCZGgm
jDvx4Crv36MFYKfl8xxURLTnafVayRtOKwINS6oEmBL5hC50yuDU/DNc6pw7WQraX4XducNsByuO
+4OZpGOxdmDnRINizAVWifQcidUBnkpEBmrCmYjRu34yBh50myLg7tfbZJcho8OoJgrccaaf0x8C
woeNaJKotsCHnENgLqdcmEsynyYM5nK5pLAQ9AOq44Sdp3y2GSqsEQtk25/TgVBLZOCCTEnwINGA
qCtwJrH1mAL9OsHCzK4nYwMUnvzhYC+brZcNwoTFEp2MiQGnw0+wSY404Bps4ClEMIFROqN4XcFG
uH3LElES798Gdi+AxTVDbeZw7lU510zeF5nCo6KcdUAwdTbFm/fPRVLZ4BfznJ2uJ8GOHwANiZmE
yn1gRxccW9NSTHUrRkOFJjTKcG1PDH+yFQc6yAMWxZpu5nIUhw40cZ8BWY8cjxi4UFs51NBtqj8C
DPkzD+49IK0buHWDou2KaUSxpL/fvb4JIOQkOYtwj+h/J+VeR2ptolE0JaKxPq5pDs49WF95IKzg
ElHLA4z91HcXLg0QnmDF+AoDNsXFnNIjFaLgjaEEcvZgfSJYWxBUmzVD7QW4uxzm/0SkE58esCbC
DwvW4O1LQ+2YdOpH+1aTyoS6wj+mEXR/jDHwWY08o7YzH/rNb0WzmBLcwg4aVviyjBp2jKar3h3v
vBOJ2zuMftjfx2bmGSUH7JFe5xetONoG4fCrMfNh6THKmVL3yEajYoScnmWFWBu1HGkSTEY+dHO0
eKeI/WiOeFfM+NVbAvKhDihE3C+zwsLLI5iYs3xU60zvaCP8JNrS2E4qPHSH3aNshgZfkpox1h8Q
30BZ8O1QwvPYMv5qMRmEGLy/KiCEV4tHRNVuTq2wqKnwOiGgvVuoeaS+jY1n/gzGb8TSxw0ggRqM
pl4Fqb92Hj8c7abSk1/TqJaB0tgtrlHTiVVSyx8jZYVT6tcmCnrdqXHqS1HqBzlHwppHmjW8uSDD
bTMs9RUkIHWDGPb7u4Y9gLS4TrorbJ3YsODd0gZ//v3qA2rG4ZO+J2Y4xLgEq1gMvh4QP+n7KU3A
WKrIfjRIziQctELffvJAUXCP402MehikWl9eW3cJQYdvk10B44SY+9G8+FOppcM+WDDdADGe41t3
YILpKRCGzixlnU2w9YlPWwhVy3vrCbt7O4THsh0SX/EhNTcHme5F0f6BnSgw+bfS6r0i3rpCa/Ac
MzcYGu5AKYT8WUD6B5v600isJNx9CJeH3+UIgMJ9M6LcFNbbglIvkY6CZ9DYD3pZgQzPAXXzNKN/
O4fgbf6/iKa71k2dgiyimcVPkbPAFRwIVsb4owv0aso8oNNTGh+C8LTyBWeJBsN6a/gF9DMQipBq
xZn1P3bqwrAlWseUJY8Xsx1JQ5Vm/rznG0BmezLpZtp9p5c7jsibakqv02NxWL2/qD9Brs7OUcE5
Ndm9FE32/LfOMexaJtHUgha1Z/LzJ7U3nRITgJ9q5GoURzw/BPAWfJJorzBZYUtYDUq7it2CdYti
NoGIhU+iiS03WvAEewLHc6WwhE8PG1VjgOomEVr3ikY32d85lWlQhcJGufpqTE0U2sbnsZUWGdBm
4xMFOMIhRfvcDhPAcx3V+yZE048E3zFbkPKyP7/035lnlGo2/aLR1PQGDqFEQRTRhllMwPERCbVA
CE6Z+kyX3D02lHLrHs+8xOPiC6QkqLU0LH3kqrGZHDc3LaSlFlv1gKw76qWfdOY+YvgG52Z+jPEu
KOC8wPVmX+TgqwyveSukrhtvYWcR6l41ls4GYCinWnPYDKeo1Qdd+nUh9kET63H9QhNaJbpxjExE
XfgF4E2/Vj9nSp5Q+SZ0OVMHYoQKeVURA5ZtOWpAKsfHzVwvJHuLYbZ5hHoKgmFrrg1Pi9aDi6cb
cO4zrV8vSPr8gR5RKuLBar/cULaATSpD+E802ifIVXBBR5BdnWtduDW6Za/pRghRSEQwt8bsrRbg
Iq2SBNnpVsUTkwn3p/wOUDXyy90ZemX27nKyivxl6PO/Br+Nqcfi1NCGGRSqznE4ARr3uMO+K3CM
rxbnvceVOZSlQ18WD3sOmnrC/YiJFYa6MdpxJ2Q5FOZBnt2VFVlOdFIcnwGSjCafYe21RAZMzblF
FBMYNttBOe1ZdhaBktXiG5mTAo+eAfH2nJa8F+JZVGxdYAxANdsGF0GMPFLUmI+P4loR4uFBcoba
aKMskq755qpDOqb+BYJJy5fKQTpg42cqu7HN9ISIBfzRO2gZTBfZY17vPcgKkp1hkFSlcVD2G7t9
HQ+CqDyaHROy71nNOqWMhoiDjqPrvGU50bqLXYB6oxC6JrpezUWZCLWvnVDcMNGGyeu0o9tQN3Iy
v76zy/gqSU9NSYVQhKMkrkA84azGSQxEhjOT2s8EjxOdAx4RebXR6PcWkp5PXjBVPq0RtYa5PXgI
DoEZM0H2jox8MXgFrooijcOo4qm5q8Nbu9IT/O1p3m+6WME/snVAy3Bjmx4gV0q9geoWqAVsZhYD
r0R/qYfXlXacMKAZ5jlkLZ+VVGvVebr0IcA8DDrku95Ll0W7n/SeuY10ShoH6xMpotH/b7XYYUny
leShab03lzq21ntJ7+YHrZExYmjOcs5KG/qcYm6CMmqcnU8F3YzumJ3k20XsOgQ3e+aobZNbxAU9
HgRu/sFmaZcmfq79BCMnRlMtHQm6V1pK8kFyXP3PMhZOqYVWfdvm+C0LbsVgPREZF5JGJ7JDICzZ
oWjxZW6fb+yNf9H6dVWywXbYSVISbgHEmAtSRUZ89Qgj3dN9RFKwfvuszmv3j5RbEPaF83wWa8Td
RnrfaDncOiftmo1dm+EReokaYLx1uU0n8zHUQ7vWZTgGwl55od5jNnDE0NeSFar9ElxEHSYslmZy
OOcY6tUg5+3sLeWvGOJqIoPodq8kgEwRr9Hjn1Bu3tWWwuFx1i/1n2hAWheGpbTSc+FAFL6AoI8Q
2czW9sWYpQoTATZdMIBW79IHswDrmNkTaQVeXDtO65JD5IJzmMYuj8gjnAf8EIg8a7ZgMb0WFHs6
x3cCLJ9E2GD3LiflUDSd5ZrUqLn7+eHkrFnnLQr0r7lX+IvmHdD/eBqGFvgevyqaSjXPN7kodejQ
EUrve3CJzu7UOC1bcej7UnxDaYC3SPfzjXkh/ZYR9T7Zcn6DxJzFSfW8IAwj7Rp9c0QWNUZ75rVp
Kd/8iD1AV74m5LkkahmQvZEg3Z8RcM8HSXtQM7HYFyhG/QidUjP+vXeNRkb0J9/wi2dC8sVE9NoB
9cc8I5yuH1t8jeJ4iTB33sAgQ+Xmd7SAWnVAZ9f8wjlpuJfOWhaApxubO+za5Lx1WbMygt+RiiJs
GGd0Eej01dnOfu9y8hs46URQSIxGRg9x33k6OELOF5a0S2WjA9s4eYhrsuuGM5twNTEdN/08Cs4t
F6MmoHEsHsG2kmg75SSmm2VCNO8iW+x+loqqN/dDntjMc9CKWHMQtWG+xL/q1PoYaON/Nf4OYEC1
gqy/vkY1yW2g2/3LjJhCkGzbjZTbbAYhJrWMf77EDknzCK4CHgT7al3KW0cPdzWhiET6nFZOt4h5
YtqhyapIErJdqEN1kgQk3KP/tkABB+FVLdu98c+gWsYLbM432STABQB+KHxK3TLVdcO3OOnjffNF
dRKz1yhAHnjx9Wp2IBGphfJei7Vqf0gn9weyTWT7PRYzB/igcvZ31nPJnCcKnYjC3uH7aZoLw6vU
ob489NXOHqaI5Ug4/oZQjuV+p/d6xoqnuUAr45kFtomCMYHezQWot3cPXRzntAg2r3Y35axMjge1
kNKYegFncPgtB/1E2bSAHylANk45DlRMVIJFnYFLSTzy93J/HAn82jbkj7VGKZNFgggLBKEW2B9j
RYswb2LL8+kAAUZruEvSuE1/0F7xfD8QzXGBdGCw+Fu2tjQHJ6lwW6Q/J2tU0TFk9P6b6fb3ow6q
+JE8N0PUBOGytW8D3RL3wFc8YFaQYHRX6r8+xXxTp/eDq1ohxNjzg/z2gTSf3h337fmNH9qILyo8
mqg71EwDPZVuO7PAxpoJlVpPt9d1/d5DoCBgaBC6voyseZ2WEFggvN2w4Ajv4xIr4s17gASQ/afO
2Q35uzxmMEN45lKzmQ7HtqLfv+486lVTqlEOl9PdHLHM0y3v/YdFZcxlspmKdJjCQOQfvEhtkszZ
uvQfh3qQvexZWsTeJsMV73tCx81LxeUxFYLmVu8eI8BBpsSLPIeZydc8yyH9pNVqcqxHFka6ltoz
IUB7ll+KYmzGI3rSsKHpeTIXeBC4GgC+0sDZMFL1sKKNIY71Bzajfch8pHaMOporq0Iv1GSLdtEn
BLVEq1C4r2CAnYl2bQE33IpF/KiDpEJPB20BLAkTNMDlmtt5BorOtZvjqN/YZs2CJHCkjfJaw9hJ
DzvYyTh03MWRP3pKvlcEQ7aiuIqiFfr+xfeQkLuIs1jQmBLVBzkFxYn/QqylpLemHDO7DwCI7yQt
dXpf5qm1oEXfYWed4ML0jJNoM1pzsGmnWtZ+QJjDAcz0Bsih/icVH0DyS7hJYZHq7VRxy36Nem7Y
o4VBLq/bk/SwZqOXTdsDhHoGtpcHKDu557enXxXLjtBkmG2QsA5kwE3s3YCBsPYXSHAjROrwf/jL
S3qgV07iebg1apceC2kLVTfhOy7mNFb8plXitKnYvtAyJaK8QkECzGPyp2a4U70pO8JvqFmXfMp3
35/tonc/zirPs4m+QjfiCVH6emN86ZRqQrlIyPz1q11FC/3Xl/2uVKgyXzRECS5+oiXkS5Zhlwo/
6f2O9mFUK1afdkSoaTaNxtfkHOJbW22QKSi7dJQ9M/wfGd+lynCeFIQ3iHx3ajQgGdncwz9UgVEH
bBdDmgxFXlj7MQBNwP4tYItvs+khOEU3XI1szolCZ5unfiihiMrfnOXWgeicEdt/IhfEBInwVn/k
5WGVRJjXKIVVNcBDRxfQaHWgliYyoL9bpS4FshAHCxc+8vNC+ejSzxzQZXRYcE9erHnX8bsifDkT
JsUqSzum+DBPLSN2/eKaqN24Rr5cQfF4nwfb2Nw3FoeHZ0VbGKt11bZOPbUyIbBmL6qTTTrFaPuX
Wpd5bC3BETt8JQAZlvNXrGu4+ab+DRy8uxPT6cL9jiOg4myH9sc3dvjUx6mK8K13t8IAu3OAJKxH
jDndRQkblmPBVUSiZcEMyrJVJRe6tNOf+ULUYfij/9ReEdY7BOkjTodAyBMWxnrQhgqvWBW2zLrA
u11Puu4aYiw3zvxrsPglIbAlAnMBVnyCWv35/hXVuINU7IMtqUUdlKScmT5T97FCgxkGiPoaUhal
oBVDFLbq3aYHp8bzqpIXsjETqzVrEuGhxru2VxDu0qM/6YMGg270/sikj/Nx3GUSkHxcJ+QvJBJw
ghF71r2P3Gy5QECrgMwhFyOLk7LT8tFA0VN2oSWf4pHPRmnKktYhULNe0LFaSCk7an+F6lABJ1SV
6dBPyOGewxEa5heDsHVx0uBISaSxyV2bSpB3E05nNYGlTexTg2JSqcCtGyY/IRFl9epjqUzwXadA
PrZqrnMhx5gNBokHD0Yl55E8Edt+2eFZ+yj43zsfvv2F198B4P0n2AyJtY/FLihHLKpcvxWwt4Uc
Nnj1RFjTt15GuVjHMamWBIpuFDyO4fg1ZJveoBpRHP7QwZeTZPo8RZZ6sb09OxDNntbPQUdpLcey
XgCKCSsQUju2JV7FNzMMlgmeQbX0Jn3xs6u51zAGFA5YWOhYVD0+RFDxqRW/4Zl9+IdkYFgitygn
12db3E9t+o0V1uBzqVw/rgyD/YKR79ZJ7tnqriqPrDNEP8pFRbePcS41Abcr66jxxJDklpAlDyYc
Dm0mi00OZCPeIizT9wU6fdHfe7A+TOB2K5C7Vv689iKLFS6wjGBH4TbajNKqkV0hMlwIAsvIVr4s
IXHbtfrUJAasZT0CZrrl/zDp+EG9XfNLOkgw6k9Cd4t+ceLSuc5WMLFqwW4WCegbTcpCOtoIjju4
ofJDhAC+oupCqLyaLYWP7OpJJrFBjqPG5HpP7XPl9BobhVAt/8fq6DGg6cQa2yn/d8AeN5hRAQkc
0Z9thamk5UBIsURug8HzB3pHUIS+ki2sc0/MeUVVXkX/GslKQTiGDF/7Kxf5y9jxmkR3KWgyu6mh
dlSgAX7lIJdIBvApUu0dzORj53qiB7ThN0at5l2FJNkUz08XFqwctFuFLYOlinQZ6LbYZeIqFEyd
98vycMPPAb1+E8/qQnFVny6JEWrnmd/yT8FoHQ+nfL2W/c63NC9ZOIReh37nBdHDoniJ0u6oCHiH
gE+jYbnsnF9TDJMYltt6Bm6tX0lSeRCHd061NWiGtnD4ksfH/yxh/K5GZUfp2RDieE2bF3ghuwtw
Q6IY11IeuF6dAd7X3+1QNUTpDEck1m5KVEx93kAeapMgASC2t5D2nWzHdfgmhrvyxquzNHTzUOeI
FoXzNU2+wnl4SGbT9tifwhqn1ZI7Xuk3I0/s1lRmYSYhJcEpAjU6zIeCAnAuTmC6ECMuYkkdjH1e
mbnqROLoxiyGd+MyzRdaxc6kiaLKuB7nX/HbE5TcCc6wZldXwqIXu15pjxJStRlheESRtQdaO1JW
oXWZEgXjjpc+JZLdp8yx42gtSQMH99xcw3th4vOkjGamIWNOvYjyRr4xYOhy1FxH+lchUw+yz2t1
9tV330qhctictppgltFJiNQQ33kAcqhtVmT1I0lYiGUNc788kZWqhED0qz6pRrgJtXHiIsj97VIv
MRPhwXXn80lO2XhuLN352nzp05URqXEt4KKY8cKlVgTYY/3aghz3WweqWJw5G1c3ajPDDv10mAUP
aRB4gHPEFWK9R9JDiMBZ7TfGRsY815iwL2gcMjMSNdfYgpoehjNaEGktFxVqRr5Rug+OKIzIGTQC
z+JV+wOxg75Ytc89CuDQt6dzdPISTiR13zXasMVF12MHDCFNQ8mpHcFTeGYxGpl/U51/7S5QnahT
T8noaf0YWkYdMFuclfhnXQVu8gU17wQK5yz9RB76SNuh2nnMkY/DKfkc0WCjmtUYiVwpxAF91S96
J4Qddoq9i+EsekEVlhS8y70csQ3N9Fo7OZnSnfidVAyPxVAnJKqaeBHCIWjbPJr8u5xASHlHJRdt
4nkXWl+owaIYOELBbqvlfwkXj66m9DDv0k7indThmS14lJSNXiHU517ZunQzIAayQ3VC3KZQ38ym
dJgKMsG9bNV730+WBIxCyMdTfJaOX6dRsD1lGvZJH4vO5YRIsZeO84+xEqWxsywM+sbRBGfe/I+h
0xg6TAsbUrci/Snb3ZcDrJHsKWgkI4yqNXXM+ku1RiOi5Qr3mheOp8Iply1cl4MkDbGOLKYMiCdW
uDg4yOO0koyxag7WsySZxjvs82go7ELTCS+WgUzUUblPL1xsYEdwO5rF/Dsbi88/pGAATXr+4SnS
6yvaVQ90LD/Of6RyHo0reVWmPy7hiLRkZ+sY301gDr5mfHVCDqzLOamfMA9/GN6ekfTiDeuysqQJ
QdKDMxGOVXpJ+TbJPUvFxuwKAQY7A70dACTCi00Fowf/5/KxX3pcW3mXSRy/X4O32EZ++0fjuQGa
sOndMNHoDvDSVsLAX1hKqumCk0mME3dQKLzxvgY/I9sUiGDQD+QsYMKc5KWpGc2lFK2qVeqjA9sM
KhBy0y7NPI9WLEbTdWdUlkh7s1VqTzuLLDZho25FetiwVMuHuTGUjfxzWJSU9XePYJuJaD/RtGxD
hg8412+06tABl8OEV5AQ48mkcFUOPzbzLONJ/5wQo3cJrDM5kJsq5tf+Ryqs0OCpF6zrcJvquXBP
RoIj7vvEMkF+5qJW6DO61wcGq/LikC6HeUDTydK5YkewEMu7hURNvKZW0+TYoei8rCzRKGZMp6Ii
vzejBW0Gc7WMTo1xn3IzqG77ActYHns8iTHLKPu79bCdBYJsZSsrJFWduwYTOVWC2RmhM2rp282L
TLu43QyIyf+P2d2ARaOK5E0Ve+R2qw1SBNsUALm9qoR+rCmdffv/plssZJbyS/PnTgRoq4DxxYHs
6X5Ge71zeO2139tNgwsvIN5waoub6v2Xb9HY4Mhgsli2LAHc3CGleeFyEODrXoP069NqdtzY5AMv
yws2l9jEIJdHgGlcGVPFPCvLysvGWy9xUB3WzX2gzsHM7jD+4R04yCKyQIrHJJhQVX7QJU83Ofzy
IqAktk/InNXYFGrxh36uzGUJYeTSvGgqH1sMxUitKCgHX3+3RMtfrJSrJ9LmECX1J7Zw6ZA0FP9Q
zYZNjq894k/tn2ud1/x06XivtaFscQu34om59XI9pYaK+s2TyIuEXH0sVpPTgj+bBWMl0Rc2LzqX
01kPkOV6YWLkQ5zxc2Cyu7es9IgQ7PhVTUzuRxH0KQe2NKxyvYFNi5RCrJM7d+idrQvEGwAZGU3n
lrDH2qSvAVWM2xfYhpYR9XxyYzCZQth67VqlihVmneGAgLRxTPctH3LwlVjgJlsqZmrmp6MoTaNx
QNLxmrxBwwZy/MD4U6rjnkT1sKM/igmqjuegNds/JP8IzgB4uzhXl8dwqOSOcoRnaDy7J6xdGIyX
a6OUXmUAVPd2I2kpXECqHYLGs6j73NoWn5PsQwNnZ+aZoIjTkI4SEzVjxb/yBlE8BkQIHxTNWb8O
UMl3W7tou2QkxPDtN9/7pLfVA51+HlwJgyMrwLreCwOrOQmWADKAtSVqb++u9aL7Hr24wfiFXEj/
/YEs2AynAZbxFXXbPrR0mjLZpfR780bO+lL62TgO+/8mhsXDZ0kfG8l2x7EuMIHuU5Lm9SGGiBBH
wQVZ8jznoIawm/hpKnCm1z530zBKMP4s3e8ynOwEpKTwFY3U69HN9MX9AMGxqU2zswu6jEtZTJcv
xfQgSG2LOXUXux3um7d1XHgkXesae8lPysCI0/qsnwtJWrCXZXgQKR1lHS69t+YqPY3X3LX4Wk4r
wAUwgZxsUeWGHv6h/9z1qDMLbvFlv1mtm286OL4AQe7Xr3LJbwyVIHYJCTDJhK0AHJr0vl3QwOoR
rz4RfXpJQLlBa+pGhjSbFbPwn4ObUnkkTjfD1W3F3WfYlkEJagYfBcOMe4Aa9RJ2s1wUr0zx2/52
Yi/YwKifB7KVXX+g/eIBqmJzpNYyxImEBIVlOi4wnBIXvD3aIx4vnX/IPBfxDcpv+ulqORI3NkFa
pvEseys7XAD2zw58ZNkyq2sz3WIbHik0lCnlv40l2yiT8sAT5yRKLZ6Twimprh6awCBOv0ObkaUe
OGl5Rg/vhnnO4ZDW5n8t8fXCf/c1SukXU+YGRrkmLW2jKD1jEFBfuZgEvgP6Q8KtESV0ITPzDfmd
GHQCiYaHgfycoVK1IzKTRGGQWNEiiq2+x27rOItVQawNSLP6i2INCmD0wTGiDM2FjmmF6KYxS6k0
6HFkTkhmb2TYGDX+xrxllia3JYGgPJ1IA1PePgQIsKie2qxiKNyKEVavRsm+0AfxAi/ojZhzAcKn
O0QPT9Ms6veCTXQjZPi7zMw6LC3ThCOObBNQgdyrVBwy7q8JInXuazHruQFZYW3I6pJxYPYPHXNz
K3F1Wjg4B2u/BQIeqjUz64HTeGGK7r8AXxHsdr56afbVoJ9dkMGWZ1Fd6bpkPbAbEWHTNzuHfNqJ
2evzjS6cftY7TOBHO4e3Yly8FD2py/vzEGmqLAh37fyKGLK1Pwfi3OmObxw84AFALPcWkfTK47Em
J29vy3FgIamIrIM1OESHYt46AkoAvpaNfvnSe9cwYWlCRxy1+bADex6rre0Fng66WqEpbtHxoBPI
T9J87nptDF7VjhHgCsPNpoJ+n0dFxlbPNjuxQopYJuJsOPvBHlS21+Y3vaemdk71DUK3j1jYii55
VhMs44X6LO6OOo8plIiwac6qj/DLctmNXTdOofO04mZHSoExpCMFh1H7DbRScCqS/N7N1Pd4CUcs
Hws6xI+lDr0h8g1VMhKfOz2zDlBhPMs9SgEtgo2oH4g+nswgxTUT4U+8JkuZLcLUH5741uWPM032
GEyZjXO28TNJRgb4eCbefTbSo0AUoxZrTEKsurj/pcrjP/uwu9fVJwdtmO1GNw18tyNOLIsqh4II
MtDmYLk13fh4vwiqymvJ9N0eUFPrzuGTncpRW/wFYjtf1naXZ3oj4DTnZJ3U7Xw0xwrVcR1rpg3F
wtSJsWfPEztuWC6HNqr+2x9BZ9bk1BzV4IDbD8218UVDaulJN0cKDxexJaDm16tpMM4fOOL5coL5
Uq97NRJM4u+8gJ1nxVON30ZAT0Es3TnrOOmrhEaTckTOiVlx+qbPLhgjkcddYVcE1AByNNGasDlG
0Q7UIy9iaMSCV84hXIbHGJtC9SS1UaocLpDTICHes9AMNwGqkn4m42Dx38LuF0Q1uuEkPQF5peoI
DVmt1yTF+vSEup+DVUTFaNpDG0srqPCQ5e4vYmjizw2/XmSbli/O1cqiJdCnRgRZldRsGPJUDxST
hKsokoyDHg12Cv9go0QrKSFt+bEWPs/IMBayqa1/nc5x2C30cRfGvzFzgC+uCjr2C9UM6B1CsB4q
Wd6roFCzQtiWLa7AClUR3eAK+tXkvCZdtuuRfkq3LOkbxfAsH5Cg9ONG9BR+CvahyWc7leIO5mw3
8jgDEt+iV4QwXfs4WZRF4KoP8Ysj0sivuVdrilKLDCCFRNIDB5rZKyAHS20/FMBTqIGp2aPnif/J
wFWIUHmDpF05vVDGBPZkoQXmPMH+rDSE6fHBZR1DFlzIQ4Fl8720+RY564kmvsIxyvMVZrYavatM
MpjZvfcbsSx1+z5S0qzom+A7tSVAIKpQ2tvbOw5jNp8yznSMcKYBLfyGKsJ5tEN8BRLDlenHQ0hk
nUYfpHlGe3SjOJBTVtXmYzMyE/ScPTVr2a6wzAonl+LW1Ch9l3VYODpKiA/axDWSVnn4Yc3fnb6G
rM4lLZBNxn5Gk34NDrYPFG6QlIi75txghTAhxQvp0mi0LsS4clkMQFMxPY5h8m7dpg6R4SwMw+yJ
CoZT2MXu3O/xeB94dy/40H8sfmRUmtr8yNOSRdOwcpa/NoQuSGnljshozUdwaVDGMT90918dQV7t
IMiBvomhbM72xflbATag9v4oqEJ4BJTUI356sjr3UxUkJI9R00GzOIbs8eIcG71Imb3OGdd806IN
sD9kWGSrYTXMD/nIqJ1HaHtB8Cj/bK6v+wC7zIKIHo+AbzGtZRSGs6hpJtic3zcnlIWKUPY44OjC
9j3nNgBnKFjbfTWOSI+d1WXHUSsQF/IZ5gGlcXeXo7EyEKA9qn8nAzW/C9gcDEuhXArpka3URMtm
6xGFxl5DqekMQ5WiNc+DqSvrAFW8sMkiOHuvP2n79ki+DFPQZMUfpHlpU/fHAHvB4F3f0/xjICe/
y4caY/gfxY4VhPn10Ob4+/rEL4pLhdE0O4ag0/IqbfMU/hxM7xrIzHkBGhv88nzhkx7rRvt8fCzm
5f6ZfjVFMeX9p0Kobdpxar+4MIbDPvboY2hYF+OrSDduLDNjw3MElHAMRfR99qRsbQWA5THwpb9M
IsDzM4BpIt90Ua/FBPS9vjUYpgL/N9o4VQkxz5MWO1E5NkoWpOWknVX9skNCtZUjOHXwtbLMQHej
Cse0NmPMIzdsNGer5bTkpWHeHC4LCoK/pVx4C39Rph7Xw0AWWX29RRN332RBuZB+Vx0Gc5tD0D2c
6SPO+YyFrBKgxrUO58yeuLbXkJnHH2uzmGlhIdC2bbFusKfWXNhdxRBBmINr3VGUuL/bX0krsJtE
ALooV6475AEgDxL+n6GKEhZ1H/BrHzhqjpUjbUPnWqqvQz4VK88M0vYoo0yUfbTMFIK7Pg48cFTX
O+oJ0MhPbCgSV8RrhqAI9lx5BDZVEWdHfV6cd7sKTr5GUCSNtHmx1+LXkMngYlYPA1t14h2KrvHn
BIcJ0y8fBFJM1hxFHxwdOUq1ynyNW8mFCHa2miUtb1EUM4HUwvi0zEVREFibQN3H9Ewk5INSBIM2
KhslDrMx74XhTm8+UCJ6cwp36LoH+YhXtqGIuHuX43rc7OSVkbCxlyb0Le+M5gLQFTLvpb8c2KsP
kCh9Bdug73VW4ewncxl5ExZDTjqda35ay/Tay9D8uRCjPDgdWGmaD7iqLyy1FiCQOI6Nz5aQxQEN
gqFQpG3wHd7oVsNM9XhOKH4nnJ9fyDW/X+ysAWyubB0ct6NUfBXe5KZUbp05Hx/LmXQicFty12z2
2/188K1H8n864nWiPTRKPq90BIym6WuUh951+gjp5agsjbj4Tndp6MbIudWnne+bbxQAhtdAjF6J
Tvt48DUiFknEn/6xuiya1Ngyg8139z1s+yXmgCYd2Fh/P2kn1uDneMiMyzmCsBpuiCYPtseDm8Ib
cyIRmYG4M8GnVMTclCz5XUHdUkvNJTh/s7p3elP9dCvbZ8vhStWSPC5ject7Syi4vbbP+ZWAtYoL
kYjMpnq5s+IODqbvMljN2oeUfTa7wTxDdhosptOy11WuEjJP3Y841Gl32RbzVFd14fkSD5u26XMC
XGGNggnPuW2vpsd3dcUspTtu3mMBj3b/MOvS9Qbly8Q6aeW5GzvXF4/MvPsh/8SNG3LmDe9vOPdM
KI8zvOromUyChJwJ7ljKn0Hk59W5sFKMbfVBvF6aEsJQ3QU593lkmfkrFqxeQeiriOLbMuFmIdTG
7p5qDe7G2L4mDDixiKuOr9iWvMMsEGPsPp690X8Sj5XfEDUC7yvlRpoS73d9aSbz6bdVbvZqiwBt
/KaMim+PiYQg4VN1DY4dzaj6maeRkNhvmHKQn0iW2h70FBU1QM/lNbikBUTBNVQf00g3kpyRU1h/
htJLcjBiEuDmDd7WoXd9vEHrfV+R1IHpYleWzNiYQK1tKW1NdTg/r9ZSJVpfByVOaUq5Qa5H4iuR
qlBeRrfj1OQ8JKPeddv+5cb2wNWbs+tvYYSRPPxB/JaD1BLAe2w1PugXYOWlXGgust/jL3okNkd6
Q4gBsyYFkxh1uRND1iMygVMemIOzeN3UFtiOzzpuBu8sP4AvUpuF7NvAOI9N++yVNrfT3usC6qNF
a8PgShSMUOIUNpuPPuemqhu2IBXjKijj8KB6okC6UyajOaurtGc1Avwopn7bShXC9+NsKqTR5q1b
PKNxSyu+lJe4EQFgDZh+aNu8NnWUX4+2Lf62HeNBCk3O7IUvJw1LgbAThVqFnQtfR0l39tXjFDcZ
dJwxtZ1V7JQfTwkYEhn1KLPmhy9fvXRtryVzZY69wJf0na0vBJiOaP4N/deKC/qSJK4Bg0Q4Eomg
j46YNCSsrYM+NYSh9vN0Dua+LUlL1OOtrg9d5YxmzZ01oxUXrwA0cE8Flb3knKXjEuUJa5TC5oRP
KC0kPpDcMJy3c3IQMyrfKc6uOjP1Dks4QWxlb9nPDR169b2BT4up9S3OMCUDuvZWo1j95ptncOXR
h6gEvvwHHr2tve/V7MZ4mEUJFCCiU9BLuXorpnH/q7rByAybJhPUtSTg2m3KxSlsU/7aHmv6hFC7
qcIoRtUYCpI6Scb5wOYeiMIfgeufFhdAEkJFHNUNtWy6Co3jTNJd2YN75uvYqN/zKBUSAm66ipHh
fNSgUd9JrmdF2lrOypvjR0NlET4689cNNi51j5jNvVXJ+VB7fAdw+o6qOs8E7JqHiiXcAqt00Suz
vnTQjuKtrq/rxFVj/Gi1gP5OskHvwqqkgpL/nuXhNN1yX/AW9kraXI6R4Ktdkx+3J/Xo7iODLhnB
cVdapS2ZkW9tddKtJejovQWHyPanY/iCOsqeICFhjgUX0UsuEiRfQbLDluP1J63mQYFxzNL8tm+F
6aVI7JR6RWsupUhjLCiAKCCx6BXymGmQF5S7Pn7O0x7WiaymKQVt0xBe6U4AwDVz/xpnIfJ1a4XS
PNmcxPPIFCkz//fIipVU3y7KZBt1IDilMCW1DWccEsU/dEPXkKTSBFcDDGna4Zvo7t/vZT04DcHC
7BYlpAqAOhs/NqVRhwaL/+qYbz0YRQ/8ViEjBYsZZ1DnplJVWm5Hcs3d0hRKIVNKyY0rQ5mOrVxZ
BttzN1784TG/QXqxEnz+our2Dp3Xmuz8crQUMHmXHFlPgDme9qaeu2cHf1YiM9k8+S5MuY7/p06p
cP5tJUdXo+KAxLASA/6xswJvNPIIFIo0izveKmSi/GIeFWStDntbty1ZMNQmYRBjqc1bd+0+DIGx
zsx2isB+QSWplmedO4l+J0W306s0IEuNU5ECH9dHkDErhFwwhetxHhDt7/yrjCGjYCSux2kwhJQz
saRAqOR4lB0tVm8qbbCG3EK7yWLpFhrZPoW4+Achhj2R+OYhDzgMH8SWymFiwJ1loTxXnSNhMyWK
5qYbtzAAUPMW4jNm+PyFKR872MukkclCSkfUl8l/mJg4iJdAhWnz8LP9GbAISR0x67EFMGA+MY0e
9e2v0uLC6lDov5isc+8OmRX+FKE/7KYBwid0U9LcLoOxMlntcx6IPAMCd1pysTOAMneVt3TX9H1U
Q+37lQVSYbRSUK7uV9OLN3Ar6GBY/4TsXMSDz2jV+8GFKXgyYgkHFTfSgUOc9s6Rd1OC1j/DTlPT
WSZWWIYdje5bCQZ/ev/Z2CF0zNkdYpUMNSTiEnrYcLpOemwc27pX2e1EM6yeLFCYOkPVBk7DeEeK
shd5CHVfpxr++KdgOE1lRNbiHWHS92U51TgFhgmPMjtra/+Hlcm+Sdszq7sZKDP1oQcd5OCtyxMf
piUiGRbxhbQkDNYMLlZPssJu7ntKqxeM9t9bMSNUlsiDuKZBSrK7vUBVT6Zneb5wtnW/dzxx28E2
VALUgQjZ4/vKES2VoWHHGv74Z2piWp12SUWu9uW8tgVvmc6T6ar7Wg+24rKiuxnqKWOc5iG5y9pR
CDn8ox8OyGMFxGzr7qWiEdPaRGPxi3XFhsNtbg4GAIrQU1VIujz/GhvsDv/daKFWiW7Md6QOw37u
g7b/AdmdnbG5GGGrYAx+zcGRfIcgJEJqEEkaItc7hQ62XWb4kXub/SmlDFlht2wzjnqsORkCe34G
ePPllwTO0+3rbWh9NPWG1ISSde9fibykq4QF1OjH0nYu30WDSkR3jIukyjBkJgMjMJm6h1BbW+2i
f4+uABI+GPbuHC4nNt6yXrLC1TS/i1lP/nTm8JCCr4tnFouv/mZC+zl2tbdoxqlD18yAjbRzDY25
NloLI4hFOr84aygTQQWJMG9/LvQYHD+QaoGj5JJAZrqhrx9bc44xdj1NjBKG3LjdhgUdOxFqHzVz
gjqwk2GmdGwnyVjbP4IYp9NqETiN+xBjwXmuSnQxyr9dAHcie0OOswyVASPG1dPbyo+3ytZdD6c0
45EH7iYaR/kH3HmxxRYIhfU8MNKZhepX7ou4Roc6T/o/ExuTnvktbM+r3UDXVTcazElIK/ZkVlb+
kDWbQIKED0j9P3xJhz5or9TE+ARElKFPpNVGr2VUjxFcXSVWB9IGEoa2AnAZ0loGv5UboLdK476/
ACfiSGIMH9Z1hz0fYF6ufDcg2kvZf8sip+Q5QAE6hILQkQK+N8tsYY8XVV1mOdC4eQrgOPoY8OMS
FhmB/uAP77wS/K27eWIH8EZ12RGyTpK6yaNT6R6FFuet0ZOWRBsx/a9yc5lNhfl9TZMys/WHbNAS
5HmAJF0AQGWk+CVq4cuMU6HOY5Hd5B4dql2rPNO0xzxhDGFXYKGNVHDXyCXokePxlOF7pe7r+SPj
W/uC9Xi/0PG5FiuBoVY5C7i+tbkfKIOyRSmPa8GOk95cDEXdux9d6GbQFYC0LGvuegRith2/0biC
SBovB8KxdOgsmRxShtD5ADMv6IYpUeGTciGz51lRaxBighzQE4BQ9oln8gSiEcW0W2HPJ0E+Q41e
7Dv5SbtqwgzaZKed7RsPZ7h/uiIGr2eZajkyAyG7YDyNNuwYsc7VRNyVuB116uh+WMrJPemNy2kP
l3IhQDUDIEQA8dnOygeA0NSZOGl+j+oYqOpehpWC+mvrKB9xOPJhrS8XoC0pvBTAzIknWfAZvxLo
esxTfBdVQtMpU2ZIVsxxxcZGbTUTUzqNoet5uPfvS+aHZnsIeKx+Cu2Y6vEhZvmmWb+u+Jr8Lep3
e+t5Tr/l2IqzgKC5VmnIUtOMaEFKXocqnMiL+e+M9pB1s5EFy6nehDDLKxt6ZWk0d3ClIKNe63/X
MbP6ywpjPEk2LA9QOYImxGVBlRUIXRhS7t11bFKTGjBBjWyaGEzVeQufztCMDAWHjYw3sJbvJxpu
fnEwhAQn7lMoy6uf+jIZj5+kNinXAU5dB6X4NK1wXi3tsanws9TQAn2kd+7k82xUMbp5++MIRUmN
LZADgfY1Z2uiEqn0KaPWJhV/JABkxGfidfCth8T62zBNQztLfQPh/2si8YJcEUBykHeehrnjyedV
G4nqu+w2Z5VXdfHQWMjGezVA2dEb1ZiExiO3W9w7dLqL4OPOpGU/hIWe7bg4tmR9JYXdcOSJRB9r
V4zO3NjCpAIWjMPjJKOWrLE8oO0rW3T0E/ck4EKUi/YOC9atOgM+Y5utDESISvBolM4KOo8pzF4O
B5D56lXzGCF8ocHRInT6yxtxLvz+8GMVWKFaer8lsuEV0bsv07AsWGm7NSgKRT7TifJgf+AcaiAT
9xIvxsylj/dONb5C8Cq1MVlzsbuonZkUMHVQt1oOLRxUEywdt70tgoz/486oO5DoDVFQYiXgUgX2
YJe9nHc3jt7TgzitSlBgzqjJuWg31FaZyWrdOQlmBxRb6SQwpvrteohCMauwwZg8pztM8jFNSSyk
rI/fCh5KtIdEZUkpfiPa7Hx0FkrWoh6tsDuCLGkHEucLHkdaVtm6qcqiFmoT9d61ELeVCYtlzKHP
srbjis2XS0MfNyXiyYXkHTN5v8lGrC4V8MFxP0a5AGE+/pDkrC8wZN73s7AhTHHLp8U8xpmBzZpl
5cweu/ev2RJEFqXa1EHywI8rKVBOwJdLxcRbcZsX0VJ3KOwA2v5l7ITiiBYT6Na4eJlwD08FI/8y
x7X5wRPTe9hojONg4b1ihm5k7EzIaLVxr7d4WiZy+B32y/nxzEtTq79f/K9zegXkgyvGqImSvP4N
U/CxPyUa64urvtrqJ38uqhpmyNxkJMsYFO7vHG9iZqNThDxMa6hwaNSAF8L8/ZLrJscb22yGTkGQ
chfbkTaxqiT6fFKsdC5z2v9ourUtsH13Cw3ajeRh81yFCmQysKaiCYZ9h2DpyKd6IlJ5hyY3WQzn
RIr8/9kJ6IcVfProvK1jrwtcqqkwivtgwuOJUdCTvvJMYUpsiAnkl0W3RDoHTZowgR/bYLf974uZ
ji5sLWxb/7DYE1e9pOMhUwfuRxK19W8c5HFpc1mIb6DxfAzZlp5owEvvET1GVNaR7qtTL+Acve7f
VFB9MCTRPEkVTl5Crr+83QTRmAsgr2poOTaNa4thb0A3424S2IJtBBvvz+K7nw/An2V0Jnh9/bbY
nSdpXm2tV7qqCOZhSbvNyiikg5CJ9hrf/D1A/uKX2pikMw+/gr6agqLohaHh22TxYi6dzSB2s1Fm
lDSVETG2q3pqVhRqeIZBEiN619HS+rKS8R039aZ1smUEwdY7Cy309IJm03zqisA43uxdHjX8Ad9U
YBEJnLrH0wSc1AzPECt+Zg6A5onbIuwhVLCRrhpfylThMF2qMAPV6aqRgy6yihIGFfeR3ni75Kqd
ZhjdKT+DqLEkkMT18tEP2uC4bHpoSRPN1g5S1pWfCqDhW4Bz5vHtqIMzsjU6l92gH18TKUUFJk7C
F3gLnhBnks1YDs3SV29elMZk99a/o7eidXvyhmAv2/AdFxqhCdmFxUZOl959V/fu9Oaatq+olIP2
tZmFo4gynEgklnNs5TBALGpzvlLmwu8ShGZMBqNIDP37EQZDoXrW4JMmr+QXLkTR1cI4bG1qJH7C
0EY38TAWQ7g5pBmWtSwhAUpz5A982YalN+3hxfHDU0Bue6J4PIfpROsHdf3c56BlxfHKvw0rKLbx
kWAgm6TADBJxs+DXnbglZVIkOinbp2kPjNHakDmS6k/71Y2laTwOAJ6ZdEeJfRtFUNaNOxTDKmI0
vrhOkIB2wX61m5cfRGrMT2nqC6BIcfHvKVXOZChLtEvMNIIM5xRThZmHthmcSE5iCJdZOzI8CxfZ
S3yvMvYk66cK+yY4/bii94lZndNCUDAMV5IrYHV7Vz7XfxddsBspQChT3wu+vMuSWRr5jlCxtdAo
BSWXAZmSI+urD6bdLCg2CmwjAWYVEsuX8coRUrA1LT2QuTrF0OVHMbeKcrPNfyAiBTWxTIHybF02
P77VvUyz0WjEd8oPGPw8/WguVG7OO1dRs0YDdHr65xjtjPtSfrfsuoW2VrSg6O2K7aOlYWeiRMhQ
7PPxiuhUagjtv2EsIrZg0Jwen5Ux5b9/sLwzOLiR5+Ok5dqbWKjhyZ4/DD1t5W/q3elhlPZ4XEEF
DwbYwTD3Ae0KQDWMXijN3wvMO/9TTdCewFllDzKyu6yFPXdXW+NzUoCY8nQIGLY8chf6MH180PRg
LMtBrfHGWoBqfVZJq40wpxI9QQb4PeJDiT5VIWzOJzCg/xg6HTXbEw4WafoiVbLWWPrAeH/8a1NH
LDLtNmUte9i7gi034nrxQDHuYjKwGRDJaQmP85xeKZFDJJZeRETup3nYOBCx6f5EtEPSaoJpuFKe
i1a4VTuA3DMcGd2QTbG6v5xWe7+t6Pm89NFgk2oITy2qDN+ZD+1DlVgfWCm5xh4IDlk4OKzhU3MM
ZOP3fBKr6Zckb77OPDRSogvtOpHTHkkD4KFNcStARBiadO7erq3o8S30Vul8VOgaM4OyFp77UaZQ
bm9QoPMAG52LmhqjOL3DQFPBqNHNOBixZLrPnfmmmy/5GHB0aIHTTHH4J8DjysIMm6R13zrrvEHO
ShoqN/isXP8bY126L0bvv8E3XB+ioymPTRKSMYNNergAD0x3Pa/BT/Fure3Z1o6rulti966k83md
aT+/3rlcmSWA4OWw6K6ByB87/kOAU4HdiIjmsJvm60nKtIUJMAgV+9YwkuBVOFVTlEY3DKwtiBMk
WRfMNrQs7NWbMwBwJh5aFTGV5kshDugW8UM10Nu1QGERAE+fZoXeMrGbERA7oQ42Aa+nraz8vQC+
KfqFnAemzal+WxXmGlFX4ezNjJTQsImrB7YeQY/6LcXjcTrxtO4u23x8lpsqTT1bagBswz8ySVnR
O2YyxRasTPHSTqS7x+ASJwINaephLI97GsPDs4pUnN3NJ1+LtNvzbC17saqm4XUO9Hha6/hGaZTS
P3oK1FrpHS2/YmA+uAPKpRhwDHSIR8n+nezD7DBtT2wv9s0WY43uPs5rioiK/tA9WdAPVtjJAV3c
5MEQoFQl5HTABQdtIBS0W9j6BD1M3Sc//gJr+cscQxMBPIR+trcqYlSrUYkcMwerqDyEy9i/UTFC
Go56VlQrdii4gt4g9nob31aqd0zjRE4J+xB3zZz9DJzOBhbVhPEmvfYRV6K6QzKEMoHasfizrBIl
YtDAmFf1dNto2hiXxf19DRosTNFwTAxMF/WJTCJ1kcn8+7Ttijl4LO3oRXQDkNCm6CaMClENK4Gn
nZ1MUKOd9MiSA8rCWl4llOU0tLE3OAn5gzRfuLWsRNpcniiyHn8Leq43TisHBJVb6xqpultwRzmX
5kaEuJl5e+fveTKJ/Jj8g1+6KDGi+HEC1WxqHuK7znEz/GyBtYVpxA1nnLJIG+dbPCYmXxRX4cJY
AU+o4avT4YSjbuZJt6TBLToUHyFeJkoy7p81p0XgtwxysoMh2Gl+uycDDURlY5qnQhqZW6Hf5iXX
l4+GfMn5+dfTBaWj2+STQtAh7qjbCjtH6yDcyOxKXQ8ha66OeF4UlBnqCRc0LAPVuclDvI6qj8T4
90K53vGB4WHGzyzHscpoxH5m9S2oAao4BsbYbLmrlA2EglkB7EbFqKLYuwPnk8Fi9oI1CrhX9+Nk
3WP/cNqQMttzjG0r/su0l4dFiflG7kmOCsaF05uMdjjRglGHUwpUQ4a+eBMVa9TlZcCeQT/BbUn0
5HzF8MB9TO46zSI1qf3FcjbLOF8/dQNuwbPtU3NWGdRAum0l33WQbBBq0qiljBybDe6tC0vEmkGK
Honi17GwM5jrsu7M0n4Mz40GnNjno6RwDh4vGe6yuUGN11aaOOWozL8VPNt7EFEwboV97mXHnAUx
vyOaOpxkBZzqS9DreRu7iPQSmYttAMc75UAeNOji5ENpfWbKV1BV4sfeQuRKCOQwlCbFwM3780Sg
zVQkzvT9rrBAKI+CwwzhM32fKuz+xpkSTKKJgSw9vxbitgTgeP0SIMFc8sM9wUOeyFr3jlwD/BXm
fLDjx30HDz61PURIZ0VL2bqIQ+mANmdYVGTiBctcTWRnf3Xrefb2a+9JfhYcpRiY3a7sD4zxSapI
YTScYAZj3ZcKYwkVuwhYKBJpqcKcENcQv5t6y4VoIpgWKDnyQWV2ja1jk83U21bb/8tYgswocNJ7
bofsNQaVfk+pZiuzFiojJDrwmzsIJXF5vkJlnc32It1kGvyJV8wNEWe4MFNwDrFlJSO1eXtUjy4s
xW57ewpX5G3QSIKUnEcBbxXlMxfze2MPX8hiJ+QVoSzXpkAV6DlEuFZOhFvVhB/cYIVqBOT66ncX
w9+NvJRcBNMdFO697uHTxB9yetgQ3mvxncuzLwJ2HVD929f+Z8N2Gn+/8oWRFrZvaxPNXCLKL1PV
Pr2Kk/huCaApEoHwK3TuY+7F1rqK6zsBXH++JCPgn+y369blfaHCtkDaAriRKwMYMOjmT3tEV9vb
8BTB/pv3lSaNf/gXj+CTkJ7VcbpNxOVJMiyN6JJJy/tF8BnbzsM2qR/NjQE1axekNA4VAC/xvSZa
NoB4GpW5dshMIa5wvGTnWD4z1oFgo9OG6XHsjkgRwiu3UnqEOtY5zCSkfQtWGqnN7nT4MaJVpOlf
vye+5cZFZaZyPxbnjkGmdA22/UwyS420yDjS1iSYZqf44OjDUu7qWca9byC4syuin4d7ZyClZwzu
/VYd8DeAZgpUePMIJlkT5/6VTGWwlK1djAVSQT2fWCGNfx8Vmft/pp/xau7GmwygcR6HeEheew7h
VbQbO82OGurcdzvpA1B9Niw5iaaNs6+UD5PWtN3zmRmu0nw00NUjmYdkaJER+UHZfNZJmkGT7RuT
iphJp2jrYeR0uT4dm0xpCAlZTa6iYr7AXvgiCKaiSQVM0fJyOPYGEFhNvT0FLmcNnoPon5VYzhI8
O94qE56VanTAwXctTpT6KjnrvNJSlsbBZfYnqLYaVzVaohGh1soWDN0Rir0CKbo1QBw9/QBfiCrb
tHyR/6JqqnkxCurwxe0k7bLvcF8HBUST3ErxzXR8QJtVmnnmwoLfP/6uYWrW++dx1j0gopjBFyNl
9da+UHjQodbqAmQckoapI64OygysYiBT7tig6YGeomrMmiOXVD1xtggV0R8h0fXU5tBo0r7CjE+V
/FBtf5Fm32Fme1EVU6efUpc3YROcSwTTI8xoxi991NOYRjHh+lmYkLUMNuxUjTPFX2L13l7v+rI8
dUciLubaTf4MMy8ViMVoiinz5TfoVaDeJJhbpRLItZeLidMP1e5QWi+Ke/11K28HvrHLg2NsO6mj
l9TRWIBiamCw9hGy2SwzpG0vuVVdqthAoohDcd9DhwH/px5V+bZDLMJvu91fvlHpqQrGFS6W5S3D
rsQ+qn7ZotKdFu0o34XF6VjSCaBZfrQ8BBwrLz2VZ9NX9/qjQeAt2KlT9IbBf9vuOS8izw7mgboT
vx1vGnQ5ACMvamfBy4vRN0tJWrx1wtBRIkL8o5Ep2zYI1yK38RT8AyrK6s1955OR9eEvVy0zu23q
7xEpvAo1+eoI7fMk4vJ89Fng85u1IG1y5ucenjp5EpkEowJhle25puyj62Tc3uMNhIJStBtSawkf
x7f1hmyyZJO+dJaHrOAc4cb9lHBrgktC6HvAGdRd1KQBIk5KW9s/xKRfTAArP3NYZf6HtFJTzbmp
unAe6KsIvaMSciYwAb5ZwnTV7CtntIfVXkfVPAb00YpLYnzAOtnMFHrGUoybXDtbLE0UfXvPegK6
c3Q4nbaaSZxr1AJIj5CQIt4gD4/MX+k+7YQeietnXrhBNwkfT38wwEgtMXnrcSU4OqsXJ+IdAQQY
UDKZXKBxWH3puHWQC83rD18AI1Uyafd9gTJBfVvGMiWU5Swc6ngvxsSXnm09MtXeQsjfJ1WEa07J
V33W/sfKeXtf0U9w/4swiyFDwtFJ17/VA3A1QHGv9VWeYzl4Ik4tn2OF08TP964dR7M2TKY9Ch1j
GTADfBSYsMXW0AumNmWDkQZE7pW4Z/QzLHkddRmMyyZhUhXf29JAnD33zwzb1dL3GKCU6uC06+6D
1MJnBWwezqUAceI30SSWAkH2fs7JGLj1kQjdfKWPHBXk4nVh3JN0IuKj6DkpNaQ4/oZJQIsS9kfW
i1/epk4T6fI6ASApd20gba2kQtxaHMZvdU56EyFvMrSGsIbgvtniBrU2Y6agG1ZMH319pdS6gdkT
9tA3odqMc25x3rd3senHc25Ee5B+Ij2qQ6iPVvFTJh9xwgUsaAdx2IY4TpZ8wi+ooMDTfGetwf9B
UDl1dbTOHBStLOgitsZhSary/rPG5smi1prIR8rWKMC+VtY1AqPGXNF+NOYbxwMOJOv4DY9blGLj
B2Xt6dUubLFHHJ8KRf7kKLoQoUt3olChnRXDhpIqeGWlMseE6aXezlamOrkR7A1sdyuBj9tV930v
BxmWoVgf3h3KQThsK3FGeL9ubusbBGliz/G18Mnwo5QL/VW7DxITmGrueise6ht8m6NdksXqzsCq
NPXooKkhqJCW6B66jCyerK/AH6H4vbI5IIaUB98/GZc/EhBRk/qw48unkoLDVN9X1AcDTH9uU5G1
+lyRYAzn7n7K7WPvjYFADm8e9IFEUi6Hp/fFzBJ/b8XTXE/MGG+kypSQF2edknidYjq5R3lefSbS
QgbX4pYulNCaYPqPwFsZbVdNPrKhIFno9rITfG0TaFJD3F6VwAkWn6XNfKMUOPbk01lRkqCewnbc
/hWWdyfGIcMJTxXKnHDpfp6t/3ORy77K0hs/tMoxjWs4mjP2vynBZzacdj/FvGZTq3NGOevZzLkJ
2kyus7wzMwtEzjnmKCWBLkqXqkTL4Yo6KJP9BOq09Z3+O2A1zMuqW9h46zWixr5OAwqLnPkymlil
5iWoeYKuP9P1IMxce/3X8VqJpW6lNaA6Hy5ebkuMqAP80dZFRHrN0LRruKbvZFNV45mn/rUQryb6
oraqfMfGccumVo0S32pzPHPk9wYrY3Kl7G+5In3ICuMQ7vbfJD/ylg85RNoG3VIe1QS67CSHzb+m
ER8l0y+BwwWeMtfX7lBLUP3aGqAu+KqH8CbGLW/yZmLB9ibrNfmZ7H6BkXnu3dUuXoq7V4KvBVNb
PJB+6x4KLhPD2o1gl8saP5hwapc9wo176mEpxe+42yXhmGkHAW8aR7DpuWWtS+afD0WG90IUjZXQ
cEVW816upN+2bXMLbEZcc2VW9lIk1rY8Sp1aH9dP/dmnXCJicf8iy8LNaRsOsnp7/fydRlCpcXDE
MmNQc9Xw6DB3/tugurcxMyO4VsC/NYFr81iZewqBLnM49d3/TpmC1VszR4FlEjPiD5okuaemq7Gj
HHEzgvzUz/W3Qi4u1cIeMiOH7QTznWCKEOB1/g7SSfciYqZEjLPIm3vns3jf9VFdzzkV6W5woHjm
KA/IVWCWJ1O58mgViuGoJO2luwadrKGa3BhlbJp1mVjPoAjihelBag4nouvPT0KZjrK44crGfwTr
i2oE8wQryfWUUfuLCOWDdZzsqJIDWuO6eKm3lM+s7A4HMB0mmElScvPL8gYFwaVP1I/PDGMhCzF1
85Rei4FhlSKq4g11Ys4OBwaNwFBJvaq/hJAn71vgUJQOomfYKkshWVDaAPlj64qUxPPGGFhdRO9o
yaPqW0FRpES+opEZoApYs++GEukUUeXhknT0V0ifHpt7REEn8hYh+TvtR4SVARAvMZ08ceICPKjn
nPlp/vfbrD1GFHEOpbz2K5PHq/1Z9gS+QituT7o9Ygf2l8L4kfuxMHGTWIljyNfVLPYk0Q8XIl4w
4EmsPGZadafdAK/YIoBMCYn2Cc+ybUNlk5EAl5XCSXEa2yWDrZMtSsLPuMyOlIqkbHlTIGNcQkYi
fh+PCdwVA2Vkj0Rz22ZxHCshHSDGs+Q2Ks4ZuM1beYl+hbSQMMTaL72DnsDbDMT5CAqanyKpNR0X
Vasz+qzEuQWksJ/kRFniKf86XvsWnt0GFgwYHQrvNdIjtZXhtzTOt9DmTeRkUUTIe/+DW9Og7cRC
Ar5YuYNPzWvJoqdLtt2iUNjwKTvV/50/h8mvMd2+kM2Z17oY7qiWV2+fQpMj1wr7FN95ybVe0ENh
Yi9bGLgDNXbc7EeChwjjIip1LB1kRfAW2YqmYyUvBx2zOoJ54Lpc2NQ5wqYZgo0sOhYpAmwfR0ew
TzVXVCXkoDGjLB1yJslMEG/l+dCE7IaRoBsMzvbjwEsL4rJx6wIov2w6KEyiNNmOED73CHY6g2ud
o2BzgWmYPVFvSaGz4DKKVuOevdouXH3NOwY91gGwAmcBJlByTgWMYSUlpAzLx/Q/aI271m4z6UJ9
rNzGQoLLduoPW9tL6rngk4bC5RDA7hdZCmNVmAQuS/obr57ftrr8SPB9bGP8iJrUpWNQ7TVACAsi
WoM2nBSIjVnScgSx24TyRQIqFqbVvcDu85FKBcRYFQyriZPjNzekm6EaIOspu1nXqjt7SLpKMBYq
rqZma9Am47Jqvs7WSV91X80gYHyMdWcthtG1DiHR8aE29RyDWvLStItfllm22B/iK+3LdsChB8oO
hsaOEyzR4HbjaqbuSSDbCvt7oxy+XV2NV30MgDDw2F9RXqFNLhz1uOe9Rpng28rL9PSIElAtxISX
QYnKhILiMbI+aXKKzc6joZWrwN4JhR8Xynk2oZnY3GOJ4FMg3FrKbD4HtioyDBkGvWQIKZJNqrAI
pAc1RrNASK7Va5JVGbI5CRsbjD4lecaaRMmnrw1KtFBt5AWODY5KP29BrGGqeqxXgiMq/hvq3aSt
59MyMvY2Wtx50NHuhq4VcbOn2EvNDnyLSy+zRqTxOCbs+F8X/CU+gHqb8n2ODgT1mHKw28iOLSOp
db1bD7yLqCYXchXOYeR5R1V4FD08jn3j8oSMP5tzgzSkDNoEe6fZNFv6VdABWhg6yq93w4RSkwv+
+oU/KGe8XnBb2FvsB4+5k0MOhLvTEr/+F/1kP9Hn3VgegCKz8qRL1HLBi3Gq77zigYnNKa97Pxze
EFb2x2brG37fTM23SVkiIi59lXKIn0J7keGq9DFijKANr4Ep5ak9fjosuTb/SPc8mOIEndZeZanV
D0IJ3o8TmtXtE6IHrfLIdlp5oIl74a3lo0c8WHTAvjP92jC/lcugI38q6AkRJA0S9LOTEcjrWDxB
83xzB0EY3mi9bBxX19Pz17i7F7IlyjqouD/O5L8belfFey6ej4Fjx1ssCde0Z/2RVXGh8KPDHW6m
OGYmYun1O32sk2DMw+QpEq0jZAnUjgZv1kORZneG/ZWcnUwefeccs0NBC7faDZ3E5OsFvUnzq8pG
0JXhbPwKZqvv9tY5OFVqacfDB3eb14ehXeXF25wXTKFDULoEFfkFzVUWbjjuDUXpswSvA56z+0mm
bKLsf4KWb4M4ai5T1Rvc/gnLXEZIUYjLT10FS9iYHdbk0Nl4PXvntSE91+hEN0cqUAyPeIVCGN8Q
SA369tRtwVU0YohU2/JaY3AVn+I5/zek4IRlchk7H1S2vwwMz0C3LKOhEBy9riHaVI0u6ga8dlDn
JrhD5QZ7KXZ2/nJmlqfKr5SvXR36DiTkjOXMY2iZfezi10umkAxcCkwnX2H8Fk/gj+t1L1qqdXRB
KoN6+VwgrK63KrmGHzA4aZQF3qEELzQWVXpelGcFfs8xesm+InQU3FbdZLTSv30acn0N/oJ/MU3z
WWKvmtyXKe8VurjxT6iuit5cRX3mLe6NTFoCCy7N4ga63ZBTliENUDKTo/hVoNO5WHiWr7h7wnRB
r7EXwTk4XfE55G0KLBIJurHhmu+45wWxetqoIQuNAPtIxpzMnzv6MXdlrA+ieDHTFTxXOh5iMYYI
pxLo0ICoEC8JgBnW2k4bOu2jIhAaZfaW4waL/Rl5MDYcnaR3mfmIAhfFfFbiEcvQXKnROslSGnFd
OJgooN/ga8+NOBeyoo0CF8vb37WqDEeaxJI3KUVCiN64r6eDMwVz2lyxJAViiRhZA97sPFPiQEdB
09NvFUhsJKGnQXUsVxzuuTgfRFTBWMju68lzFXYGGQEl5TRAz5khS3zH7lk5nfAwDsyQMoudiG+8
tr5vuiZDFrWjtXL7cFiKRpsaJFyejuFlWPn5s/WamD/wN/Ea7Q2lZPXVl85/VMLnsUJEcW5rwTsw
Um/eGx18euQwJCZrCm59UR3AqTptCNJwP92oSVPbaNQOjr3gMYCChe0knnOlmzI+titiZTptJYsc
94mRdhsB79Zdy6G9+vi4MKetCgtJGLWhFljeUMY6fha+ZG83PKih0eAcsoOCuue+AhcvzQm8BYev
JsIJKm4/mX6nM4Bu9XQ09ggr+cZiDV7pBtexSpDHtTDWKLpxSde8T6Ksq0VKBXeZf+IntAppCHzU
wTdjViGmKQOLGEoCqfss27JSH/4noHd9ZgbUI4zTsqEDTvkbwtd43/CXwxTLYDviVS7/4Hh0vZ02
KEcdNK99cMOMlp/xYzsrtVYiNyk3R0VS/C79j58C7WZ4pAo1fML87UZ0dlky+SV7yo2FFRsMPHIP
DYCyCTGBoOjy4iIbiJ92slT+1VCUnqU7kX9rukQSRK22Dvx1OYRYNl65Q4TddUw5xSbtW/hnPzKo
0IsdzwA0pEvCChxpUx0YGOTqsiYYj9GrBiPLdzER4FLBEXOATo4kAYpkhanw0zuQYLS1B4vJoc4T
kxD/qxryJd3Yg5r8L54rb8MTlYGYpbJxbTtpomUR3TuX/0y2sit5TUNAzpJMAQD8ydXDN2TOrNGl
QA/ZG6APigA7ux4g4JE8UJEKjww234V8/m0auE3NaZbk384N+YPA37ErOSeCqkGqPwEc4sszB0/2
r9RHOPvR/fh1AAT+JYXG6xnrceacwRzAFnrhCBs0KX8DgOfovryolYFmUPklQobD4f3qYlpNdgVi
END1YXqUeZmhM2expDyZGiJs77jqx2IHOmNABSNLlxmfrYxzspQox1yOe0aE7AVU8gIG5NkkqSrf
UDZfxMjGW0F4jfI8qr8neZwWqXY+2XI3Wg4oTI9UGCr/L5HpkbYQwpXbEauTUM4uwW29/RCt9tFo
UhMbBL0NjSJo9KuQ+LD3Kh0ZzyOy6EbUNEk/ZOaXY/d/DoCPZNlzy1EraoC4aZYoVdSi1n+Dpz7F
UwOwMqeiUpUjj2L27FhFJAjc/tepoJ2GtV853XcEWW+emVdWzdXWLZgQSd1CvfTRVu/JcRMyEfAj
bjYRcVHru6ftFyOQ7cqqfw6Xzq8u3qnmzeGKQyg/EZlDCkezsqg8zQ1PSBjuQ20QSGmg3XPFCvPW
/Il0iWFuhHpWZ+pZ7k7cdB8/9rZGMv3M6pO7t5IDpHY9kJCfFGHrPaLXy+8OMBCTtgSVzUKGhN3h
67PQPUJ6Vhvql1A/NbYLyUhZ9o7p4ddZshiL3xFHUz6cPfBMKPQgNfDdPho62xALoABcmC3XzgAj
J4nRc/obELAvF0v6Qa1L16XoaXrZoBbF78abC/TzAIBgTZEBgR90OZ8muGPxFOLW+ICf/cNEe+Ks
PJIf/hNYmOaqZFHcLQxN2I8jDXzkeAM11B9S9Trq0UNMi7YWii1cWtGVe1Mky5cFj4lGqEjk/FBW
PRyymZ3wxNAHmc93/bisdTvFc2eelu8R/gszSOj+nMFL92tuA514carU8sTKdd/n4dguLjJ/ndz8
Yn/yxnVsL5vn3Mo21ihCVklJer98MH77GznPBcopjIFaVluxDMxkChSudIsGtvRZalxgvagZu6p1
sjPw2z9kOs6sWufB2B5bX8h4IvHYIYKYyUUXqik+NRqL1QwuRX1fMtiXLDj7too8stm0UL3wq/Kq
Q4fTffv4nUNgKX9ZNcyhOwoJ7CKk5C0XFaOFTStI8E2mP7i4kJjIWj4axNI7ehV3Rs3Qk6SS2QWa
oLZMhdTVA5STM71HQfezzMovnmATDlFScp43LBlrRcIjgSzFA3xeHKH4RHYlGeRII5IWEoTFzsUc
JzAqtgH2v+mOY/emM7tG1WLTfIAELSyhPJCia0o1xqO6CSqfrbgvl7S2MEws0Q1ugrApGnMosFGw
pbYhjNkRskLYvm5Me7yKGyjyHrCKTwAabLaSC1EJu+UcSiVgBmaz6cZdm+Q7AjB+ugeUMc+l6EuA
e3pntCEDfdBi2N3VtoGhNV3Z+PLzpXy7+HFG+yVAesuA8gqFCaRy0nLonEa6WGuDz0pt6wtUADL0
zziCzqJ1IljUNHVF3uvrqZQZtvAQqvQE7Fx5pqW1p5vv9S8Ybi3qwxsWIlilCSBODUX8ZW3x5NaJ
EPah+nSF/zUhdI5TMhbp4NrE+nVvB5ufFZlLIxPWXfwXE9DrEAqpft+/+gilGg4391/ts1XqUyef
dq+9HcKBy7w7GwaVqM9uYn/I3fe3dhjrCR1lYgHA8XVqySUh4jJsB/990DPQHNwRtmz5nWH11Wrm
bAIswBHvqeK3BXiXVIcIRpkWLFlBhFPcStK1tEMtMI7PfZ9H1z8HP8V2WFrpwoXbSSFbxIrYOdQz
ScBVdrHnQDy+K0IkKe1cBPRbo1J8U6upfDi2zf9V1qZ4GVjdGPNC6Baqeiy/Rl6cOVLbMHJPySxH
d/0pJdkQI2STAAGuLROSc/ilHKZYpM2TYbindSqe45vA1O2Q95boipLqqVjC6mc0l+S79vU92bWY
5OMw0sdawqrztczQRVymcqUeZ23JHqns2RlvYrXjSny/5FlaMe8r/WPwXh+XCsPyDfEMAsqbEc1z
QbZkbOeHJcvw0SSPQ3JDFOTCHJIaloyukS+Y1KsgKUw5xUbG8RxRtjGV01Hj75og68a6Vsqv5/cW
HtoUfeMkPBnJ09F4kmbGpCYmXcpjufpnzJn5I+T3IWNYk2XRuRcixv7sL16zotY5SU82/WFJV6sS
kuV6TeiZmgyxphTTuqUDKNt9UHnOxGW4Zl0TU2yw2fIEmolMQLQr75CgB3WKfPAoy66BD6NV6LHr
jZ8Sw3I8UMjCbZ0LrINY5V7GJdzekD6hXjqzgx2P+IZ6LKzNRANlGLRISm2ZdgTUsVZFM7pe2qJn
tfKOqWDRdzPx2bAF/Rtioulc50ujRF8ZXV1/vB1F8+Jn5bE/wJzz4JAYJyi9NmXRB2UkS8cws/R7
V6z6snvnpxkpS0zctaOfAdx1PlTO6LNNXB2ybA1ym0bqvLvL5WgFXELu9/Mj87YiHkzNdMRDtDhM
raxIumNRrLRYgwOzBitHbk+e7jgIjbYdwh3+ap1s2p2shGiEgwpklxTBxIGbIvu+OalthpCqdKlU
xqJhXKgE7PgyngJKpJMU9flnMGlPlxabOoYfWIakc1kT6OmDghxS//Tl4mNzTlIt2gNhN7oWJpLZ
Of1Ri+n8eFerDToTkXfwPkrsff5AG8G1CcF48YtRCUQ04ZMhJV2s69d5LyHDTs2Sc3Tw7G6/Azhz
EGAk6cwMat3kMKXh2E0Ycsv16VJ2RHdFQfnUkk5Ji2FVsk04KDi4yj4+Q671/uBqAsfYZriWAxj2
gEWJNusTenXDMS9UTgxSTnu/b8wJ4RdMPd5/RKUBMhaDq/fyp4Chd5uqJ0JOkY33MtG8yLgg9EUm
BlGSnYxv02IQ8NCYkut1oaApVR38n+lCSMudjqnE8thFFBImYB4bYfp7OXwjpCuc0FPmkVVY00nT
9Jlxq1aDKBWxil5QQ3bEvldHB+1mmpS3t4QML6s6F+L5UesmNS9zOsbZWlhsCjxm70Z6naANAE31
rcbhhPasx1qAE3z16RkSxURYtjf/gVpNdiN6IF4v1kbaa4+WG0eGqbVNCEuJenhlkQ0LgntPcdrE
LlxH3PzcsfO4rz6zL6vyIK9V0slrbooEMqjWh5zJwDwQbyGjG5NsKyuU3SyNRR9neT+3p5QJ1H6B
uJHnIobTcGZC0WAz6KmGQv2hZwu4AiHi2jAQbQ8pw2t1F/bXop1CCJBQh3270Fqx7WZ/6TmPLmCG
mYQA9lB1YP2UIndIOvB7JWzggLMcPFf3AejMYqeYZWI0DoD4NsaqvdbZSvVITVAc0DUFwyOo6LGr
TABSACww9uuhXu7rA2MbKZW3g3maR2SMVA67ay755IEMwmaEjItMBG9vdkJkLKh4bW4YKcjFtQEO
VTfwQPZb+JFz8WdvlCuNaWVGmZNcx1FfmmDlT/2sHDWD3lYF4uwhUy5X6vD6FiQrCQvLdJy0aeNR
JBcySK8JnUnLyRoSXKdhqVzz+gCsZNM3lrLoVxz1QOoLUXCG9AAjcrqrsXmM6clRJzQuP6le43Vh
Baf5Koocwc63D5JLnEJTvFIZQgfG0/+kGTunZr08yCUq78aEFSIRAJBYtmY5cyBHd8Yq/RczA0z0
+CD5jfpaQ58l+d1/qn+evQiHxRBP+xKapsW4P3ElfIGt8e/aHKAqXml7/uIT3nYxX+PRI+JX9jol
xFk3C8L1aEH4BCEgsMhbbWAYxj0Le63QYf9D0GhSLDzNiOzMD/icgfTh6AZIXg1zqEEpw3RU3Dks
SuyIybgo/qIBGl2Rb8M2skGdEaXn71VtW/8aj5Q4sbiQJxbH13TBdqd0UGQqAOmgyqBSB34ztKaY
EuYiWsWZi8qkE9rMgOsLtCKxr6zN8WtNdt5qKJVboNxIakSI1jW+7hlK/wwc6hwEHZbIovUpyOwv
zDvxmJc++7jXVZzJ4Ll7hT4/GLwYpo2lJTEE4XbhlxzgBNyPdcBspFAb1xVEe2zlH3Cd06LG975Z
rmssYc8bCROn8WyUPR6Tl2k89sp8KvvD+NGxLXIIfALH8DHxYlFmcTWeSa8+tJt3drob9vW4cUDH
6M4QRuajwSBwvJBgJUau5EXIaZl+sxGHmqMFK8ggYDoqxLkuigZTAe6pur7TTLIsmYQfmUyCGlfA
0t0CshEsRLQnkAVU8Mb2hfmdwae6yiuvp4FGq0Bw+UTHbrRxR9ZJ8yD2iCqwwqC1GhyQ3GJjaps9
xAWxPS7QhaIVKE2TwR3zZo+KmTTzRn1ou8BMNtEVvyK+SM1NBrVESBLiWCWou580dlACctaDWsU+
LXJaVvA6UNbRih3oxwZwAMvBcq4XiT3LQp7/3EbMH3L1VEFteheFpyqttHSTSKnKDIPX47uTR/Aj
R3KGebm7JPdqYc9sopYUK6IY9kPnikUXRWe5L5oL6ASz2ZcpXeVg3as9wRYwCi+FsbwR8mqw2Ztg
sxdF5K7zE1BdqSBAtpm3rEUrsi0UIZj/xxphoqojRupAByGrj3lPXAlWiUf9Ny/ZOwjMwj/99Yo7
uO+0MEpNsAQaMzrE1Um8ziOpqHQSf9x0nwi6X34V2KSJhxkf2n6oiupc0m8tWqNJJ9s5MKIU4f00
n2BWS+dzUfdcgs9HJukuZgbY0rHTmd+NAIo5xVRfV8F1Tis6fHRfMRe94F7hZA8ih0sJlbJVS1ZZ
iOsoSkbjOs+Ab8M0/4rry9c7DrRZzGpxyb2P99GyfmIL5umfUfBzkqeKNHlGkSPE//a1ISwflBKz
PpV0+4NX5P4/ZIHW6NzCpgcYgG0PQMlMQbrHrcSUJjM7P/HzrCAvoYjXHBwqe2xAPoB5fKFGFy+k
y802IICDwPBMqwPnjkidbdIYyPIRmzj8lWNyz4Ylx8DguuXRGzZ1Y4FiZbcOExGbrtKQcQASNxkz
fHXCsEH1snFwnDUQwpZGZcrz7wo/mc6Y9I/BIzmdMaBQbvU1pstUg3WOp8ik4rMkdsYSTzKgddfQ
uaRCdoGnXymCeoK/eU9+rriPnOAtc03A6B1y69jIoYBlPdrSYKvUfF9Nl5eDRzRWK2n7n3f9sIZk
mIWxt6dceTEkwS5Bx143Han3ybI+MvoPWqYCbT9VKZKQkw31hho5YMilqEHlW863loyYh841W216
Lub5Ugeex3fG4LAdZrErPu/5TLYiX4ubbbBCdPAEMLPrAN5AJW6ieTQP9EVgbXakFOKGHuPmlrAz
0kKCmh4m6VD+3BmsT4ydgZpuWJlDkYaarH5uxhEB0hvTpc2eCOb/xoZ8vH6qsB0Xsmtgy0/M9R00
pf+RjRX6uz+ZdtmqZgEXeePb76Ca2NxuQE5tsF26M3qSSC9YF3OfWJ9urynTD5ktXVzstJcQxWX1
QtfbjY8o3GgitSqoh12VVfHD/7jRUsht8aiGfa8GTHtrHCWszK05Lp8RcAYn2dzc9nErQ50+DyhD
DzYIfM7s8Yik2wpTv7MHmC3B1r0gcCxnPzISzmCj5cchZbQITeYk4qn35sOI9NyeUafqzy9R8qO/
waDyTtKOXJFatB2ZrC3rYPVSxYDmGsBhmtu4cdpf1Pg8hHbV1gLJNb26GauprMaU1C44geLep1FB
TYctzcG3G5VK+2Ka3f7d9HEbWcSthmLD/YL5dFbw3dpZLy554lSfR/Elb2AzejOrve6iIRVsgIoE
dbewPGpI2W1qo9whEFLMJfxeqIR8cRYJheZgvY9bvw13FRVAQf7mPXfSX1//dGThro65BJCqGEUS
0LOeIVZuUAuQmoa4II/1IKtjjbPCMoZndoxbsZnY0bis95GDODi2DB0lrw093tqzkOXjtnaHe8kf
LG5MyYJCpQySxiRKXz5+RQL9Jc/N5lzk6LRvcLip9+o1gWn0DNXsD783R6iqg0uMgigQ8SE6/Fo5
8NVgIpB+gIxW7flMc5VeRvXn5qPgHv+S6ngTytdNmHoaX/EDHk/FxJQm6cLOkt8opCqcdkl7ssGx
gpZ062dwD3aYKHO6qUmPK3xe1oGGZUMka8rh0GZraEwgvjcyA7HBbUzNhOGh0EIuONC7moSsqNHD
EQ8GCzTM9t26sJxFh53VJXYtnQFEx4ozYiaEANjHY0cFvn6EuNkK0xZXdKDyJtftKiNSkjcT5/9A
on534UZ1lvvlvHAq+SmROrQo8oQBedCpFQPbfwqkIXSkK93zE4p3bJhboOYMAO3igKzDNdBbiPAu
bm2Rwv1PjYB3VHCTyZ/Pw8ElqjH3yASUHzb9PpGpGGFVMB7hmJMPDizRLo3OW3QUZwgH00ZQ2BgN
CBgoYs/L0A2spsJSDi5z7bBSNsbMFrPwIfgKLid0pxxrR4Gb18QRb1clFOHqellVaQjHeVxjhwAz
kvC30aXN6xr3xktG2Y5Sh63wVZEiwBhmunlS3Frug1ltfWWNGOLeUBUhw/doFi6GWoyaWjh0vfVJ
f/+/I9oLXmGsIrlqcd6KuW35u9xFmZxoYh9kvSUiqfUX3Dw2EyluuFBtCSacIKZkJCRt5A2Ss8zz
ixJk3GEQYRtj9CavRO+PvAZgWobie/c16dYhO9ooimjs811h37KvsogClTAd5S+uJN1DA2kq8l/P
dgq2Ma5D4OMfF87sstveH991tAt7j0cdly+JMQIW6PjN/UsCNq38obluaQjse75R3h57/OEYgLP6
nLyr4J8z5ygd9P1RhZY7Dq03Uk/rFpTmUujymQJQMHBfu9omByHdv8ZykizWQvtGooS1dYwfnflC
wXxwUhUWY1XxBBg/Sz3zmvoWbIYiJ34j75kDeg+AWV4zCigtke8yzYhozw6NLP8RQNQLKNM5gmPG
DZtwIDHy1zLC1M/0BYFJjgsOwP94JD0G1gDLaLhCy40Dk4YGwSJsaYrejS4ttAgiiraaWjsxPxJ4
+GOCtWddS72PFUPovUUByIKmBLCfAPaXVl9GUs5qffkgzlsZ7vX4yaHPTJGM/d4g7Ya8KhP9hv86
P02R/x8rUmSXLi6y2Ws8Fa+R3wriaj8HENb3cnAOoDWFwm9rgMEt/HOeyWBuWXfNo/LujVSPBPmY
+fZyjL/xeSbsbDYAU2yoil2Bv+NINaaJc+aj0IoAZHp6nYCVxG5Xd67HO8p6fA6zPEyJtDwuBSF+
BSNzfIXuyPX1EPJjv7y+/l2H09BJlFCCepqRhcCoBUg+MvsP/JC6fLSdx3u8tuwK1XEEtIDWiI1j
9dddLkpCSS/z/oqmsRCLjGFPKJeZKBTFm3a1tGJY6wKk9JRqaezOEeWR2sfIF0XmNhowo3kXwAQh
UeEchaY2dh9AX4n7Qi/o2Vq2+g7FoQv6UhaMfZNF4BPp7rvko0NJrhfLzT7ZMhX/yPVBKWT3OrRM
EFNLanSF4UhjDhOVT6clCxIehIZlj6lzvMjBdPkhxvZ8o5g7K8vl8dmzFh3beTZwVQl/OAWqRZN4
vAu8bSku6e/cWrZ3ACUrguzBmz+/FM5EYj2OWkl9M1UBUWoamEZmpkuMrp1do7PkBdqqhim3hx5A
ueaR+JePbO2BJ4eSpoFbC6PaOQ91wTS2qdtxSrlr2I/vRP3/R5FqBHX6DT4vMA13vnEYVfSgUMkZ
h+d+QcmqiNR1dtLBjWirIRoYpKWmDL4dI1UU/BhRo9Y9NvN0LhqOcXkaYn7alKd9IPiEOAyMTlhA
CKwcktIS01g7IfSAQwmtpRRQE0/nqktu+g01FmcOwHK/PB/hVDoXFkJ9Oqt3uVS8tFEJw++/INzs
hrkBcKxihOBvUCJuWa7Df+JsTq3ikFX+gD56/TgU4NsDPSCYSUoNTM+5nGfCivp48LxbbhStAqZ2
vhBEVty7f4liGV4Nb0uVJb71gagKxwripyLcpwc/P4eO2et8GxrubHjpj38sEwdt7ZtAujeojAPw
xZtPXYcsP+I4HW/ke0E2lGCpQ0pS4rABZ+FBez7QUOm7N8eg72yPIZTjf9wRq2alT9FibaUAWuZk
o+G62U0Ed0Bjdf501gPAuYPc1xkZjH3avjXJT48jnGIeeikfU0FUBoPktL415q2CXlSD5+5c4qSC
1WR4t9pydeY2Pxjv+S47yBC3vrIvYlmFosfwjc9I6PWjJl44x4QbJ3vdeGhVGsAIR4AIFaAMypB3
7pO9KqGAyFgsxtNg3V6gzW2TjS8NUiPPY5o8XKhv+0Qjn8Ljlll1qQl5kcFfxTFrR34asmNdR17y
4BrUKsoF0pA88tSMcF+vCWAht5skpyLQqXi+2a6t7qrRCZ1PSDBk3kNB7amQPy/FpNis7te25oSG
cNyMv3M0eAXGwGhmGlsRLB6lNiLkVPk6jyBMgc90fQpiCrTaHaH9zDF519I+7YTJkWxeacOTgtKo
79ccfkiG8VsK2YaNyIeFdcAZczGgDicidGiN27cIoGXX+xwQo5dK+Q+rGm0hIMH6994RhjC44crB
vwPz9Xil7zHjTv76dx5oTqrKn4Veejp++d1wOJc38LkikY/f7MuzoV08FCbtGcWkZ7FXdse63tVs
n6+h2jGxfftPHjilBrwrD9vAA59knicle4zV9kiKlJUWiheXvpcQTKsUKh34GfoHcHmqEOwlFt4o
pjbL5lA1/w+6g4Vo3cA9RKs47ICxjPtaAK2kMg583cZBeJ+LOiNx1rwk5XgAT6bbRsiJZqpZ0MvZ
bpXQqcfqDCXnDihAI6g40IK2OBCUTIJsc/YlF7K+RWicUQekgF6R8pcLKdJX8Cz3yz99LfNTEPdk
VJfykUMH17/7fXEGrAeK10yiOwR0JYq+iIhu7R/5jrswe49vt3s5qzER38FGBdvSzp82ASd3x6JN
QfJmxKJ+pTQSJTNPkLbdw4B0FZYgHGdcnjPZGEJReKyyL+LJZVQQBqzF4va/3vEKHG+5uLP9rT5h
TMthLpmGUr0ZKlZcW1UAmJV/Qf4dfpIDfcFFiRYzpi3/DjPiWN+lZFAqrY7wi2Hxp0Tk0FKY56fs
NStKoQJYI8JtM/TKqG+MwVPPfUEahPxLV1uLVoC7S123JPhVqFGfy/AzmWfPnbyYnaDfxONe7lPt
qztvn4U8TARAOMYUZd623t0PxxHUaZvGId08BM9z+3XhVAMREY5YwWQk94kg9aUAl6upqQEVbQKP
rprqJ2DqMkwfjPngFNrmVE7/cG0cYoZ3unTW538fVkRAKTjL3ilXG2UP4VQ8kvsnOlkmG+Os4ffi
FUbgUx70QPljL03xefYVE/hj+MLpvOc68uX+54Ttlv7yrFao3cC/KzCI8HRhpn5f79GgaDmHTjjU
mtnLKr//BsS3MdQf34CjjKbnNKVIuRr7TKG43tmmArHSGq5XaRCkFJRkaMHi37JWoZ7C1w5d9G8D
/WorDTptms2UIVLFfX7zpPNMW3BdUb01s64cTrTIFTtmNIjPP5d7SUZ0WKIDmW28Y8OJ2cuG7iAN
jvtROuXyOJRTHLCEuxYYbRqmnvEGUwA6kImy74yC5CVR816fcM83M+l4p96oGSw1lXipfFGVFePH
I+f4mh4Th40dCsxGfOoCwe7CmXBuOdk+pdcejIlYAGfx+Jrzf3E7dwfkvRKAf2WE3yCy9Vp2IDrS
k8xz+XRV33Yfb8icHL0CfDSGWeBWn6n5Mn3IHjsNwI8E7osdHqMNbv3DTsS1CBGkPp8J+WrEhw3U
hd/PlT4kQVm36EiUvpukcqvo1jfLkh77/vyplUT/rjpgzuuP0svrUzbgfhmc8yHJ8q3cwfgJMU9s
xOFp4e65W91s32IIy+GObUKCwKTeyKP2VA8EDaD1M9Q0On5/3NEs7DlH7+sgFKnnN3lZZK2HK2np
xVSWplmESjF7P3M1ygKs3VfHJ3byh3hFED97gttvZi0Rx+xRXLh0EQccJLHbeKAdvSNivj5dzTTi
484I//DMteRrf4ArPtabgzIhHY20DiMDODo5o+QeIdVZafOf5nxKauFKrD47sfwzJo/FdiCQ8o9/
npSX/ZudQAhgFUwhJ4ERsvWQCP77c0z/1g0tnrWyuBYnXKovesSURAAmfgYSAEGibZDBRnNAV9BA
IgJkbzdC7FIen7xpceyhRS5/O70h3Vvx89PzKaiy9aD2hLeYDTShy42T7HoBwCyrfG3qV3XvA5Ap
dqsZ22qKyrdi2ElIGhVF+TRx9kIxx6Jirq9zobATa/OZfbn/q+JV7UlpBrskOXwhiiZQlXH8Iq5S
oaJL9WevUuojvlnQMKJZwR7i6E470drgbUnKxwYLVAc7iM42GQhedutDOrtkiq4CcFD2ObTEfoSX
k85yygQ0X23axD2v4Uni0BNvJUHPH2qP0g4sBI4CxpQlLuLzALfw3kjV+w+ZefxK4e+XouL2aZRg
uPJQY3NH9rXz6Bl9LrUiSp67wviG2c/TzoZ3ywQLUZJ+YxAZAjfVI2S4MrUXWdSDJ58IyY7lwhri
18VqcqB7lQCIPn62cxMhaBDBRewTpWjjwpb6DtcQhVYk2rOOmqY2/bdTdaoTSJ4cGhiGaZuEnfcn
83IhwsAj4KeUhlloxZa3uhqRbRQRTDOg6Y6Yrd71IPnPcKwm9illosTh9vLjVLUFD+NFCfV+vTYR
ApLthk6OgdjL95FBqKPZTwqoALf9TS3HwC4YE8sMqAejZwGPdl7U6+RZEGd8MJy3+5jkivEutV43
ZNEYCqWf2u6+/EdKgcufEDkWgpNyzEUl81X+1yXvtEEFnOv6BqcBFjUmcKAfjnThiyO4aLYo/Hsr
/PtTAPC2xROoC06mnlSxhKCX1Ul8+7cayXjHI5pM98AfjxLu7Xs7V79agu4JxHcDJQ2tflGyrJSc
iIKdqsAAilh0lo45hYNw5p42prsFH4+2NqEb3Nr97nDVuqyysOeHe/XSjMgWHgYNoeRDErB/Zyo7
tOjh8l/ZgwQ0+sGTcStElS+/GoLuksnfgnU/6Ay8Vp+v2ZFXyJ9rUL9DB+1Ifed0ugd6bD3jgUbN
zptLa/MIs1jDaTBlg2LJvwOLQBqnOVX1chc4M9DbdXHINxo2JmZWK6tgsF8hshfmU9iR2GTGZRa9
Z319K30US/6f96TF2G2ptSW7iaNW6FTCS5Gatb4K307SyFil5XDu5nn72k2v/LAItssLj83P3chT
UKFxjVaeOyVd3b6vI45hGeiQv3ME0fM3VWKxLCGLfTVHRK4YR1rkIB45IQkZMhpIJ/yFVPmluFkT
nGugiXNIcciYosE4AewMahY+EiehqYLNAlcqRoQ3kJHLUsZdQtiwP/g42Cn+ojJGVaTX27KhUU5M
E6XloQh55paGqbgDHIn7m3m/Li0FwryFEK0hcsX2uBe8yPY4SdN9S7lW2gZdLT/zZ1GCbeGsI1wD
Djwy2PCwwLz1mzT7D592INJE61MnIjhMzRIIRY7qVMlYGiHTGC6pRulekKc7bE69udV/qfcVf+0s
BBnsANG0W8l3AvbEziTxSBiQEp+iF8+0eCNMMDmAvduAdi7sJBGRkGGKs8e9xsU/np5w/Xr0/4x7
SAC372O026lih4eV/E+KZk8oy+7f7Mln2RrJ5T0SgqJfPFCeqQBB9K54ciT++v1cs6fbO+z+V/79
YHJWqmwr/L2t/74xVXT3BLbcT6ao1CSSLv34I66oLz2RTMX+krFZjMOK2bPSWfxtv43ilmuwkVuY
MGukBx03lbZTkB7CWuLta7E1sNi4VMJzczvIHHXYz2ppfPmPXl+aBr11/dZ58/fSqWDh194kqVCf
PHoTgERh+i0eH/zbJP6ofEeub8bP06fXl3eVSnEplKVqpiwRVTChTBtPbpzsgHDFq3YPqDi0OOKa
mwjzHTfCdWiI1OSG5ognMzq5zfWvoxxJ+ytxHGo3/L3mlONvte7eZZJw6xwD+U6n65+Z//gSQ1Nl
z75M6RjZtjeUVzT5M+0NmCR/M6929IzZ2F9Kv4n8xtIRj/okGeeW2DUKm+8AhQSKemuhwRiH2iB2
S1V5AGoMaFv7C1sg2IQSXQR4IKeJb+gjVNv0LBazXzM4RBwquO9inR4rnM+htAbY1SNc+f78AtT8
zuFT3g5rU1jN86L2D39TSmH1C5SAWvFHPfiSrx6j9+kJdmkJCYDoJW2VCAU65IZ0EH1XAqS34dh7
QogtCwr2ZjVqcfubnWrs9pXyk0duoZ4KMk36WmWNvZSdl4KVFhRGXSAqKyVN1hmuD4LWuqAxBF0u
AB9jaTEMPFfpMp2mV0rl8f76FnRgRD23IwNDo7+JIkfD8OG0UIPifetsVvCwVhwI/V5Pllywph9X
sg==
`protect end_protected

`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Soliton technologies
// Engineer: 
// 
// Create Date: 12/11/2017 02:09:19 PM
// Design Name: LRX
// Module Name: iodelay_n_metastab_chk
// Project Name: WBLVDS
// Target Devices: TSW14DL3200
// Tool Versions: 2017.1 
// Description: IOdelay configuration for a lane has been done in this module
// 
// Dependencies: edge_detection,check_metastability,sync_stage
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module iodelay_n_metastab_chk(
    input           app_clk,			// metastability operation runs with app clk
    input           rst_app,
    input           riu_clk,            //clock
    input           rst_riu,            //reset
    input   [15:0]  ctrl_reg_16b,   	//connect to 2 bytes out of 4 bytes of control register of AXI Reg map
    input   [8:0]   cntvalue_out,   	//existing delay read from HSSIO IP
    input           bsc_dly_rdy,    	//BITSLICE_CONTROL.DLY_RDY
                    bsc_vtc_rdy,    	//BITSLICE_CONTROL.DLY_RDY
    input   [7:0]   lane_data_i,
    
    output  [15:0]  status_reg_16b,     //connect to 2 bytes out of 4 bytes of status register of AXI Reg map
    output          rst_ctrl_reg,    	//reset signal to ctrl reg signal to HSSIO IP
    output  [8:0]   cntvalue_in,    	//new computed delay
    output          load,           	//LOAD signal to HSSIO IP
                    ce,             	//CLOCK ENABLE signal to HSSIO IP
                    inc,            	//INC signal to HSSIO IP
                    rx_en_vtc       	//TX_BITSLICE.EN_VTC
    );
    //STATES  
    localparam  IDLE                =	 4'd0;
    localparam  LOW_EN_VTC		    =	 4'd1;
    localparam  WAIT_10_CYCLES_i1	=	 4'd2;
    localparam  COMMAND_DECODE      =	 4'd3;
    localparam  CALC_DIFF           =    4'd4;
    localparam  VL_CALC_ADDEND      =    4'd5;
    localparam  VL_CALC_NEW_DELAY   =    4'd6;
    localparam  VL_LOAD_HIGH        =    4'd7; 
    localparam  VL_LOAD_LOW         =    4'd8; 
    localparam  VL_WAIT_5_CYCLES    =    4'd9; 
    localparam  V_INC_DEC_DELAY     =    4'd10;
    localparam  V_LOAD_NEW_DELAY    =    4'd11;
    localparam  WAIT_10_CYCLES_i2   =    4'd12;
    localparam  HIGH_EN_VTC         =    4'd13;
    
    //COMMANDS
    localparam  READ_DELAY		    =   3'd0;
    localparam  V_INC_DELAY         =   3'd1;
    localparam  V_DEC_DELAY         =   3'd2;
    localparam  VL_UPDATE_DELAY     =   3'd3;
    
    
     wire    		trig_iod,
					trig_iod_re,        //start iodelay trigger
					trig_iod_re_dbapp; 
          
     reg     [2:0]  cmd_id, n_cmd_id;
    
     reg     [3:0]  state,          n_state,
                    clk_cntr,       n_clk_cntr,
                    delay_addend,   n_delay_addend;
  
     reg     [8:0]  diff,           n_diff,
                    read_delay,     n_read_delay,   //delay read from existing IP state
                    orig_delay,     n_orig_delay,
                    new_delay,      n_new_delay,    //delay to be updated
                    user_delay_i,   n_user_delay_i; //delay requested by user
    
     reg            load_sm,            n_load_sm,
                    inc_sm,             n_inc_sm,
                    ce_sm,              n_ce_sm,
                    direc,              n_direc,
                    delay_read_done,    n_delay_read_done,
                    rx_bitslice_en_vtc, n_rx_bitslice_en_vtc,
                    reset_cmd_reg,      n_reset_cmd_reg,
                    delay_modified,     n_delay_modified;
    
     wire           error_sb_riu,
                    error_sb_app;                

    //edge detection 
    rise_fal_edge edge_det_e1(
        .clk_in          (riu_clk)  ,    //input clk
        .rst_in          (rst_riu) ,    //active high rst
        .signal_in       (trig_iod),    //1b signal to which rise and falling edge to be detected
        .rise_out        (trig_iod_re),     // output pulse of rising edge
        .fall_out        ()        //output pulse of falling edge
    );    	
    check_metastability check_ms_i(
        .clk            (app_clk),            //app_clk
        .rst            (rst_app),            //rst_appclk
        .rx_en_vtc_i    (rx_en_vtc),    // in riu_clk, to be registered with app_clk
        .data_i         (lane_data_i),         // reg in app_clk to match with rx_en_vtc
        .error_sb       (error_sb_app)  
    );	
    always @(posedge riu_clk or posedge rst_riu)
    begin
        if(rst_riu)
        begin
            state               <=  IDLE;
            diff                <=  0;
            load_sm             <=  0;
            inc_sm              <=  0;
            ce_sm               <=  0;
            clk_cntr            <=  4'b0;
            cmd_id              <=  3'd0;
            read_delay          <=  9'd0;
            orig_delay          <=  9'd0;
            new_delay           <=  9'd0;
            direc               <=  1'b0;
            delay_read_done     <=  1'b0;
            rx_bitslice_en_vtc  <=  1'b1;
            delay_addend        <=  4'b0;
            user_delay_i        <=  9'd0;
            reset_cmd_reg       <=  1'b0;
            delay_modified      <=  1'b0;
        end
        else
        begin
            state               <=  n_state;
            diff                <=  n_diff;
            load_sm             <=  n_load_sm;
            inc_sm              <=  n_inc_sm;
            ce_sm               <=  n_ce_sm;
            clk_cntr            <=  n_clk_cntr;
            cmd_id              <=  n_cmd_id;
            read_delay          <=  n_read_delay;
            orig_delay          <=  n_orig_delay;
            new_delay           <=  n_new_delay;
            direc               <=  n_direc;
            delay_read_done     <=  n_delay_read_done;
            rx_bitslice_en_vtc  <=  n_rx_bitslice_en_vtc;
            delay_addend        <=  n_delay_addend;
            user_delay_i        <=  n_user_delay_i;
            reset_cmd_reg       <=  n_reset_cmd_reg;
            delay_modified      <=  n_delay_modified;
        end
    end
    
    
    always @(*)
    begin
        n_state                 =   state;
        n_clk_cntr              =   4'b0;
        n_rx_bitslice_en_vtc    =   rx_bitslice_en_vtc;
        n_cmd_id                =   cmd_id;
        n_direc                 =   direc;
        n_inc_sm                =   inc_sm;
        n_diff                  =   diff;
        n_delay_addend          =   delay_addend;
        n_new_delay             =   new_delay;
        n_delay_read_done       =   delay_read_done;
        n_orig_delay            =   orig_delay;
        n_load_sm               =   1'b0;
        n_ce_sm                 =   1'b0;
        n_user_delay_i          =   user_delay_i;
        n_read_delay			=   read_delay;
        n_reset_cmd_reg         =   reset_cmd_reg;
        n_delay_modified        =   delay_modified;      
		
        case (state)
        IDLE:
            begin
                n_clk_cntr      =    4'b0;
                n_new_delay     =   9'd0;
                n_direc         =   1'b0;
                
                if (trig_iod_re)
                begin
                    n_state         =   LOW_EN_VTC;
                    n_cmd_id        =   ctrl_reg_16b[14:12];
                    n_user_delay_i  =   ctrl_reg_16b[8:0];
                end
                else
                begin
                    n_state         =   IDLE;
                    n_cmd_id        =   READ_DELAY; 
                    n_user_delay_i  =   9'd0;
                end
            end
        
        LOW_EN_VTC:
            begin
                n_delay_read_done =    1'b0;
                if    (bsc_vtc_rdy)
                begin
                    n_rx_bitslice_en_vtc    =    1'b0;
                    n_state                 =    WAIT_10_CYCLES_i1;
                end
                else    
                begin
                    n_rx_bitslice_en_vtc    =    rx_bitslice_en_vtc;
                    n_state                 =    LOW_EN_VTC;
                end
            end
        
        WAIT_10_CYCLES_i1:
            begin    
                if(clk_cntr == 4'd10)//cnt10_1 counts 0 to 9
                begin    
                    n_clk_cntr  =    4'd0;
                    n_state     =    COMMAND_DECODE;
                end
                else
                begin    
                    n_clk_cntr  =    clk_cntr + 1'd1;
                    n_state     =    WAIT_10_CYCLES_i1;
                end
            end
        
        COMMAND_DECODE:
            begin
                n_read_delay        =   cntvalue_out;
                n_orig_delay        =   cntvalue_out;
             //case structure based on i/p command
                case (cmd_id)
                READ_DELAY:
                    begin
                        n_state             =   WAIT_10_CYCLES_i2;
                        n_delay_modified    =   delay_modified;
                    end
                V_INC_DELAY:
                    begin
                        n_state             =   V_INC_DEC_DELAY;
                        n_delay_modified    =   1'b1;
                    end
                V_DEC_DELAY:
                    begin
                        n_state             =   V_INC_DEC_DELAY;
                        n_delay_modified    =   1'b1;
                    end
                VL_UPDATE_DELAY:
                    begin
                        n_state             =   CALC_DIFF;
                        n_delay_modified    =   1'b1;
                    end
                default:
                    begin
                        n_state             =   WAIT_10_CYCLES_i2;
                        n_delay_modified    =   delay_modified;
                    end
                endcase
            end
        
        
        V_INC_DEC_DELAY:
            if (cmd_id == V_INC_DELAY)
            begin
                n_inc_sm    =   1'b1;
                n_ce_sm     =   1'b1;
                n_state     = V_LOAD_NEW_DELAY;
            end
            else if (cmd_id == V_DEC_DELAY)
            begin
                n_inc_sm    =   1'b0;
                n_ce_sm     =   1'b1;
                n_state     =   V_LOAD_NEW_DELAY;
            end
            else
            begin
                n_inc_sm    =   1'b0;
                n_ce_sm     =   1'b0;
                n_state     =   WAIT_10_CYCLES_i2;
            end
    
        
        V_LOAD_NEW_DELAY:
            begin
                n_ce_sm     =   1'b0;
                n_state     =   WAIT_10_CYCLES_i2;        
            end
        
        CALC_DIFF:
            begin    
                n_state    =    VL_CALC_ADDEND;
                if(orig_delay > user_delay_i)
                begin    
                    n_diff = orig_delay - user_delay_i;
                    n_direc = 1'b0; //DECREMENT
                end
                else if(user_delay_i > orig_delay)
                begin    
                    n_diff = user_delay_i - orig_delay;
                    n_direc = 1'b1; //INCREMENT
                end
                else
                begin
                    n_diff = 0;
                    n_direc = 1'b0; //Do nothing
                end
            end
                        
        VL_CALC_ADDEND:
            begin
                n_state         =   VL_CALC_NEW_DELAY;
                if (diff <= 9'd8)
                begin
                    n_delay_addend  =   diff[3:0];
                end
                else
                begin
                    n_delay_addend   =   4'd8;
                end
            end
        
        VL_CALC_NEW_DELAY:       
            begin
                n_state         =   VL_LOAD_HIGH;
                if(direc == 1'b0)
                    n_new_delay = orig_delay - delay_addend; //CNTVALUE_IN
                    
                else if(direc == 1'b1)
                    n_new_delay = orig_delay + delay_addend;
                
                else                    
                    n_new_delay = new_delay;
            end
        
        VL_LOAD_HIGH:
            begin    
                n_load_sm   =    1'b1;
                n_state     =    VL_LOAD_LOW;
            end        
        
        VL_LOAD_LOW:
            begin
                if(diff!=9'd0)
                begin
                    n_load_sm   =    1'b0;
                    n_state     =    VL_WAIT_5_CYCLES;
                end            
                else
                begin
                    n_load_sm   =    1'b0;
                    n_state     =    WAIT_10_CYCLES_i2;
                end
            end
        
    
        
        VL_WAIT_5_CYCLES:
            begin    
                if(clk_cntr == 4'd5) //clk_cntr counts 0 to 4
                begin    
                    n_orig_delay  =   cntvalue_out;
                    n_clk_cntr  =    4'd0;
                    n_state     =    CALC_DIFF;
                end
                else
                begin    
                    n_clk_cntr  =    clk_cntr + 1'd1;
                    n_state     =    VL_WAIT_5_CYCLES;
                end
            end
        
        WAIT_10_CYCLES_i2:
            begin 
                n_delay_read_done   =    1'b1;
                n_read_delay        =   cntvalue_out;
                n_orig_delay        =   cntvalue_out;
                n_reset_cmd_reg     =   1'b1;
                
                if(clk_cntr == 4'd10) //clk_cntr counts 0 to 9
                begin    
                    n_clk_cntr  =    4'd0;
                    n_state     =    HIGH_EN_VTC;
                end
                else
                begin    
                    n_clk_cntr  =    clk_cntr + 1'd1;
                    n_state     =    WAIT_10_CYCLES_i2;
                end
            end
            
        HIGH_EN_VTC:
            begin
                n_rx_bitslice_en_vtc    =   1'b1;
                n_state                 =   IDLE;
                n_reset_cmd_reg         =   1'b0;
            end
            
        default:        
            begin
                n_state                 =   IDLE;
                n_clk_cntr              =   4'b0;
                n_rx_bitslice_en_vtc    =   rx_bitslice_en_vtc;
                n_cmd_id                =   cmd_id;
                n_direc                 =   direc;
                n_inc_sm                =   inc_sm;
                n_diff                  =   diff;
                n_delay_addend          =   delay_addend;
                n_new_delay             =   new_delay;
                n_read_delay            =   read_delay;
                n_delay_read_done       =   delay_read_done;
                n_orig_delay            =   orig_delay;
                n_load_sm               =   1'b0;
                n_ce_sm                 =   1'b0;
                n_reset_cmd_reg         =   reset_cmd_reg;
                n_user_delay_i          =   user_delay_i;
                n_delay_modified        =   delay_modified;
            end
    endcase
    end

//---------------------------assign statements------------------------------
    assign  status_reg_16b  =   {delay_read_done,error_sb_riu,delay_modified,{4'b0},read_delay}; //1+1+5+9 bits = 16 bits
    assign  trig_iod        =   ctrl_reg_16b[15];
    assign  cntvalue_in     =   new_delay;
    assign  load            =   load_sm;    
    assign  ce              =   ce_sm;      
    assign  inc             =   inc_sm;     
    assign  rx_en_vtc       =   rx_bitslice_en_vtc;
    assign  rst_ctrl_reg    =   reset_cmd_reg;

//----------------------------sync stages------------------------------------
    sync_stage #(.C_SYNC_STAGE(2), .C_DW(1), .pTCQ(100)) 
        sync_stage_i0       (
        .src_data   (trig_iod_re),
        .dest_clk   (app_clk),           
        .dest_data  (trig_iod_re_dbapp)
    ); 
      
    sync_stage #(.C_SYNC_STAGE(2), .C_DW(1), .pTCQ(100)) 
        sync_stage_i1       (
        .src_data   (error_sb_app),
        .dest_clk   (riu_clk),              
        .dest_data  (error_sb_riu)
    );
	
endmodule

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Qpo3AJT/cKwgSuEvbp/4RWbnB3sjV770kHb+XXi2uMhVZW3uQU1fOfqEow6SjKm7ePue+L1kNzUt
PBuo9vAS3w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NCveSwNr/VXXcn4TF3W9pn7aMafXhv6qIlJ+QomdzYQidZ7xp8Cpya3GfvkFBs+5BEnuunoxrizJ
KRpMONwPu5Va9XcFTHCq9KQCsZ7oIUc3Pk+/YRFS6Jk+8kIhQbjaPKpufXa8qNyxKaYmgGt/8Fil
6ktI0A7aFF39EYblmqQ=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
A3W4kzxyVve3BBoYMw2VI7YzWGfguGkOb0N1x4EwpKwnfY7UsAXOVq4t3hZy3ilOFv/xzpHjQjg8
5G4oZfoZsxiePAz5x16ZHPVYw2GvtLAk9yA+dwbtwzrnVAXImM29pSOGwD9e746RhprsoPpIy6wL
nPspC381e/l5Eu0ywF0=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CcsIEDN/mmn44yljCbnNlwkLDonAulX6jak88ukqQRYe/DVzmMLOhttFc0vJWQaTu8vwxM8VIIrR
0hPLWSKELygGWFZMmikDyTo++Y/ZMpP54c7fzKvPUwswlotX8DXKa7hNupAp3pzAzfPpmbBBp5SE
7BseC+8l/ARw9ao8KQosM2Z9jLbFzGhhtZsqN8jsjdF46ad+elp/2yoK1gOTqNq3EB017LiEtE2v
H9f0rcT9tYESd2yRZ2H/u6j6mQPxg0djUkCtUObs3Z4Y+KkF8Uow2dMdW8orV2e+tnnve00QdGrA
pb85iJT1+5sB8b7VIjShJqk7Gc0yPPxQkq9CLw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SCeLnLCJxqJlc+H8i92PqkoIMkYBjH6C1nnHWwSc4X6XM0TCdIwnOucilmxUuywfSxrZXYf2PmpS
w1Wy5+QOdHG4mOqeK6Pdmm3y2yphvfzivf7qCzFeYPrVpn0Hy3bioCXKb/RR9lRfY4ZIFTj7XDen
srcXa1PBaNnBGbYTNFMCCWo61UVIkNPsbzkPTyzrlqiVRpPGmCszoNiSIXGYjMezDfAkzKvQJclt
fUix03YVA7iY1o++BNau4ziaETBdp8lOm9LeR3uvJO161WnIAYg7U+PEQPwvonH8wwx8nKX8UeFa
h+7jLbz9DodkL226TME+T67lyN3vOgSf4rY+Zw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iFk68b8RyLUljyVu4Wrn2izKMOSr9l97Mr6Sf28ViOgVZH8CvTtczGhoJ4JChfmX9/GzxzcmlG+c
vBMyhEg5w6L4cZcvLD05vq/+D1fbjOYz6l2TlDnbhgYxmA+DaqAwU1ALhYK5rJJWzebY6hT7vxzg
H9ULXBMsADfipi361s8kVrI+OKPcCNThWW2Vngkcm//JlfkBSNpo6pB9zbh6L2sM7eaVrhYWMYQw
UsUnatTxkpJn1j/Xa1GF0XTupRb32B/bIKq7q4N7whljjQGhX5FGzt1fjh1xATXCu7z2xAUS62hl
8zWvM/1b/d3cQe33qWZnTm5/slNRqfn/kuUhcg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1051216)
`protect data_block
YBNVUnfApaCCj46QqPsmGHHnK6qQeSTTmIPA7gx38yBEelpplzfxwysi1un+ULlmtdpsVvKCeKNT
8W57J8ITXATIjoWdHesAS7Bxthxopc8v9jdixiNG1jtO/j8kT8K5SIt6Ff8AhN6x/srQfahLobMs
m6Pu6nLh7hqh/iTD7b8FF8WNFSEzsFf5LApfoL5j7kNRYve4n95KjqYxNga/FrhWD1WhPMNXlqyj
Z1x6rq3QGqckCH78kaipJnBYHu+OqPN7Ss/MAtjH5hfEUSnPppyaGXF0AoCHoNRI1GcpBOrYkYRv
6SMD10or3qxI8tArXg7nD1Lw7Yqhm+2W/WEGiyeyYUDIOCmdjURVr5piABT/PUzTKS9eoUF6wbT4
r/g3TDU1P384f3AsR2+X4a4Hfzp8L877h/sRWx8fxClK7BiKJt63IWa/gn/Ul3AedRRF4aey+D4U
ZSdx8+ZUH3G5dmwskZmQoFk8Qvpq/DEHOIqY1b4jSAo+2YZtEgbFe5tkTaKnxfQGYnT+GAz03Gl7
DEnshMNoBQSqSctkavcNW38EKq3xf4HxU4EoMmzx/wH1kcb2lT13bAjHpGMjuk4KkYP2+ZVZZk6g
W8RQAK1FY88lWrzBzpHqE+wtBKvBTFDDvtgSAPTsrcA9mOxtHIpgG/Hwpnxx22ZxRjrDf5NpXUy3
yK0PaXzrkZX7qwmz+qR2A6qtcaN52cTNCQ3h7NZQupRZFqTdaSvLxR965Tyk3inYnfT2JV5NSTZJ
qo3qjwbyLqcBhhquJLl86NSl4LWA30o41Z22yQRM4VPQrdTFPrdNsdKUWAdO/dHQA8q8oDCfzTbk
gWGDbjnhygn5aWU0SIfH64Gq1DEF4v1Qrm6mBt7u2AR9uMm1O18KOiFV3Km+gYacQ+az5HgSfMBf
DwOL4kRQXtvwnIM2ao4Hxd54MebFKf7KFA/9ppYURq55woM1nOE5zsuYu8p63rOqNiK2cN/H4sXr
OPkg6LKHFnF+ZTR75CRXc89VqEPYSbpfljAPGgYuV7jX+bQAXsCN95EsPI+R+D0eRB6GhQJrHX5O
X9eAaYCy/fvJ9nvrUEAUNPye7Yktj21CNIGhZ6VDSi/7WSd6YKsFK88tnz1WrHvptAVOUP/Uj0Pm
lFMIiXPii6tZkxhVe8cDKuGtzgi+HWjHCgIofTt4hoEa9VBWkg75M9veQH6CTpVQkYFrwVEVz5OJ
ieGBvN3yVeb8saH5h3WWxsKvwlr9Zav2l/4Ryt//Etm6hSzRrFSc9WJlOGUbyh5/MKnFF2z+h8eX
Q5EOPL/fssn215KPsI9sjof04VW4lZnBHj+0+WPJzKPxWlNrlt8Qzds5NTlQI04GhyK5LTGMl6IY
H8829YE2Rq+fdefDomr/IyWsB7fvRQjCDs5XFMTp0cW/8NGtTO5uf46oeRy6Zn75KmDSsBKRiZZ2
lm6+yyh5CXVgO8ccd6ZAF87gJqvAbkD1dchylKS75VFMSX0EvytXRWM/gj36e3YfxR0+Qghw3ESN
qemyfsoCAIdTVloYhKXWukexzj9pUih8a01OZ9kER8E3DfQXs9a1/XOe8NmK87MNYE8ybx9Eifg+
k9FRx1AKuPHim9B1+gEc1LG0u1fqRFXdNDe8PaqRROuXp/ti7PSRCIxc8nj/yjVae+ipGNaikOW3
LvCktK+sirnAu1RI9Ebs2RaCmrNpDujsIA8dBfNnXG9RG0rAReLfEYHb+ZPJrb3FWVHt4V5b17oC
CmxeAZvig84A2ERMwkJy1TrdrVtdFUbh8aW8ereeDRCM6hLN35uzZQh2dP/ocheThsOT2hrCFaj+
WzXrMJ2Cm86hoRc8EjvdLMPtUe/CDtb1lg4R42zj1IXOwZspLIHPMVRwpK4987OjH3gXWMp/QFRM
9YFoQzro2+xXUkvQsCqKiqxYbKOg5ocPDH4iMide0zh41l0lzxntUvSCSvAhrJqHUh7JoVjworVg
mHGTSzvWAIIiI9L64BIt+Wu8Uy9B9/lQoO0+FetW3Iyxd1mr6XklT/bnzbunMzJy9shrkj2Xu5bm
Sbqwb16nFxt6W1Sl8vJTcsP6sx5xsUBjhApeg7NbJs+RaNwYYFHfm3UCnAwwvQz0oHnd22dUzm6j
aQyIXxPkpIZuGm9UhmMy4knlRErTebp50V1yJBZJQqwT6azuxqwPrT/k/R86GULFauGUwVFzNzbB
xXNFceP2LrjJJvN61hv2/IN3uSLKGgYTsjDrccqx7TKNxmaBUI0aRosW+NG5BMLHXyglEivlJr/B
uJKoDdFBqkiy9u3VkUFWrKJhCBIJss8tBlC++9WXmXLxcls/8i0oSVYRPtzWxqmsSCZ6Y0gtFI9r
pcR0yhiYZLJIQJ54MODVdESS2IFsxHbhHpWFkiZH+l3InZhSUUnjpPL5uO1SJxeFzE5VYQ2a2/Mx
DCmGGsUJ48/R/zdcO5hE63YaBctbTLQEDhQq9hZySRc0XQxTtr/QkPwWv9jg/gJ3BQhw47TrB8IQ
gv1k3xpCWdHGPFtFLQEFY5iS4UoVs3HO0u4zRvO5seiimtRvCmQPATFCl92J+Edbhe6FRv/XrLqh
8ATcfy+SNUuZqmN1+GjSk0nrQCKZfPxro/nlaAwDQHwDUrBnLnpEg2OUcgRTIfgtqaze2+o3iQWa
CA/1mJrdOz/5mGSJi74P6arO7lK5A/VTW4M/CU8IIvy8N/TVbK14xRzcFuZqBKCGGAuljuuE5ssS
JayUYkDxoe/5hucC8U3gd5otlixr3zdThfFnTr92QtNL7hE/2hR27wiJ1/BTQ6g+3ULmeV/XCfxK
WU2Q5ydfoiMejZyjIH0bEDEKhE+l8vhCFq2f7WpSvMn3aaRqOrstCYQ09cIQWoxN0UryO2GMrtYt
cNr1Gpzf91cNv6muFdQbov3LiCoM0KHExqgRI4zXHi9EAXNywyfl6+fUsGHyGo1WfpfXJCtw8evH
fNrjjcGb5nZiI98uldmEQBZRt6hNMG3lPYCKriZO2etmRXszLvBo2wl84eoMqTD03lwUYMQnw0Mj
8+cltuqPAKEqjhKr6oGVoIKOoTeuXFCrq/er2wE9ncFvzkXZ9i1sxzMrPGFHXr73T7NyaMUBzbJd
qOqmbN3VuH9H3TRqiD+O2YalrjiJGvD3J4uTcDauZ76N5guDQLx8BU+7UCS3FxDQ27wpl7Qqdl2X
YgGaPrxZi9NAypZykvoG0HnXRLpZ+T1M1AfKR8alhWyjHyeuIAs5axObJufZFUOiPRw4pQjuZf4b
alMeVX4lWS86LtztK8cI8/T3acElwdHti9GB8lyOQYw+kt6Ti74YNYnX0WI4F+YNZQwFFJY9zWnz
vQtZ1ENZujVl91WNiAHE/ifmiyk4iHDf/AmoHLxJsLbz/6mPgXGayFhfGqTtM7W3AKYj81J5uFkB
hGBxsn5FhUOfVh4chT9aZTKgd13Hy+cY+tM54Nojv8UsCe0sL8R38fygS2EC8bVc4wLCYAheSxfc
RDd/dYDF42ynkvvvmkximzHGAKk3nZgXAkZ7ztf9OmOBkbtBeojfAKHi+6XU8PojJVCI2AjKQwNZ
an/Gkt8viH9JcniFatyv/aWfTkDxIi/ig32fMwO9lIbqp9b7VBX7huHFdsfOwCVSL8fP1GAqZOkD
51mR2a2JqoSdEIfsmn7JmWwed3zJ7PuYhzzmiJQEh0DUeQ30NXsvkvVG5by+rEpSRxT04ZVGIZt3
OFXJktTGfrnHTED5Og/MTmGjqtHYiWjzzJiHCcokrMw8miVC6yKsFgWy1fW578i/zTDOiqN5W5Yq
La6xQ5qg55Q/5Q2hnoDWXrQ4lbxpT97H7hVLcagdmuxiA4EQKSrSc+Bs7inxmtKvS1lF0TBDAjap
s4J2KTjsneEPYcc7Y6yEy1olicmHV+KYos4GYna78e6kl8CBMDejaf78fgA0wELr3orNqFt/bOgd
/Yep3ErV15RBCM3cExQT6xxST4WVJgOopGIkRGjcm12k4Hy4KVrHi517LsOwLoHxPi/iV8LI+Zv2
gRdhok/uYohIRd+2uyzN6UY/jZF0NBTIW1ByXMvAUM1dOfFhwaevarxa2Zs+Z5g8AWQpc7W4I9xB
rnmYuKvYsDB+vyJwMROQt8CNzI1BmXiFN5lN4ByimY4N+mHOBIa9UeSaMCR4HBDnGcMH/Jf1aupv
aQLhMNIT/R4IkJG/wquAD5xG8YC/rrlvJIVqAPgSVDffdLFHUToPK6hofWGcl/xmDqAgx3qwMpzG
PDXSAxwBTn0X5H4yTtyMRxnYF+qoDinZMNoA5NMhNvBEOOkeDDDdx7rKi2CPuF9O8tA1rpqQbWyw
rXLalP7DjTTie877kgWWBzdgBPH+FCvYFjn5yszeK0i8h4Gy4zY4pnO229rRN7NZHv6zdbpNaUbp
w6seyQvpilsIcThmn1mGmprbQW2k3FvAXuHvVcAdD0NXRqSVRe42eCoFkmZ42CCos3T3XfRIko/P
c7ElFLj7m1YzmPnvi7HKJ76phFf8sV1A2W/0b/wVvlNKsV8U8m6dvzzM2gg4wCKB5+IoMHO0nT3c
NmTjQrlW0yU1PSXyJ6GaBuvtmmxrusGc4sSv20kNFmAG/oMXj1rG3LZujN+g5tNxNUcdvIc7YP6c
CXftLpkqKT62QCANqfWwEah+sNobjj1kyE238I60iaOYYd05r878XlswuN3smgkStJJeIhTh4qUK
vN/giqO9ekmCJ9sNG1K9wgXlXpRvK5BkmS5yL0vZfmBA1Q7zT4bft7aTRPMM5lkhBnnGAUD3xyyl
k+EmoZJIzkECzj6aHchr3FF0hAoxmHT4rhv7e389dl63cqUh5rNYpCQrlsZXhpC8OMYjsN+RvezE
qwpWpE4KmIme+f0LZ+Eq+Nt4+floUJWZK7YlTN7OkWYZZoCXxwkM+Gqzv/9+I+fA2Av5qNIqus4V
NpuMQ4bM7RtuvsNcR2yeHAmRO0/HTPbfBbwW8XI5VzUqnlLvgC7SUj5gB+rZ4e4bfNXXQtFKzzXF
mjNmcWRBwgNTVFeaO8RPDY2GH96Xd0GzsUOku39Cos/4j//zcicpRM35rL3cTAQo8aivsUH/4ooy
jbiiE4yxaoTrQttAXU3QGzKTmo0mygGctUs7/DDTu8Pb3a0LfcNtK4xj6fVSJkbc7OKMZU/nzk5u
2DQcLXhhGMe7Pzpjs/JvKpSLKPoKYNC76M7HWKEiNyj5vbsx86MU3JgO0ycVU2cYFexRnlU8gQtV
d8f7j+FklCcSYPZ4arDNSeLaoNQqty2L9ojd0gqf/07WTqOhl9ui7CmIc1EWZ9xJBXNEaDBF+He8
pmAGtjvav8qLBOerozPKb+e7RcqysieuI28le+R3AyfqrRJBE3NcrQnZGDMVs4oeYBIkP+53/eZA
Qjzd/MgpSTldJNLSNQXdYp+Xa8GIlKMPR2rZ45rnIUSnPwiL5rdaxasNKsQ8UYUOqvTUmJgsTpXX
S89qgAeiE0W9LmSgPEqIK3TI7wktqf6JKz8dv3kD7iasOPVt6dyD7eUqJhYbDBX8AWF72+vzS9RA
CwMNUEzLYzMzCcAPlBGuVHFR7hX2n8TMJoyFKXpO8/E1avgqCY+YsObqLHn6fO9KG4vXZ/636PgU
J4DJ6UhfdJxooL7jxOapwW3leHnrGvySLcuEGpvvkVi7h+Uk/GWZCIEfJjtPVp/3hz54x9OD51ZN
RseIvoAiS4+v5uXH26nfUpcrvLbnL2LpPEIMj5hDJNDbXSLrx0B8QHIP5LlAAMn7NYnDbTDs7s5p
MEOA/KNtbYmNaQUVRNXpCZDB/34EFdITQA2DvZ+Affaf8a3lXYFGNvT1QXErGlSxkofywoBllta3
ird1NpQWbAuE+h6oZdBNF2J9KzMHkPfkLD5XmLjz0ZLdf6U7SrNiziblEU3AhdOsJvpJFaMxdjsU
ePUwn50aEnRCG7ZtgZDw4ydKspx6qLhbArzMbdaOP2hwHQWXM+Zob4jQ+ODjYn6zfvQR1sm3Ix8w
wsO28xt3IxB9E9T4BD87LTDYYP+BOIpyZj8VBdBMRhaNyMecHzBZJFGoezrIKI+kpGwPfrgzdFcJ
8a0oLF6D+FB2N41pFI6MPabOFus8NOhwyFtlNkg9ot3HQn3GlBooZGdVY2v7tyjXdh2mq13gAgk+
7zZ9XNUukEdmrl7LzAYF7Pa3StVwut1NKptVBuLVLOHYAWEcbTSlQG2iQYi0Jx22SL+EMWYNmWTJ
0NIqVdjpStk3rW93c2hnnusbCipBeyq3PjrZ9QRT1//Hx2elzbXF9u1FQErOrSVxDAxWOe7sbEKu
a3Qm1vQ1TT2rQEFOgoFWaE3TXJuUXX4VBr5QKrCgI+wR0EDV6Ri2N5S1tXvxJ3dk55xR2KxvkewL
/bpONz3SlrXDH1sFPdyxz7D9/01di8bWhbkxAi/YppB30IiPi7yDEMnljjHbp5mjI86NaahrbqM/
bqnt0T63ZgDhFgUDixXYuPcelxyuDW3w/WMDPIhG6bENRgyvRZZri+LOhCYunoGIEhvhFgJit1p7
waCIZWP83cikW2ona6580au5ZdhkMfzXxvh0Ldg50EhoL/x8G4sKJEivavY6jkDw8aObgSGj7uJZ
ozMAlCr9WXOmbhtQZXthSN0HVaEm2kr1xks7JYmYkEvT4P+3gA9HjoY3Vk7MVMUAbRpBogoPywVh
SexNKTIPYqvxHWk25s012MVrY9Y44dzcXC9OwSINEAIeXZndkjcbTJ6OnTpRLLnAo5UsoFnzTD70
WFDChJI5CTcQlGbMWDFQsEnUFjieAf3UP8kwCKUSFdpX0EO1ddNHIatHmjM9zqNzbU3OKCyTzPSu
nmW5RQIbGf0ZmFsGzAD9tXZLkIbpcBOoeaO3BVxHGlknSsVujSgMkWFo3aTP065iwg76oRabvZbF
djLMTGilN8159z9yBZauhHKytLB0eqwr6MIr0Oql4xW/Ie7PbSpoYwP8cdWSgLC+2QjoUaDw217G
JP+f9jLNNWZPGfQf7xG0ff7Olsan8vNtbSoNJCD0Ov60pDrIdakG0e7Fa5snIbPlooLpeH9zUXOs
dgYxa2+1lcRw8m2fGD0vPIJLPMU/ZstkCEDAEuRU0R8BF1NV892s5ASQzvhblAkRtQu9mB83oonQ
Xqu8YDcvPXsLxeHlOfHLU0HvJv8Po/ZsR0C9M61Loots66oOLkM67fdxTSHaS8c0LfIZvlcmhZnv
EbztWqc2QJ1WXIE5p3I8GMD2t+QBOto2b5Ud1975AzgzaUn7FZB5kFIyeqg1aqlTIyjoPzvoJ2mp
7HTuHY50Qz2CHwqb2nbWg6n3RGMjuzE1YtFLlui5gVqJ6a/yg/wwpsjg7iX81M77PwJJ0T7FVEGR
S/I522WClWBDcTihhp823SycKkumevxkvBxNMBcsk4vufghgWxY+BmZ4uzrBFijRJ6x0NJqxtrrO
ii7LKMXgZkgKJ2GA36gSo6vfFnFTp8rrpR0UZUH1pciBgtZNzcyzlp5U/qQAkPXgGqOZriAPWS/+
sNY6TX5zZZjhYfo1hZJe0v3je+zi9aBv3DM+gUxAMN7SkPKSbBRB9StvFGubOO2wcIlbD2TuxCgx
1BKYQqeRmr+JBF1EhhbrBjnlZVFRlbpqMX9UquLhQ7+UJ0ZTP6ecW1e8N/w2x65fo/j5lIyzFX1T
AzsM5YFXswK9+HOzt6HvijR5K8kh9QNs5mEVs1bQYAcCBUrFv4/9+J3VEEihd90mhVsvKtj9aZMI
tF/2YZvzO2lC2wfDDoNcR8XxjTTPaaqqN5KEaRpg97JELyPn7otQUNQFqK6bmQDoykDzLap6kTEV
uwYM5LXshUzYRtGmEPqFtKwvKUkCs0kyAn2TOWleH0ARpX3V4Ed5DMVwNYxhIIM8co3y+TrMXtH4
CUFNnjCWdcNWYi7niwjsdwq4aeQsQh9la5P/gsAAtN9QrhrwwusUC+D5ICww1mTYBLWEWIGXhtgP
g3ajwNVlG3NBpUxAh9w98iJbyVyW76Uv2+2Vy7CLg3VVGBDi5Kaa9uDJav0hFD3q5kisp+IezP0O
UdJXS/2NQdB7fORvk5wRZ7tjqYwTbD+19sy6xfq1HdNEBoXrEOfiK25x1sGfw5Yk6BkaHQ07TmN5
CsJhJ+AmuwCC/IDLPWm5J2o03sqBTmUxDrS2dS0v1r60fxdLjyPZkeCAJmw0GtnOaO7MONtZPVMA
D/3pEsq6yAmWmh36hLJ59N7YFvZzUmnXX0dz7N2xH1UUP1ae76RZNaL8RLozRd3B1YtVmJCcbpTB
qYTgBf3ZGdpv5z5JlU+X52ggIumn59IZZnIB46L1MW+qEaBiB7ke3MEf/MBofEsDQZNaWHPbrUQl
cqpcJhmKcK5QKhCAfdNE/PkthKkn+Ne2MabA2tMJzX0DahXwl42EqeoHprNyb5q+vPNhDg5UPvf8
ZI/l7lAIjRTdS2i0pu5iLANrucfbACwKFk3VcTCOzfjqJTMPT0Z30eBlACOoah/wcp652/BKqaP2
WPBAJk5zFRo6kFE815J3WPkR3rF0gQ2BbZK15V5A1gCYfKtvbWkU57zr0rfpHuVwozHPTKzfBESk
mRiH5bX3uz91YrxH9p2Q1LR47kEPjyihyPXXwTsfQvAJazjBzGx/5zHklD4QV/53H+rzTaIvN1SN
rCW+Yk0o+6Lu3KpNi49hqQToOo5gTIxCFnv0Ikw+nwP7jdnU6HQuuNkNQhEJ6FMAG6HeFk2jlZJM
DSAOdC8t5zpKIEiYFhTVB/X5digvBjXiJpTK3cy2bfP51hUhBhqUUitHa98+RxEPcroF38rF9CVN
ymb71pyFlkg2iLSgzw8bh2s0IIxF+AgmKVdZgrO1C1FtjX88VHOy/Id6iSgGwjfqtmvBOZ/vtKFi
08mGOZWkrmEiYX3rGTcqvmteH9E0YPzEmTjYWypmO8n20tNPFmmJbP1GQBFjB2KVSEK2TJUK16ei
pCd5E9OeB4Z+MRqwQdZEr+3mAKeNAPRrEWK50Z+cSpzJw3VqOafU8DgkmM2ISdZ0mBcOAvwZ9eJV
ZhNs/yZ1PjGs8pW9QINGS9ulAWvvPuCl59o0eFleE6CesPtPJFSxCRSCAwqiC7Wb9NkpU05IEqdf
qnfz36HHzlveqtc4r+kC+sI9sciotu8WmwyZNw4adix7WmRFMvheWyNa9RY7Q+1T07Wf8Stg98NP
MOiO14M/ac+hSOAMluifoOOMr300gh9jC1clCYhDzwU+McBWl/6TAgZliMagiSFmMXIYegqkM6ax
uz7utMvz5GkOuPHtFDLbTNtLC4roILm3JKPLOlI4OeQao84j15XvRgzWnLtZR+yFJGSH4VPTBS9J
Jxu92i6hGgQh+N140gN5kftczj/Hw7OUfG/404icySbw36oWpwH3KNVXeMPpj3aW8/W/+kEHZISw
vB+JB9USaazTots4FWTdh83gQo7a9tTlSMxkP3GlgI4LpwT98H4a6Ji1ip4Vf98BvFTmvUXyrxPo
Xv/6Y4jLasMbOERiCXxLawl+W91zBvrsJuQurKj4xvYnMFqy6H4S2qetwK9QqS4ohBk4XLPSKgeO
BQ09yTeD4TdYKvXux9cSrXMVOBEtSvg9p+NPLDUZEPmSNsE91UP8zxr+yTvo8VdnNPSzuLzv+HcZ
KSG0l+DoJOLNCshnIoPDJD9XvUU2jz9BGw4jODTUPZLfrsXQSxNP/h0dC3+Luqq+5S6vrfOnF7Xt
80LhQcqBUcyINuSmv3mUa7aVS7Tg99eew/kidO5s2scp0YhnKvJfTqyQ2qA0jaLSVW565J3nfBAm
Htj6eeyYh5UcjQ2IrSZfio2HGuh705NRfuUkJw5BDvmCpC5thqcRBx3Z1iwjUQUh+lzlhRxzPRzd
7ZkKsFgBSRc05bJGhkcYKCXeiNpUSGYFTT6fhMtpW3kj0G0siNQKZsAhx9JDHNG5l5qDnbBoYyIL
H+3lv8cUb8cZ5/dbyQ8ZfzlIBWriIaMi5lqPszvCyY3S1WO5j8XdJzCtERWfz2f6qYDcIV/oW0Zo
tKrehUIOw4YtEqTSP9GUGYYlYlGCLbg9Iv6YSGzCg90vN+fCpfSUlVuDO3mgjtteI2WXDedPBJ8m
uZuovH0YpmTwmPMPBgfaPCn1jfeqZ87FNMNLhnulEtsUVSheM5iQDIjiykF8d2O5Lu5Lol9+CwDq
A0F0ldKHjyarxXNn3oNCbw1hNzEWvalbVsc8EvF6bsPfE9ij6PlSPQ7qZeZclfUYua+LUYqQl5zt
W8k7QmM7IadJceOUwOTJActoRVZpehQKxPTujSavWzpyveKOviWSIyiydJXbNkMFAEyTnsGweMj3
uyNq6ntK6Iz6cRMnXe65dtlxHiXNlwsnq5dLAPyHZmzMRbWFUV00nE6MJfn9EWrfzvqphzykWA0C
ZPq5fiVh22YTYg1VU/AQsCYVpfF6hsbCBkVntimVe93jTYmBhUBe6iULAXVZvQXfuPZdtR05JzG0
iEKOXbArzIZcDZ4v9q3/BLgIM+A7mBnKSGO6llUoq/14wP/hRgn1l5MUc0bq5aGpZdfNfW6wAgNG
XwCHlgpIn65pHN8qaAX1XInlKIIA6hno4we/8wkUQI+7gFHUY9lF6HFF8iDi7lU5HICnjShoSagA
D+nmGfdcBlDzknhbb3UKC6hFeq0I38zcNjmNxIHoF+MMqjrAbUibY2/E2dwz9VZ5O0scNWa52Coh
w4jZJ6Vb19sRlyOk17TiykiZkU+ij/BUSQ5C2MdyEuNSCr9S0/04uGLPVlrWNW7E5TGcLo6TxFkW
8aHqszPC6w5JPLVpZPhSyqe+l8xzcFn6WN7kwmF+yFe/QuddqghvCU1iqE1arczXI4b7kovigx0d
ne+3CmO5kGQ/oslN276xuf6X82S6yBmcI72dWWOy8ZILoZ6BMqQzl/Nj9ft3BNj31/55eP9CfMCv
kQlClAhHi9NDxSqTjMQOlLRR90ieJZHav9DrEgc+hXuGgV+MEu6NvD+scaX+Fb7Dzor/MeWX1hcs
OjpaJwQHjLe0qLhetSyHWwvYDjGAH3UGD9/4YdDDa9m/13ul0IZKuLaS+NUQ1OCjDgIG2n5T4XPb
0bMuENniI0deHhYDK4mxmfKT53TXHy2Jk+cokaKRgwrhbU1IZlaDH5YaowuRWsFII+W8c705/Ywd
7IyD8tjcaWc7Q/9OCX2zdmzVAUhWRYsfV/81em5nebIfcIuoMcq2ae5z3IqcOyGk2Vv7kv2m+DfT
7+eLTj+ydE5Nryps3azcPbASu0nY4sTQGtPktmZ5RCSwmbCWgZPA0rugDGkUnbvBq1pd6mL70OoX
149/98WJSgXluFR2eXtdrc/1QA46evx5ELLEQw8FbX/kgZqMehp7H7kKWUOZ4Tq7CxdzrY2TwNfv
A3tMMWxV8+La1O1K/F8ZAN1LMHaejsUFdW7rqf3fMyDLtb4gfJmV78ulxMxsH3CSzfeJO04lT0X9
hMlrdN/mFC41w4RysPc0B8Hp5hVbBmxFPeshNRrjB0tIyTUpM1f/d++1dyiVfEM/myLCQfMmucPB
sBh+G3ty+bt8WzgSfgej07lJv1SzrkoOp8of8zJ7Jail9nnxOxkJOX71pS3Xdtz6LO7hzs/W32rG
j0QcVzUXhGa5UVsg380vSZECWR5/qco19q3ZUwFXi7PWvZ/s5psxuT2aKn7oz5kvFhYRcpNvrrv/
Tj1KMCu3s6/b6bW1oiraVCCjFB56s8wZYVqlGkosjBrJb8noHzQzACYLqr454M91i0yq1BL1+fDv
YjlfWyo3eaGDrwsKZWZwgkZjKYz6GMWEv3wm2cajvYIB9TieHN52f06nOshUH2saoYSv09ge/FTb
BgRfZ5fSoH3/kZRUUU+JJJlbge8qLzE+uiDWvYyo/rKRfFm95oFzX8oufSe9/3Jj2/O8hwyv5Itn
ThxO8pFX2uqAV4uX1kqcQygeMM8zuD5YCqZZtKXSPUIQinR/ICs1uxHL8DXwSqgwJXi+MZpFqZto
q1iABDanc1Z1106/FqpfMq+m/nUWU+A/9bgc1HcjAvtMCWyeLZRHkHZJC4TwDu6a6fB7V3ShA45P
v+ygonyS+Pf+zIE0hvOZ5NijlgBlA7G9KgFfAQU+u4TIUiCZCby1Mt4f7XgxKDEQ5V3x5HTvr+tY
MOFnOP8K9VyaR5OzV4KMt4zgAsJBap/Jq+HlHKTPCLSUMML/CNazDiqMwaO2qjIugD7rWlaISVgX
bO2Fbt94/YHAhOTqwlqIB/YCnMf6uF2IPZyF1NJFbP2fAw6i0tMZn8diYd/1pIvPQ2UAS1iOuC0B
OmlcIB5JeGHPAYMi4qFQC5titDrF63NB4FpasKZYu5cCtRxN8fjO+9jSsm8CjE6KYxt3pJMmbu6X
a2PsPh2TszjPbJC7wWAL5Tq/W9jnXGBjKu+qkevScqIwVKYPuz2byafKFWoOUn2Xzr1TrP89ylYb
brjsKvWEHKHAFmrCUzJGY4nhvHMuEITTX+8MkeE0ikrd8zDQji+ZrKoAyQRnfvYd/wAn+Tp2moj+
MLxuRiKInMiiS/agWuklUWqBuAiOq5WTOncp15gWNvRZrSi1xgl1V1CUcdk4GoGj0HE950RBK8EL
PPuzMAhaXZ+UNd/0kXztA7c+c0WyVdvOyR/TRhoh9e6zU2qUohY/Vnl+kaog3XKb7792i/bHW4MZ
FvzS4og4Leim2l8N+9ieGNujGRviwuk3Kb7ozO3zW1eY1FUhnJXKR+LAOPk359mKevKTATT1BcyZ
mUbNcN6ta/SxaWYUIIGcLwq8utixF23PMWsOT5/y6jr9BCWAEvi6EpdHaLgKU1M4GCTouZyptkmv
4VIsyibXFp2nfQWMUAd04jo8WILAcQkA1Q+tMtPhbIahiVRcL8DiBUmXymEH5931SG2TEO13i4Md
f7Z4EiEVVP667oT90r7byUSyKpjEQd4UR9UINM4Djn9OJq5aQlcvgtMmu0mmHtYRxezgCLSN6qpJ
nMjeiA/4toHZ2FN+9rDKfZsI0qOwIJP+XxnrJtoQEnH+U+ZnAku+l9/eco9uXTOUk1vo2SOceKuB
iKG62x39elcNup1WxuCBH4+mHKJvD3zmSlVbjwEgbWwIHJ9fiE86D39DN0PCuaYrpXYb3ZU7qhj2
GRwpyL4HU5HXKiTDsacRvOEb7yrQVSqah04xWzDUCV2n6Rm5rElN5XgqitKOkgGkrX98tzcclUMv
1j3BUgA3TzrxAjlzFFvOjz74VMrXnB9jAyU8Eek41YDsjDkDWGgk6Mtmi+E/k0z78YQ77q5uYiHp
0lEE1BTR3tSfzfnK1ZHByWw2oDcbThvQOl6zIvR5MC0IWeRZaHTKDBLs8WjFolqrhwXnQqsQI/Hh
lXzESejAhTsZYojmWq8Q/Ixjs7acJKZaN+tW6QcHHpLBu6tp96qcSYtsp+YT+/FIoQ/qqTdv1WrA
Pidr8i7QX6N6X27ejfwj3egMGcDU57z5pjiTiF+g5HeQcrRWgq6teeBKHZYxBLF8Z7HfsLFN2XaH
l2KvFPVzTgeD7WeJi+xS+bxZ6iVeugjSKK8yCJkMT96Wf9Soj5NpQU0lUW4jeDFtzRcA6Y9IA8MI
snH1QNUI8eERZaoUOn74RjresqPKj/BWtBJDO7a+vWmg9EZNYQeWmZ+zttSPUzltwKUqSq0fl5UP
eSJDuJLjYABPyLWAQ0flZBwVs/Rshl8wvIWvV2lbmHnbKUD7t/z+KrTTgzmmPOA8p+wOhHMP5k7r
HA5LhLpMugzkhZpg6bxcntLW7w21YZ2bx4QQKvqeIU+m0D/XK9asUMPUaTmNXabf8YdoEoBRqZhG
36uAm4w5oxqhW/WLodu290bA4JX1O973T2ion3LoFLlvUnj63ZoOaWzbUPXJGZXxrYcAW5Us1tR7
YXcHGfC19FVrXR80u5l/tQOXzBr7v0f9DUM2dVGxsDK0TbSGeiC25g3e3L13UlT9mrnYlic03rJf
ofJlzXV+31d4kQyJo7tLttjwaaKY426CI2DIbDLJ2/FgxD82yM99s+gRUZwu4nlE9XG2zEYMeFvi
4faCV7L+bS5fJm6V3ZSft6rgMV2DKY4DYXmstrpaVRNU49nOoGM+czwdyfqU12p1KSKIks4pmjGs
ryBo80b1Hxzpl3es376BMQhniJ0sutKZ/mKFT0QIFO129hyCm8irMcq1xWXaiv6buGN2pE6bKylS
jOuiKZsat9KXqMJvRF93BtxDjwXoavF7MhPH+8GRmlQUYd3tfOxem2Uq/s0/FPJ2hsmEnHrGlP27
dPleVZhx6jqz3zBAa+FV8K+sry8jlYKnbX2ds1fxQb3Xzsqc18b66oF5JrA+DWA40eBR656jWX35
EYc3knRoOsjpSaeNuvF9/TZhtW8DkJFhOqz3ABWVqPRT56nFyqJ7Dv/q07FDltWOcA5OsRMyW29u
rMuC5MOQGxQsHV5DgWbKCODUUB4wPNcKWqa9bWkCAGLbv2+/5MqQiMhEyaH3wd1Z9nzV3YqepfSV
mYCdrK5cBADshWkqMtKAIynHLmF/GOGGwYLVCCqywzU4OZmfTzh7GUBukdtRr4bzUX8M3x+cfG0f
B8a3AnhDkR4aCs6Gl753STHUgvs5aIWh8e5z0NB7SiVffTz5qmd765aisMrf0fYAA6EGjimFTfz+
8JZoCZ5lTaeAyQ2xiwMtQt/gu0jkxtoD51vd5c8YKAPnoNPxzPE3gBuREmCZXxTUbEGY6qSYlue0
uQ02gX6Ajv+sXAwkwqA8p5ZLupyACPe3sKqpmegQ4kPjhbV02R8hhSg5YKCgaYvqQjbsUa2+ShWn
01YrXEm1ufons/CNxPpGgRM/VE0mFILB8R7OdvQuTJT4TPqBHGLw1DbsGtL+O9ZmAFhUFCFh44Mc
HJb/QJ9Jy+Nqzc4bqZ/YFAJWCrPTd0kUXC6rrrFW5iJHYfyX35HJXU+ohy+1YJmuQzpJDMjC0wYe
ql+grdTh4/y0vuEe4rNeUWvAA92ZSFOSonTgVhQlUn9BDXRglzudrhZ15h4zJlaTGz445FMuCCe9
ORbN+M5JauOMLTCKryA8OTcK05c8twCq+for88Du6mV9JArhP6xaXKeKZ9CaH0BfWAS8jMZmQMw2
cYbPudn8LYzi/VM6N4QkXiqVaCS8NK7Zx0V3DSsHXs4AyGLDYToiajgJ5zG7lJ2KZl4ww/UvSsZ4
vGDJJ/Sih1rACWUn9MfeWAH32smFUyuZQNvE1eYkbSnQBY7PR33y0eojV8la02HtpBdxojS/I1E3
MkHc7aTB6NZr3aNg2pnib/wt9uIIh2RDWs7ivaUoNmWwTKYH0MSKS9VL76Wn4030udINvDCN/qTM
0qlnD5NaQe/6UwF/jDD7U2TILvlicbweMZp+RvxlBYUWL5Fu84F9WUHGzBpSovGIl0CsJ6L8AD6f
VNNj+/cOpJ5ujWmqtVWugU86NTfcwlNkTy/99G8up+dusmu6WuqPPd4ahBo9d+1+NcjvRlpiB34q
s6PZhD5XdI9yh6WINx0TurWpvlLikkbqr+xlyTf4oezB7xjtA3XT9tJhuXXrFEnm968zFZxwJ1UK
XRzAXGeKywsPJsbNBthL8QZbu4+ACBK8PZHdumkeitYlPHMvBbebR92QiCy1/3tU3WVqlU+6fw2O
W03kjciaP5u9yUfAmFLTl5FIny0cn5u8kssqDwW44VCa2fNBChQMqOaTMXs/0pszULlk9JFxMA2H
9p48x4ORIKyN5HmdFs2oCVHE/NIH+tFrEUT5OhoRW+FAbzqUyUobbBBDTdFWwdrjZJN/7Fmhd2Df
NtMlCKDzz7ixKsKJIjwKpRLOafg7KTQyovQbzkdZzxGh7MZsjvOFKvysk5iAYjwhT+WFXAp+VRMs
6ZDt07J9koOOdBPs+puLjhU4dLydTYu55/TvsRf5G12D4Dp16fpOzMMncJYJYgBNtqTTI229xLCW
lrURCV8bqiAhVSKetDiYYGAjN6nlsrmRjsATNeWosY3DwqnDm8BRuPCr7UTwdrIBN+bfbMyd5MSf
Krec3I86c0nGT/8Xx1B/rxBg2mU9dzIRUSCJae2gm8s1x8lFXgDUYq6ceNyMAPvKi3N0MJaQKA3o
+ux9kcxH9zDjcKThxyDJHBtf3KUDA0ydbVrwq1CWviKBBC/HzJp2UQ84GYjhpdhs3mMyJpuqi+B1
yxxb5Lj0A99FtNwLzcBbgbiDIzFdp1s6uZauyM4SnUNZLLBNTk3xmR10nbcF3G3xX+Xc5L8ykd9A
8MLBxT0sJdjETsAyWcU8NuPx07my8b8dc11uoGTqbJv3mHgKY9+aa0TXmEav7PbVcv79DvOowW7s
/asXTaQ2cTzOFlROG1xBrNdLHrDjEMhBvyfUO4yWX0yBUG+QXASSHxkHIVkDHcwXZIbzAAz9OyFp
c9Mad4dVHrgo7MHWkqPEnBxeJY3KV/htf2szbjWAZu4uitzUO2Hvl0mU9uJZAU6PkGhDlw89m+p1
5xlT2I4qmac3uFWl8XPDWgA5dRIG8HVYs4fAfAMUdGvGQ+Pv4yYdCsqNUqC8vjpBvR1MYI9lbfyG
00nmKww5nyDOwzhajiIChEIEQUNCBWHIC+bbSeCUr/XaUz53pVd3wbvEE2t13sYjoXOEFsEVGqii
cU662c08h2NlVJp5NUIHQ4gn9BZMzec1qK4+JVQaLg+lvzh3BuHG8a78Y9Juj6WFcBzC4oG+62ef
eJdZw3ijlMAy/vGmUgDG/G7xxU6HJF9aSXfmXR/3McmfJdne3wP6yGV+zG/fBKL2P4ck/DRf9UCc
I9lojRo2q+QJf3VHDi6Z3vj0bPfG6Dqc1Ba710FQeNrjCeuZH/JVdqtzFiC8ZCiy5uGdn3bgfOu3
fVWgG3iOzdPMmHh/+LV/lDYIwPDO2s/dEjUe/F+R/Apa/agS/of7w3nmxJNxgGfmw/DRdI8F0hid
1P5DZzZfnT0CYdN9GnnKCrM6BEsT06XAr+CR+/erQcRBV6ef8HQg4LiPmiLZd0nF9dI+Fs+5569d
//TfFqj4+BtvbXdzi5LpyeLmegGu4z76Xkda9hfiWZUDalSf4jYRykcsO3DQB4N363EqtYLqBaYK
8N4TR49ThFxUiWV8X4WhpaCokClfdHaZDnppsAy/D3MMex7cYh/Fs64t71ax8bESE5pi40c48gsK
r6BEnrb2vbjJxYGiIlw1XDYCrl7IwrTZAgy5XNhjLTNq9d4IWK6A4qVCNhleg6+KIGg4aTkYa2qo
6O5dAFCZWqVlgbkiH4yBjOwXzmfLrRhvmEypT2GS2QHNEfr0HzCCY2IgYDjW1e4uc+zWJ+gh8EcN
0BM9zthc81S2IMQqZ3chJCUF/ViHqycRt9bxHVbTb4XgHaxjPYpK1Wrj2s6i9OGEHahuGeTFrv7T
ySXS+2Cphi67t6pO8KJLjYepLpREM/7KiWSxZhkyVw9t7Oms/Wfm3y3EgjKTpS8hVLCqIM0Vip9e
7BAsNmukY+1JYvIB98WBj8RgxqQs00DM+5XkDNxXujo6lyU7/NOBbmUDThDSmhrd9WZ17UZnH7H/
tWfT37HYvRw6xUqLPzXb4s7NaXxwrTgqKeZjgw8dpBzUWhbdgLUGQBwPLXkW86AV8GSq8KLt9LCk
tvrANiQBXrBnh74j6qUxgb73+6S8RMQAV7SAa061/W0uq2WJW2mD2gmS8cbFPQBoGv2op0S21q0r
c87Sebsu5ymaU0KrBzEwwAYBpDSIJEAfPW/6D+Fzxw22O4kOOCXJb/WL9ThRmqhbHg3JzA8BIwn6
ZV1bKNsQycUtN5ajTitfSmLltOroKZoH77k5XeScBg/6av1aiBxNQZqJStP83Kn3W8x4rXoclV+s
hxAEIY0kkSHAKf8CdChZCI37cTSWX3dtcDLB0L7kG1lxfsb7L6GbZ/6S0qg8l1ByD2juSNhUjjE8
b12bg1REiMr0+DwwKR6d+5vsFSM28BjQY7fWcqGWJPkSkBw3z/2tm+7I67yhWQ1rGEd4y1Q7PmKm
D7wHnJVX1hSoVH+wXdSZJdayqiYVaBDrM9/EePQj37RUrE/RFf0zrlAeugnz7fKeim1NGJZWDTKZ
VDhv1hOIWMf5inQ+kTg6iDkxl6YNSCBQ8KnB9mroARYWQBkgW7XhA2HkFsufK4c5Cvv5KUVVEeXQ
j3l640g+WKrH1OcaWPbGrk2Dhu8/eYBkzXnIXtNMPFMunop81a2OYXOHYteBrovidVLRVtjX98UM
XMyeOphZRFEub9vP6ikTWKzjkqJM3IPQFwQh3+/BNSeZmitELv9vhf3WCSYLBHsk7ukjH+ux/yud
orzBEkj+hFKeAtVTZxeTM+GVJhoT97kxF6jImDwGjDtikOQUnGUJEHFg8AehJrDmwz1h6f/ppNF/
m+sU0jVMO14rRtE0MU9DO7d2XOkW0TK9wMXw+T3Fz6YdnlsrxOv6W05NCqYexv6oKFd6omy7XecU
spM0ZUhS6oUFBLO7TUUpCoK1Z+uzRhXOXx0SRQAlbALMrhgoNxy2VGewup22E1i8clcIxEqCTFnL
hBmOz2tNQmFdAzELnRklYUdR5+VcpA2fZMkKdEuhr1011TV50qVqAx/0liIEsJALgvMn/jXVfXEc
/StplVWREdH5Ms/veV7tMvnc3qJP5UgPIZ4oO3Cfw09SA92n8+FA3w/76+Xr2qvu77n6QczzmMFO
waZ1+fV5LFQr+UCX0zrQNhO+r3LDJBxkT0wjIOCSuFexTG7KyouGYwYkmqE+ajyQLHPOmnWK1ppe
Fh50BbFt5yUEqIvCBZ0WotigxlxZb0wOqUGNdY88tz72UD4u5SkQPg/4ddZdMZ8iLs25nwpbxFrC
NRi/CKy8y8alDOoAp164UZmPG2UBUdCszNvEhJ6wFfMoG1PRZExXgbj9Y8Y/9TUHyUmHdEP4IN/E
78mSkltSpM6o+cucl1ZCEo776ufMgL1IDY4KxfwQNYYt1zmVQynYGLOch8hIlXGpoK8EB7z6jmea
dNZo8+kR9HGrNcwylU7jF+e3LbgJC7tzHyhrqfdaCLveMSFZ+dsPGPC+rmyHhE7Rm5szp1+GcrxG
sQgp8y/rzIcEGZDkcgXP2yf/772JXILHeS18F4Rl3badqcaEqbGY0uoAlngTQw//eCMoI35d/bzw
1o1gHL3vcGM6t3zRoAMCEjHO3K3BOOFZjYeu0WGarydT8Zc7eSRVbi87Me5xBYVPJrcGBeOCjnnw
kQxiisPDwDPT+3ArG44s8KTc8oMGbz5u1gZPpCoYxoUlKLjnwbz+jyYIznvwuRE0uloGrTalm84e
8l9NuE5m0i3+xL0WmlHFfJR0soxBgEwJs3hNA/ZU0yMFQbiuAGfc7eitLVlX7QrN8izMWrL9bja3
qoWlrosIj8j9qkJ9cgzhivxtTCV62MbAGH6nL3/oJ4wxahOXXrbVxj56w6EY1OFBvEL4IYWiW4fU
1XYnJyaP0058qMLDSgje4ao3dbaJ2xHCJsNnNGauaNMaGJpE5SNFaPtsBpUI5ymPIYkBp1yvD+9i
uPi7stbN5vzuPBjcRtDu7KkHL5k6kp3E6Aj1PXs3FDydv3Ystj+sl1wfJDqk0DQLuoDAqOoftXr0
486WQGu/p0bKOL/+jGRQguaVq/7AO1pfXdT9rHSpMD5n2RBr31Uwyz7a5s7kG9pCGBs9mqlThgfH
T/JNCgA8GQQgIQsl6bzUsv7TNo+g0eaUxOOss57+RaRqCRt4Nv4XccDrU4Z+JosgEMaVr5Rzxlt2
jGxEEeIKNLuwLjYtj8o6WO8lkbKTKyG2dRtNJaBtHQPjWOJva0QYwCKdkJArYPz3X1NobCo3UI6i
gTzwEdrXgavvW6Oyn75rGp61fMwb6Q0Szt5TEErXLVmQ5kRWp4KqEwUCYQjf9A4RqJ9qIrx5xWfn
ViMibyzCwhVE9gPVVc3ui09PBs/kXT5ggE42kLYAOWoVe7Zbuph4IGjDSdZS3XCP5eSwtaxdTHN2
ebXUVeo+WGTSmOsENljvqfbJPb+oYFyrlmJloEx5r0suiBmxKA2ACDyZa0Gcs3CAX+vEjnyxblS1
9LFaum4Ycry1V6HWxRuLZh716KS56D5oNe48dkRbAFJfG2nWTziWjTSszyhPwX2XvPPAOdhcydPS
ELiqEVUeseUYdwYNoPVDWQUUDWAxqeLdosktEUOLZ1LXxZZ/me5gcFO5HxdrlJAGmV/HRRpMRJlZ
cFGPNGmAvo94eE3UamhHfnIrdQyCrbiX2oXB89g2nbkxXqthJPrXwkbBYy2+abKHqBHGZ00ItdUz
EzYvRCqlPb/5asAixfX4T8RjmDpB9PNBflfuVVL2tQsG0lhbz6F6la9wFE3yIVBcs/Eaz8aon1lk
PzuXTsyEdvQFyJ+jExVPenHhX6JirD1P3zIWrVvPTKx+wwe+sjnk14QolNv8RMbe4BeCXERtl6Se
svUMQ+8+fEHeFNBujGsl/2AKQ7NBAB0cmXJSnDu2B3/Oz+YHlOot/Qmuz6iH7qi5AdLlN2OBqH+a
TQEtDsrsVUWD7TtSL6DjXwMeMo3FWABtLS9f92KWjR7KvFFpWJsuAE5nfCUeHd79mnG5SFCJUJR5
bYy9M+hpjoTX6o++la0iuuS0h0DyfzLrqyPThpB/tspR6wD09cFq7Pt9GzeI+uANQXuFgd+sEMeK
umN+GfchDW/lcSc9x26doC0VMb0FrGVStrd5SGrEoXY9S+iPPwAlEYJy7pNH6K0QylNKQvJrkzwI
2tmMKEIXh/i3/pSmJ6OiAZvnNLOBw2ceRhNLUCxLWmj8tR6yKd+aoarS52Q7NREPIXsm8JTbWFVd
Wj+KbhZ4DueHycUeI8qXxbyJA6sWuEfTtu4gAg0Hh2VIB3SONjkiX1O8Jfo4f3XKDkwFxh8NGCxG
iGpgDwSmBxTmLwL8cC+Z/tdK1PUgTEVwnglCOvyy3D8qK2RuBTitd/rQwjK+4mxuzdzLZgF0aP5B
aXrlq+7SMtXW9KNkVlSA9sGvQmF/aVeAFsAJwxtDgmCWMsrFk8QUurxPgAna4DT+vdR1e77Ste05
15NcSf1aLGuhRY4rGFP06DwoJYsCxxR6/wDm0pRQfKxi1hWo9Pgxl7eTOlAhrT6wzZAXiDETbiN6
7mc6yZ8jkMKLFrAyk+W/oEbIzm2upzX0uUcwy9R6OP5EKyQGDlZqo23T+kC78/6tBzU3FnYHP5fH
ipaC3mRi6nr9OzeuHBMSGtveeaYW3T9CaN++JzFJeU7EEynsLJN16u1WPkcdz+TfrcmTQr7YfsC+
b2tXf+FduY4I9h3B4Lc+Dj1/ZIsX5cb/HeJRo5+JFqJgIoPHEGFnJCshP8flOKIMjYiJWtT+9aoR
9Uzfg3Yt9mJHlndm2zTfmja+ue2/kpMrtvJWgYj7GP/Q1WdA9+ATL5T87NjU7dL+LJhHuQpihbyV
DljMltpPpiuhEiSaLSB7rtaAFPD9MPkHHbxTlfELgUN23BfkOhGUTnoQmT4lj1BBZrCyxC/y8BKi
aKjiIxE7n4zuLTENpNiZSBJkPfXCPkYr6GHtK1KQooT9jZQtMv4EoCmbW5pilZNzEw+F2pA/+2Py
RfVmgA4cvJTevG/+wgDT/GM2Oi+1vK4J1/m5gNUQSJ3jUpqJWpcyJPLClIhaWauXgNfkzfqrGkTn
w2ciqWgoL7EqtQwUfGAAr7CZ9mjEsSyImDdh/fLtr028zwWfYsl8MHhbN4jHP4/Pdixd9FIC6Z6Z
Uu8FCea/tfqNbdrk5zG2R2HF5qmNawExl/z5vM+lHSXk+zXXLUmuxZ5CX+Gm3edWG92GfWmpaydd
J69T9VUsbePIUlmzwcECHxqpkS0AFsyEGTOIRSRq9JhRF0+C5tSWKgIdVHiVW5r5d9WA5ObCkUzj
V8YgQsUJfsI6k8jdJ0vUc2MrhQmOUTAPyWx93N0rFVVcTgz/yZHdsw9i5yNQxlq1cLyz87xaCTQj
R7X1VDs0m/jkmHGxu1v4LOWRpMZgHpgTIDDNxQEVS/Bftl/r7ktvriMAT6hb/Kz1W6gpWIq0j8b5
ToZk3/tOIv0HW4Nth+gjSJqjY/GAsraF1EuFG5D/t6188HjDSEzJkiyUnxQHwdLeSiBaonxBKOMM
alyXhSzlLWUAhd+fzPt88p9w/67PvSnrjXDEeHBSAYS5erNybjrEjd/4iCPVlxetlLgtmMYpaPkQ
h5KcK4yfZ7elLoA6DoXmnoIZB4ux8nggGIjXQntZqyyH8XrqkPO+E/2/HqyMucq7AuSRHxtMVe6e
qk03gt6OvEi6Jf/C8pIgjrQVnB5oGU4qNJkOq7emJuaaRGsTxNrjogPDZ5lab1Li3UxVNohADEVh
IkRMCt6CVUB78hXqjoFDSX4JLxoSxqZ/G0Umyg36rh2uCX9P27V03SrT3OnDtoz/gQxDxubyAb4H
cmpiO3N4zxwV9p6fAJASzW/c/kVmENEoOdSw9X4YQuDs6EH3J/cB8F6zCIiiV//8+5YIfxKUU/HQ
pyTy9OpaiIBeblr7uR5EcJNz7jUEoMamZxfpTAv4mUUxFMtYt07SnVu4K8fxqef59lLm1FZOPW7n
2tOFZwMlE5Yb3b7OGa74NWRYjulo09m6p+nSG51dYBxMTb5rKrboRd7pY6VDzu70/57dQ+lhJTsA
Z8BuEJ0bFNoTzXzNL/RJOfujTJjRnkJrz5hZyOBS6e3Xguxj8tljGF03Lxo8LXUNbqC8ncI9obqg
4uZBbndsOOkkrNrnv62DNmHlzzzgMvpIS4G5RMk9XBhbEi8o4FdaV9C5akL6fswNmZrOeXVWK2cw
qTWX7xesPdU855QiVF29pQVyMV6Z25BsVw95RuYBXAqVcikXvjtJBp+H7PBG5tZoKa8npy3e3Z1M
lf8qbPNOqIdHSdkE925olO9cmRvGNHrolVIk9eIcRdfnb16sAW/MU5NtKZeRs2UD4d+kEBD/0j3m
eoo7swD1TgfwvN8RcD4fYW/I3WkOJeVbvqUTTFBstW9dRWn/2krtdqu8dxUaAiVVc2viRfUse9jU
NDSR6pDwVD8tpiv0lxALwuIs26DSc9Cd6T3R2vV9jJ6Q/K+TAYM3sC0Lq4uAPgsRm5loPw56V4FB
8ILhpeiNfYgegd2XzJN32Uh2qDdi7bbGpvknml2tCJ6OHQAOB/t8sz9jrrBiH74499oAQfUIRm21
BVbqCqMAEuEgiu64Wx1CpSH8QYAtJXFr4YCx4Kb8MlD5ce+l8LUZHvaBhl54/UKzeitk+PSg7txc
rV8u4C3DUWnd3JthCw4vse7/ZxKNa0lrGO6p2at0sB3amClgigGG0WNk55u7cdrXJQOTPsXfLCYA
qN9a3vFBqu85y4ebNj3QO7VD4w+MXrD0QwJM4IHRVsz3dWMh4DIVSF67aYtJMOvE9+xH1TSEytY1
m5YwiuTpeJ3163z7PCYe5VULz2nACMjN09FyiChmbe+HoB5qwRnaJToGegOgvMDotNYtwUBe83mz
5VX4oL3TwB/atUEwin2W/YryERHb3KGclTj1k270fvJip00kv37FoO3VQ5NFCFmVhmLZsLVvgvyy
3yaPMRTU/1CAGyKovlDmQRHb7RYs/xQ8zjImh47o8yKErqaKSt2L2SYaJ0esHUWMlJNJqzRj7ecx
2UZJ7S/lNKz1cba8FURj+cRSGGM1mbaPRhpZi45Zb4AYOWObcsPLN0/Y2n211SUMcZ5yFs+xFAQ6
kvfhZ02cF8EpDNGo6HPjPw6oyLdpZxJu/IIFW/f52zm332ZLVBWES4B8kqUCagfSCVmO8R2H1qtg
WhkDLvK5vDL/TR2kEKKv9ZOz+M2wiftX8rqbHOUWm/72xY4sz8Z0n9wrAfbRvSGO+njyb7ZNcAri
7f7cLYLALvL6S2YNr66pRQXHSXy/IKSmPPdZ9cZ+zi7ogP4DFosH84cCNMvyWuL1Z6qbXfBWvK3T
saNw8BU50NcWX8YusiUpUMdn/ZwvrK1jer+WgldOmlvHKxxk60TWMS3yZ+pqZZG9mlAcrtbixlmw
MUZyk01WlS7IZncp6ZWIQ1E7B6yiQsA4Ulc9vu2Upt+U+ERpfOHU/SBbxXqrukH/MikfDMb1jXlb
HIXOVhBz0U1SWfgzdSo880tvlcqHKM11r4rGqULiYu5Zu2asl/OpQKUjO6Kxh7bZc1M3aI+jpiRZ
ns9PvdzTX3TSQDUmvEaggCrXL+H8NlawSQ4s8YbVkZ9uOQYuf2wiZywxW74KXdMtydXjkn542/Xp
yAmqPYmmfYY004x56PDShYgnQSPKX62REBSVC+vw9YyV70DVzIUuayoQIXYR67C2vq5lVWVSb3Ta
smrJjfQz9Ko/opJ+7U68ihQW7Gc3IgU81P2whC4rnsqj19lDTi4XL0aEZMM6vup2oJhHpyBWkMno
1strMJRDRwQkNbJPo7Y2kSTo83BQvypSUia2p55Nq/Urf7XpFUGdJslc1m/IUQGYRiEqRL7VuGus
khsbzJIQPQv1tw2SseFFk2AY9qKyTfxQmb2MF4K2WydOKivtd3CEiB3WfnXQeDGPZRazCvi1bIuF
JOX8ntzZX4qzf18uF7CaFuJOvgtop8tDSO3bdZAtol4/tqobDcggz/8yJvHUW2coBRgBKYEjd+z3
Z0bBH/mXiL36yLCx30Qb0bQGDoxkNEZ1/JLW4fgAOxdObLMHAEyv2enInZGzHKzc3VS/ByHgHyCL
jz4ZS+OXEJ1XqSury3N6v1ZT/zre36VwkBVUMsnq+0rjkHvr3cC0Ms6q9BW5MEIL7BQT8eX89JEx
AY9aJdh/WqrB9Hgtraz71AE0ocDxBt6LM8On8U470OPFcRjJsUGihKQqxxEr5vHEkguQFHZdtXY9
MQW0JWh/ce2HIzzyEKR8QzUIxuLJzbSGSeUGzr5PuqcOIQsdCqc/N7m2gRptcf7MlTYoZ5H9cCD2
TXMbELhkh4craWbpJUXfdYLKZAQ3EbqrNZZKmkFa3VDjxC7zeNEigOfykTn4sVUgiqX0xdpd4WlO
r1ix4JWFtiQsPZB2sQfttJRYjoPk7G9Fj+5DDUyYx6Ie4Xd864Bkqrp5Douxn9U2e9Lq3dI+nAU/
WaIEJCX7iMHNKSwmCnXeXh0N76fTqYKWba6xkk4Yxz81DzLgt8X3h9Fe7ZyWj/CRYT4D60FFT6Ii
gIWh8Bu8suRdFdcflyCJPXMJUbhN1zBtaE8bB4asEzHvYhmexTTmuaOQ+MlFO0KbzV+NF81Blm2r
YvMjDcrZlbptMrh1zJ5yklp4qwRQ4GRyl+NjuGlUgRLuJuxSfGdYVt/1P+3nj8YIHg3m7098sPim
qtUiG8c69kzq41QgRomTTj52YNZIdyrLa3GF6UU+elfzOCwh5232bt4CLhlePKmp2d/k7+y/rZ3x
hdtrX/tN6uZad+OE6a3DXj720dlJfDv8uY+PBTB4DYngE3EZouPcY2ZKyfeEKa7z2AOCl7y0TErw
B4doodMCKbJy+HKZNSj/OSEGxCmJsfJ+jg/wj6HWN8BSMT0Uv3bIGkU1HpnbGmczoyJmtbAI/U2b
NVgbIct5Yjouw6+XCERqMCqmVEyNDO1HLBEuz3/0UxB0NUwvzZgVqlGwAchSci0bmFDRLKDOJzen
ODTscyUEEZY6c1gpRc1HdkWUKKPf7KY0B1ctgHWUrOYpr4oK2Trtey4De8KD9oCSsUO56MAy7r7D
EQNtWZABA8T1DoYJBQAgop8eEYPPeRPKiQVfnxOHRkmHd5m7GmTNtvCvCJq0QXTW8p41f6IYa4GK
C1iygYVZdguU+XHpzxQ3XIpzcuFgBzGMQS5HOj1qdgZuXriwge1c70zXrceMZc5a4Cyp28cLXJ1/
Y16CpQm128CFo1D/GjauYeSwUPR6GoX3oAp1JQPOoVpnutx1QWATMAVe8WTuGKRLcTXGmMUQXz7X
d6FtEkPSLJCiUM8VpF4AnBaTn07a12f6frrstZJJQOcE9V6oeli9GslKHZ6LMAkmWd4PyrD/EWPh
j+G262zmcNTlTT2RRixefvUVRIZB4DXKyDEhGvA41Iq/w+0kMdBtFQ6JG7H4dmdJDMrIPNwxwi00
c0Dcvg/ib44pTOiywkXOR0mM/Uls6yL6Er+AwB/9Lrrebcxdi67gQIcORGVhZADTyTEvg56t5n/y
rMxXxBlSr6Lab4J2XjDmcnMzq0hbXrSAU4x67Wtnje/2eIOFggvI34m09V+7RdTW68IDgrUvndHs
RJUNHWbVSTbZZ5FkHJzPUANpGFX8YjBjSM2dzY2292b7Ql39PBmSxfAtGwLyLujjgKSIonx6EUUW
bkBGCh00ZvB+8aFOXab1oNmA1ML6hUNkbP7MeOCWWZgE0S3C26OG3s9MOlCKCf3B3W5RxMwYEYkc
TozAxHbG+BP9GdZeHkteSh4LD74UnK4NWDLADhb9T3B2Ps1GCNgKEf71kjlOSUDJTV5EtQ8nkNtW
AmD5Vn9/tWcs4FHb0XbWgCqstHxLINEKQcHO0FqlmTS44gGdxeYkpMNsW69Pb9TrsHce/j0z2myr
5gV+AyQVJ/ShvkqVtSZ4rySUONm2C8VGPBFlkZ0E5HUGm4XBggGPbKch5jkQKOuOYQ/uDrSEI4IN
k+Yh/b8cSYRW2mWee3OBkQLZHAVPLjvRxd7U2INi+BsrIgdG2MGgyXJ2OrSowCEzldwseQ4r3fql
KHxqdFYCn+aYLtnzFuKkxSLGBADtlhjDoqR+sexECyI5XmCw8p8PjWeayzFAsOzbm1B344bPCVTV
VIF80M+CMDwfv1XA2ZBFPsIrJVfzVGf5eHKLBYwK8VwznXcUf9ZjYWdaxBDAaGpu9OlcDdeYfd5Q
7aP/T8NXY8voSdoA9+ZwiJ9Awatp0/V1y4c1uihh8i4VILOy0hf08NsSeOZ1Jw+1qRN13S45svAe
g7FN+XsRybWCwaJxkrghk7ydcaCZrXY7LlHc9i5Qm7zd2e93uq+OXRhAiBimDiM6Ip00e4BoQgsV
wpYiHH6NVSmV22QCws7SGP08fxvfPNofretPXGS/Kj7JtxFtlB+zqSxuBEiTwqkkgCcxl2Jvi3yR
a26P02T2wqNO2nzPJQhTQde5jL7J8ACFEG7G+/AezYUFwKE4LEzaW6s+pH/9dqLrjyK/qJTnKYPE
KNdog2IVRscHwaZQNYsZjHomqeGZg0emJO+g5UTrJs3/pnJEMKCGxl++i2jf/MqyViBkEeaG0eDv
jFyD9pd0or3aEvA/AnOQqKG2rzOEzwtzGYCXdmiznWX/cBL/8bFZcbycIyTCgsWW3hqXpJhWFv5x
ezlN7dXE4dY3K/0JEkw3AfwrsLI1pxtKNWmEWA2jhrQlFddsWSE2iZ3aKjyWXt6R1BFfIE4qPzec
kvL0qGMBuyUYf9Sr2JI/vl3fiHl6wOV9kw3w+REqYiojElIdrHk0Lx/1KDMx+uhOAYaZsTTXwZbh
Mp5CrL0nsma0GR6hEHFY/QbbLOT2xMcEm09OdK4l8vOnhGJGx48K9Tpdey7YvzezuvNwaeiUNCJW
LaTq2byx3u2qr2RqAeTdiMtCWjbBp6/PLK3cH5QuQv/bT1QL2RlvGFYCxGijdwATLJCIuLuVNDly
ck4FCPxeGiCsgz2zP1s23svPZGdhKtJS5Cf4WG+WSWaVTLwzdK0ii42bnCO9yOv9vtxrL0f7GoqT
L2Rrp9lDFcasp0sSrAF6owgyH7p/8fCwuTgGqmzSa4UB2xie4SdfMWv9U5OaQGABj7qoyvAbORVq
NDOi6/QYXWzmnf4Q4iV7Qh5v9fwza0itTHaWkAhW7CRksKxdgx7UM+X9xIsxSrWSzyxWWkWYVTsJ
XRUNw4Nvk8OK33H3Da1Ut9xw7GQZyaqQz9x2oHlzu8ZPvw8a+KHVlzUQD/1oFnUeHYnw+MhUAtGC
y95ZA/LyU5JfI7HeRgHnsxIzr6VDQYS1wZjZ1gfcCc7QLcFA/bCljjcqVgF6JYmjLJg/q9zufz11
/1WipawZsAff9KIvFtjPgIlGIHz4/EeUkW2OIBh6EEgiIeZM+BUAOx5F47MJpYgz+I3ZEJ23Lr51
l6mdrn7ZBdr3TIUJfc5+uH7UoW8fbn2pcj6YhukmIIAMt8t25r8S+3QOTbH6htoC60hcR+mgSrGL
UYjYxvwJQJtjUhGX4wiQCm/BKOyLG/itQ2TsKiCYibxvJsTMAq+9mqHvcabOP/3rfiMeyUxgz1l6
GKNgIYaSLytD7Iwi6eLKiSlApuGBhLW+edDfQond1Ov1p9VIMpa5BlASJ3A4zMwajEK6lafzi0S6
ogg4Bw3MFkH9tMMdEqntHc14fDUZLD/fFuAfP2bcXvOjSCm3ZHYDROO2TuvNrSJ8PoqyGHxUEsi8
fC23wXgVyJXGRsOFKmBgbRh0aMBIszT2xaCo86CDrRuZaZfkEqLZIO0DccFSuEXvKBXhZDnKg/Tx
BeCQvJ/G0WSA5roPcueew2v2ToL6rCsMzhu2V8ykaZbvqGvL2SEH6Gm1hMSrTDRNviTr/QXEzu3z
jY97Z0XmeQV55EMZv62tQUfpqKfCJWEpqTn6AeNAvUMsFh4jMvttURRsOQIcWenB1rO245rWC0/f
oMpTVf+KG31gZPBE0UUKzhGtkazrqTa/A2zLdce3FFkMQ2vTOYL4zdTrCmHasCmEC+dz3pHp6uaR
bOfKjJqTrnFnykAfqiuAxXAWGWf0Ym7iUGrYGNYABetUtRTskR/a/bazTJreOSxvtkUFc6mNikkb
218U1+Y4z1bUwO3ocZ5DQTysJ0Z/bQspZCjzJVGVo6z1+xUbSb7MsvYsH4ftKrRRe+hJm61ZR1Vz
F0GU3pHt3qRPUjNUBUs8xW92L0ZSWw2GvxaV/y4Nqoh4Cm/iypVJ0W1oVZyEvEcze0vWKBwcl+cW
LyjcUbJKchcYNovBTiCtEkJQ5yM8fl7GJhsfuDhqCRx8pbnl8IUoQlf8WSef70iNQdsdtEDhLUJp
fSQJ+oPB++kERqqg5jsTbHf18iRhhClsAX1j2zI74p7lz9c0b/8OWjNneZtrD2xGc6OOKKSsgJgm
v0FcWYLGsdAWDsuueWnRMFX/MMU+oJ3+yOuDzh/5TMwkZ25TWQmJjbV/2Fl2fo6/6nuIe4OmsBXb
Uoj/xKhL2DLnmKOmQ1yzINvw3d3CSk2p+j//S5EtM3cVw+FxwN4ntj1YCBELX1Wdw0sNEq4r7MhM
jKcV0shHVyx2IDG+IX2ZHRNnK01AG1prM+nIQfEe8O+IeCBPgm5cGczW/C3SoWCG/a8MekuTy7UP
MaHwJmuMnyIULRC90/CT77yIaus8XZ6aM7Rkz6C+yDf/BS3vNoJLmJeX9MR91BpJGweUyk56YzF9
Bs7KUBfAg6vXvNbdHUsbbQdbOFOij9j67lCuEBtJeZ/vrE4GG7a4UocXJZZo7qxtabunlPQdVzX9
GSpXGBAIMMtfk8N+2PUV/zvnKlBVKHgcdGjgqfZnAN6QbcfbDKchXpZGuZll5pyjHkeYNZRemPCe
uk4+vrin+2EXftesncGi1LRq1MW8VKnOjt6yhcwFT0vGxCGyQyuISO3iqTnHOsLVtDD88rpbxsHf
RwbUIfGRLhr3LNt7YmFB3FziqUccSTYaW3B5nF+vmXEbd7llnFwlNFP+1JGLV6K4h99Q2+X7UHBE
ny21trlGe13ijJEgsS97DYqIIGMMo/r1j59UiHXSK7fBpInlc767LFokY7wUJWw0admZcvRIpEWP
ziwPmJR+d07OFc0aOQHEv3WI7/I+s3j7MVucf80htIn0trb6z655WnRJau7B1/J7oxMYiYnegxmR
uTbCEzs86sysxeeM97EzReoKgZggaOexUpd5izMD6Ravj+rTL70b8g4Djpm7yUvc5kNTHleDIkoi
xvDXqlyh99GzZZgI/g7eBwUuvXmqQfk9WP4ReyGG0nKr1jVxDN1IquEZICb4ajHhRdYLACbaMnRe
KQ/Zc8IQGpJfVrD2kPefV62PBv8kNeWOaTcx0mOXEjryFKNtv3TOtNOEXemHguAzZndxhJZhEQfr
ldeP9PnMN+o5SfQlH4aOM7fjbkmg2OlE067Mkp9R7S7x86v686UXS5cLh7QKwb03EYuHrnKblS11
EdjAzc+y9jZyxperGPWeUpN1RnLobAG0wknTe8AFlVSmmU2v67SRvHdrjC0L81OxNZ7PRjFLN4kj
vHNQRMbIhPDa3jWxrDmIObqaGnxWiqkvoBuOeeFfbmtlHJhjIE8JFoJejQmMuo2zC7dCPSJ0Neao
71b4l0ge+szaxN9SMfmB1CnvjpiPgT+kR6YSTifABZ/JL92oXdNj7+CfMng2XtpoAu5184xZwERC
t2SRuaAk+U0Y6vg/MboP6vv8qcYgNqd+YcRXxkEcdI6jgXIKc3PJr8ZYDDG4OaAgL/1+VdnlOV2U
WnvMG0JqGK5bGnDD4pPVRokYr1W6UYS4D5mWae0IrzV84+DjpWMpiNqgu0NZqKDf2Bs7nqzs96QQ
ye+0Z7oEejWBBMeRooJFMFsIbGtmWJSEzfJJgiCCCEdsUTjSuQS6lDvjfbF1g/MQSfxoMzRoy3Ko
p6FugVaEyGcqCoQFzpa/jA1eiLNhOOzb5C7fY3io1zh8hO2P7qrSkk436IVC1l5BGvKTj1RpHeAD
FZGZ/HyjwAvQfr70jXZuZWWAM/ri8xcrLNtnEG3IgYRq87HATwlNKF8ZN233pzK5976pHsLEiIOw
zh6ZIKN6lIvwGdabMH9yaF/48+rJLRVlj9PbmjyA0ab5gSOcNIKerUJT+r8IA+E8pqjP6tlMy40h
6Ke8yeH2c06We/1saWCRticlH48QyPt9x71bWQ4frJtl2VbgRRFMBjZSvq2IbN0/6VGY+hl5JUgo
rfCvwizOAXBZ3GOwVNNkFjiGL27U27lU+Qr7SdYuIhX9ieDiC9rfOxK2nHuUE7cncW1gWd4bJKaP
zUTFcnNE3+TsHwos/M8F2sBKHu5Cn0VOad+BMyxfxlgWxBZCPRv9oO935ZHghsa9SAz8p8HoAfNJ
NoM6Kf2Izqciel2gjj3pukxL3DYKO86umliuiIw0xXfux8exPHgJcg+r8hXP/0ZNG1W07vPLcBFE
jJg7EGxOwflmKqOGIcZbeTmdVScrKxZ2MqgLv95G+q53G86jQ0YCp+bciubKYc5Cc1ZwLkIbvw27
nwl/ZoO3/yYj8sBACyxZceO7zPvuuQ+Vj6jaT8nzabA+pGjtPsArm9wyqSUnm1SAbXoCACiJ4w0K
6joFP3dkzDBaTj1mOM9RdVPkR3D/DAStXenseAQTXRAOGEyJdtoFPAVAsk9RGYhnr6g8eaxbiyAd
WW6DMmXaT43Dy2CRyXKujTVmtCmpeFIQYDhseVhB8dJCBgWI8+DEjkgul5Cb7CUXt01rtiWMzMPq
JztR2kFlIoX9rxq6+wDiLTx6gVFfjG+At82IBIfS+GBrnVZthOOyNHMxsAt2Bqj7MzbmcYzyfSfX
wrCAv7mPzXXEst99Je83ZmH7Jp1zDNgA2z5gmRHhSpIea/0a14Wh7hVF/QdG4zUUF4uYkEy2uPWc
0SsbWAd5PGqv4t+kXmLJGCOcHJizQjeqvOx4u5pOMGbryKID9UeH6mhazZdl0OzOVAnM41aBCllG
KtZ54GmdVYEptpL4yDyGKoWl1EUadm2r52BNkX4KnQhJQLeP3px+jokJf0pwHbl6SsRIXQNYrncs
QJ2trOvIHD5152kxCR4PSWit8cbR1mV1RRFejvaI9N0xHMnrGoeGfFWekM5hXeeD/c86hlxiJ+1Z
FJLaRcFQviHcu9Zs+dOk8OYGi31nbVkckti/MztojQYRfF+E2Ek9PVxGhnsI4iRS15RNzki7cwb9
dxDsdQxOZW/PUi+HAY7oZvwkR1fyhP1xYxoZfjRn8dl6PPg94DrdRQ4KvtQC5WreUJ7q5sfj72VT
xhZ5aFfiINxGbpwVr5rfW1wdTUxZTMFUksYyvGnXGPKjHxpClxQxJXOl7P6MgMu5GTgsRd/NaKnG
/tuT6DUz3OLLuXE5apEuq+F0EeR6OhvfQ6jCpWQjuxeA5CJmiHtbPPcLv3dNNlMe+dy+KNtSR5q5
zd8fqH1+7gdRL6+Ag/B9q80MFqeRyrIoJrG+95IH3g/qr3ccmhZrNDR8rBl4JhMgspO77pazVmV+
CFyr3TPKQXDaMRLPcwF9k70evCMMqqY3jcWuLDAtTKB3ZCivgcEIkUw1XOhtAHE3DXwkhFXNmMSZ
oSrS5lVgBRy/A+0i550u1ZjQy0/RlLZAJ17e+Y6PBGtYeY1pYKb9FET5arTbAgD7czVAkeiCoXrg
ceGuI1kOKXWIes0/X7JZ9DLWMDO3ouGVMmQjhzU0RVP3NH4n62p4iqb05KeYV2EC9XSz5U8VjUV5
0zGrOFAAYLm0GFNQAEQm+taEBGDa8lCeNgniXiv7NsKOQy54YSDgew84sF207MEqYiJIIBnF7xCQ
WY1VLuDUY8uHfScOZmwocEId/QwEuw1VYeh/TdMwX6+w6UBCso0zEomRgIe2f+w/lOk0CB1rHx3p
D1wzweh8meWHyQ0xr00I3qPQtp6h2IClchy+0PwlBhPzfldHpQdAQcfmIPN3yACGAV5sIQxEpg/N
tpI2gF3EmMCYFNrIIa9ME8hrtQ3EuWHCDkqf/6nEkvFEuWMqFuPF+iKgJwUM1zVjL3Xpjv/8GTLu
HSicZtSf8NxaJbA908dDFCy1pgtbF/REzaEtUiWU2dYMkp6utCHX0xex+QqIna2vsy3+OHq92Q/m
6JPa/C21+xyBYBEe7Pm85Tj84rtphrWOq7iBououUykIVt29KSdQG1aTdi34ZGhtpdgyqSHB5Nd2
Q1ZSamIk/pfTHlcn1jyhFfw1iNRuOMi0B1iDkWAABK2b+xPh9Y9zLyvCHBcxHWff198ncr5KT5dk
TfM/06YIPb/5T6IFMdE7O41GuNLMKQbvbexPPKoihWHK2fMBOcil39a0vxibeKC8T2So2vQkoYLk
+DuVl08ax5urOOETPYnkiMVZszDcNyJ+tAWlND6NLhWfUfI6sFBFt3aD1vi6YaQJwjH5k7/qXqoL
x5CcyOf6iAx5naT8ATYTH0XZ8NQxIvjq7mnuJHcRmmt3Jcgf2bvVDME5j0F/iFKxRoEgeWAhjhHk
xDfDSpQzz6CIlcB+N2FldGll458zDm0c92COl8jUZphBRKoeM7658+m6YoZ6ogO9OHNU8rj0PNW7
KG68dXF3YajX/56xdchnWYg2Vjv9udvTm4ESrQmGjuL32/MwQBBg6odOMexN/BRXhf/I5x1oK+Lp
UWpvpfInwpnVvHIA8xIcL1u5ErVsabf7gL195OURLz+FOexA5iQDdNU0XwUrJNRNGZeGGPl5Dgtw
ZScQL5jVpp13AM6hRf3QcW+R2WQ399kAtfcXz2x2D6lsOta5QSIJD14G6+Dp3CF9tDW0vYJC2WWr
I61YtPfVJ9ayNQZ4JztOy4IGKcWGD52h0GxCkKTA97c64+4J5Wa7p5XxSbWwcAoNFd8PQ1UyMtmv
8hNZN6jc0PmFrUiQ6ot1k8KBgVIlhLpzJMmtGjtJQEl7bX3O4vli0f6Z7bdonk0TCsRsKtt3QSq8
ElYJPQNt3aCMDeeMAhkeEJXsRO1tDsyaCPEJCFTRpYSUEEBCEiMRcYZp+vbS3wuwNxhm4U2u1Pdp
QiXbtbMiPJtCIe7rJgY2zURYGl6DU01ASKw0L4i75mqyXmjZmX+0AXguhKEf8+ES7Uo4Nl0222Dy
Bb1+qKvqySjSzl4A6Y3MnkTXRHa7EJeK3IynH5vFE40iJq/77Qmq4fhdadzg/Va/Qfg/CyLL+F9P
p7RzTES5K+YC4Fdt5TVPYAPoPzjHfzW0L5M2916wf20NHyqF0BuaI+uNWI4LXQ6yU28aeIQnwEZ1
IkNJxAVAt+q3VTsIg9il9VpgZrTfzhMtdyu2qU0NH7q9hFztvsRp/URljlCa5iZVkCcLil0+aorM
5aU59pApa2SaD97ScMCH3fyfw5ftI96fjXQdUR8chDCCnSKCoRsDYe8u7SB6hlDE7g/nWJ9SXPCs
k1030aOUNNb06tJD182KmN51K+FrNmilQ3FtH8FXTqyAe7sxR3L35jRC1DwRp9W/5RY7Abz3EayW
11KfsZGZR9bioSBXFeWOD55YunHI99SkbifAGqkOmt2axZVY5RZXRhRpAPP0Yg2/NzxtaipfNM7e
mnuuXQlGdwaxi+Ffk6uOTn6flNfjCA62PeO+8C8JfUnQm3Vdu40efI491qUTKMe6z9dQ2zGlYi5h
Oc07ayb+E9jwmuaPIONQZ0uh/5/oBXXNFCuHq8MRqfV+7lRGnPtdN9oLMR/tiPV6aoKRzixtVWlt
pIj5xhy88nitq69In/+DNP5nHFMtrJIG0EEgpn7U4cKvEuEvb1W/ff1Y/VYfkQvm/lZJaRNRhxZS
nqs0PGhh7RKnBwLaYXCW/GwJMB7s6hb2M88XzK6oT/hH94qyGOETudpvIDrMSkfSpm0imVd/2vWV
/racLFcD1ztlijdCc58oV1BLMQ2Xajf49Az30YOwfW36HEYZJg4NrpDh/aOB/J/iKx1je9dTjcwg
t6aKonwpLvqW6nMcCqs4zEeGAIplIjNwt5s9K80x1D77tUsolz+7nPq65i9Xdj6xeVZhO+4EroJc
f+THCIimq1HjlLjd8MoXeiC3esWamoyVIFBMQ4KvdKMo1q9miS3CYAjY+Jq3CzySpTKfg+GWFnSV
ek+DuiiaUVAPTJzCZ3uYwxaCySwvNm/SLy95O3e2veSyWR4JQ4pbIJvOHZS1nsof2wRkfUXHXrRs
5FnLOpAwOuZxeabo0pFdhcqhnqKGR/WCLWh9ml9BHsQC8sDMUjvPfFjmxlfhdIiTD75gxD5YNV29
29YfEl9fbmMe3ZDFLtxxb070WrmeTe+TcfhwEcTqaDzNC7KPh/Pteb5IDBVdPXkPmwBrZNLf/cOZ
xkGYQbIwrt6EAkptFxAeCnuNrwF1QOKbNf1Y9gekXfQMa/8Jk+YwWLc1i/Pz0lpHr2+21Gp66Dtw
hJhHaaaR80Q/1NpVMJl5UQYWPJgn9ApBZqcr7tQYWlXbhSymw+5pPtkmfXIgzcJ9hNEASeSefHvm
gataavLUeQZ+u2HhLxUnDvYl+EsVefiKYpqi/+uX9xKCGxZVoNqvmJjNnzWiVGhGlv1VAKGbepIB
46q+sZGRWKyv3SlHxB/9RcVvV0a4LtMQoDVf7tayyMq/2d5HM4n6AXQqAX27E410+Zp5KVLgOSo2
9yqo9aofJfMyxpNWkyB3Ysj6IeM9lW7MpJXQJsXmwWifNL2Ai22PyJgRTPftBWqMWtZnMle/o4OT
YFMHcJDc+8XWu8bIIiTCx8qkSbOX3dE8JoRiBW0GGRjU4H8gICGHNGK9VfO42O2XMc/5tzPEZfnL
3ccQTG1uWmqPzqZI65VcQAcuHeHgJ+7Gpg8W6WuZLj7sqhzG8L4bDDaNjiMvDWCrrb1F7HSDwpfo
1mHnJp1qa2oIgr8BFWMUBioDfh+lLpT67/E+ij+iGoA3AWCFSXZ4EDE27H8tet239VRSW8ePO/WZ
dTcmivKwTbTipAba1DYmW32jXLCiQpuwhX/Q9DMVpS8ioKqZw4Tynl4XRh8WeMpS3ZEcDu4OmcQq
x2LqFLnAcB6e9HN/z4lTRANv8EyPd4rr+UiMsNeWLqR1q0Duyd1VLjX3ow3cDWzoBZCVXUwu155l
ibsiqqQKJ7piyz8rnix8lWRrEMaslyR4msojnTbQ9QhDsfI8Nnn4aHL6ac0Mk8Cj9AijqYoV4aSO
IPpQG7QwuXAZVgxlgjqEisb4QpjLGPSBSQjKWxOa+7ZUMn3PCOhPfRUYKT9agHISlTatTmBg6zrv
TrMEyTRWIovC4Ue9U1vhh+eXHm3gbXf/yzbdQL7vh9iv+noJf8P+ogTqLAAI+zdW6xFsOt9pRhLv
j4/0vhhU0XzzDzXAtGzbDvPn3ZH5yDd9TvTN6jt8C0RBoNhzFEBFrKyqbuKU3uKlZhyEeLSU3SVn
cXtAqxvDhOq99SuDj91gxmR3wSjyy8yaYiO+tHN6xRgFbbHGrbFkCIEMCwOEQ98xQEJm5kMJ1shn
pjs8KHTVkZKU81D0UkVmCoLOpwR5VKIT0bsCDBotCk/3DP+aIF5iKoV7ywIjtPw3ERkzYAO6Oaf0
y5q5Nt1GR5VUkosvy44Urzq6vZT3/V5FqhUJf5my7FJkDGjpAihQm2A5llEZePgy5TWnYiSmpSa0
vk88QOWXjNU2jhWgpxuASRdQ39i65dqBUy2cewXpobHlwmA+27j35pRV85fWQOnqVVxE9g+sT2+y
+lhHZbVAzD3djFxRxB4LF7+9Qr6/lorRW25JMdpM480gEorb69UlsWp+sCRxOJudaWS/MDmik66p
qE8zPc4BS5GSxGi4h0lV5gMFIo+S+/lQHeDQsWbutLDl/J3RarLUiN+85YlKrEY64XTonodEmxs8
4NmL7LR096pPcisK5XMXZjXWMU1+xGpnHt94B+f7r0I16WGYtLZmq6xnBJCrqZMcbc3HnGDDDLRC
ie0G9NUkfvCDZ8X1aEMqZaVCMjCEftVnAXedxpCFcvBGIeHvm969cxxbHaSmEse2VLwIcBhT+0Km
3PeQynZyp4WdeKEmhSgGjyZ5Euqb8HvxKUHeYlV/cZ6I3X3eBctdnZ+ci3ELTX70u1WB0am79y+/
K4MwwF9AeUchrmkPSPQBPHXrBBTqHBMEC9hE5g80BJwsnZKLKxhMMUXEOiva86ejHuaLkP82IXje
TnwK7x0aCPpw+3vTnDQQXSDKsUeS+EreW24jtwFhwGa47haGcm+BEhfEGZYHIzs8SpfjqtmXiZ15
RpQex2iz7U7fqcNRTzhGFKFlM/m9/RVcMQSJHcQ9+4vlASrDjqRmSYBmrWiJZeZUd3sMFv2dF/ee
WLAJgwp0WfE8M1KFKH4LmLqLQBLEJrhUtAMZ6ImoOvtixvXKh6xCFw3+wnQWn+prxX0Tr6y4uolr
BNZyIkvGKIaug/WjMqD3NFM8eQLs6kNXaNP3cRVhaZ+wpZw5qeabgc+OPYiM49cKWEG5av2fDkv3
SPz5ar4Jk/3So34A8rsi+Em7qzcamgI+QJH0aZ9iMwS9yt9KxqwhiMlImM7UdPlb+JqJHgEasnWA
dOFaSFa4yhK24ZnLZuL3suefXS0A2s3RW00neJBb6ocFz7Cuy1fjHs2foM0MCYwkZdDMQzHfj+68
kJtyWCjc0DYSVY3hFVwTBO0lK8IEoXlVvAL2ZL/TAzvq6+4YvfSL5IstcrCEofQXncFVT4aajlM3
vcxEJGnB4eBR4EVPFtPXyfbqSwiWVzjdMzGCqxFDFxlLi7fBYoXYk1fTlPTZwFQSd+sKQ4mszvTv
gDy9XAj11efknv7hhPNuFSeluz3sSzPYWs7m/JXtMsVyb/bfU6ig3/Lcc2I6GGM5KoyyI7DkXXMI
0y9lhc3QCKQqREnQb+Pl4YPH4+EDP46JpzPu0T0eg6KlZ5Yx1AwBId6cLtpZPU+w7ZRqhOvg52TE
RSLCX2+7C9mYt8+BiqmHeRWj+LoXaHA5fGUnbu6lQyQhyqo1H1/CGyZwaAl/657uklqR5/12fgIh
o7KFIc2pG2REtDJ8j6Sm/t9LFBSFccTCVqFwrFT04f2O2Fp8JJjYwf9XAO+g+LidJKCj1srGdulQ
lWACcN9LpA4cheP6v5S+BoH++jACn4Ugzxjmt8NlJ9zSmjZtk6Txe7cZYw425cwYE1unMj1mpaPV
JlAOdRkAwBP10D/1TuayA52WygCiUs7V54eDIm5zm8HO/KMLZloJaesoHBRiyN1fhNYB7D367YMf
sIDuQDeXD8rml4CPP1g8tffH9OYEGTxK2ttw7lq6lbVpXCMLcboONwyGS7GlFUaKv2BlEP8X/RFY
CDGNKQQ6KmGNDAJLCSAhla4w9JnUgEG999eU7kvEw+hD0XuR3xq0/hQe7tCedv/iHtv/JDUVpSLa
RmR1QbtX9Os+dCcdlsJd2pqjNSFYnZD3XnDnANqPTOtk6g33dZu19GT3JPZma1MHifDLHEE/bDgA
VJ9ci/7SVODVVw3wR000gGrwhXLadzi+ZO+NBVj/ZXW3byc9T9NydI45pq6WgOKjRq3v1jVbKaU3
7qfbarVUL7fWarURvWb8HD3plr05u1Ul4N26GxgpAJ8kXzRuHcm57bjkt3N3LnLiBaE2aTysA1hz
FYxl1PtlGryYeJ2zAhYpa3rpqRYUMMsZCXyBYi1nh4b1fUThNhSgdNQD6g/mKDuUaj5QG6D5i1KZ
yy0VrPuZ/1WG6xyghaox1LkCwYGGsrQsjkxxl58PN6KltvU0Z5xCc8yi3U+0KQ6YKCvA2kdOsleA
53VUYZ+MOCIOk2HmOb8I/UIiYdjv0Mk1SVtSOT6VseBF1FEQdCpA3+LbYh+20M9hZrb01y4PegXh
HkBJNbqVHCzD2JSqwR9Wch5rjFp3KC1SKXuRoTuanIBNi6/iAft4XivmQn6TEPW7ifV6k/2TLYnB
kabdFkRnRQjA/1MUX9fUeuLR+dUUXkDryoMmJ1AsF8SJ6UZPqEbFgCj89ubg/IxKnrajzDKBBz13
ew8++OmQPr8WMZylrntFDNp18L+xPT+deob+CluFJGlr4qLvGaW4UxD7vSKoUmEzYwKTGIA1ftnJ
J0JCeeSwCrlj1Ar57Vq+EtG5e67tj3cPpPi4cOzIf8OPkOV/2ZWhrsmU9pkCLca85EZMw3BOTkfc
0zLw49QjEO+12hJOxC6ujByH2ZXmLVIwPZfR7s4jDF0XZAWAS2KnGeT1I23phFB0uVkIZRhMWWFb
Z0X9LVCzu/Peca72n2saNc9mQFT0+21PIN1JKA9r5rEEsS1ihfFtJ/QfOxr3r+al7N1QW08b9PEz
VoaCEf7EG8Uo6EfF6jxul12nDjfYqQTVKBgbgNIHv/WBYeNpMaKBCGnBKyF5cEEdJCOoIRbUboJs
GPhUy8xwH95BUyXAMGaovzDuz0HtGor9IAz/fKIdqM/yCuY379D/gm0U4GWHEpebEifaHwGy477E
s9MDn+xA9fXHGeAUPGxo9EppgjckZYfTpdlMpeb+cIy4cNs363rqhkm1dAi/nggsulHYcaO1737E
MbAD05llh5K2STpNzp/Klc5CMFYgXrK4AfDGIxVBsgohga8YBMjGn6bQIA1ok4mCU4bE/aKbJLD1
EWmJyWoNPrgceFwLOnDELvQ2uBsx1c1v/cI4Y+llxfHsreSDciBMA3+SDbYD58xwy7hj0LXh8bMz
l/rQknyVU/SVx7ewmJpEp4kkl+OncUkAiGoalCrn4cPj1zUpXt2tSZ4M9Kq7DKA1yNB/Lvr6VAXE
TD2JDDDn0Pu3Tg629hwr1p/+/8YCZUdj7WZDaEBpw3y7JTXt83bQag8saRuyeEpUFOhOcctwHk1U
o3jw0cpjdALypZa3YfeADZWFYAXaoqyk2UywjzhyJ47MhFvC5OqPHresiA9tqArtDC6lFbUGex2j
030O5ZLZir4AvQ0hw6UMSB+q43SpNL19FKfSUZo6c9/Rva15EZ1SN9PhkEBKhlfnGVRgUzdVS6LU
tNp6xgBiq77f9YfJWKjr0hLZdQxk1m1FaTsmKpqVU2jzSjk0tI5+bgkmNYNGPAmP3BDzhRwWCebH
iX6FgceqOs5YDexMnEii7c9CShas4aQpJZJm3dGx7tnBtvlT26sHJFtdvs9zC8Rz/vWFRoKXXs7l
VhZdDSvO07IgUaghiHvTQCVxfAboNCuYm5S8lnOtPU1u3oDdK11TK9lrvkmWvnesMMxjklD5ZV9u
+uwebope5Zj73pCusG1tHveEPcxs+yJ1FV7LFckzFGz3+rt8aowlbSZ5J8bmbUd1PGv4pyj9J6kA
eqvE3vBUhaS7sxOYDd3y2WxkQqLhOaeofuemRSxvNg5QaHOJgN1bDU9DqbsYnfstmlj7jM+DPq1x
WFRazVLmZgV42CsEEH2MjQibjisxeNSrxYx48b7UzdsLUqfordaeNGSRA75RPcgj9mn5hrHXI1fx
BtR56U3RsMTxDp+JNIv6s3N++aFCll+jsYikKfc76B3B59Yf80jPX/IxVAuy/b0SWQbLBibMcRNZ
8CdkT/vhiJU6Umlw7n98/Bg0DSvSgn1TJ7tiLaYLNOkKa5/7rvV2ksODpseEWF1gDgydkey9OS+5
jLj2XqqrZcgz6viLVkbh6eQULUEqSuOSkccLFbL1d1NCmmRrlWHNJT1KNd/RUQw/brx1QUVb1kCV
bAcD2J38BYv6xqUHBOPBqc8K1yrru3c0eclczqIC0x4ZKikXbNCZ4vlEgjAHmaE1Bjc6+UXxcwrJ
37tLDnGpkCddfQgu7SJv0vRKPX0gGCRE5/H1itmo18G+q53qgmOotVWJUwvhCdYTZ4Wf5Z/NNwYT
FXwkMj37dOm6XuHhJkzczW/UOBrMC5J6oAcAF6JjVsOd73G36kjhWLMRj3VNY6OroMeOLgo4DJSi
pKf2XoWlTG3knlO/GBEPq49jGeZuReCHvUUbiYLLFNZKq4R/fY6AShrClbnYfT/VcOZsuC2DzGqX
2ASzyd4n0ncP4POGMZOG4J1NqhSMoSVYuWAlmHNzu7AOnEVlhnslU/kRWdAxgY8E+yl7eGau2vN1
jewlfD275rq93Hi0tXvTWZ2dvvxQbFHUZbj1la4Lf51WC8jHmQM3FFVBAZZ2xxe6B+y8os6KumMG
TR48L/83xvK0J+430xNpK7OuwR/CNrxBAV17Xs1/uKaNu0dDBQPAa1f54GEAuetPIGnAbLvsRENA
zpG1PbXkZfQEo+2IYmb68q1tI91r+LUNAy+Thv5IM321h4io+6RcZNiAEU5LmargoqZxcW769Y/8
uCbfuLHp86clKwvGHc+mgOPYOZZbbjvoFDn9PHnXoZuejDgvUNkmZkTXT8inbElvPy+sQBZkAok2
RSKuSusMxvqtLNS2HOEq5Qrf03oFxMNoVCIda9H9CW1Gs9zs8H01W1S7SYfUFrSj2Fnn29+iX3Rb
3uLhzLdHdpSrRgvThkLNoCPt08vtEhP08KvcS0eX7sN4PWaJJAcSd2iFXEmPVxR7QR7PM7Ezzr62
HYV8vQpRSdMk7U+JbZT4T1RbIp3GjxsDIHjPmRbA4aB+6meUJUclYKRSKDz1YYhS4UDHjJBViQP8
eRWX0d9e4r1rOzl0F4nq3/4YGtFJK67BrK9JgeXIXhWZdNHTqn17EzW8v+oyKycyEwztMpvpmhw1
NtFCNHrOCT7rwoa/5mmYTww1tjYuhxGldnG/EBAFLDhoLpfaZHH4AEesDrTBZS2UIFDv6EiiCJ7q
THZBfCiPKTZocYlWNuptkaf5t6UsO4HMfCF7kBiF5TeVgN3IUSnfPqhKp2QK85nm3WYBlS63aypj
xlg6sdTjJWxZd4GPK7CxOhb3YEDQOBylKuqZVOCx+GKQc+nBwVpWcyXyfW7hoT6dfM8dsKfOcs/P
6Ajqc6I1ZR/BSkOFjcRJapfr8ixFW7BFX778zRtCm27qMVNwilvhfpAYZA/SsCylAqLCzv4psiTq
EJvRVpKkDA2CY8G4PkrhX6nSus+UmNVLBmYPJMhkX7xEe80v1VSdkCTcRgokvMXFPYuSnz18faqc
OsWwWQL1RE+qcRunuLhuf8hJZMDG4FSb6zuV2QOqVDQXeoLp6KD42q/g0SmTPLUtCO1hEkIM0ezT
oSeXny0peDLrk3i3ql3s/2ZRkVOj5eAS8WF0+hsEvRmp2TadkiEZVp4lXPPd8JgIUgL3/K1s9V18
oraazK6KsI/6gmBCgkVm4YaRFk66JU4OOQwRBZ5ZI08MV59Lt7pYgTWRwH9iunoKKpFxUd6s1Yib
THP3LjF1oLL7nj4nS801XDh5KCteS4QXhc3RE1ErMBg0U6LdwgPWku720zxQexOnT7G6NnOMqzf4
zkYVoxBjFn0da2tzYGN9sf2W6Bf3JV4pLX14T/1tN3C35kLcpJngw3ztXoz+xA9zPKEBei8v51ir
aYBfyingYZFGXm0A3sTX4qmbfw87HvYFazn2ORjIzERZ0wabuxS/2atMpRsEkDvunRiCsHVixmHG
aqsDv7XP96Lps+ANeDqa3qZ2fjFJZC7VJixujRQnaSPzu89C77C36Zwz8z2CLEdRGjv94+Ci1MXQ
PgpQ+tSjMtJtkruuYQcHkAOH6a2a1Y3AotcJTTpqv42w4ll+TqcsJxT5B3h2WGqYDjmOq0nGeuBG
0LrIgOQPfr+yAmLCDEu/haCFcWZZ7XbY25Ch2aUVSYWtpBQev2+sdZTyaQbDYVmv+GpYOiVDWaWu
Cge3MajHMbwb3NkpCAIxCVbiO79LONyFP001rkMgfEnV3bAcPsfYE98ucO+plu3SsXIvI1KKGfqL
R3LPSdkCX6zVWLsSsGRCLUEpLN92pnQYN4iiY4Z1TkEuepzpSxCyJP8rahrniVaX9oFp1bvJKXW/
/Ky3+CoztSYjT2HmiHOwhEPGAwSFH7VI4JOahPJFbCheIzkJ8g+Dml8RyvwftLW7DMhWaalujAQQ
/R2slJJc3a7hM/v9Pn8I4P8apiFA4TBJo5NhIanaO9s4uV48DwXtoXbrKAc3bz/QO5Xp4FpiZZNZ
gTGgu6pROnRgAN/LEV3cfqPLfddwMFVOztdop3bz3k66FN9yRvoMyKgNKw2oBTMO3A0xj0spmUv3
eei4fnjd9AyuekPxEC50nsORmQ1OaqZ2yzJGntAoHVnQKrzUWlT2kkor99QwVOxdPLRReLe4lOXc
+IwyGCe/3L81YQcOOw1yOtYwW/9Yyx+5TnOcoJIQMxmBL90C9YrHpem3/bnRlRapwUqbfep8JxW1
avVvKUHc6kV60BWai6Ggy3Nk7vaZ8RHYelnKBZfycjFZzTejMvFWCq0mMii2c/wl9gN5ZwHLU+aN
fq4KOq8DU+5b+smL5xafWp3MKKth2Q5Bgy6DOEKgCJYu61oelp2yY1OC7aKhmsUovZeQnGgHzUug
SygM4ingq2FmZOhxq0PicsDF1OGFKa/37FYTl+fOsVCnwsRZM1O43wbUKwJGIy46/svoSgF2T2rC
24G+Z1D65gGniZK/p0Gd5rsSFx4hU9BGxNTAUfbcXAb/OYqzcK+omyy82v+/oQn1y7007cS/+1yk
K0WPQ7MBEftm7Prb7Egog8DW3GdeWruuIw6V+J/qStXlHMIYQd+v1FJg5mKOBbKvWGoRCfAAdypf
sBQmHVr3lpDRebYZeABiYuSfqEpChNv7JNT9pcK0m+xg5tr73goKkg9abI2pIiw/DITwMA5WxMXs
GyoKbJosqmaEE+mXRouI6g7qAr8Plng1jP2fxCzJquXT2nFp/7JXdX267rF2DAAyaSk+7H+UWG4R
uHCDlkcdRSPS5hWgE/hHdjxQP+vx1hx6IVbepWH603OVOw7+/GX4a3IWtzTHXC5uWSwzwfq+guYp
t0XQXYnQcbux72XeVn+KlZiL94KcLJYYxsTrysPbYgRFj+vCUVnzDlgaKrosHNOCd8EovswOatZB
0N4dBDibm7jgTwT+pZKg6jGfxDHRdFcL7BP2CMaicO3odwQ1hj9WittXaEk8/N4aniCDQseylmni
M9O1R1+izKmDYZuGvb07PHl+G5K0WRsnq88ztYdJLcnvOj4eVP6yYN+NX9fAC35IaU/YWxwy5b54
zwkMqZHhyDWEb2zxNgcGpA1CRS7bknwT1E7nRypDPXHQtI1TQ6yF47es6F1W2wRVH9B4m6MNCbHB
VenIOx4YTcMTVttEBN/4SJ+elwtqd1dx6S9mgqRn8zF6aeIFAmNCvBZf2Ir8MNksotTayE0mv3tU
Nl38HtltrSSL5rFNgrnm3VifAmdzexncg5cbuJOzXJEZFp/yvmQtsuw3RPVRAaNm3VGJAH3gD0D4
654AKtRnfsZk5qVWH6LrKE7quS5We14Z4kkJo6if+zGuxHIXxAuk5cPVeRgcK45KFJ4BXSjt+Yv2
zSLdXqDqueQzLpo0HdYif5+4vcRzwV0fQKGEFc66k/C5jj+EppdzFCiw2rDtTdfWm/bmmDemAyJ/
4+B4amiSP+HvJnGWJCfaHUBFYNR287CYg0jsrwwBv8hZ0zp7LvuG5Pqf0DJtmA1AIM1dbXZ6FC1k
EzC2hbzCOGZ/1I2+QtFDyruwUD3XJsemt14N2OhLMGPCjOXWOhf06iXGBgUwoDxJRgf5KSd58oyd
PQt0RufXk+IRyDBe/Dyup37v2LO/iQcPEFxm7of2HYjRthdNyHyEYnDHQ0USrY4SVr9n9GlYiopz
2A/F5k47zX1Euh6fMKxXg8+XeUGpQJGEB9vYABk0F1xWVnlYeQ09yB67n/vvbrWLuUJSM5k9lM9T
5Lj4wnM/YitpluPc5/8oU1xsJiXMq1rFE0qG5LC2jrlR+Dkguk5gpbuFSRBiU68q/TK3h+Lz6L+N
bXb3TTQWFGKpXNk/IW7QTNNOCeGNNEutOjQ57+RTyPuX8oFCzxcfmxKLrZyIb7qkKjVJI4D1OA/P
4FO9UqLhie7jn0sXmL48r5eUj3KVb1/vCoV2GwJun1BeO3FwdmC1y2L6ZqDo7sZMymG3YtFzjkvy
zZBULs5w6l21AZQih0B09N2My2E7+TyNclMXVa6TY1Ga0bEPrwg18Z7+AEwhHZF6s2CdiCXHRkz3
8k+1C/nRWUppkgDpLw4KB2JwJh+manhOD6LB4abJfq65hrpBAjj1/nDBIhe89mpu7W91IRq74X9p
QjC9IW5vIUrJk5MiJe/kCIyWyPK47j6iTJ5Ai4Ys+6qzJ9WnG55E/Xa/Az9nfCCUzlFwVT8ay3d7
Glx5gltJqAZj48jUMST1R8LTaDoZuMvfqXKMKBdsLH6xUDER5+g4EeK2sCEtdeo9HnMoBs3UDnAv
2zGaUE83EW/HuUKjcVqiWeq0oeVkGOOuaaBEtYGhXYhA87kdUlxOupbwV04EJrid0/tVTptT8gUs
0XKuyREe5M/Df4TAubG5EunHAKkSaz2XPBfjXIEkPo6wtwg5mRoJaWJ6+ZvQfJa2pyBrCidA/aSj
YG64nsMmt5sguhPSuvN0fcRJOwGuikqx7ZIeRFKSz9dLOR1/qtD2ecclQATeaMmiAfh+9S2ccaW/
mVfKy2dwLHI7FhX36cDQyFV0g+nga84+fMzPHKaxDFBiI3yLporg0oP/bvU3IuM/SRKVFNfRdgnu
TZRIGo0rq1TuGi8vNrvZqQaDYSmw6kGVsaJmkZ7fyfvUgGHqiNJOXPVnZXzNbIebx4U5UYfB6stC
JQYDZaCQmf5kAgwofzHGSI6kP8cDz4ciBPY9eiWxPjKQq4eny2stShKFWfv7iezGegHCjip9yHSo
lk6jK3J5OiDR4hkeJ+aHWNSSxpdrsw9ZhILJnXNcu25HCH7Us3+BvNjSkP80xP/U7Ly5m8vYROIc
saqDeQszF3ZLqzQD3Pq1ZUzjQXtUloxLxreNIE0yiGQkDh4ff/CfRrzw3hc3bSv3l62/KfiMmi4O
qNIvN0HxwsgjmrgIgc9lhGIYbHatNfhRsX/g1Xbate6HboqQKX/gsqgFVgv5IrkXN4TfaQAq5QMx
mm1b6bY/qvEAOP06tON7d57ZVqkyVCvtSD29tldGEWL+r601K2uP3ujP9hG59BLw+/gCh6oIYKtN
GhrIEBSxbqMnL2MAAKlzyMq/OUKWZIxS+aeIm7PDqnVHX7Q05giKhzdhYiRWFs28+c+XlkjRs52K
ihWV0NGFGDnmKOik4EQzeDdnjXh/BPIezDXcHZ5r7vaghH4CkELuoi3P6DUPFPGQnjMjrJH+bZcU
deQfonxl2k4DsALLwrjTltOshTJwB7sOEfcGuDuZP90lj6OxJh6QnCeTOy7wtEXc8gKgNLZZdNDT
cGgckbQJwMv7hD6mP9wQ7u74dMXDTXVu2UrnKTqGAVEJ1f3Bci8Ez62yT/ESodn9DyqEC1RMmTu/
SE2Rbj0uLfh7nJYFTxZcNZd9XgLnKCf1C7RwqLS6MIMCmW3kqZd6ATTdHxIi9GmLv9JJwycwwOuJ
sCMfIfK0UN9+DCkFTPYHQ36umQwzG6KSHLG8GpFVdejb8ArX7EBLwZDscEFBS/3bbAqOyrFwrooB
RU/ZLXntvvWAXdmBEY69/NYdx9F5X99nW7kJug7UeGvXmFzl7IGPoRdwCpf50i8VRxmzb7gPazLZ
WCJXulmrFsibmICXO7SMnPBmHEdfYPtgEyRPtMI1cbqzE2suJzwh8fk9tq5gw2EiM+SsQVPCa2cz
JK+IYD7kbjPUyRfOI0S5Qw5DEfLIKMGLrTxTh4SdahjRjVZ1w2QJdv1yMvcMf0yFbGUIh9gPrTEF
C5zZdnhfG1nMCib9329rU5RfNaHj3vijtVMDJWCpPLGr21IGZ+lMRH77+OFdB/LfEVQPNK54uprR
qE0kLlKBdwk4w6j3KUvnF+jnk1JeEi2uvyhtUfZQRzcSoz8eNRz0wrdyany7+vV7Cqfg3LK4Dalp
q976NyXZy/YLXLNdmH85PAf7hHHYwhG3YqHOgJyFGQbw+h17/gwxIsTwasQPSGIkM3imV7amGRrF
lO8WsABDH78mBH7SCsyLeN9Bsc0mGjMZ+ZqfjTmS0VQLnkduoE3vvbuoQKblKsN6alU4syZRVHlL
lfVOOGclabF2hX+VfrMkXaFajskAL177zaPpxnnuUpFcKeqwsSLJccJfH9kjn9DIL5YDri6mLj9+
JKldlkN+qFYjQA531TRMWOXL35cnz5G/aEENgaeT+Nsu5ayfRwTDG8zqAAStL1TowATwss5yuo16
j9PZWbk7ASaJryQMgE/hwCvBTJu4NPiHdUTI5vLPLki5XcsXyb4lbdUCZZ5yzvSNUvsenkkX9Sp1
FseC5RJgyAD3tMvOaLEhNDz2/dz5SaWLmCPmALMtIvGUjxXS7utfG8b2V70xdc3yIlaOZZhqyRQ6
wbK8UMUdWxaU1quE9kYcC3Gb+pQLx6Hm8VQ+GpPruByvcN/THiQeQr/O10Vojwe5dL5JZplXezlK
D4yMbtg6XNomzFnztWdwPBuZj6m3Avh2SIaEZQHYipqVykCxz9KaqVeSdaCLycK3ano1pOt8t0zm
WdPygG4UEvlNhFmvIUaBI9SNJcmr0setvfSgdSAJOiRrn4amcdKmaLzV1IuOHUZ0BC5DPMaHMU6c
12ea2o5IzyoPPMShcwEWlswIx4Mf/ljsAGKgtEaqqwEzmF4MwaZX/X/SmLZMA2NJWPJIps9h+u04
GRIC2qJifeHHCZMPcgtsk4S5vzpB5Gok0NHOGiT70N1oxTLk0vBuRzoJQDm88oJdmuH2hxh+5wqf
0fZ9wY7ix7Sp7zsOLawXp6RTAXfHliuNNVDiBl/xx4gaXfSinqZIxN62dy8TfPaq+p0CSuYxxCfJ
0E+OVh8TMmE2IgQYRwVvYBdgJFsLWLms2iGzgpGPO6Ny6hrV061K9eSVuAjFVxU8mpbVNOLcnofg
qxL3aB72dulZT/zheHPIAp+AUqTz9xtgP63bkB31cl8wjH2eratFqxFEOuihxnFZ/DVoXJ9pnfjt
5JBIeIDDKTtnmHi+wTzfvM7sYKS7AisbthzymRuqupkhYxODIPY+A2+ZPChGiGwZhN5QJCX7+MPO
j2N3venOCsrZVq0ZiKgjDUODs3lMkvCbKdHWJ/kcsTSq/HExZu0pDxtBmwBQe/bV6RR4tNqcvO2i
JGVEYvUIbFbbzi97Uoub6nmap1nGvTg0HJjYKkPbbS8QHJ2JDTdLdE9gNcvjXBuKMHFnXG69JULR
Scjg32RfmwkQACY3TeSqYW1SZrQazCtYGSyXAsVTiB47Z5AH5dSySgxmDfT2OqGPQwGYuHMtTX3X
VCyKfmJpj2/ds8GbbaTWIshtAPYzkcj0JhLnIEs3DXxvcwlRE040T/3a27ya2h6UN2KF2xqYscD0
Jd2ph1s3jrHwT8izZYO+Kk+gZdrju2k5R/39DRZuXMk6Df+sbC1hbhI+Ga2Y4xgpJr269DFmg5BY
d8SqvnfYfJg5WMGWSjxfz2I/+z3stRg4Qy08dv+GY52YDNXQXOCId8kKGM2D+qGCuFQnqzu4rT4W
EyEG/Q36oNKEQsTdscNOZwS1zd9OjLAL+CRpHnt4L2HA490Ih1UTvRs46qizEBRvJ7ublGfOyZyI
+cL8kB6NcqOC3tCH6pK0JhoYRYdt4q93c62QzWfNAf2YABCigeQt5ccMVh0zSY8mljUl/AjSzEuZ
5zZZ0ezeKVO8v1wlk+61Sp4AzhN/EttbFkR3xjWNQ0Tun0v88Qlqvg+QTOsui9lQpjyA1amQ9x1W
xhdhAOrQj7CxH9O7XcnkTeZsGxHAU8iOySU+hsDc/V4b+ZoQLOzMjLZtJiBbnC+PbKl0t/LvR65k
jn88P3Og5Ff8TuWAhRPa7bL10oJh6SkqHmMv4qryvuQ8U6h5ynw6V2wUZ8WCfpnLOB3yG48tdvrK
IsSkZNM6b2JhLaTZV3kE26F0+hFs+5AOAXJ6sOdxF9zMDEyqmgAwnTLDHedCQNXVeSO5lbyEC75p
Ix7ORRIheM9ChpbAXfZAoEe0cZru7e72WIes3x+pVg0GENyJQGUiGsYCUOAD1aJqwUB39JUvpJJ5
m/J7SUtpKGlNTFh7hPaUJ4JVzU5qoXdJa3jdESQIzZqFlw2APSrw+iy8bScONm6gWVoaT/63jTsp
vzK2uNwAw9x805snCKKhWzrvBJFsjqGc8pci/vGjs9MUyf3dV4FaFK58YxKJDN6bEdo7gIjWWMd+
pH5dGcTGqsj3v4aB8+g9Jl7M/PPdOtS9lsAV71ozE5Eo4G9ByvA9mkYaKAWarKignTtzHuctjmNC
ttkI81CncNjpYQosGWITTU0rMp/XPpfF2tIsaAXfgMY6c/AjSlkhLMjkj4EDWqQB0D2izgjKOXhB
DpCaDKFhl7rLSyLBU8Bz+vJz8JuKcgTD4vjxvwoOXPEJGtdonzUKD91ll5MX7VqmvcYLN8CbeNWj
RpPqhY69M9GideWNDEyCgHqUGLfBgQKF9aBw8877B3ql/he8G/sh66lxTnn/lBx6QxFNk9UJWp2l
KQq0jazJbISxzlHqF3M1Jsz+FJY1HBHS5T7tIQCkPN/y56f+aHuqD4bc71EGR9cefW30LLXGXHMl
Jruu0cFzXSAQuxvYN6IOWJ+EqL3vnwmrUbKmCEb1aUGab+NCa6sgfYlqfjWcZ+nX7cgLwojP9yR8
w7An98LOcRq5aF3fhdixkGa86hRjVqEzHRzuzk39nTeXrwIBixqj5Um2fS9HDUAMjCTDTTQIbC8f
W6l3vD+RjSQ2WPk+rjZxVp6Z00Vuzle7WJ6wV083Jmkhbp1L4gyyMQ1Zt1jeBy9KEAEd06TiD4/U
4IuAOkePO610ZDVaMoxHBZHjZAKoqxtnp3RweDZ6MQP5Xv3UlAGUmTMZxQzw2bC0I6lLOlQGnWS1
mkPAaRsHtCQD4njpxZLVYO4FUgbriafWdGoNU+hTGvJbLh7EZTkWGrsvmWek9tg9k8YkpR23POgA
XcYXtMuCikxLrJTECw+pEUIlR/jRHa30F4Bi8+bVCNtF6ulRhKU5yzhYm/3P/KMcH3gC+N1qbAVo
v0JKSyGo1z2FgB8sfOeAQlGczfnYB0toZdxHmPWKApDk6KNy/WM7Q5kL9ODgr5vr9iAzsPTYYQhC
qs67YBh5FJkWKKVi/nJzTUyW8UB2vVy+wbyfjyZbbamzqag5vojFeQfieJ9eP5S1feSifHwiHc/P
pfE2k6fGXkvNu/pc2o5u9IbjeGOmqxzAKPyjxzPbcSgWLTXrkLd0Nz+1IWJFTMHjc3dN0uh+aIyn
+oVnBVvn3muh2QJY4UZEqVUX0zGJ8jLTeQlBPQHgRVR1G1qUYznLbpFRMRDATXtUWlORQMybM4x/
Wf8FpnxRV9fQCbguZCeHFJW1FeKgtOpmMhYblVCsYz9qGrr62/qFKj7XMTVViqej3VhZu41lRRuf
sqsSZvqRnzKFfxadXE/mCHb0cHQtGc0q1loaDPBxNM7C2rri/bH+ytf8FpUGNtolLLO8haDFDJmS
ZX4k6rU5JCfq1tZ628EkJoJrHOmFeneV/fd3ZU4qDvP4jTvGnYYk17xhjXydczhrClGPa8xTpyEP
ZazasT3gckO1H9OG+PZuYjR74OYLKCkYhYdx+oo5v28C/o0j3IRMVirqpB9TfIIR0XfFswPNPyJz
nOOKetTYZzjyLqh6CAKmP0E6GZ0Weta6Fq6oEtNvWknH6JQe5B/GLWfSKDf/Xvpdsx7MLPQzk4nw
LTtpmkn2v/EJ8un9cOu+dP+8ehdanJdWpC4eNGNH4141icwUd6fXcgbs7qyhLdxxbHtXXl9Qa8t0
RHlazE8kzckoAbv6yX7VCkoI6roNYO+XxOj8LPS1FVUOfpQMQeB19zOzEyLnYIo6HQASZnM2u0ce
W382Y22dN/LD1DtW70sFef6u9j8dHNscO28alPNvKn0BVYxhm5jmAvLXeCSm+uqutrHOganLFAvJ
ZFbKxJxSkTWMBtciUGS91IBJpT5K+GjHHo9qswdIbK+X0p4GMcHSJ1Vn7+SdQX/8Whp8t49kba8J
XBS5xGUaSUTlxyzdUVtKD/OeKS9fdGm/BMLtkU/5626ioPSCSAblo4FkZ5zttX2ZwWpXkJxVWy9z
awPAEuNF+ZKLTy1b1c7+QJOlyjJmT6v1n0dxGdb7Fx3xp7g4w65fpNpcuhgidYH5DpiIV1bWmvOA
tg2oI54vYSw6Z+ULcTjfReqAINWmWcAK681xiooHdsDjabbAyaGARgbKFqih1Z/Ie/Pk4OLJ+URr
/YHbqoC2IQuD27AHxV4QyIGgClCy3JBAwS7oL8dfgWhDkYHrBfGWQSIOiYTczCcdIsPZgDAZx6Oc
noagCMh6yiaAlzqWn12QqqNecRb7RRBSHwwVZZrCH9MF1cI+dNHrmlKQEJZ61G/cxhlrrXXhFep3
JXaINhXwQ+uMIBo5UomclshUM0bQmjgsxVIO1Oz/+dwZf7Ls5eMGHhDzhFXfeW271NfmB9fgXjFw
2Amx0hNXzwgfmYFOLzIHcb4ffYWBbY74cc6d2zIhxXU6AaZJojyEYYZ/3Vclhwh3dl+SjJigARiY
PhIktkqYpIL9d5GBiJNWEIdE8eMSyOs5gYiguFcEL5LhQ0eXasLcUuY+c+hp1WXLCKU7S991nXq9
3d4iakWReURbT6vumd55aRcVrXIB+LhepGmNh2BQHG+SnJg6T2DmlMrPQPQpWYZgiI20jsW2qTns
jPjvJ0PHXsAMOg23GnCZlS0caIDjsFBPd1seZA/bN8kpmpYBYKX9S8e2z+5lr0pUM7MiCAOcbOMD
nlUFwNhnqoqllENL4y56B8UiakcAOHkkXTFuTZ8wckmjzELuFwrW2WzJF1Wb3XzzB+cLFQxMw8X5
bYJiKHXfsvEfQwsWX3X3kFgckd5ogaLKUw+CV2CN7Qk3PvuMm5MJH+Gh8MlNpetWGuN/D5X3tVdQ
/hfgrxbvSuPKgJMuLfT71p8Y4nvb/g3Km+stoNNqhS/4Ioj91Ylkg4Zo1ChYhR54FostTNZ9JjSb
p8bqJxZrXRg0fN1tV6y+xDYuOjZNsEzi/sQ60VanvY6ezvLax7un8108AQx3/Wlm773r51eSsLUf
h7fy/PWQuijU9rg1ozlmlBQRlvK/4f6esR8S9JRs3iQtohsQ3naQowwCqsNcAOMrBvfgL+0HgVwn
z7bL2U6x4T7Z2YeUTVM51Sdg0wATbzSaMOBk2zjHqr6WlmAQqsRxxYih9dRaSEZIcz770Qz1Id/1
jAuE3DRlW7NKBMERjor0pu8LDFl368/5p0k1lvLbkoCswxAa+dZKHNvrMEfaTqYgm7D5ggdQK4r2
FnhdDyfU4c+hIkv4XDSRsW9Hclt56BXtA78jx0ULdPZ7bBbNt1G4FnqU/sbOMJ1TmkTr0Nqv849a
ngqdp1C9RkZBpN51cO5I2Ufm52/DHXJ7n+ap3sNYjZjnhUuRpiP1938Csrf1ZtKn8l/ntZywJt9S
B/hedmycha5GWO6YRPXZPrW5UNGbVaJWtj3P89F+mbZmxdKSOwYUMHOGWFdEwULjML4+pkQ0gCqu
IuBo3np0EuJIsXkC7WNFL0O65m+Hj3MYT4rLA0S7WPpLndKk5eQ7RfZ5rdoIzDsua1mQoeBUwuhN
oILNZLPiNDWy58DqCtAX3qVCly4P0YJ/4Tk9YBRAg49o+AqbDWmJG9+jmFrmm7e1hk2ifuKWhEp7
9KF0GxaNcahA3WDSHsPvIYohwLATIUoBdzCu87js2oFaGY+4SQPjkgTPjgI2CYaz0Yz0ULNddCuV
N+TweTni/XhSR+yb8PzbN3G9ypplO0kFI6AuQjCmYHkI847UQZyiXwSCPRlTRq1OT9HNAiAvWe7s
gqYELclycAIVME7uIkXO8PE/Jsju+I28sgfemdf9lx0h8J/y39WJKahkP7JCMOqCfkHRt6Q/3ess
P2tBPeiyFN3j07XKWJ8s5iNdgUKtVFQqrAYA0iZ/fdHV650/tIcPttuiHVL9L08ZfFIZSUSNXj5R
5GJI4yXT6XQG1/jhOWNwM52lrx3d8UtDRxw2xQoiaKzXLi8kz4lnxBCBFaIPvCp/FOlh8hlCwGrb
3PNDIblCDRUHj7L9ZbiOepeMOL30elsLp3/aYm/d5lCdTG9AeZIBofrmLkxOHRC6C8/bvkZV4MWY
/yoQ+Rvl6M/esInM6YHQf4XZMveqni1tWrjKmco++FWvFPx6kh76CLzQvKCZcy0yvw7XRndDe9NW
ughessBC+BrsJaTd7UnJ4gql0xeu6Ow2CO8XOzuXmr32e/ZCBcjH2r6Vpr2Uvw3t9lNMzQAbbtnL
NgJFgGAHGrNfQdxJEC8iRyEs0NGjY/2arU/VlbZ79IMqPCsKknATplS4B+NT+Ed21zsANGT/6pzS
oUqqJoLzXKrAYJD8ffJREKTGqLmXzNA99B7BQM1ooiBW4X6u8RMahf685mT+AB1RcvvR2wE8wGl3
EYhpHIDwQajAkfLN9PXjEKo3D/K7ZbmJRO7+ViesRVdTkd6k4eMJ+4QiXphs/6HPkwE9pH1QzLDB
EGhH0Q4IkBD+3ojVCZfzCYt7mbg0JaDu5MxZ2m08Hh1RmO5zjj7LRirAkbaVZn/ryMR9/G/m2Iul
niHso3h4ZdWUp9DLKgC7Zor7kKnHtvEdtT+3IH5YMnjOPojHS+/KUYnhdTgbdvnTYxM4ZoOHdt+a
wJEqqHaGjku3l3B0XZbbQ5CxeQJrXtqcWpipItfzpvVFfc3k2ON0OIls92M8DOCAxFSaa1XeMsoQ
vOo7xLguHiLM5ciKAHedVvLolsB/a1TDq55ThmMvPKnYq6G2uAx6khMFYlLIKKtYrJfT2TUU4dlT
jmR4gUyyY8ZeOrc+74l9TMpvyCrXBk+3TncadhtIefhIoRiWCI7g/ln1fq11i8Giwl6JayiLepYE
mMDYyT2poA9B4SIcxEOJA0bLsB4onU/5O6bjscPqTJmcJulhVo24RcJGV1BRFMKiYy/631yivLdn
TImwZDVaD01SMUIRNrOSZ+nSRFvQd36NaS12fK6Qk8ORgGDvVR3lOPPpUPHKWXHgWgmTywHiV8WT
lWXXkG7MZXe1/g9fpahk0XvpPVFpgeDIrz0CWhIqp2MUoBcOWuooWDwxjbcc2RXl0r+8Ouy5L94J
NLjlbHwO6hrNtJaJve9plQykgf2uoWrnX8N53lqOmougYaVXsawa5Q2K0jo+YFTb5CGedhqaE1uU
uectu2ihiwDgTMIsIDrswsV+N59afV1kGhLORKFDYxnQiIrE9qheM3/n0bbFuoxw/8MKqsX+iwqU
TvbpaNR/zZRP3r7Oa6JTqazDRC9U4hTEGi9vyu2KA34BEXARgiuMl1rTGYbIWzQs/UQMRl3mN99E
CxTzat8u1vu57s0Yt4b2BrCXDZj7QTsQ88uIgjmsg0H2Ef4Kfwr41UXdSkDqjSsQUBRHsR9BAZ4f
f0yN76T7hKP0+8uDXXASEf4Dd4qW2VTRVAgWpgjb4h6WsuiZDqQXE8c+hbg/iyGVQY8r3cAEBGoT
f1+Joyk9FeoGmd+D3uZWtgiSt2d5hWMBme8MfxeGlspbE0pTV3v7TG4mzBeVwFuepp2/4w/qk+zm
ncpv3c3J2YTLxDjj9uw+WNs3d2pX4u+S7JX9XQvNlE801ThsF4U5U3Lk0AgxuYjoxO7w4yNXmhGy
qvRREGcGWL4+OtTdwtrAF+GkNwDhYr2ZtXkAzwEZ7FwlHOG9TXa6xm/w7wq0VBIoxG162+pJ30DO
LXhdP3RsVU9KZ/Ay2BllDr+IzgdqoJczG64Vf3mIEHX1+Xmm/zwZq2bEFQBWz1pIZscKehB7rNZu
EDLI25lqyOhmkN9ZGzqKu0ZUpfXVd5a39tLnlnTbm/CdTlEv4Rqg1zIMHvZWlsdYX5SR26rnFWkh
D8NRS08BWPlzK5nizenoQly+5Dss69xwEszM4iD97U2iuK/qnbUW3cqncqWRRc7nRtSzC30NhMbI
gJDKy1cTD9WiSdMeBH3gCGxwSQtARj1mN4plPVo+LAnRscH19bUh0KTkU0X8oTTu4OmvqwZxkTUp
Wku6QQN9C9I7+SVYnWRn7nQFriDJfXLowds7s7Dk3fa3Uk2nGLwpyZLvd8mDP/UFKbxmmJJNOO4b
rbhZu3rSvo3ytEFhZZXtByU8Pw6RFdG99QmD29csgmj/8iIBzY41+i4CI/YZrtbr51dTdZo+uet1
fOMeK6qrtebtOLr3d88nrSsORPMtaEkLI4VhMcvtXsvmskJapwTESPigMJ5xweB9x2nKRvFNhomq
gHxmlxmb7uEW154mmzZQi+Xcy4LM1skxXKfgVitpvaRVkSRGuuzcXVEhTuGk+y3VD1oeWrLhoXYl
HWI1iU5mDJYfmbFM/QArJNJYRT6jyf4j5W2diK/6pIKSjNUUElcw2QgfBcb3/gqovFtfIkLkC6kl
VWlQh8RSlKbxxbQN+qbn4j/IMg8PbU9Wp/XrG+NqFKs4WaTbYbGD/rjxKNAaS0m49HcKQ4cu1HI2
O161nhW44EOn0KjCjfJnAwSRFHQohMeKVfE2v5u77aIn+HrtpAjLBL/YToCqdacjyY896+hWJwkz
IwOdWu8XQg5Go/K1lUqG7xGSs1R77O2TS78vngFxZP33XglASzdZjcfWA3OnF9q9BHj4ml7w4EFr
KPXmFOrgt0btRCvlSb5wDve2KQ4yq+ls5i3os2Hryj3q8yzzcJGjeZWqaoqVrNYfNT18bt+yIiiK
mJxCYyjrt0rO5ZbPn3tKqChgJgCaLVg/lxvaj8Ev8haWMYo8wQn4/YGDUDoyM9c0wwkxk3AF/ajK
uR1gp7JQKZWS1uCAN37YH1fiawzRl7a1dKs6Q16Y2H1gFML90viYZuwtMfVR/bg2NlaLZksKCY8a
+yVn93dCorjC/AA6pez+wQE2ahKVpSuiVqTFaeDtPLeL+t0jvIAPotWviXcmtjp3y/lsJs5Rnyzv
B4PJwS5OPKfgZMBB39NAA0Ed2DhvtBqREjGXV+X/8ExMP442D4vzZRszlJdKTG4vYGJNSnEeROnG
4K74wW6daDrhA7i6XQ/qQue533vnnvTM6ojPuYMdgewVgQ/5VTdajDXadnjCHI8XmU6ieywiHoaa
wDXSgHxOUsstlLNrRSgCkXgN2wGVaDQDEywOL4hzEdaKDYDhRN3shT9CHjGnL8+dpeNsY3ciYeiu
daUl+hxNmi/scXjMFx8ZkNcOF4gjTqzuBfbr49B53WXYA7ME0duAMu4hSKsg0nZPQYnpSFm1TjlW
6YuIdQCiP9uOUgRy+vIkPxZVkg+RW4Guggupdnf0XS9EsQ4PQ2czqSXkn545zOPm85W6PajYYBTQ
cySiHh0zBpg+BeCeDNI0C78k8FyT1+gbjB0jDUKKmmJ0RxvH1nmov83CZWukFmeEbxWtAtHij7UT
WHh391qVYAjnW4snVzlozFdsddN0mDXhFnE3lhS59BGW3UrZE5ZTEaiWYRVNDKR4WPkqu9P9HhiI
/ggKpqUVNEQCvGMb7u8v241ynYbRpOaiya57Rd+yanTcDgcKXppQup5wxNGauLfXmU+bFoxOogga
+TkHSU1B5B55zHHaV/dJA1PG6ilIvlFSICl7AmKZ4sUTidJE4TBg9Mb3VJFZj0X4/BVCzSyvz9jC
oFzPmCRQ9dZmdJkEUkUu+EIRgTWDhVSDfdL88D81AVjMN3lCnXjg0J3+e3JsVPRjCNTzn7jp8oMi
VBUHyxyH55Vq5CTsQE68j4BTHkTI/JolJtPCOhYb7iXaAK50stGsLfsKbV5UabOL3tTE/Z2IUwSu
bljVBwR2aYrLKa/zx1MFFkfIdhj2ldDqOJET3PHtTWnSsBi55Hg7tL/n/vsWdI/jAmVBjHKgWQWX
zEeFr4LI4zwIfrWJrcBl/MBcp9T8asip7neZRBrhqbcGHtJzk8UKSL/J1zANTAzwg30W3vV3LyTC
SPeXoOceckTTqI/WZHhSNdg560SmgaQb5M2bSWZyMscKgj5uMBcBjmxsvR/+V7d4DF2j8OqCquh4
jpQA+lepGjttpac6ToK8sUEGJjT+iCZ0QHWNIEGpVHarkH7NczyLmUJGwR2dfWSpc9RRjyH6/ECq
Bp+GPoozRAeTpiw4QCEcw3y1HSb8NYMYMe6MMqtEM3S6XTpmVrMOAP3L7iUs5A6Ocma5BPIb0Hqv
8bjsexVv0KlAz3cIQ4zyW7jc1j+vkidNnQIHAzDSOL+DxSI8ey6MVyLrEv/qlSYt1bp4lG0foTJ1
Aj4UVY2f7aI7hbPrmzUAWTG74URVhW2ep+kcn4RqZIoxx2am0HGcNAsCOQhCGoyTCXZltzufKnpz
fwbQ89KQwCQ7/C5m7u4v5BOzmL2z4MwMMMV7/ucBXcLzi6k7IeHqzFWOmNOWNHsGfwLil3KQxitb
VBiNnam0/nnTSMTPPSG39Uz2z6isu3D+82kQYJsse1lbNN3tTR6vLWcGcowXB4PGgBOxck6uEBkT
yPRmxpElyTKJlXdehx05jo6KGoOZtQZLzF8iXZtHiMBnBvOAj+0ed1KL9Ryx2nSbIRxtpbBY0gra
TJ4vF6748UG4kw7V7iorX/HEbA2id9Gj2tz/ZdOKT9UbK9XZHGjmhsn+PS7feEAtwhCe49ZRFDp4
tvUnbOKSkjGS5BMKIw3KLcnAZbWZ8aP3qhkSX3EwzDNXixkPmlaNh89ade+dMBE+4WOm13DAYkoj
HmfVFm1lY9DvBic27MM9HgkMYNiNtdq8++hIOE7s01msJTJrCbRQUFv/8myiAVYrDH4GMBCcWyDE
lL20nY/ABd8DMyU5a7TTiL02YSGvftzrL0oh6d0cR/fai5x+xlx/3kFGD2V5Z8A7R5JBN+dWIxKv
NTF2t/sti1+UtZEmO3G29X2B4zHGmPaRDkiV4XPNF2bfQlGU34MYDs9co6KQfgH3nbk65SVNajoH
3DdItjqJDMEARVm4RLQN/Z367s6SsCJCiZfdWcN3EvUQWFpbiG8B/LHb63hQ2B3VHm6K7ODDsNku
jhBsRlr0bihmiBfe2mSAZGtoGr1pBOox8yy8wI29JRUSFbXnjduXYw8HPlqqjEHMzEc3Ixb5RY/k
KNSvwpuDjGN62jilv1ARwx1TnSVze1tcBqnJQAA3RHkQgeWPjmI8cqwmbhQdMogmKbtxWZafk7AD
9Q0z+lbn4Xzf1bGQAlBJHp9fYlWthbN4UB21Bnv1GxZ6RvBY3TJ1kB7VnfXwXSbDaPKwHeS9cMea
DEvcy/LojrEO6yDAFeSCtCPY/Ls4mW5Ubq5/021SjZLpj6kmkD5uJ4SEq7GsmF4sBlzYrm5HF+LG
Xz9V6YNSkAvZHxn8JPAsSZLOB0zMtPf+tv8LHa0RAOiXLTB17S2FtDaPED8GRN0ZT1F0TLT4OFF5
zrZIUGl/W6bIjc+zSEU3D1atWWNvbkqBUkA6G/Q1uUzhTBC9np06bWAZA/4Z5wNW8psOOp8qLNz8
OaIqqlPl7pwW6mCq36abBJTYU3e3sjiSa+ZGMEESC5kCEMCaBjnCzpggnkY5w+qcIbpSx/SEbjTJ
1T+dhoV5YN3erGVTQJfUgFWwS0I8QOnfZAdyBcoiIa4FkAzCfLkSlyUeNHZnb2RQ3slSVDrInJmQ
nBDig4jQWheb2OGNuAkDLFINJG1TatytH4aruGIBAvNF/EUmVjCB1JYEjI3rGo5wYv+zen9iHR0r
r5CpcNUncY8DMbeOYkWtKbp/grdxlaPjiNDyKAOkHmFCVTC9H6RK03p5c40wSwPn7wnLPV92Qqtz
4iIc7Td3vS4Nt8OP7lspBRPtKYLekaKapEC/WJhnDFXrCadBUAe2kBaCUH39yoFfgISDYEtNTI/G
oDYN01SEuT+ICmeapbw+7UzjbqI0MTFyBy7A26l6Ehlbu5FUcBAnUD+Rq2jXGIX+UCphceqYEKKh
KoVny60A3lTPggHAxvs756F7RrsZVxrT6flx8MFlxtPQ9FTMD3fzHb8V7TD51OCpwRRI5IG6g8un
Y7UhkM9yIC4GKGqGrnvvri0m3GLeLxFJeNhgGW4KyhQUjDBfEef1qUbc8O/RSxJljODi9aHHHbY6
YWZjms8YL2YUJ05SDx02Yg679V/QYhD4dVwMdFpQXtzCVDLLbg4YnXchLWwEnFx8A6miz61yFU7S
8QK0/hSuXBkLMxVJJoqV07fdBIOMWr68b+yq3EmFYNegmBKAE/bjHZJZH/A1no3sNd5S6cQBxK0q
oP9cGM6ecri/oc4uJIlaAnXCDfeCEcBdqpXIA77HshpnkAyDt/Z+RWA2pCzNoBfLmilVoGt7fSVE
I9Dn8qv7urdGIo4OepteA3FHdST3sXLtmW1DSteVMU5rz6iDxZzHxwraqelBW+XdX3aGDDt5ACST
WSDvzqADrAMLNXbHMBjNR/QhAzrDw6YKDFQH7Ro5CoQs4SMrEwgW3on/9eGvNnTslHgAI4+TAJkS
7Q/XGhGTSR+zTVIolJul+fFRpIdnBjhAQ4Pue7Mz4pZaP+LEXFUpl+u4KByeqbeyTxW+8ZgsnLKn
FMHUIKsBLAFf9bMHnuBvBMWPvHLe1/FJHc4gvUbDV7JQ2KU02Rn0VjpiHvu2oAz8muR5mvPfIv0E
d7Cr/G0YqM5CDkWvoSebMOqlXxvX5cvbgRZZ51uGrewxV9V2dfswDF7h0/3m5aytJdMcgapvKZJ9
ku3FKWBKq+VwL3D7ydojWAuRZ5qOscfS0vL+eOZOvu59hozaSxy69VXtxPZ2cRF1uXjx+W3BXQWj
MgpbnZ2nf7iAaU2f5K2zsW9K2uU3g1YczGFbJ/5eo+WAU1F4ckbSXmVw5z2A9PkuDFtKQUFAVjGX
ADsSERhSvoySnTJqYtjuZ+i1G9u7u/f6syQQaOIft3w+qFrShvqSkRmUcyeYdcauBqIB2Hb9uu06
Mp/f3wvkd4cSGFNyugcexhh9NQ9JARB8L3egW24jKnq5c0RWxOv9y36cP0AFSEIsMXZ+L5CnNCJm
Tj+H8COy+iBlY6bam5XIHTISCp4yXDGitz0MIVpllHcd2BD4on2aQOpJMJ/f1OEfenmIxtSNpd5B
lEDE2sa48Ydo7CoX+4NvGkv7C6Nlu9VdoXO2RqQQ1z+mtIc1SKfFo7CiPdCLj7GCTWCuZZT9yyeJ
Y5BU1C6AFeIe2wgajWQpbgOQ2EN3N2RoqCM5I3QsvM/jkMhZhCY+hHi4E3ZjNxLR5N16YVfggd1x
q8rx7dew+98EZLOYbtKMZzWrlRQELldchwe26i0Dvqja+WecFM8P105MwYjLaYv51zkvNSgC1ZcW
PmtO56nArtW7u5Kbkznozx5XqWAZvB1PIz2JzQrsrbl3FiWgwynf03mRQ/f83ItmCrN3aYT5xsdv
W5tLNmZHzUaF1aetfD/XCLRB4qpPoVtEaY0B6vMeKGrfxuLgv7ItZiyZTRR56L0uGi3kaDSRjrsQ
a+wQnsSHAQc5JHxXHQzburd1lwMmAm0snbAJFuXsPVGzUvj1Q9E7tms2bvo4QGCQe3I3eNRBRII6
QdEORwoK2qDnsNWn4dvxe04ogCf3um2ZA3Br6AxQYSd3xjTWl9sAADEZBj9ecATTppzm+rBPE/y/
lhvhIWTbNt9V7zhochmPE3xhjyKAgtVBuNX/j483cyN6fNkJdkyVB8Y+vIv/G3GQC3ArfHxXaQU/
5q/9DzzjrpHOe981hb++dnjPSkRV5ujsGQrkmr578dgH2Mn4dXnefWj5tX9Wx2eKAYQ6hmz0uZag
95JmZmKI1YmJSPnfOkLtC1GzW9l2Q2YJ8iHNzKDMuFkm8ilpburygWZpMcQe1co4sDQfMi/7odiR
iI3nSeZlZTJC7/7eJpJkluwlvWNud8vwwFEPhrVPaNOUvz1jE67EaTKtIBvDoNdKulxUsgtiy/9p
36K4bTYMXQQI1KxAB2qXvTxNA1K8ZLhH+1EZxGSTxa6Gi8uZtNunMx8cwXUXW+f7xytRRfF0LwQT
BtaTEZh9hS9F53wZbwkc2hPp68aQESaPy7Ir+k4pfXYgU++5AoxqftlILQZhrYiD5ZhsSbguM2OH
NcFTay1BPKv49gJXXF1xk3XoBb4aq2jT0qdYhpyYS/MT6UkEFMAqF7No70nEi6r4Iuekg3Fy6zaj
baMRUqoObcQj9E4eZsHe/cYPzha+ZDiWAKtZcm9KgWvY2KxT7mRLJR/46n4Ur3tWNCu6RnBhkFs0
5Q+qmq8okDHmxTUbI2f6o/ycJzHi2oGonP0smT+40KrH8WrkH5ABZ9yRiqLEuAjHk7QCaGkn72+P
0r5pPi+vmGP/OHRmO9/pQ/N8CGMkbtjhd7FXMk2yPPrkVvect5cQmPeyxrYb90+1VbO+c9cR5ije
8cJg7pde77UIPyI5khriBFiKhyTN8LfzNbWeQSzM531wLdbgXgGBIZ82Zva+9S0l+1suIryUokT1
FXHeuYg02U0xlSmw+fh5RRqb0e7YQM3t7QtDsfYfJT7lGm6OC96F6RZinnljHRtqvan5xTYRhEIV
x/ncOjTReqmMZuSuyHVaaJV5/sFvQ5L7u0odcNTuRprUI+24CqCA7WNKSLqnoR+pwR8Osx/g1O8x
p1AnmQ5rpIfS13il6lny2tIT/30gPeR3RxMm7Q/H4vuaVdFw4Y7ZC9AXb01FhM/2kYyg0ta+laZx
M+Ej9DccpBYn47n1UmiS/GBPYoDBord9BCccJxYDBhFu8vtUJmTvUtFiVcyciQVw/sj30SSnh6Nt
kf5RUDwZ5S2ZuiQLke7HrPnw4dbhSNkLaXBsPa4UZffuxusZicb5NVJZ3wSlsGJ078lJtj/6x1zr
0YkHatdEuPkYT/T8PoVEsV4AwwQAQu3mxUfRw5UnnzZuXi9/ed5LsPf21VkijB8tBFnst/mQcOXk
If/bhXamjzoldOjfTYGVNGAHDE7Ij7/q0C2SglIy4AetYjFzOk0QEQzNqqK2pWKHH9r63WJ9YsqY
fbMSIdIQ9wuXLPYc1Uzo32lWTVAj5InS7Nd3XTFVl0xBRc2R1TiDkDQqPNQ3QxxMPlfh0V/S4PBc
s/6iCemzMfNN8MqK1561eR8fLB0324wexaFeVT9zg00yNR/CT1e9IzDW3fIdH0PvOr2DMM1tAfZ+
FidRjhNV1KyCbbPkiZhOh79yThgD+OA6upJZOvyulxbNSTDZwVUqISnkMBQl1Bdwnr8oGnn532Qm
PBrGKSnR6AE+EBTeNLbXbF67R002QCsLJc4eTF2pHuvJI50iGlkHj/LJlVWeHmRz49jHKb19qlCf
JMAc00crux/fKkwRYd0sIbPKU+wJ0klkfaE6kkCpwU7OO0/3nirPrplvR/b/n/bjPLBu2DBoCJCz
hrxh2t0kCHUxZ5K9M7mq/hUPWnT1JZIVhtP3r6z8ADPp/L8vd2IddJYJMh1FfTSmVP7ZlCCBLBOg
xk8EybZM5Ybkl5bwNjIdxopdzC+voOBee0afOJVMYfNHLNneP/YXCI60DHRJlJF66P50hXYFme+f
U3Zl3aeflfPm5jyUh+/2Nifx7mtN2AgjnzlmkuYxp8NnlON058bJEW2HIZPFlxOqsCPCuSIw50eO
TMR0sG03Ifd4DV5MkXeJ5Di5A1HOOwEhQLAh20Z4XevTtNKq+FAuB1Uh23Rqc8NV1GOGC4CioGh8
KZeIXT0StUmKGfRgZsijNp6i3luXp6Nq12KiZGCyN2koVCxxaPHq5zYIEl/5wkYbBpnqFj43FdAn
k6mSlE44A/eWbLKuXuhBIkqwaY9B3f9yutSzqZkE2f6gUMDy5EmuLeNCgY+pn7cH1VqWh0upIyrQ
41I1iBCXqUqVrFK4n6K9h+qkHYwFapnBxe/a446JmIIl87bhLa5SX21TeSW3haLpIe6gLRi6/ar6
AQlfjqGSPXeSU5kskCQfCeU9zviTKStRV3hE8MmfdGEvB900x37cRY/HHodk3BbHX5ZXiLwgZYMd
kbZ1jMcjVncYCIswDf3TnznA2BOwki+JEJddApxmyY0CkbVjqMiNSbtuT36gUZTlxq1hygrplDL/
2EJ1MK2DyId/o791LffzocJSb6aH40okAcgVUgHS8ILfjIm4FN0SRv/LjU9m+OXz74WanbY8OueO
cFULT+cPJr4i4WoqypqF7oFoiFFPFzHVNxau9R2jGIDqIEEkRHm64HNZQEb4Gj1Yi34Eq1etsylZ
xdiSxfgUaE6jNUGipz38Ycf0/b+c2Fyw+NDNbnIsQfh2TwVH8iNxVsDnY+OKgIsM5E+jY8SpZ/8A
yucADCksEYmqxisOLK2qaN8LRQtAOckHcvYcDEIGtQNzKgZ+2gLr4aYs0aRmML/YW3hT3qHH285b
GHEpVuRZp6VQKGPGt8+3k6iWILfYN4O4n0PpB5arnyHd2wZrONKm9Fc0OvtGTz4mFSbQFYQMMPdQ
Kt2k8BOxM60+vLrcm4HFgaN5F6/engxv9cGUWG3YF6vTdxog0GsmysAM5vlF1/bSjm3GhhEyLcxW
H26KkymyGb8EZhptz3pcsbmvLR7sIhOjozmnAv+XmyC7Fr4dplI6wbkoQlbkXxxsSqwMT5mAxzuO
GiRppcO31D7ITBRpodANCfp97xPrdQYrBx2u5Xqfji6uJkPUtnrHs04vYkO8tqYug+AcCn+tYbvx
aWkYuP7iNSeCr1EPy2vS+kvsDYifmHE7oLfrCRoPuy98PoCr1FcUfKmn6OJvgEk1YhWztlu+3uYH
UjpeyWvNpFHwgC7r17uwZvwdUqRidKJrXImuNTB6fDEgvHQoDw4N6LhL7sy4HXDs5ejcIdFB2E8u
jdW6oVMN52S64iWINKRn1fOd/vZcZaA4mZ7ZRdXGGo4EDc1PqMbnJhJdLIBf82MByryg29nifBHE
SSpKdF+jJImQ9We1HI1Dn0kbZ0PEPJoHaxAU1xyeBYaNAlIddMZiJ+KLHyIMo8cMHgIs2L4q/dRD
kGLitscgQqN56iQPDjHWa9zK1V6GNynHebEXI9vX2DdQm0AUC79bmpZgPx61ZV4V1lhuNU28Un0X
jxNs9UXQAueQx5EZeCAlCvKVqpfkAor7MNc7FmPXRBuASjBM660dEzVIub9aFixxl/vQouUtRt5y
l5MrEiJv2H9QvQSwuGSCehP8mHWCYk0CVRS17W+VYipZ7feHyZGZNCQzB0dTMePEzu9RYtDHJKhB
lLVJBle/VoDV9oe1ov9B/xi9sN9L5Vj3M1atK0ErA0ML/jdjVqMPsnFUMGPT1ahxPuQ8m8w5vtKX
8awp1EVbovq8N3qr5p8yy968wBNl702ZGrcCiaHeB1Azsg/Ozn2o9DP5SkgFKvd7IZX6kNy0dY3c
1gleioUyqmW7f5GX47DYKZ8gPqKaslQJ293bCbkdoUTOUTdQ+XK7vkqH3oqgUNpYl3oJIBHq4ULt
SSOYj6BLP2+oQSvJUKxb1yeaCto6YbYEy9Vq2vIMJJnD4KJu1RtpxBPPmVnERLtYoTSsegRNpx5U
8xrN76aBlYXL1Ok5QURdbJ8E0aaN1eqVhPl4Ue3JWJmP5cggK1br1+UqrD8hqEBqGG8CWGGjglqH
wh7LLnWtTumWDftV1stwZ7QO46elR4A7jUOvfQQLcluL7f45TSHghG7QKajLEL5M83Kcdip62C64
3J86ABlD3DFZGH+puCtEHtnK26UtaKiMcKOIsYB4RzO6Xok+wuR8lJR2AEtNcqjY3BT633kSqPjr
TdlwTI4go6mykOEJsnAPd3u/c8tKzBXbuQ+CKs7KvuqtNmID00cvEAgEAteHXARggQE0Nnu+l9+4
D9B4gO98Ouzp1wSDSKd2SU+GX1eork9ECw2rkuk6cMHDDWFGMvyMe/rjoCBDgQKqGIl9isxg1htS
Ku/lUUctHPT2mkS0Gza5b0Z5vonFkR7eD62ZpDlItZ9fJtU3K0b6Mr/XVzito2f0EcpoWUYZWByV
1wQYzZ30tWxf89ZCxEalYe6F41OMZTYZSg29kR4+YIaCJkAS6muvpb3Pl1ZLR31MHlcejd4IyfIb
SNsCPB5yNwWbl8GClESNxuHEyPhn5mRoookiNU0YwhOhE1EKGPRe0GMJkcS1XZgq5emTvfcdRBd8
ZLjJ9AabP6bLkV0bHlY92Ut9gv+OOKAfmWUHepss3ZVu8t0LN4fArewGSB5zY7yKmCEU0gu1XaJL
KDW4kPhlXFGA2xVL6ra+3Dr6ZX5KSD6QPt9lkajrNB+D2fuSvkUCcP5m0Xdan2gQ0R0Gv7DMdVN4
1pg/iNTVgtoaudEyf8ZgcyzTz2ZU95WD0XALd9++2O4IVJYy0iFi3wRI5TV6CMQwWruHRqHmR2A5
V6qUk2oLz3GvYy3zczqH3+1febvk3+CdxbpPy6dtGsnv0g6RZNvULm4MWbldZhE9dKyeNMWhWPME
p0aiJ6QbvjYuZS0SNNe5Ujhrdq4eqTO1GAItMUEr8qsdxlPYe2/UT3xvIo7xTTo0/O537i2QwPDd
i5DVgffOErqyeOJYUbUijm16JS7Jza+ASvduMjww5erEE8LtrTa3yvMqk9846oQh+hWqYoYlLzWG
uow/q87dp4ru69CcYV/IJHXw5mhrL0TMIJn7lWZKeXk5KccvCXr6+6Pzr9G8Ui5P7WlQog3ZJrd7
V/9NN/wX9DdPraZKmkShrFr3iXi2SuLM0U8fs361dEBKDw+NCvXbhvcavnPl9amQAdLny0Hfa2l9
Sy8Y24k7cWz9aDhI1XhW+X5ApmCi689Q4B980sYNShH7mefGdR5ylL5v577OJeLWcu2hJOuUISuj
J7KxRv2Vs1z45ltQ44spX/eEEao+bc23XnTQycZ9k7AHjK5G6+r57XA8vkEa6GlxkIrMugmVLEKe
xgop64EVXYjz8Oys1JV+MkMiC3vTGrguFSJSJR8x1oO+G7gkQsEAlr9I5UNvVNLUkjOlNVNyVfCV
I/8GJfLVpBL7IvOKUMfnoBog11LjpQs0tIRphYdpty+IxKqSMejqgn0gS1NxL/Pu1adTh9FEWtlJ
c6s7jxpMmZ7EmOe+WvVHNVFww4eHJE1Kp8UQsR6NVDCiaGEkuVkzOLxyQ2WGQ4vNO8UFDqpFzr1i
jB10zdJIfLU7WENKAIbxNFdw/cV4wLQrXUfyRuJbmjqwLd/QqQx+wyuNggYdOJlY9CSQe8hRNm1m
qvpT3iG+dmhajTsM6jRUEfi5oaM63h7lx575HxWWGxAuKCYJItCt+dKDK4bWyXnxyHmMyphDerYS
lF2U6GECnlaz8xqFAEO7aFb/aq+GLG32v0pOZDau6/HyS59xrSbRtUmPGF9n02uu14YS+C1YU4E5
FW+pQWLPrTqggzFcFSpk5GhJqF98lzFmOtGvnK/ponjOSOpZPtaDWnZZKpnd5MbOcaOK/DNSYds7
rbJmZwHaDcOiPbVbAyQiBS3xNS9LILWHkyxC77e//pDpV1aKvF8PXeYjBbcBOGZFkXVenNtWYJ1I
4PuvCqdYz+2gWaIp9xduoCIqSqX4vntT+SJ+SIeVlbkYRfAmIuos+kKCD22W5PdwoL/Fss1x/4Xf
JZQFYmB6QNrCdWpSG63G8a502dm8YC86NYu2SBp/2o/PfjVI15o95gae+CMtJ1SRIhDuuA6DU86A
fb8SMbKZzLoiCilro9tzk9Ly09CzRLfhA/p15sGpXXdK/sTnAGcEKDduy9IwearwjHGGJWqfU/m3
j7jUKmuPdIses5UmwWPqEUIip6E5LjJUy2YVUa1mK5WEe7llh2ik+G48QyU6GRtmZg5t2a31nKvY
ZLg9uR16N6JEwlTEhLL2H4YmJndTnEmFZ9e55Sp+ZvYAMNoHzcmk6/89gnUCdSscsbeofzCvUJ24
h+VJFDny1OVlKwSd6vyopw6M3ZY0TJorl4MiIDnOXMQ2gyjpzIM5oA4veM5eHv74D6NUwepcH3/M
jL0/XB82yNftlPRCPycDES1BG5rWhmshOISqMzwyqgqfH+7uDxzskx9dFZ2B6yW06HlnjsftqBf5
4DvgGeyJOQslixdPEkEddM/YoJZsSEum0gT0vHvZAlxdV8HJmczElWJx3OykakBiPo/p9K4JJ2lJ
H+Zh5isUXZg0vik0ce8+GC7GAQWjwdjOBgZmGv1n40KDV9gdMyZo+wnveYV+onzi+/mShG+jmuKB
VgAoTLnwZ78oCzc4wdawQ8ZrBBJ64PwUvvAF5Zs2S4/AJPabCy0uru7ZYL0KKQvo9/MBOrztzhy7
Vcabc2DKXi3rZzwGa5oEampS15YtKO7m7Vd5GCuVUc8l/Wy1eCv1UhXgEzjzvjVbAh1uKX2Vrrb1
iXarM9ZfmS3k9ubFF/2Ak/kiUDJIwj/n2XeOjNspsW/qkXKAmMeJldEI9HT36C0mZLnKlq1NoBvf
+DNFCEZvscoiCCmZNMXkrTBYXCe63148npk/wBgph0MG7DmQJ3/kZwcyCP/uS9ynLIjHGvd1ue0o
nFaFxK1aot9IgBdgV00HcSpJJql+8enJKjS36g3DcSKrJoxjsqsMRH82OnnDk3SZHqgkCcYAXk4K
kf3RPYQ5/v/uy0zY2gT33x1y/cofzjgnMqXFoMnCFsQAMuxnJOYcFqC4X3eQxb38/1zsbasxRVxU
WuZkOCH/rxLTYn3ncEf9nZL4Di4rYs3llRSPKQEYFDJKC+FDxUq5PRyTF5OzS/sIvTA7UwbZAHX2
dCjAljoHpfgBY3IZ+ipvVju+9lkPjZ0kRwDzZhmKsfyMzsRe0n40frh7v3u8AEEZTPVhZbVYJa/t
w2p3Hct9kc22/C/9oX/iPmT+hGnoPoAvQ6CaVSuXW7cnFlyqY4Gd8mDvb4lDrDOR/uSC8qrgI3V5
7b9x9ui0WM3wmQ9qpoETCP7/N20H6tU7m0l8HuMVm/YrBFuwndvn/c0SLLlVGiCJAAJ73fTUH/k5
CMxTcbIpVuxD6XvyCzEaIHiQtYNzB2xFAfUAhXQ96G7X9mD7gfOkU1l46gjo+A0gFMKAeVWYYo5c
1KZAm+nqsBZ6oieHcu+IjFn8n5GCy6eQZRbHpVR8HnDShCNCZ/blJpuGpIk8YSIvePoI19VZCzaq
VChBicAVLwFET2esBk1as41mHOCDnkTmYIBuy2rgkHy9S67DLuyBbQvuDSTZ84PfYRdEIlFggfFZ
bFSDD3NGfAf2OItl0yFs9GgX4trdrFnSMVFUNRQzt+mmnudzgjBvHpjmQLnO9P71Ei+dPa6thehF
QTiVh4/I8cRJl5CM0okA/UPJw3ic61MWvuOu/1KR4elNlJJK2uZ1u49+hx3X4Sbeewyo4YT4SjJM
aew6O8VVvkmk8gevCaSvGENcLJbI1/LQg7NghZ6KETm4LNC7snxN1DfsRt4xXk1U5t/us/qK6E+c
ZLsJJYLTLuEuaDwnXgcYxU8CPZwyRtB1cMW5vfUt8gwrPoBBoqKqqya+btsp0DTHyQuAJzp5+Mbq
G8vVwFRskV7idfsqLNJ/pDb2OXxVmWLFNmAZYP2MBNariOY1wvJZIa/etqq4zjVUPmZdZvbTEuxT
NO47BOR4sQwS6W93Yq1Nw73bTmYfeRo/DIcrPQfvqR6V8W39V7BMDV2aZvsE+TfNn7KvsUmIEX9W
YoIW/zS8P6K0aCvjcBJ8xneGoE1oFhQxbMEkxC70IRKvSXnSXsXyQI5fBHhFb26tMd9tY4QLHDwn
LVToqeH0LcI3vtKAAKOVX5A69+WdydU03JILqCgux0GpIUVBefODCAykbeFutf1eLwrr8WWKOAcN
tX6dyIXtTvVONcu7cKT4Yfx+Zax/Pv/ksKZnoZVUogG+yIfVAjw1DopN41YWwX6nME41Hm5TUQYU
/q+7SMNiFjxnVfM/+XPtQMBc/pbC/6E6JhDjXlTnAFMoHq8LgAdAy6IMpIFaxDGAI3Dd0zJH0g3r
sC8yzfKM/ifLWSutnMgp3mJsMqIQmc4SqSaPBGc4wdzzwgI2nHfDDhwdIK3yjmkAITBqvn5NRhBY
gLhul2HDlIYJCzbHeUrNzShNHL4HZrqyikhs03Z9RUG3pr9G/T1A+gRF6tjxMnMZ10S7PmMPDs1A
OtgpiGreug8H42NIjuNfRBwS1qv7EmBcCj+Zrx6iIeMhJgejb+c7raEOEzgvYshu0BSWL/iOB8tY
fqRYUQCJCCTPCxoDD3axXogjjn+erqQbAOLHoBB+6l6xNWs6gi4CHRpMvfFt+/tf243GnfDjv1Z1
Bsg9Q48M1ggGYjLcZNvsL6kygJTxfNIHcBOACr1Cn8ybNx0nvhhTISo2BATiytciUjtTB6B/Ix2/
INrtlScLgopZ1yw24A+R2OfhWzGVa6oqJ2MWOE7qFx+/4Krd7T4vCrBBTdZOQmti2U+EQH/+awfr
Lun0Z4hzVfeHb9Opfd53dBF2QAVTQs/X1qMxyowKSGAkJs824wQTsqwAX8dBCA+AECdcPU1BiohC
6QPp+MzSKBW/VYli5OltpbrbFhMe+RWloWPaLHW81a0mHTMqdR1T71JuStS5wGQr8ql3OY8ENlOe
iLXpvSpcPZccCH/Ie1vC8bbFtWWzfodTCXcBeLle+aknWXErKQPEuSfzlmUouA2OGlpoqPXSeCP3
dRXu+aI4jcMDZfOPsvtp87F7fbqlbXYr8YZytjwlx2Mlta2GqEs0llmuLQYLtBD6NIr6Xzvrdizc
Xo9vmnxcXkjA4bZSud8FSazNrK3VlYH19/0dBE9AM7XaP9UTm4WOOnDyGaov6/8dxP79GrS2EYhM
09aPHjIuk3g41sR+5bkqorWkYioJZeNIHpb+Rnpx8bmtyNm8QfgmvIcCyeJCvcpNxNXhsbI4zX6M
CwH5r2vMa6NmrdWmA6cKSCKUC3tok5bk1r+1MFyVxlpwRTg+n/xA8gQ20aQD9GfXlQ+7Ec3ziVnB
aW83+Pfz/7+lR/kOwdubYa4i5Zg+u/rTOgng+iFGjq0dsRFeEJhm2c/syn+cwImiLMdeDw1LxDUq
HHk6LAT/QnVDSHGQDWyJr6CBxWbDEq/3xX95qqDzLsv9BIDT8rlwUVqnwGfeOeXWNfEMVXRx7hI4
Cj0nEw25GZdDnk1PlwEy2pPKH3QPOpEW/zQUQndwtMh33qLfU4gy1HSNQL53AvwJ2+B16BVrXacN
3kxdO7Z6gAclo2oMnf1r1Rhx4BnVfB2pORzLtqTPwvU/lS6Ra2EZKpaF6NyURW2yAtB84isFfda0
BSR7RcHn2rpgC9yrDPouO023pnDs8c72yOiDxe5/flE8qTCwKTjjsoQCkdQ/e0LRVlzdlYfdSqxd
wwYgZ7EpxpnMLWH5OPbNhONVspQ/ZzD3NBkKhh3wKMZu4CpEPzH+O5tr8exkUoz9w7OiEorueeE7
VTIT2JlefggOX+TieCpbvOtw1/gu3f+r9TT7i9hg4kCuhls84Kkf5nXqdT5eo5HzgsnOgMlnt5p+
+DWxHIiX+xqjpWp3DJyHE6X8Fs0E0UuYNY+cOuigLmpy11nmrnomU06VQbcmlaRVpLklCtV2Ods7
Du2QMy4Im8uKhPm23HLRsHRn8aupSieYPaz+36cOVfoKkHP22VuFcYnH0sXlhDrxssuy6vpWjiGL
mBti9Tay7YyAfktbd0XRiKEDOLfQHaeESYznDIpVXwlbxeGKSyzIe4AA/W8YSb73KNAOhX4RPYyy
eRh8miO/BPaBnRjfi4qAMDYQHNnDsS3BuY7jtf0H7Mxuki05XbssZtmDrv2Cymuwif7m4QQNG0y/
6zNckmfwY0LoAd9+NZB8RJhmGr5gd42/lwi42/mO5dP+/i7msKBysCKAV2gCbIfdVFq9B8t8Afnn
nX2o0slLR1jBFGemxDkv4/HXvu53boPuG/SMJHJ2bs5iBJTtP8Jw/waNUjNLIpsifP1E4oJpsZDN
XQdCJzZ8yQaHDf+oFrhzL0IENDW9MGEJNLm4KZDkZqPxGdUAytuozSCvbyvUZ7+sfDNSdbNzH3Ha
3xOKrb+sS7t3ILM7QZN0Uu9cN25GPtxIzGfDEzEW++dp6zTb9Kg4U2FEJo7SMqTL+jIevIoMNsv4
7q4fY8ZcZcHE0QzfR2wQUeR7YfQ3iMvq9gj7fTjqHQCFzgVfyj9lbyk+R+dxfKBtF2SNSrrtr4Jm
bqt6AEP5c9XXLZxoyQ57S3JnDLnFrnT8+OTxO/l1hiKnnPoNJELTgTwbjHiNbp/WaZxP9oiJArOr
i6FdZIBynpnp/RsOcI3YIXHevWJocEwuGPB2jEITdlA2vSKAemfXCllRL3PpwMjvvn7QgnauOTAC
Dtn4riHvJZJ/sDYLvKj27FbQSpVZbddjzQ+CaTIou2AjXmbfwD5UZSnu3SsHUuLgDJAg3goKNHfb
HxQZBVIvFHg9XEES8Phh4ZqNHLwQqNnZQBc76vt9I5dErTRbz5THGBbYbMwmjo6yOxxmm7VcCUrP
fxOk0lJ+ms826igd9XVrSiwUZCDGeBQxfiLAQqh2QgHpYQXEX13uyMh2PEorClP8EnRL1tzk9Fnn
0FB6BDqdf94Eifs9+QhThlWgl1vGUvkL5eoQcq8Gkd0JfosZLAuILbEHkLStbdEU5NhvylrGmqy8
TxXmyEMQW5IgtB9jRaNbXGo6yAijHJ+5FW7QtikmoeIUh1qqXq3lIEScIHVb3rm1vkmd/yF5fVgJ
yRMTW51J1vdqQ5WDVOJDMD+4yqyFdOyQbCKMNU5I+6MUTNM7iidjd4ltZ6lbB1fa8fOFu+AtzAND
oXpfMJOcAT2+dj0d35Dd9HP1fYEz0PQF1Ow0lpq22E1cYZ6UxsSCL55jgkw+xfjn2ac0HvBd4Tsn
58epIReaToWMhoLUut4NXtSuCv7vzZqhpWYFapS1BYDyijwWrIsQ3dXrCm06pfl3rTjhPu0A18bk
U/n6GKASC+zndjhr3wSnwBjkMOyZTdkiZ/HiUKbCbxypmAAZwLbR3skUUyeZRhhOTeSVM/nwP1sA
xH82bdTj/GnfQyUBfEc5SfCBzw9iSOleCrg44Clc01+LBygspkxFQxHm5yRNA4pMGbVlB6aPxick
WEzt7ma5qgLeZXJg0kPD+/RuWhUfIiCrbc7XsUvm9Vq5QxiXtsZwKGxFO/Os0EV6oadebEIQqtVy
8waeviHI9Cwbph82+Gh/MprUIPg+hh+aHNuqQwaaQlXvfwKAuMQRqhsfPMkHeR0P3MTsC8ShEOUy
X65M4fSGrSzoP//4X3oc8AmyciCTjbDHTTJcqr1G77UKqIJcInhAJNn8Fs95ii1x0PH67xuQeI88
z0F+Gat6UYaByn4IWgSNN+dDUNkTHemm7GlP0iVZKg8BRD/eJAE0Sryamz11tsjSw+Li8MmR9N3N
X/r7RfV7RS0ZXXH5O+CfofNVYezfXSoH4zr1wegPA0LVO6kNF/mCIWhnqUbb8cUD/aylM6ROmSM0
dzdsdrBpapR8gB/c+O/xtDvO3yze3SDs1ExmjvgbRFaL5zxx+WLtSNmW6Chj0fpxBzBcujpuckh4
w1RgPvpajVMddlRZPTV0kKmpVDCMTfI1Ac2qGAEqk1/9A/pBMWwSwqWQB/l80ZsKsHbvv81/i3QH
h9rNem5UtV3BRYMycVL0IijJvfYoepNyYOC22E5tHeiRhp0NCgfMvpCrroPPKHi789XTpIbBYXho
3e0Y4U5kxEy03O4shi5bjnAUicXH5zPpaW0ualsXEvxRKpU+UQPrjloz1G9Oj8/6m7MBXMqkoFbf
Zs4fSVWHncsMkr/NxjHJVuR2IT315aEeLzxrZDMOlcpgFt43+1yc9jzITW3M1mWHEcozGxxByT6C
JuPVs+z21feHfnOt88vJ/eOto7ej800VogrQxrWVhK8N6iJsMRsFpkPVBkY+17SBh9pkayGtiS4W
rStcPZY1fixgDPJnkONW4ZLV8vwLKWEJ4tH37Y/xREIa1NCcb/hFuctOicTxwVr7sM5iz0kGpkQf
sAvUPeYiGqfc+l/y2GRKrLld3JIN14v6Yp/Zt6hO6UzCxIq7dbII5sNwmEIa3pqD6bQuklru2Xx+
lsLONLj2X6RiG4LplqKb0i0JqCUEwEGhCTMCWi5Znsq5jdtu+uTgX2dZwiL1bHcerMXKfNCb1cDI
bq/NsThPOT6RKNLfqgynkXHzCWi6Hhjb1OwYbYxLXCdoyClmJf6Ry7M7qa7BEXS/yDicdTXiLmSQ
z9QZ0WZVHrbR0emNbjwafcxRI85PeR7ZXx7NAzhhPlqFdgDBM+SD/2caUBsByoCOWliZuJb46mWM
5Zi30vd4XFWeVAg3ORElQY6t8swc6vQ5zKCTW3XimABUJrOtoPOB0EqU6ub45HtJldCB509cE+C5
V1XvXdg6Y4RBdzfSRGEsYG521NjHdlNyuhnGTG5kcp3+X7uAQXQSSc9tVOfIxcCJWMdHGbGOnM1i
SbrsgqJcz+BEh6R/h8S/hA71NEMiJvsbBJO/3rG1a854+JcfvleXtN47DXAJ3dGOAFxlWMKr01G+
P1NOCjLXAJSBCTQV91+wsl65hxei+fs1yaYT4ge8rvtFlQ2L0EcjPKfUIhX6AiuUKEV5z0m0t0xU
2GWty4Jmk2RBfeTGX1ps52mwTxzb41qONl9axHY/y7T6aw8ZiW8gKQbB43TOJdWbbDItM/lCW3C0
hrqQ/kdzADrkUNRGHnZUMej8I70vBmwXYmrZW2grau7FqzkGd7rwghQKw4RIOepIBrRlZo69LPUW
fr4BpRPKYnEZmNCkfqQ65jp5loxv+nN9dl/6Wp5+qzNZUKI+QxRIc1saKKWKKgAs9gYa0HtMQgOl
9Y2ZgdXCBvkS+NimcjPjTwrGAE1PUec5PELmk/yv1nnegb7bz5s4D1LFa0gbv6U8HD/HqOYpzKRJ
0+0AeWXymJ4VBpMfrwVOAnuGL4gGYjPAPMgqEPacSCfEb4aDshs3Wp32zv7CpkXfPVSMg2aKV6ia
+ZataBWjw694WWsQW42PYbukXzu5L9dvOXzCeg91WJsuvVAA1nKQRzLJxu0BfLR4aVSUGT/ox9Mr
q6PNZmRrY92YqDXP5sxv/nqvBinvB88uxqEsRwgZIp8vpcN+yUanEtxgI0z3iVMr2tPRv3/RlTDB
Xo7++8ghs5tWp3eQV0K5jhRvOkBMUohzfO7zmob7HTKJae2sqcZkSWDvKcOuqHdoL0i3wJQVck6s
hFr+7LDnUdklW6VXmQ8FHJDPUZfVZxf7POmoVBOU3qM97t4n9zvbABgGynw+xdHXXmAC94DBZObO
ZGP2VfW+62oCwbZcBvHj5yAR07hOs06FDxS3M0id2jTm897OAXr3aS9DNbf0WIp5YWZdbpMBjWhw
IRWyfxS5fV7uHmPCqeluHdZjNzz7zr840CPLjf/dvCA20LXXlqUNsTwKRZFVBilv2zNaoUj1mVT5
KDR6JcE7LqilHJnokI2ELg5iDsj15PajjMDSY7JA+yJbP736qnE0I2FvY/N+WD19/FDuDMOTvKgh
qJc7RWrAfKVMY9BF9U0XsVQmN6tXz1hDS13qYB3Yv59z9Qv94scfJQhmI2W3qyT3oloyPSqMVV6+
GPhZISAlNhZChTufrVvdURvb8mpfQp8TMu1y4CsI9UtZg0OMNTAwVCOSiUdI1LjWOBTw8ZFZXYIO
j28fzgKTPQFFsJ2RtedrfjBewuAveF4aUtLz3fEe5P2mm337d0bgru4Mhm2zw8oHgMcuWNFaZZZn
qAWeHImvec7ZsdY9GFhmJge+eHiaUM0K9AO/IXJ+sJit+CcNBvEuPtvJMAk3envkKAsQ8HXP72ca
FfOSNJ0eeDFFzStAmyxprrXmty5NgW5kvzPAfXAyDuUz4Bk6vQImguFlMcJ8Aeg+KKsxOeB1Hbh8
FqpBlstqOVyAdYcIS/TnwmvP/8sRm1moFmJFpJPtS4u6Bq4QFN5GmaCJF3WPxrF4DKG+VBFtsGGJ
i5u61xVbLqNA5HtIVzgrGKRvaNvPPXD9tDe4qbr5qH5hjUj/lb/llaFH1sxFPqygQuw42HbfQr3M
D+3RMkefmpjTPjuLcG/bTE8Hkf2cKW8bcxTf7Ue2L+eGA6BjDwi+JetEcpsQ4edS6HSBYafRtMWq
CDUN7pIxyPoiACNEiXzlFq1ruDgZ6swZbZ0EkIuEKoIeuClq3LW1k0BDClhZjv5uf9vleGogV1+M
SkzZ6heuJqhuMpblU/7b8e4wLiJhgRP10YW4kikHRp9MYSzah6ZhGslkZopj3npQ8oTYg1fEOHUc
QbOn69JFUJLFHld3bLdWRguCVTHnI4eNVb2SeP4Mue6ElBX3hU9xflTD71VjknJcYmJFtYSlMHfI
4r/uWiBQoH1vtmwI1ZP2r839T6bQmdr4EQuHdgmx3x2rkCOLYdLmR4p4BsaEgsWhDCJIuke2pMo4
sx/XfQdKTZoyAfPbqHx+m/nsKREUTS/JkI4KO3VYQtruVBD6UYUyrU2+NcFCkHXDLBuInQQ1jbsZ
F/tZUGie/fTOlF3MxClLczZlSvLdfjiQDNIGHXBaeEfOMo3Y5cJKWn479D9JigvLUPjP/8Cx3tB+
VD/qUy62cdVt6RLc6o/Q/ENKsBqsdnyaVqgfMM3x6GW/pRorVvxL8G7XPt8nlBgu4S3Qw8dhp5PK
O603BYlmCcqVnt/3WBg9a166CUlNfDaA/pzBWlBJIBR9e+FjbCi55p+dviSJvVqwUb4tyCUQ6leX
wukiVFbmUqim23CdCtLe1nv8u19U7wUaBg8wJbG7KJTH0H8mB+ibz4FNew/2SCo3/oryS6WS7CXN
MWDxBUmcstfWEMcb0cDyGMNG77CY/lNSpUfNZOsSjIoFyvHt6IrhcZGRhKJNGkaFH0YrlTNb18jQ
rtWu1zWYfhTac2fyHQyAn6og957+7k6U3gCRMDMJq0PHEZh5y8uDNWjYqQ05+GlN/zo4kxZ30xhC
GtZcni1zu1dcgeDFnYvBr2KLT6swmI5RUHa7uXqTYehMyxDG4FzryT8EGEl5/7KzCq4cuC3NRyyq
vrIBwx7uJXWvI5r0XFfCOkKQl0WbH5UeJL0UC92QfSuHYKN6dvgngl/UUBP0MxoDdrPTjBIC2YiL
CQrbGyUjAeMn8SRqfFdx2Zgu47lgLDdzl9rli7XLNheA0jaZt/p33kEnQ46BJUuM8CK1q9gWKP7/
zT7/F7Pn7IM4mXerioVawfd9605xhOq3RT7ctr+zD9uGKZjsfWpMOGHE1w0s3zlbUtm4cRFz7o0J
FxfQpX1fL8EW8o6D5khJQWymSULQEc5ASEPjzBmBbegziJzgXp3KC94J706NWdlm5Va2vJL1fOgd
3cUMhzSzEy3fPPaLmAETQ7Y473rp1sFCR7fJo1kCV6/WpczFynHv3I6t6maks5hWr7WIlElOW9Hx
2tuQ5rgCe7SZAZLWqYnKTljPjkO9Ae/O4bt3fMxAPIaN+xs9Bbe6iHWJ63rPfICCp743gJixztpl
B94pC0R1bxarrjphr/h120r4j1/ko+NsW2vPtZFCEkIUd3a2MTaG1K5hN8QBSvKryoB+W5bDDyCt
j//+bN3aFVrRO9ZtaFTOgh0JXyJJ4HIDyM11tHiisck968T8zbE9KLaCLUPbJlr43O1CRnWE0Gpd
KI/6kjEabSglngrNqUB5EFKHXzCInG20Qm7aGoxTkPnstuB65lsXLx8RPymbaDXWd0sYPAOpfG9i
PsA9e6J/pDfY96WlXZgk8vc2ovIuQUpzFePaqfEK7VzjfCaE75XZM8scTOBp6dV+50Abu2o87khf
+t+aY1c3BS/LMOSGcRamcOG9h4XxpnNLNH0lKhqg7sdIq4oz+st9ume5Ixzl1RYRg59pfKqdBzDk
qXCKzEz+Pg29b7F3dn56s6ZePxAWlArj+MwSbQC6sAhnEflv8BDqBWDOVET6RLEZb9j/ZmiJZaQU
JX/d/gVL54qmIMVkAH1YNgAVXYwG3W1sIb7u7ZuXzeootEXamDwrD5VNizMt4DgAYMBZ1FW6Lh0s
NQpW1vMy8v7SF54qdfWAb07J9UWdlG5JsUirJ9UA3H21HIGdgm+BLWZEDhjCtetq1puT5KBumw51
IT8HoVY8lLvQ557DNjCuclQeEYWGmmrw8Bv+E4IjZQZpCD9Mb6RqIDv9pfXNROkMFL5ZwUWV88mZ
J+lKnhiU2uKsJkHvX/RvibVx2+coQ1aH5Wj68663VZHIfk6LGpo/Qk3nZT258iSbeJZmxx0VGRP4
15iz6icOX+x5VvWYlJi9GhmRfN+o5y2dR8AdBkuxReeto2P0AT4uXZJ6kVjvsddah4wTtaPzA8Y2
3DYpWykxXGSWeGV/4tL5QLAw+xnPAtaFG3G2nGwIR30cf8NLuGqc4O5KB0jI/lDHaZMxulQZSOnK
m5vNDMlTct6vmzZ3Wf0UKASbrSqUdK1PLpmuXuKi3VukrThkNQy/iIgYvZTSmezjme0La0FCUrck
E0KtOmFboBrk5MMNBho+cWZOPZMLSL1hSAilmBig5qOXfqESlc7nHQVrboUURmDAnzLtal/x8Vlj
eRwQR0oTHOeOt8hgDgAP+pOp6ORmVM617Dp7BrBFifo90vDaSUnF3VuY6TeNmNso51i+j+2aHI8o
l70r5fXM4oG6qyIxDAHCqz6CvgFSKW7hVh9hfmIQEE9eMbnUJEzecqvp53Q6QETMRIGkqWdNLWvk
12Rm8QNZMxH+WLxL7RKsu/R6kzpbiMnNfNPBcOZmWZOfB2vtBIJ8BvTHTpNbWfYSQVZsS/Z6CXTa
lSXmYiwdTx5KLcZkXVZathL/sUfUHTlEFjD9yNXSdSDiUuq59J/sPmeU2foPKheciZmMjkIa8rdG
tVKHJyqHo8EC7HL1y3yYvYJjUQCiXRNrUlj8d46eYJpgqeVf+gjEOpWvxQSvVzmzu6zqjsjFcPDk
SeAExS2bQ1VcGmc2ErAxolzXgeWg4Qr51rEs9VIom9a+ntrCLroxhklZfE2aVoNIcc3FhxcSPVL2
6TOa5+vFHTEED5nAU2KnE7r6VOYofRXw8L9/zDT4H560aF1UQWuVnBzrGsaeE97iIr7Zliba6ejq
/LUB77keMGO+KdNd/T+Zo/n67UEHCJ25MFqcUkMNQtTbm6+TAb2HSMYmVEIhcS9duPu4TBd3lHUG
0Bnlt+ujTI+zM6vZo+HLtxIK/Has1bHUvv2u7AEvTzUU4+DaX4+fILM07paEqpQtb43AomtiMHCy
gSZbfzK/cvvqFmSH5NtLIPjVY5T+D76LFW/tcw11p5T+PCiaIzAOawu10uG5S7P+VU8cvWxRnM8t
EJGF6LQYGFnb9z98HYjjLJjA/I4LcePD8R/14chjqJD2wyf0TCKDxPHbJefzrrGFnmeadH/r1/t+
uObh/TLgGA9rM5zS3jNmgFaDwNxeDhH7pW997+EBoeO2UBvbOyLnuC31xZsG8bx5XidKUfuk7ezV
xN/8dmPTK3Y5wFbZ9PKulfRKOnAkOc73V3XrwNpp1GFHAcY0syeMN9xPNYMnj4lIholV4oJxfjfH
yJd8495rQ7CArvDoFF4kP1EaCE5nmk1Y3C0OG7rFskfnLHmlBhDZeJn5XKh5dc1VYo6HyS+usSy6
gFdV0xys0lYqAOygDSfwhJQ3twVCiv6/MFPzTWEh3/DDiXjvhVVhDqXshFdyXAMgAQVixrpzYKKn
YPDRb7yQS0EDzonee39mO0tj6UBdk2sPTf3Ks+xFOhRkavvltbGzRZB9e4M6LcUwlL5fkZjMfXjD
mZZt43PZ3204rJysMiiUD8LClohGt2TkhjD9D/WW+/LIHyvR0mL7t/VHl9+KHWkq1+o50isel0kD
b9/fdqSNVmaFNyMHfWjMP9s2Bz4GDGOCcnqYn3Vgxis5M3ii+lW/lClvE2IhNjcGXgAjwdxC2XZb
kkXq/eTb3z0udud0MIcCJvE9gR+R3kF+cS/DfUeynvXMLh9FC9NOZmkVn4EywKCIvPLm0OpNfKPr
eaByj6BA734Wt8qq6qFiOBjn43T83z7wF6Z/uSS7d9FqdmH1OCoaUTNa7ME7oIf+eDXJw/zpdTCf
O/DfgJG43a3RQIgC/kU9ZLRq03ZbVSxFlmCul281XJNwSYqL82l0k2WgRzh4wWKXDx9l6I3o2uXs
QHw2ZNPDC6uu0WDD4NUwNwLr98MD7YzMShHhXxUs7ewwesgXQxLI+7dPVIAxUMgm5BOuj7DtFKU2
rnlYFaL4GmjYvCC4zoxzSn4uRL94z7SzreqrQq1L7ZqqyG0y3b3BZajxUrQ1EJFyB1VRupNsKeMK
6uGgc45lBpdc3Cdon91MuREufFsyd1psGvoM4LdCJluJuy6dFDAROo0ypkgLmqSQGh4Wk5r7Ct8P
eAcrXN4uNBdG6iNiDGQg7iBnxZqgGCgnPGu2OynELLl0jkHcOqF++pQfdB4XpgE8aT+1upZz1CJg
iQ6Fso06slaA7v82Wrn8ONqObICz8V1DUV0Fegap4pSdsg4iMOPECQ3HZJcvKe+ky2ZRpX+HL2w4
9QUiaI4ujoF54wAu3rl2kH9UVC7EK3nhHchXZM+5YwqXjgA+53jCnj+J1nkdOiXYsyuf0eyLodjV
3rBAQEVMQTnoVihV8f+PO/2WTL7+MipFOO5/g+RvFFK8wBSvsFySmorcEIsfs8dN4h9wnJDctlYo
jOsrMXRoPzyEQySgAg/YUBAnZYMztPQDk6GZGRwjpp/UOLLsVDrEPchmRC14XdrfO7Am3k50E5lK
b5t8G6uTaVGDvKi6ExD++/hm2nD8PerqulNA7/Id4y90y1vBEwOvYq6lw1nAOauHLv49MCxhDBNC
I9JQD+NA44yil1kiUR8LzHWlb9mMlO3EUxMI7Dj6+nlbQqN3twutts7iYkH8UvwUHwUIETH2Riko
1bDpIFi/FVbXWQyTmV6YQSvHdR7sdABLbstPAmf8R3TIhHx4Jf4yfUVgjyvG9KWkcK/IUWF+NZdh
F4Kx+5ZNfPkiPSj8ukZmW3Tgc3E26YdSquWTPgCdK5REym2yEneYNK26A8vlfxH0LSQdrSkWDXrr
3f2h/CXWhaemuFiPedwfQYOoWb7qSC6H0vFn1ZO/4rrfjMcBad7TKqnzuXV1jF6fV2tViTcy9osT
smDJ8780Cr/09Yn6WgNTpInWE36ztemqHErOYTS1XIJGT8cdAXRAlEV1iBT2AF30EE8Cwp5MopZC
+NuUVEcYCRj5hVUUTvTwX2/Avx+G2DXDMHbEhFKf5eeQdlXnPCz4asKNbx2PqYtqLMgBtjtffWVK
q6zcnqOLp/z5OGnSbfoXaSDeHUNoKFlHU/LoDQUiy50A9YRQASiX4yfDPb8F0U9hMxJdGOGjMI9I
f4ceMAafzIi+BoTBpCSkrt91R8uE//MKKvDmOVWPtgiQ+k6B3Roh05NlHT1u4p+FGF7XxEob65bu
1tU1bPv4TbhkwWEkE6hGixoeCRBWppaiRF7bZdOziFODhh68Wl+PEaj1IJlTuhySDNPcTN1Y+4fk
jEfcqjfii8PSOCnnZf+VxQpUBUnr2c2EBSJL5thI5SfphXMFMOrAa/1XhUAxKDVjvj4DMRPDVD1M
n55coW6pzTx6E5B78I7O0BX1lc4G/XeMW2KlCI3c9XmLXamvPffGJ0Rm4/DjRoP7DqcGHA31vIsE
vuVJHYyxy/N1bgGuYUaJe/ziXOBAdFSrwPrr/0sr4sujHxNYtVPWeE3jA9tzNq+Qwx27khtTmP4D
Y8n9+zCteFmxZ5JyUIrgncYjMYrmidFEeUVo8OMIv2sZLIIAemHENwm6/0tIL8V1gMEUzvwY3yIC
ej0Gcd1kplap7kftiEx37IBwcgxVhnKAQ07YT/pkrLtmg3GDq/Gpv1tjXc09Qkh9bpU6A6aPPrCt
YmpzSOZAhB0f6eD+GEx0sbSCZz3aowkMMucKyy9z6aoFEeP8yOMjiDhBxRMXgvtquPCY2gET6yB7
3ealEmjetc1Y5PtugP74KP4GYTfQVn9W8A4UlNqBf/3U3UfWsmMQnZX6tS70goeksBmEBrxayy/T
KitglommfuJay05yUbyDAhX7fbmOXnBoF2O2fga4QZmKWgSdPFK2Se5L1utVfSjWNOjyAyJLxvFX
Dd+eMBzQ/2h/3QxkiShbjzXbHN3hl1H5yucxL/3HMgLdhykvzsnlCE+a4WqgNHxu5TY09vfez/52
EY4rRi7+N/BsWrcPla+X34OdRcffk5UMm2XahNWlXvUIm0qm10pZ3zH1SQHVMC8//UZWzeEXuo/8
wWx4ZHetgm7wzNR6MJpYKRSdH2MDBTak0t3UIBPYAhJx5ZTBuFsrOQMZP4tG4Q+rkWuh9DUWGTyE
zJi0QnAdGWHLIw63v61LpNQ/DAEPFmmxKln4F3UW8xNZ1XVbHzQbmzoAvV2UDDpN//Cxc4jVbdqx
Egt1GZsF8Oq2lABu898+slwYGyCd+lU2EAoyfHEMLoWwzycOnr30T9gNpK3ROO3mqWmsX80Y5C7w
rWZPuIgaRNScUDqZ+Slt0MZXqkrs9JoN44WZ5ZtO8h5C7Po6zyYKGPbW3j3gyOznTsAcRefNe0Ao
mF7mPn7eGgbEBvnx4QNI7sFwQNpSOwoje5IiRXhzdfZkelG27peAz1xhT16iZqU0W8XqFvIDn+Lr
j1E5LDuaVNBqojsYnFdtAcACV6RMocnb0gx2t2XHwXgNFimYA4PV10yzN02lZ6q5lCHsX+HIfbbJ
zYlt/WNS/Tn6Fwnx8LcdgaC3JYRzC9DisUA2ZLvU+bC+YNFzJI2vw6ZCBKE+urRDhp1q8uDOztTm
Mg1Wo1AsGx5fD05unQWpbc8LWXwQb69Rqp6dkfVVxOvGi3MwZBSFuSWkfuIIKjCGnjLPFA/R86OR
HJWuPJl05HVTtvDsNL+aUBVlu0Nhhn/492Mj9wuRnibd5qNqwx6SUtgIB+IQGG9+Mc1qYLrIAo5w
klPqK3RI3YFAM0IrFIywut8soOj/R+RhO3V04ZDvwGezMkoUVfVr58hzS7VrtShbgnBrYg5okn84
1ItsJY8sURBWEqbPW7WZe42cypZLUTo6ssqoBXT35InwcxbEdfhCo6JzLZVepXfQGjqk+KezNa6M
6SwibKXaPl0wXIk9gL9xeB3NYh2wdxPHi/41gJwGsds5WOQ0XA/TgQvHcrM0ct3skVC102bHZ39b
uxbyM6dVLyvgP1nBTJDZ2iv3JjAplMRwEvWSy5Ay1vv4qA5YSI6Iepx4U3nZyDfmRWmhUZua31u3
LFEr+4+SMSOoXFIdiidRCa6NT8xvBKRakg2seWld7X/iel+OQ78tMDfpQjJP9B9vjLOpRBEdp/jA
8OSRaICtvOxmHu/R5vNLRzliWrCAgUMRibA1K/idK2fiuEZ8eNACMkbjj7APuKCCwUnZdlXXkSU6
D694h8pkg9rPp+BnS8D4bMdOz+ygt11SlaDm45hC75yyK6+utUWpsB29/HHgpMeI5JlaLu8mTZXE
DmsP2zxdKjEC6RAO71Hr5NDRukWCGRSshOgoYzxqxqOEMGGkwZ8ZT8GuHgGwipY4gQO2QM/TZvcz
/upiKaSas/qCqZblBnGMh0BYvHmguCQzr0XXKIAuGWGGQoJL5QQ/SI3jGFcUAxU29sYuDMpSUzMc
OhR1ZESQbg28FRJuEgokLBVcYcW/a9eSgJBKbHVsh+veX9umj0wPF0YXPa1YUyOn4ewuhK6Ub8HR
ZgpAlnDc9zWCuChxNjdFVR88Bk2HMNTo2TEW2AntXOh13PfrjA2eVsxDSN99TA5Xj1CgSjyY3vmc
989KmT8khveflYUJ4pF/Fkjd3L7S8AJOP4mchhm4YbHKyynt+merFSyq+9vVGCEgUcWfMdr2qvob
US2YXxDBDtwrcZQo+gOjFTgsrWcDK2btkl5hc1rK76NESQMz7DmfuaNi6C9e0RbFmNaQWiZgEB49
ODD1wHvAXH4PU2JTUyf+FewHyIKGGtWe41rdb/98P+OpHm1S+YLkFlZtI50BcjpOV7rXpH3aR6tr
cDw5w0lLFKlj1IUMe46UK9fLZUUiEiougNM9h9WYkzF0B/tBupqj97f97suVhv2Zg8saXcSAjeG+
m4t/RP2oerRzyajZgFhVpAfsIyfCmwZTacIp7SxejOexqss8jeAVEzjX8LbyTBDFwVes0mZXUydZ
dfyIU1KP6rjkJ6NXjSjs9UW4sZnTCCatWmN2kxgsnVMJbaowk4T42ksccImOqpB9FTHFFF85x96E
0TOUhlU7Kty1dq1fMF/hM0DI2VmJ3VWMS1QDBpsaIfQEoC2R0F6u+ws0/dcckH+KVV0P6efxvpUk
QJfl0FNwfOobfMxfF2nsaCJekK9iHLS+iKwxURC53xhKVKV2Oo1k88xcf69jxOhLtvMDrxY42KS5
mHQgFHA7ycqgscICT8K1pdB4ciAHGLM1XyY+pBH2XgNpllZ7XpfKQA9O9P1IQY66EvD+2yGSU9Dg
P1f3IZEYGK8DXGMjCGj2WWcsoFwTa1KA+YjxC1Zvl9z4FzsYFkYHcA0p+xBaVdKDVuzEDdTNbGQY
YL3j2kc9jmekIHf9oBnXTEyU0kY+Xb+rsSiBKASAqDqVvR5BRro9qpjcm+P+x54UhFdE9d2SWnJ9
DTW57M5hf1VIoV+6WVJpv8Wx0qJqNp/xlKRJNApcLbgB9S/yhvjT+MHX0CONFf/TQVIIThal1SKc
IZIGhAKglGcjsh7kuy+lt3QPDkS3iuPAGUa4lc2ppl9yx0gttC18xpOVHf2wkUCz8LbEGFSKIQuY
2E5lHHXUgCfdMVJPKT3++AtmW/ZHzdAis8Ja1Rsux78hr6vb6RHSkY3eRkhttGQal/g7HMTZ0hr/
TJlyndbQesmvlT9v6cnXMMLXyk9cllyHc8XajvwvhpTsM22599iqPTxCExb+sbHItjFnQTJNs1Zp
llxGov7nTermwMlopQ4Nadbncmm0e2N/8CQ/lNyBz8Zjsyk9guIC/+SyTTtdfeCDDUWLlu/auVv7
xYF4jUjkv5Hu9ujf1ZqgeVwkfDbrpZfIWffWV487zbLvzXrMtX38Jrt8mT1X3IC63kFsKUOK/UlG
AUwmSRn3ZhZoAYVBWVDdS62KVNoPbEs4WGpNrV4GQ2eTPfg3zi3KQ21Xmo2ypfNoHoDXOcdFBuZk
4cjYgtNkACZJXjTwbBJOeai4kKiKUc8u+xFn6cSpvowgDtFgDa5CWvoHzEj0zxYSyOnu5wDEWCcz
EzlDnJpq8NsnRamaMV/SxiNBZoXwLI587Re7Rmdz4Rybvq7+87XqVSncv29mqYiHRYJCIbfdrQeh
nmOOUHXF3cplFYVJf9MYnI2JXbVB0F/zPe2SAVoGXF3bik/HluutzBOut93CvFow1vbrZG8WSNzD
ILXKpMEcR1RMxtBTfwcTxq1mrIxfQj6Ci+L+9Kl2DFcfEyB5RpPhPbj0dAorSbveLfVRp6vhWghQ
efsVuDo0LVgd0iCjYF9SCQsd8S/LZqlIWSyb+INy7XO3V4sUaTZFbAU5ilFC2gXtVFZ4sru0xRSS
7EIMKI9EVAvbUtkogjxFvXy2wSzZyvegsmdeA9B2206SSdu8R2va9e3QvN+aLiiwIpzpUjXQdRrt
YmbSy6Zp0uyzaTKAV6JL7qqNCPYx6FGcIRW1xsNlrsq4d1EGimbPKg1IlzO32A5dP7Aa/oOhWNyr
tENbcr61pVmdD1RuBV9ah0oo6FIvw2ZaC8BnJmvxAX+hGHe4aroVAScmJo4RtCH7HxJecKPrkf4Y
B1p7UntfhRw+r+atc16PCbTnkBeDzBH2DY+iGt2PVZ9VM8g2YIGxGw/4E7RNs4fIEVgO5rzP7MCs
YaEcP/xhI0FCmVjFmwLru2IbVQaBoRvNp0jgr6vBCkmFGvc9kFTRmrzeMtyQDDuBNwD4+fUFGLPJ
92rLPWd8nyH2TwkHCcnc6yminr6J2oAw7yrmSi4HgcknBVjDrQ0vIpMwpg+LQDAYOvgXteg49a75
LXehMio1e1YBydzIKOp+nJi3KVSpFeN3Um5o+m9Td5emXQ7fNf2XxjDpoaAhzrlPv21fAGnGU1Tu
05CpKFnZJD6WYGiCz8tHWAcw3YMqs/qbniBfyuhK7Y0IRC0d77ZmP5/QfZ7Lmt2jxP5cpsIRfGyj
WCHyWvsputgue9K1mso24263r0i42WPp72mZTJAFpggc5MqwdL/EDdy66m+faXB3w5l83kEkZhe2
tQNe+vzaZ/qFajdtEp0YbLhZqmyN7WH1WqV9t185U4OKQhENSnyeR7UgyfmUT4LIVwaztXeSCG4M
EFAdOcaTtJl0AXRXOqaZwl4CNGR9WPZUYzjNthqNuS2MYkYwqZLQvrYrdVTCggORyjQS3PzjZYnn
AaIeZVAJo4MZwSNv4ltA3DqiCr35ZJfyWW2iz4EtN/cbPhAD6rrubnCdBErNqnLvUd/BYsi0K05v
i3ybKYaDBM1eBYHeE5n+R1UotDnRL+iQk1FLpZield4FFkV/iJ+I7Q95yg3csNLzoB+tdPfSShcy
oHk2cLqgBXgAfM88jCjqVk+g44Af2xxNrIB25S19UEmQ3NOhZzCA/BkFaCpMQXIV9WXcB4R5NDin
4u8GlSm4OCW7JsILJZIezp0NIi4HjJd19NEFT6VdqC47K/XdndfCw+X8SilBITlsqeBHE8qXRlgh
pv+92GLrQUyUPG0/0IvPUhSPrGuKYEOXWNh7aIssg3RTtH7Ldp3RPibsK1VEYuMv7PbJR2EqYi/Y
nYCPVWBHf1vbdCYhglSGNRaHYxH6ADpuuHRr+k8HmMCtsTA9bsU3m3tz5VjGm59m7ZBw/mZEqRaS
uKNM5tJU8x2v2THm9ASUotW/jAGZnvIV8DKv83z3B5UG/st44t/ZwUIdf02xovcv7ws4VYvPtK4t
WNvdvLQMiEckr4Llm3gosRwioWU5KKaDg6bQhNv505BYk9RRWNFSkd+0SCyvM0OUIBPhq7L27pdN
D7hnmiAZn9e1zbw85yAkhNXyeuMXziQrA7m+xFw74Hib9lRaZYHnwOzZe1qNivJOMwZDHUT6f8l8
Q5ET/Xh92FEEty1OLd8PsD8/+wgNBCjRaFnLckhAKwfbHOCf3OekHOJmTF5j8KkgIbgcJkl+rKb6
ZAFqOLO55y0nHfLiUIk8JlUOOGSF89gnMJrFDc2+5W5vsLromT1tjFQzZty1k8WjRUMH8CTKIllk
ci00SbNEkZepNrhor8orYcyRSHpyYjdgcEVnARnLiHGAOwL+MA/Yi7bsdS1H91c8sFJ/m9WdSGuj
yrUeDolvnYNciVLZyCLMKNMNvNRa7qhfupQu7VWelTeBhv1g/AYZ8ds4fnmJXr/fHF22nRVkiAKg
Q+Ivcmxt92ZADKSvc5rwL/h1nQmcoahIttpsVNVV4hCPXMrum+T2y+uYBFBgWg4utCW1Tn5jwJUs
eTZ/DCg937YSdYkG7P4l6NWgY81rAihJ4MDpyenVa28YcLiLOD7Y+EQP4h1Xlilmc+foQMy2kmWm
RYoyfo6GjeNsHOZovVu8ELEeZaLwY7aMebfNsn/UIwMDzl1YIPEQ7wBtWlp6K9ardCk2LirMgRHT
y1XMUE77kIQag/GdCOXF7biyJAwZ1PYKjHbC6C/IT0/vFnMYaA9uqtVUjR13RBoNfDvHfTCgF3qZ
NX1kz6z8U1N7GgmfIcgk7zIPyAtqy34oFWuPCh+lFm3SaOdFSX+xxs9WyEmHwhjW5crl9tKEwcon
Sx+ocnk1RAC0DOecEy7UuIeObKp0iQle1GBIIIiy9LodWKWOrq8XrUDBQCFdiT11E2y4gFTDk2H6
QFzVXdC1Dld3tpcKNqKA4rLBLKRsnyPfsArWd6hMknBY24HZx7x6/omRz6KwRNqtpk4NeOr9IOeB
XYJTjWUSWPJ/HMP3sb2sEE+cqdaTQUrY9LmJlCvuQcthTO+Tz7IVbezsDTTQMb6x7ktOArKm3nq4
hzxaPHmNQJ1EcAohOUNlprd89OIfqmY7BTA+gUon51jA8G/eNRAQWp490FCotuuyEKmJ2tophDJ8
6mT2o3Kc9Yw/vu0HNo4kgavcDpgkp717//0yR317kB864eDJR7lpREQJnNIXfWZDUlVJZGvK5GrT
0Xd55yxhevtIZFXz7Bv5sSHkc1KS+Bun1ex0gT92eo3CuRoD/OTR4p0aXXPi+oCM8sAV0pALLGUR
h+fW8uPrYSGLiZTGFj77jZBSmC/AR6UIUQUcvAeRZ0SYWOR/bCpV26UGk19FF4FtAqm+SLg3jXpK
sGzNOdgdnXQjArOgIcPYIjbLdAwVfvDJ2hiiU8wfYhIZ3YgvCblQ1iGHUmhJB+C/p/eDhpJ+dWP/
KLznQQ2PsrfCp7yr6xOGE/qKCH6GW7vWHAS2W12q8/kGHGmdQU480NWao5kHqtFrt9dFmOBiayGx
JQsVoE2YszGXApX7ok9UyXc0J9C7/5nKNn7R22Et9kblpi8D1rFTAL/Vk97BoxVcxV+EXtU8IUHK
a+j0Vt1GdxBs7Yh3bGgnFOn6VUN/OGjvcWE3H4g37XGNU/gdU2+k23hKbIMxUZUFHdNYULYV36Jz
fGxH51kKVFVxhb3uW1ePYL0RGOBe2Cg7slJPsXK1jGhakpd87IGUyJw8AcsBnrNNChn5QlGyM0h6
A2bFxa6fEaj5pMnZuHc6k8oWzgU1V7Q+yQk4Os15j8N93+mSpD1jAI3yIkPAEAi8vlt+E/dpYrnD
rZo4WPNWryoEQswuhrwit/+XcqO96ZtoK/TLcPSYoaAosHh+klYe02gxEDlNlsZw+z+KjKgfFyXO
9c2+WhiV9tG7ghVlA/ZcSUnzG402VmPfMefqGoy1nVQbPxB5oLw4NUDPcqBcQxWtl/XnM2nR/AtW
iWb4fixixbmHBFoAOTPhtcEgauFIaovrH6he3lcRXW0tngFJEwC6dOA94vT9MhbIUnvZAWacr0V/
dsPJYEy2OpWl58sTZPLgcIgHLH+rzlsp3AKKE8UTWG/GzSc8NdbootA8rXVZw/IqMUfcHGVImVY0
rdeQND9qxdAoOPLJM+ewn5ChKo5v0IBX+7umaMoXRLJxU8ubG3AcUq96NG6CBVz5CY+YUUAt3zVn
vHoeVfb4qzm5glmSS4J6ri7a2RQvx1CvWKZL95vyDfFD4gTZbNRXpp5K42h6h6DMSPVu9frQgtd2
eo0RAn+QbobM90NOHKBGWNjPBIUXLW9/Hh30Tyxdod+ig0sCUPaXetkvcOH5zPiMyS4ifyAiX5t7
yHTIK+kPgpomKxb9gWCAmNPHqGDDI05UMsbb4njcTISUaAcdjGj//6Pd9D0RkChFsPq52UUQUMEK
7BW/gCuIcO8irmOe6FtNXYzwnTZgbJUQ5JV0F33kyLE2u4pqCi0NbuEr5jAqEg0o9xzLgYCwGA7d
V/J6yIpApRA1XEflq2UVNAjDol6RR8G64frTuGb6BfnuW+gyPrLYzr41nSF4OFG1SDiQhIn2Cjyt
a37043WGcFlyY45m4/jgr/2Ewj/Tl3jzj86Und3jWyyQPrI+x9ISe1wdVDu+mmzbY8IUNc5xuiLH
XkMbUgXPryM8dZ+9osmbraqNw481/imCubzmw6gbF1hXK6spXAGIlesSfQpcA0qvToB/SKCy+tck
FHSMqU8v13uu+fwuxvQZ9B8wJj3LVGUQrWWUDbrXbIeYLtgxP6/OLvNqbnJLAJLk7OPfepzzieQE
gi7stVVezYjnfbEUS1WMihpVOLbB3Sr6giYXkyYfaOPoFXb+NyW+D/yNHAMX6BAQQf4iQS7HDwj7
fIvUnuAqNUASZUiffQzmTY62FphVtumKat2s3IYloxIk9Ga9ZM1ZMEQKuQrSJ8kWMdthUvKENPr3
SWjfKaBsfvBIzH5SgggFhIWEE2O/YJy7xmVIwAt46j7h1/8I9YVIzglKiz6xoyXpcS0/ZcZvXt2B
Giq0h05qpTnm2AKSFkvuFk6d6LO7PSmk5tNJfkIGAMmw4l57TVP5tx7oI4UdN5DqPBePQ0TZwb7q
xQyvWyf1Y/D91BFZBtC7MK4KNOGxFTWfd6ZMwcKC3MDa7c1fIrUBkaCxIXn+akFAyErrmcRdH7XG
L/S/qHs+ufdsAquuHv1ddTGnLZ1lFqHP9m2fzcD4s+duZboeEtPqhmZlJ3soBSgmYbaHhkQNoblH
g7HzCiXcInyd95cHcTTUnMHB5M4vqmJuivtUW7ah7wYLIVAOSHuAW1W2b/hXetKmz+XHDVxVvqHY
3ZH00S7PlrUcX5kq23FTc4BVWKm71s+rfk5rCaXCxC/atnuKhtsFTB6aciF5LbiY2SeQ0KJnTM27
F9hf0ZZNKqJsu0rCHsbWDHKSGcqoEaDJGEGFCvsFk2o4qqCkyj6vb52JcvdTSrpMyJRAhrjqGjjX
k6sW4IbDR0xfb3Q/7PDGuspjNAkzjRL6uaBiPHs7eeiWLudZh/wPx15AyUj0LxEaPT6GHii3D7PE
6FBx8ZmE+O7+xisqi9NqHPtDvjFXo6F4q4L4dY0IC91WJeXaxCx2j/nnwqy/hw3r0TWbMPaWpw8u
DJ4jAIARRpFrCFUNnBJb8TzrSBa9Sz+oyuiO5k2OdVmHCQKJc632WuESd3eF2dp4O3Y20+OJVqlI
M+mM/wRPgolMqOp52uVNN7tuabKCZ5HY+2broY1/QOFh6fhJhdSKNaFYtwxowJDLIQMRTNkKUahx
6+sRKtJ3wzo26bbFdb8XbwoVWYgdLHP5/WpKRxyuZ9nol0YJ2ovHZKwU7ZKiG6qQnXnXKGW5hVQ4
oBUDHlZ1yTNyWVLnlHWZyLxVU16CTbZ+UnlGY5HbgQKrfRCTf6AR47mmQD4imn7mX08lf0oDyUgu
gCSHph5TujFDO81kgMHvNXy0V/tgDmDt6x43wg7KjP+BB7HuaQ7aQ71YZo1Oj0rcMBluT9n3PJpt
Br9Bcsv677W2/7oC01qugmN7aCkx5i/kQpMZDWq7Ze3aJZ2UtH7GmXS6oPGD4ZRnr9SwsaoEn/Eo
y9D00YyPLnJ6y+xyG0CTlX3XvZPFg0LGH4hYuMTxkWHVzTARFnsXcD67CIoW69O+oYX4sSKGtv3Z
Vg8S1XbY5FNY7HGWayCzMJ8e+R8NrdC4lmI0lEKNDLi3/iplQBwskdPO8Cxhf4ffVzZAzsUMbiQo
nKJFczhtCEVITHC2Im40BEbSnRm3M9tsfyhPzlSe//XR1gwuxpN0xJZR5Jm3Rr/i9JRLfPc/4gmy
5dkalGyQ3Nu9KLbJ33iwVTvjRCsqwOpAVcHXPlF7FfQTv40E3EDSsgybY359rN4w6L21ZkDsLyLw
zideOkJXwUzp/+dcfT7NQGkxuMbl2sDgwG/xS5sqDCUhMVzw1wlSS+Z+mdOGwGXldnGs9KnMOyAa
5o3iktmgo/RA7CkQK9p7M7gRv/gx5bdHVUQe8SvHZqBEaEkmfGKd6R8mi7N96PsjyUbNzw2U1InU
x2/HeECyUaXZy5KXSvtr9nMFd3OCLpEM2FcsTZxuTLiCuv9QrG/w+yshkFgRelnJOV1n0CA5GGmP
vL1DXhbNdl48cFhMuvoBFNqIJrQGM3e7RyPmYTepFzUOy1eikqG662ZNHHWkw5HwfhNfH3exI6IE
oo3UH0FKNZB+8p+9HbTMXsrEQ6AYfaWWIW36WthTZqqNoP2awEeTKd0D4P+ICg6KySZOIKCNiLYd
MQ9smEpxJm6Pszd0UnOe9aUJhk8V3tfCWQ8GfwGe2WemwAm+2eKOK6qA1yuVUpQvv9hunmW3ahH1
pHgkvNz4vD1rLBJ39AuebMJzzm1jmZfheKMtmay4+QEYOvsK38ltLFgpBTVeInOcEAnmqB2XMx/g
32Nr8F2+3XIt5lrxnMMswkrzNrkZ2JrdurE22lvxCskaS89HdG6hS5LFwvqxfs2deuWI8aWmdWZb
j//mD6aUd71xIPgqFltnU7y8e55T0Q3QLq6bfbs+PWQg9xx5OGyPEv5ktLOEp4dfdofl0C58oB+X
Zq+sXD5C4ZmvYHsFOrACdEIYkg+NoNrYHX495/oqMSC98sGqM66Z/WzclxfGqu2sOCvHCOmX29i5
AJkM7P+RObZQaccXmYhyYSYULAJDQTtDs9BFejts1tWe1yPAgogXKdwt1A1vn4nLF2rBd730WNx9
7zmbob/qks+ToCkk5YZdM7kgTH6iLu4YmiZXA0zXdK7hC1jlYGvRzGieraADpwHzltC6vlFvQhyl
nZK73jk1JaitqjxfewmXQ1fy2mXS4DBn+JEX3YeT9FJXgfJFyCYzh70oj7TyY+aH6ULAGg/ONz/m
6a/XYX9FB2l9OiicmJLyA4B3PWJbuz2Olvoap2x2H5UpoMz0a8xJDeWQ2nvPqNXhclJSGxPGw5Mv
Qn/cQOASNknzFqoVtCkFCQJ1E4Z+BIfslXWiL/QbEEgdVSncZB+gLnMeQLBRpicbMVT9GAoVy/SB
5KfbF37eEcLnKwORq3RLQzqvUGzbiEE8Pu7yFmspKDEp5vKFAQDGKznJCKxDjtZUrBukrdYP11IX
pzZdx21iV+Phcjv1KSoMZfA6pynl6WbG/MLmwbosiyDVkerTrgVm87eTZJafwa7XqqkRT91DDb0s
NiOmrZLVOuEfgvtC8B90+gkFIeMrsW+3Bj30TnarmjPybBCtNvRPNpwKM5QHbAkU/tdymIvhMbyg
yrgy20Jyi7Ka4HinNlQB9I/C1iBSfmcID96HfoixTmhZycYf9OITAjLH9PGLrkXWiLlsXijD2mu+
2z6iwkJLssIx9XZ26Gqhupm26LIJVf0VJ8dY3HdMFzRT2li4e83aD4MXIxzibt3qzadi4KmP8tfX
64nOdXovitao8hQLS2vDw2MwRDxbLzxIiRcEldAckTECtHaEM5S4p2Bb3UEDsvlpZZHBJrzqvzyb
1AtGpJNXOEVNc/O91PSp2r6PYTVRYboAKf+hFsbo/T8bpajoAhO7my5YLu/FoLH7lJq5J7KT348I
vkeoHtmhUvys//vzfxPA9rYPs5uzYDtrkRSaLUD3voRIAeTUY+pS2NoZeGJ1uweHa0D7SszqvtkF
AUuXpJjMom8fV8M0hlKOwwpuGbRyYQfaxfAZIHGQg6W7j0Hg1y79sSZ5jyIe+EFjO1XcyaYopIwt
eB2WikxXPRbNXoU6RQxbWRk97dqp8ZhPTyWONprMEVY6hBCnLxXV0FggeAU5hQ7IKPsGnMDsmFgC
RZVYtwWiPS6NGUdMbcYhi71hSm2KeJkKbC85qbG+eGNskCswEULSLsbwGFw6KuG7iHHXoZ5HToRF
2I36N9n/eBtxdjPej06+Sm1Nxdrna5+bkOjOqeVwio/QwNoM/06XPPaAnEd94xsad1kbILFZ8uJl
5fZbCaKay5mq7ny1RWN7+OYSHPqVsh4TWQEe+sgoBz96PUxYqtQu79ErvGsCKmKuuexSFrYsvNax
dvc+BTrxGlIEfL/bXW3goGot1A1s6WEKcv1UM2txIE0S6H8FqIWKtN6yO26sN3iWx57+fPT6cKkI
TmiN9miFrN7tMeJ6dsznNuwFJiRArVYpOeHkGqcCTyuCBNfo9gUaVI3+NV0Ll+Wf4Pz+U/IOwGr+
JHwKm1V1cDLGxtayY1zRXjWn1ufdVHrqRdZDhpmzQElidkt8DYH+1WYduUlZUvgpo82Z8Gy1QwLD
03CggvWNNfRo/3221yESJY+jm1AoRCbxScn5S/RXUSNdQyKPqpRGGxRnV7i1k8nLdbq3hcX6uwN/
J+CPEKBQq+awYkDruMfQPYtM4uVjQR3GuPGBhYG4gJ9mkUJDkSAKUAeoe7ITMV/xIa0Z7lynoXCs
mGaD/ofzDFapxPAg7Dx/J34BqRypbEHK8rppBuD1JQIeNYIzdUrxCMs0H6e1ND0CVFVGcspcoGqm
v6rpbeX098MY+xaNvEqJ5p4axnT7LWjif3aGfbJnOx2WMRZdBX6h62/cpZ4iQAPDSIqGQZJUGQ1/
hiAi+XspZOlJVQrHP/QpgyLnfVVRC/vLKYJFaDc1lCMwm52Qk0asnihKxrGOTh541BWVZ8ic4Zn8
dokQA8kWbBUgsJeneZrpP7bJONlCt7Km7BcD7xXHFqXFcQelVsNSqPvku3ZMOHLtHv4FaIHUxFXd
tLGzgXsXui7ena9yPOjiyHAiPfSvnlOZK/t3oj/7hhMVsQcYkBBFb/kHnjVw3c4HauY+KAmiiZyP
pHkPiA55+9gms4llwZkQjiRfKHjy4wcCTf5BBzlrskaHIRuz2UygksYKiZexsGDSzfoRBBUJThzM
CDZW+uw1DQsU7g6p17oZtrcmUAZT8foVHZctDiCRPYzydtX534vu2/ULRu30ujZGjOlRalxEH0Z8
3q4rVV3SHg7vNLgN/YyoNeHngaW/HqBuur6MhD4NeehtOwa7rgazQ4Dl1/sLdJ6UgKgUsebYOQj8
i9zDlm5j9A693tzz5WWUcU+bTsfBZMYLyeaJdA40/9ToBY6F0p+NTlq806RwEB5cc6WcKYz+2xB9
bhg5V7ns/ieRrvlnpXkb4lOZdmxN8w9wBF7C8mU/ZVqT38TeFjsz3dg5p8lM0KpTeBM6PjcCN6hE
FF0Xo3NPY2yvI02xp0Z3ChWKMYmm09ISv/57p8gOKWYywxHFw/w4Hy4j/mmC0N8X6dlzUwhzLbVm
5O+cvEGxnS4RtH+a9s0Epm4zrygwOiR441J0ynPgnKQfEwtFIdcpNIDPfpZPDOe0j9D4DFgvBNoa
hqEmTfjEsD8P6dg0Q7gjzN3FE7O/ulpo97+p5sEJtZB6dCIxANSbM6mrqyZpnLedmg0R1BQPplC9
+QSCunqWrnEK1NZMnJ3/e8l13ZGFxvy10CMUDwiqWgRcVezrGVEEN2rgxyFgqb6+TVkZ1VN+/TDi
iRT0H+nt3n3KP1oSL98iRsN66U3vML+zaQkxaUHC4MSXvINyhBd7A7QepeEN7th77xYon7q3PGXQ
fh+Jj3kYkv1HvVHuQjl9MTCDBb+G37zo76q/dKLOgAc0yDgeKA/l1QUu+pglK8tvL+2Plr29T0qV
Eq35Wo0exCYNIKgQOizDLR5efCXkZnSHl3y427RFCTN8iLN8xxA1vgocoC2v7/rspN9yYU89clmp
2/RjcoT3OyJTzBt0Z1dnYEe6phIbjlbdfYeE7Du0OeBe1J/G4Xagjig15+dX6V+Xuamoo2feVoms
kbHiNGVUIfdfvXI9QLHMy4I026lG1gkxFGf4z44m+AbYNHjWW9aIYiXjdSS2y6C4sQSUMcFB8mpe
Dddlhow6nFHGBDuOPQ7Xfs9USIikl+X/2zyjbQUD4QAbhvQcshInFQUk2/cmf8+/XST3Y51bPELX
G0EENAXKrLAV7FHqrEeL8T/MEgRQWqWKO3om9/kJoGd3L4AQwR36H7tlXHe8MsbyPM6oprfX2bY9
B7R2ydV0yU8bjZr6P7wfBgkU1pmYGZz9g97SjD6Two18RktNQQBcKhl0NUhOKyLpzsiFYOQHjHVJ
DBIod3GBEujlgX3ZiGE0//68ToI4duzs8Qg4u0bHw7QKnfqs64GqTt7QW8IEqRGmNEzLmce2h/2J
8o62LJPA2UdTtYCq5x00hxLssW9Qxoiy2VkE09yNLEvS/37mqfMsnmTOH78vwk7ENJWFXn9EL8Xn
FTLaHc/b52miDGS9r4fofXuZw50CV5FZzhtL5PdkqDLCR9A7ICT4MgJ2eJyvf3cCWPPSKMgabSPs
T3UTeFepzaqOVub1IfnulXnfuHmeJrxwoanjXSZ9F9bHTVIkQykleBe88u2JJu2NBG0MNAIbCRUC
hEFiKdT1gnlvjrFS+jagDxESJgHEMbe8qcaAv+rZJm12s95C47tUfwZ6sEkqHJDXsf8F/vrdxLdD
m9cFNYR3m91b8Vs9lA6FElZBOniFp7HetpPYc3idpmgfTcrHTvDenGtFQMoD+eP8PxkAb3f26Uzi
MWoBf0MLIKFD/ZKahmcTc8XO3Dii35xRJFaZnQ+Tefzw0AnX57cz0uTWt6QHiYHKHRmbY/o43DQl
6dEnr8Pq2wcRDMFy4jaMlxoHvlLZKjp/C/loQuhxkj9/XKGQqb1OlF9pLsqDW/wLCGUD705b3/K1
LiSeEiKilMvlA9l2VJLaKpTTHWFWFtPU8VLdr0xqw5KjW/3FYtMlvpzxDPz0Ddzns5xnWYjUHjKY
xdaVO1n/LbuCglyyYavBRXaCu5pYHSU8gmLxQwoG9iGPgTHHbEmgX+pRNpaqDovBOaPNw2NhffdI
MV73X8tl0T66+URK0hwlqMP7s69gn21g98dPTy4Mr86Vh2oSSB5PYAD9ztBVA3yIGantPW5GXx7Q
3Gw1to4SZ35TZZC4xy2fbBXe7wbXIfXFEtvYhiurp9USIOcBMXQBat8xC4QL6H9rsoK8+r8EnzFx
mSLZiDGyuQqU89DWy7GiehXaJo5E2oBSYsCIcdad6iNT/vIi6IFyKRAXuLScF1/8R4dEPredzC+T
29XludpAQrr4hRVHoXPhVbKpZYcyFhg5RuOr18L89Kzfj80P/L/FzfryGORhEatHEYzuO+JWGflL
1xGIy9eAkCfV/KqTURFv42TiQYX3I4BmFRcPaytIRVmHsBOMEzQOUF2JqWCq5qokl0pRPoKQOvUX
q1dExDm2VMG2k+tEX9wvxkDgNkpPdCOrwxt+iWVTMUxlOv7FRK/0U6LqGZncg9p+s0Hec1AznUeN
8SRwY/cbrNOSHdGIec+Z6Ehjaww9rBIf4xy9eJcul/g7LzV23kq7KTEUu7K21SdL/Ekpmb+Bq0mM
NMQu9W90lP/RSKFK9TkKUPUupJkcw2S6UqBO2tQxSK7IEth6iAFMXfFDSEQYRfMRaj+bcFgc1nly
5LuudbbLuuCCGDrRn92ezbtYdqLL+tez+PY7yxi1KH10K1rqrzARLHX2tw6Dj04MJma6jWs0Ts8Q
zoTxOQiUdFhvQYXdaiWvNE8gr82jMENWJygu/jcJNht5OwkUSML7Y5/RCP0OUoDdn0Rs65rtsZHT
vtxPlkK3tjUdB54duUBqgILxHh1w3rY+qWHbfR1oT/qHBTZ1qQ3FfXzvSWEd4kuIgk+l7mBA/R9C
dygA9JFH1HFJf0qiVAbbc4akQB5wiDS5drDfXKMADkkxDzJq22ZamW7mHgCMlPXGVrFnqD7pASU7
knd/ZU5EK2D0F94ZOplpG8mCcjm1m3KNAhLV4m82lxei2oL7aorfT77w6qf83t08wHmW9FLYEcpD
eUzM4geowCZzbJWjs6dVCLlfyGyq77mfEUkj0Du6f/4gcXoAEUV2oMLk57HomjCKZM46NAh5GGX0
/SCR6TX2M5qe2RUrZxIqE3puvMr+zxUAJzMjSBKsNa5WZZEfILYAGHojqayD67r85xfBfQ+nF5Nc
kPCoYGA0E+cta+jlk8EqF3JaWFgd/eCqNiqpl/MWIWUAE8L4phTNQpXLUjv9rw1DNvSNaGyQCKcU
xpMdFr0Xen3SZ2AAtKNFqllvN7Wyv57a8xBqLDgaqSgzSH+hpPZ19lDvGe46e5Hk+HJDWkfN/l7Y
aLbunhS9i+pwpZBGzEVTJ1383NTRTpsZuKFMa2I1kfPHC62NyJ1bdCJQNI9irmTTDNrUxrGcnT9I
+xb+f5xuboZK1m7Ot6v8nrSBShXW/5SsiVBD4XjAtSD6KLo7fxY+ETibOevESO00+mMa7Bq8FIPW
qaM9nA2yI8rYVICi7rw+KK8yDImtHq64j0ViHtFrxLjb7b8+5rmog6tun2XfuXfk8UbYhwXYYxui
gzRnsUmm4Jxa2DOjnjbAIA2fH8GUZlIuneYE0dL3InZOkUQw4PmlV+XXXXC95f5+ImQnlfEgKUOL
eVv5TiAwzeAfFFP6JTuOHPVFGK/fGAwU/48AKm6LgQkp4y/YikQxSBUIIUpzkgW5WJ6CzuPWRMNE
YGWDsts1EXq01Jv26rLkTN/Sy8xCIIDlxsqGs64AqgZ326fa0Tk3u9OgeFAOnYxevXOKYQ9E1ORc
cz6m9JLpqn7UR/E4iE7HsFQWa08Zzywj0s0UHD+jWT/J2b7e6umSj0r1h/qL6fH7iCS7xXFc3PtA
qRBIquaeJ668Rd/4ywTG3c45KrZGbpQ6Hpmhmx1WFl7vqBKf0W9VcA+pYwrP/f/40xF/Cl1i82yG
eAvGOz61GhMRAVspRxlwdDuugCIidSy4pgJ5qQ2mH+YYo8yFG5C5l09fo2nYVS051blACe+6oyEW
kw3B4Bn+XkgQakAIFshNXI+DaREtdUU9uVFUCUAF3/z/N0P6JZcaFwIe8WAHCQOvlvF4LzGqGL0L
LLeBCZR832YOwJM4HdGJYAtsVcBPk11AFSUfjyM2FXIpLOSInXYcsPp7W4MYgzmjrI7+u5L9vMha
Y2sAK2UxVv3vvdogkb3NHIF5FsAG/0NXo3O13D0olk2qRWrbgIunRe6L69eWnpTP49DWVIFIPCy5
dID5fCuYE5rWmOTxvMG0IbtM24K2pYf+o8HN/2bmJXg5Y4Ve7CvKvytYnLmFr9TiKFiYCvZAyJIh
lHXC19qrFBINh3Q1KtLkcLfkWFFA/SnlE/rEv8y1WSsYk+TD8CldDfiuwuFsVBRmzm9fzBJQJos+
OdNX5cpUgCQBYEUJBmy0g/1q2DVy79m5+9qMFIHVPn+EdeQu/fb4ZH3Wnjn0oEdUBjM3JBtPgZu/
1dLwVW0Au7+OJnyD/nQUzC7/Esc3RVzrKx8Yzi75qlyxWEPBg1s0nzlajf+DcMWgpmav0JGaZU/o
xDCMzsHHoS28FvBlL8TN7qqQvaP7YeszZ6bdu74HZU6Ztj+0ae8Vurc8A4HJpvxKV4lmETRlRk9B
vSb4KheuzuQA/FsN9jqNmihxeLYjTLoQRo80sM8OueCpZMdmZqKdNIuXdTDN/TkrSgr0E4iMO6nT
oEQ5TOL0QEmD0G+z8/7U8u8mZv9T1hMhKYmvBcYECPj83opB0zdi9i3Hw8VvMEWBWHFxzkL7JeoP
rTWJQxu6tJmfpuBpAYbUtjvDbHyAds7uczNZsvu1G9CHtger4oiJzvEAR9F+ZBDspZOANbTkWfOz
cj6GPlHtueK65ehkLYXT0JJXNrWcspeAzQoZy7UG8irOyBhOfDwF3jH6JlhDhxu+Bo8uTTKRYS+X
7ACo7z4zSEhVGsQzromzitObgFcJazsWRTDpvu8hdMyygIVPndp7h44bB8FjGF2VLrGOYjwR1kKe
ilqbrOSFr9/Gx0hVKVUk0nMLfSwarUfxR7589VSt5LNDy6QJgRrWZKEspGkOrbK0OgJCbRQSs3iI
TY+7GysYFOSWIOpC3H2jh6Qs9ZtHyCK5GmmftUQnH5DmNdvRFcL8qdkXTJlt0h8WB9tHn3WKU6P+
7SlLXFXvZa3E337VPAeu+2ifckcKMsFWWz80rylyOdWoTn/HRlphfceL3p4ppCo3+MlTVZ3R3Ys3
z/JUeSgsz+Sp9903seTwSnvC+mMNgX/mYBOjNC02Odvcq1IGw/HRH6w7rtBQF6/QuE7IWiZfE+rl
SayB5bwIQ4u2fsOLWRul3SZlWP0Fy6a8QzfPeHfWTOvnZ5bM2DFxIJc88FC+BTS2nO1JPXzmg1rk
ChXwcs63fhewsC7vmpUn00mkFtgQ6I/5FKFtFuprINYaUDyimpMnh3ZR7H+e/cTEi5AcM9M/WHxG
aL610vv43Jfd/JFJOkibWONn3nD015XFoB+ICnl/VtKUskjFwfR4ekJ7CfTLazp8NUzLfUa8E8QQ
8gr6V1uIWvwf1BRlwb65wf2ZCFLDM48cxvvyjWQgn8vUysYjEv6yNj8z9x42GpT7TTrS+B2SmaOM
4HRn2FqPp9ijD6uEqnVxoLhle2G3JDmcTRgb8e+XhNArp417gKnz+2/JOoPSnvk0h3fJ9nuIZ5r0
YeCkGQ6wEUdStlJ8qH8FiRYZM8m0ECgxHMNH9AAcYYsqwZrFuoZ3RyHUtZNdt3Rk0x9zfivbI7/+
5PVplG0DJPPP8rt7ns+ENCPXs6Rr2knuAcsnF3F74qBaGMkTeGhQ8vH0t/OTNPyDDS2ghDrbandA
tYA9xWGYOpshXdCNneWalQ0XrX2qt1MU2EWATvHc4YuHhQn3D2joDmSBEPDf8itv2o6o3aXfo5Lc
oNiDGm34G34SVchMURkB11zzRSBf1nkh4PaD9CQ2+HIrubHHUW+vJipxI4oV5n4DfCgH50aeAbA9
7i+OwlOsnyFbKvFxBw58udc6g5vNjG92iT7bpNLmisyLQdwjAKlZdDEPAk4c1QcVr5iwiSNJAfsX
Em8bH6pUAsB2PPj4oEM5nUWLwJszS31/afhCxgXii7h8vNiqcnQJoDex6jncojkqGTx5UpYIWMNy
lfFvI+K1UurKqOC9faj3FFW6cQ5OhcW9t4f2JCIMxiH9VI/OvX2xEUoxO65lDqVD0C5PG751qH2z
u1ZoJ0fNzbl0s/qTwhdo8i4r63YFb+EIX1nVxteFzba8Zi5nun5fFQkwL5xIPNHgPe6nyh3HXViG
4+5X+vmrxWdQsfsPyh4QB2DDOLk88v6WvN2D0p7dC/jRjG6DXcNeD9XOU9qCO8Ez0YGkm1+/aCGd
lGhLdpAOhUTyhUTa6B0y6akerxIKjlXD7QYr+38jnkGJ8OUi532SrKOKWCylC+XelxQLFT9+Nz6h
GhNjcCUBeXmXhEjb4v+pHSaXHJ3KzAhin5NBzn+fwhpj53YSqOT51lqaBrqMEB58RhBhhRHE+HYd
u0AxILAW/7AZBA9//G2Es0qdMx7p8k2Sut+jjVXXQzg1WXi/OKIqJG5GrPKm4ULsSKCgzC/W5TCe
ByPraf+SJw76vRGhnJ11uh0KJvjLisjIGbswVP5Sd8yRf9uv6u5nkdP/2d9ntfjF+xSYIuWpMKya
ybmJqVPxVtDX9JoFoWsVrIvHvkbW++UnRqh13xDxyx4YsNtwazYnScTAY6OtAPWp+RyZaXxq4wOC
dLq7Jpdx83mcacDIun8kBqXZfCvjBlzcQj5I4BCIwYHfUBjH6QpNh7fs3RsPPODQQd+8Y5Y4vSo7
KMdrSZMq9q23euqjUlSbVEp46dZtWV0wQ0xt1ofx94UAzE9aZLntYHeuWg8TyrSSNPMrtv4ah9AT
FVljr5UYNnApKAKW406gURqw3g8VOD475RGkgvpzKJbxv3tmNygf3XQwRBQQELFHDJklJWg+h+mw
7nsM6ydmq9nojoApR0FWINryE9Ruy6fY7hQRZKaX6w4srRTAsP/PpYOZSncZ5aGkRlwFAYVEkJUO
ckgjqxFMBcnaARCdP4jvv+dPtRMp/tD5kEG20v7PchXpstj0dsGyn593edkfZbh+Fk5C3j1n7LTX
ZCWS7yLfnWbCCfOEdNCyx31Pz2QD6/qaW/3ygaRPaGimafCXUlmmxSmm6kqb/Lo7RT8gjTkAr5MT
4+aqvReBsgZROSuM/fYDNug/ga2ViLwNUNQND6BLVkoInCbCa59hbhjLHZSi7zWuL/9txGjotbA/
8Oaw5hCG+7WoQi55onC18eNDKuwmP6jgRnRojFBmRmfHm8qNeUJ428Jilpntanz99ZO0GZSY3GsW
zELferqmkt7QLAX3vRBQmvGL41ahzKMnMymsZ2S0ka6IlRFbdhqGSveUpmxP0XLRzDDQMSI3TzVp
XlqhB6In1Dka0MbBnAPwwiyH9403Mqos5ai6FNZR5xFx6a9brRioap/pxlKzzLmr50H+VE0SNBvW
IpDhB2zShOQOHlvnI2t22xZ7v8clMr/Q4rLTJ7W6PvWuicGdEoOQRMRgs9Sfau8U40JIXISeMAUX
c5IS8RsAlLv/db+2ORVcIxXPqlZ1BebSZXZM+vt4s6481aozgtbYeao8SBvZvsgZIMVNMVXWtcRY
V2J4GiKq75AHuC7czi2QJ/KyQTYoqjeP007whFR4ih49xRbNHtkPDKr4Av2XEGC3gzH1YwxqbpJ4
6jpukRxDipU/lODedAL/ZoHWqsI/Xbk9rYIhLjfiLX58XUuC4v+uxjUD+6Yh+e77nKY2dFBrhsnO
AWBOjBPT9NV1JrFnVK1/XgHxmplw+k0KYH2NOiGFiRXaOejcWK9rnX3IvMaqGX6V+5sG3z9EoqPC
oQHI4n78tb+fje6aVCm907dQjtOEYxhhsofadv9x5kEDdPagvvTaiiRbhJ9RDrrWRCkr+NGnTg4B
LnnPcnsEEJhQF8rJ+QTOWyiq2GHVN6pHxRfgaQw3goibnz6TfNleWk+/9CaglasBvkp+4DqDZ5yn
Ds4mog+nFIF8JwqKLWzsaCbWKuF4RCgnAy4vk4lvWy0pYXurQMjipT6vEBw/ekeEbm+gPx3caV8g
e7SNxoauWTrh+erD4QT8vJP5gxUa0Q05dPkBLXwbZyjPhHtcc5FcOPjyywy5tuuMG83K7/Ghl++V
masMl70AS8Sxq8/OfZ5KM6z6uPWfeJURN+RqbW5LM5+dMxmknIO2btn/VEXUo73yaM4mazSQiCXc
6hO3ab2PfhtqJf24Ua8rx51KtpQwKaUmZ6EtNjpEs0Dz/PUCcOOO0VBK6B2YC2GZhxxHl5mZdPgL
ivXyl0AwRLSq0ogdFBA11NnPuVuvJy17HapRN3LBfdvQrKPTpaGOYe+72+PnykdKNBXuARAlJNGW
BCBErWOei14fMato1avz2jTBZ23xxzVzJUDiRrWZOl2cISqGXM9oRaRhI+N3KcGV07EXmVpy31DE
6vJPSnk+GdGRnuAQpa2x0bo4ylGIw5WToPF0McbszNqufUnR9Qd3isFD0J2SR6yusQizXNOrBeYd
e9pTJ712WDUvfnWa16s5Uo4Q5FF5hBPMpgD/E5NFPPyXx0xCjrGCJBnFfS5XNP59HFHrvEvVhHhV
LtdSSuBnMvRvCNhUgNqTAX0BbeTNIj54uYhYiZs99f2OD+3DwpKaxHMqkg2dUGAK9PthjauoCtmj
25ZTDnBpbQNqoFiu3Ot/PXMMQZaCT0POHjoxqefxhzmRnrEutmLja34hVe8vvrfeaNNiZVHjMYPi
rAChdGWOcTC7TXDaxcjvBQBTwG9g+zn7kUxRtXC6RRcDJrH3mT8yLgQSn0I0PqMJfSncaZXuuvP8
2+MWMeD0IKzoYo/X4aGrTOVy6QxjrL+GowAgPmSaHwqean/yEDLVhW8SKuUQ2A3I59mPMea3+SrC
D9PgclpnWMzWE5XXaLkXFWhTLtNdiHjtLgY9hF4kt6DMBCgFHF0CCkluq3IvMus9P1LM+aLb3nkS
GT56cNxLkNAjHX3U2gpMlHwmAn9k3BkCItnNw1Y2LaKWpPAbzrp3CJPVhhMknktgbEqbnozq4Tw2
lZDhO8OLmokQyJgHcQd22v6mHDybykp5ZIJdO8YUpRyS5BejJ490T1VMN3q/UMJTnM0tJOMSXgFt
UDa4sZnB5sjV5haxlUPa5CoSMdnJ/Q/xsdPAUonGwI2azRkTe/E9ld8ngZnlBP4Fi3CHLeb7NJHT
Tj2/ex7A2IiHyanCghxgGnC+f8G6C0tHX+O5Jj/SAelXDJPAKCXVk3CpKtKWYcOIAqNABPA2j7aw
3pYnvxYb3/pHs2Zsyuc1RPQwjisShZy7pgddjJwFjnAVEKmL6DDM5qR3hXC0AWAXj3R59X98a++H
ppRd3Wdju7mcxQ7BDZ5D9mCESO3Jk1IY6k9exvpn0d5N/j7aNFzcx4ZSzt1kJoyySRZfgLUM18jo
OTgyKLF+ordcVL3XluakUEcO8UQ5CUtFdZc8uTOuYQdBfN/Rj9In8YXv2r9tXS0bEiU9Bwic+3D+
ZLiHRkhv+uhDO8n3/Cgdge+hJh6utCgoVE8rct1HHyc0LXdM98XkX91Ov7wdHd+cPT5xw5goe3Lw
ILFcQ4uMKK3zfxXHyRlnfPo/nHVZRBbOI+dQYA6bnscV2aSu/awEzOFsLpXzmh4SkrwwOPm302UC
B3QIg/6CVtkzNsslFJmC4bsR2jvL3IrCiBEPgxqitewv1tkDi6MPbBdd97DwLOl6Fdq2YnUdxBoG
wi9eottiq4XE2pwRDjd4EIWBMW/F3yaU4BshOooSh/TRgiMc56AAT16NVuRFEGM8Pzlr2LgMgs2U
JQjEmxLo626dm5jlveysOpdT+pJ13dwH+vzdxQ/DDgqUPMax/IUJUtBGWR4tDmzzqnXBg3Q203fQ
Iba/g5D23D82dwpopPlu4O+2KVSVzWTGPr/ydZfHqN1gBhCARirSsarzLUP4FJzBTtU9GYYTXGcI
xj933van5TWa68agsx1+4c/9XIawa9MQ/TFPBQum4HeFP1L/0MdDcSgthNu3/7xCDxQmfDlshcU0
NDO/s9gSunqRMkRl9m8vj8RQYNUUK9Jpk36NdPoQIh+3aHgh+j+PUY1NZ8lRdwt5qnUAPbvIFuYp
Ql8gKm29UJfKePWsihDSMiVh8YPN1MnjHamR8D8RRTPtTtNYD/2kWTdhMqEWGZq5fJoESi2jSNdT
Qw/z8IDefOEa2s6fSMYn9/CtxpSy+Cl7qSWx/AVPuTWNfaRIno4bQIXikMPzCd7QGW8o2IE9Frig
/3cgDH+poftXqwg+ig9YpwZDJXBs4YDOCv7S6GoRF1T61XFp3u/s+77GUKPLM2MLkfPcg8jaRxOo
CCjoOFnbK0x+nY9uOdGAtw7VSKIdGyLkJ/M1BYxnMD6Abb7K+qWOnVmFi3ztCIx+99uM0OFAZj1Z
cSTtNiWLtIivDnGkcH9eSGYyua7SCJ7pYS4bqr4Jpl7BPqNX4OgLLIwwF1jAQuz6BxqN+t8Sk4qG
gz9+/ZfxMYprFfkXU33jo3mr+K2vTB4AqMnnwXxVBDCebYNG/H6voGZZYQDPnYE3CGZealasC4M2
jPsZ6SKA3H6dZaZm2TNCu5RQ2HUqDHe3zJpkDeL4z779Ii6LLn/TN3Lz1OIXNq6QZbLHDhHK+RL6
UK/Zlc6hTcthnCemLwi0uIxxcXmUGimE+RzkzBDC7GizNtK0kssgAqkgRIuKuWC4DYzRScgtGbxz
LJ638nMREfme/WJlAZbitNDC4mZAKk0MFZpUocTlDBDdddwERtZAF4dhP9Lg7etkQvrkJi3NN+ze
aszEBsD8R9DV/QLZmlJh/BAJVFNoqDePG4Dt6fCst9IaamU71UTw74lbTYbS9qLNx6nsdwUV/6Op
sFPd19ZIjllHoq/zr+y/KYNO7BC1u1RQWa3QzYIcO8kl41ksi1xospSyS/jlAe1g/+eTR+a8UGZk
wPBdcWzBrqvpUwpFZMLm2DclrUirkZhPZtiHEmgKu3M10p50JQvav3u8hqVW+Gesv3noR8hvoqxD
n3nnHahfbuXxIOwxxpM+iXbHo9s2JdVzEY0/LY8J3JzyVVFtYbvYtGYZoQtGEHZsfj1Gz01MxYSa
xpqfd8oeAuNOwE1A8YtQ898dMPwk1mUaOeSW701klyqF/IXqalLaZOQoI2Eq0dgjE8H5SajQFi+Y
zt3+wOzwDwwUZ1AzUc4qMUU3KSvaAjcXae1eXy4ZwrdWuMsUnApskDMppdopYNEBKQ6Ox/A3UEIb
LOWSlGsRsb8ya/5BdbRnNMB6TL8agp8NWOk5WAg6MV2VwIoZqE6g3GPOatgjZ12JGXnOq5Dbb+Yf
iMRy6ekrw71N9q4sm8Fip8UKukPPo6ImmGqjTCp+byyzKsU2w8+7b5xmgFByV8VIM6HLdKuNBDir
18CpEV0k2QUghRuzG05JMsf1E2SiSAcNBqk/AJR2/r7gVGcKviAF39rqmPfLGSXKjtdy4DonCxYA
exM32DAxwPwlrPRccjyNFc4v/zcfGrsh6p0EfeGUa7UFXIgJ1aBbQ9dIkDNn+GegiULPvnhLWhL2
PKGTxid1quCRvh1lOGjaOKXe0vi4oXaN42TfJEdma+ORbufKJqpM3/ZWyy+d/gMTmnx4E6H5uNAe
2qjOqGSiSMveQYCoSRBtp3rppQ8YbfYe6B16VE0YffoI2s1HBusq+Lk4jOcnrhZ/ZlSzcxop2znP
EnXtSL8XRPHQzTC041EplnIdtdgx8buiFqzgTKsbxGfpQ3hXBdeGXrJkfeakaQN4doFz36APDqvK
rWIfYT0P8LpXxfpmvqOPCU4oIKTOkjCcMJGNLyYwVIxxe+Onp1iENv3EdgZuRgzdrTOICupf6lfs
ztNcY4s3tnT88FB9btJggOGcf12f7mUpc9X/DLiGTyiUwtK8e3BaDGgVbz+Wx4JR0Gfvz/3mK24j
UNGJDezW/WZIdRRWY7rDoEw5RZxJkvziW3gJXeatFMSZ0lOh4GoN9YEOh0TU1L10Zd01X2eUJ0SN
ArrZ8b6I2W+fdO1HjgAuap7wTcV3ckZfIXNmKDnc1o5HuKKkNPya5HDJrU0NEVSPbpDXJ+1EPrMD
UK2CIq8iWaEVMdvaarnQPhHqwLiocrc1cYReMcW5g2WZGNsmxN2e+OlpZVv3421s18wZnhUspWm3
kp9yHgoV5bb4MsocsbfxD6h+MkcC6wgue3aESsYDdACnNz9xHG6sDWlUViGfbcV5RfpZnv5AEthM
YfHPE+J7GesSEvRzH+rTz4OPmGQvy6nL5ZrglzRU/EnhuO2U/IBSlzN+WjfWQ50Jdc2/PuFcr0NX
c1b3VGLCVkxhPEUP36LMmZnzVROVrOJ8ArLU1m64iaIlqgho0PUh6lzQnvFfLBU/FKNn7mKiAg4F
O48h5SRub5mLbmEqeoxD2K43J5CYwBwPamDvvm0f26hNfafj4pmVJy1Y8x9rh/ex+nDH/Q0LoL8y
QyFURPkqRALSE+wy8GRiIRyp1N69TyyLFgBvGQX1G2/p+KQVvzHirnxxzBkTjeHriAlOUsDzJjpn
85LMRtpNjSysBUwDgyiIcbmEB5IeiHx7buwChrsor/5XOuBa5qeAdmkLd9JOPw0FBB75CnXLXPs4
OEfsJpY52S4LWu55zBjLCRed83Ixelv3djGxMIlLPhAVujhltzaqV6J+edeU8IaXBiWZASQbMKdv
qbfLdRYocldYThKuhTlwEmRoXM86kpbvqMXUqMfzl496LclhtnBMOZiVJKlrkcdFJ3Nw+7cmTA+T
bDBsi8wuff+Ev4/ZLhIb1fg8cSCo0a+pprPnoN7SyrnwOtpPUOrS7C/FlLhQVgNAo4aUEFK1xhd+
DSS3ZMYFmvfUcyLsF0pGA4tCI/wxosPs/A2IVKKSCvm/1N8d1yiuQmvISjCWerM6WtK9y/DFZUZZ
vm8LuaPAmT238NPou/Lf5uuODWwzWl5omR7fc6nGpJNN+2H05+GJTgwB6LbhvGchCmBQGunWCImG
x5G02qzlUIBLBGfkqZWW2hRJsPb4IbCnwIwEDmHQzm/yKUgCq6TBLlFQgM1KcilmOy/w4HehkWpH
aYoty8htYpDWdvssKvbma7kop2MkMsoNuiOEmQH8qJIZHPEl8ytr05TqABG5LifKOQFxjxxyK6bQ
z8c2LYiEdFs3iVKLAJDaxAEjf0k4tR4RNSclxTfxbRX0ra4mLIkFSE2Esc9h91s8XS8JpcxyNrsD
eOk4cfMEadZRZpSZA+If6RKjo1t4N2wmxFPf23sDZyO+XM2aJrydvm3iSgj/x8uDdRWft6QGMyFs
uwDw68AZ5DHlMmUxj6WQ6j2/jRpVKfIaL0+YpW7xWLIeFJGL8FY3jolIuzdYk6fN9kuP02RroBqR
GFGmJHPbSL3zmS3vhNvUY2conuMlzr/C15mjWjIte68pnltafTRA6RnhmeUhVurrP/fKIy2ooiAR
1fmnyN3fVh/wwxxzhlU9AkCTiPbyZIYqzyFBAnH2GQGrx4Wakaa6V1NY/TpCJPLbUVliJbaj20/9
vTqb27yVYgte4oKu6edcF/5Qvf1KHucCK8nMIyz6EUhDZT5RtyYz2RIBRyk0pSR/doAr6cg2FeW9
oVpBLbBE9GJzA7F5AAMlrB0WPMaK7QmpF+i2BtSZKV4ziduhWHP+oOGmiO0BDsr9ZqaW3EWv6z4x
4PiXu9CgwBn1nnRQBybdO3+mFeG82x0LjIQdVRtkBypgnczuDM2NijtWoKvcIh4dB5GVb6yHUovy
u357FGSZX1g1ffzKyNVBu2T70TmNiGO2PI61Jgt2PYKzCRrqi6+E3Eqw+VJ191OQnnZpmJdfZjR7
SgLAJ1ZrqflKDbEnNiSdNU9OVSxMtHBqYxs/fBT4XN+PW+RYThLcX2ndGskofUEKFfa4rHarPwzI
yx6QvvQ7Uv//mnenFFu6FRAH+jdvWyMdkw3jgpBc+L+7b/nnhk+WPQlovUoqeq4LkGc+wFjm+/SH
cn+RNGkGHOM8gvz1PTf7akepthy0cRGCWM8tCpaFhPNg0jKiGGdkHT21hOuLqt4t01X9zeSefvVR
Fe2NItumyCnty29CNJKodwdCwc6EsOrIQghmhvizdA72AlJ31tNabLnVd/5hJS69BJkyWSxaoI0B
4TAIXgLdf5N9kyJsrXMWjaO4HbzXU9O0UaEq2TLnTJ8c/nlyeLqhBm+59z15tBllZlPxujfFxSkY
9Ifw+CB+be22nY/872DD9VChGz/qcxnxfzjwLRdUIgUdKwA7CNYi7ZPypeolD/mLT+dO7XYkduym
s4+YsHu6QdItBI6BaGGd5fmr6DQom1aJlSKy0CjlKb4DVBFMQ4YG9l6V+5iRT/Lm0cEe+1ZbBmV3
8nJV+uxEBD5rQSWrUskIJqjFGgD+4+tf2bSnIXxS0VNaFaUSXjDcW3EIgzMulL9PGFw+w28iGDia
6peL3pOAW6xbaqUzhmsdmIh1efZoC12Kqe+R1yttEvNvkUyFBJFnGTvXDvUk7SXKHzR2dNMY5+gc
CN//SIFJQM93254s/GwFXT58oG0SKd81gIXevxG+CnpejBVCcbGNXN7t+XFnjztWreyuk/nm82QF
KLjRx99/EAFXR4cxBY47+61koNrN/zoRnFc+KOAdbtRutZC+Sc2cGxGaEQillqYJfLTdCh33glFX
Da4WXdB2mxnsRPmhyQuxg0Lw4o8RXwVytjxsr1LhR+JMNSVHLxatlKAXNYK8XKycKGc95eJ6qCMp
fAe1KvCSf+v/7eyKfi2NdHWoxvzZWRJITETS9r6CQidEtyG1vStTaJ0HOOREsUfliINrLXrkRiza
v1UaY5jLqepOPEA51QDanxNGPCX3WD/nqNYVflfKKhyVi8+V1FezuDtE9nNg+1Mr4QmPahvH07BB
qtVPn0iuRA3Q2HZ95emn3Ik3bgSm8wxSpmY1TCnctF2wgbo+8d3XCCl9HQ8Gxn9Z+FYDTAM3yPXi
Yqg4AVd9WvGeN3dHwp7abA3IdJtFu9/yMlF/hTywkh+GpN0XScmS5mKQooCW35V6RjxkClmMHh+Z
y+FLkS98pB3ej20/+AxUSix4rEGa2Q1U+RUXQwkHAj+3mq/BXE/7m8NxXPimZE/DLIDe7UuNCeRg
LWg2Bm0gH0I7I7WfB79m9RlefEk9HuoBHIz02kXioIvYXYodQcgJWfVkmUtul6Hbp4JCydtw4rVs
9tLrt1VYhvNdFiRzXFtlhuOv2GI1DtiO29tOIK7PabGMB8lpgWZxpOZODAB4KM2AkwlYH6RHR98t
Pvo8X0HtcmefhjLGFz4tbrlNlbCeznOMxp7fEwmFcN7Kf/saW1Bp7eYbjPINNtWDBi3bAzrGWeJJ
CjAd75rQINRdlKKzKgOFuMBt6v/WpMS9pbp7NAmll4vJZLggEFWsDqEC85mYpNYN2b++Q6sRL1o3
qw4/ZIEMKD2jXZnbnSpW4T6YrZWeTbFDiqtjqPiO1csjfOJKL/5RE84ECiji6CQWFLXRXnB9vTbc
Y+V1O+Y10tFvJdk8d50Or9j74+uv0zQiGrIqEsLWXxeqQ7UnFtY0ch1NhyVMPEqUk4B72Czf6FDd
rkJWhJTskmZtoF4td5mP+Y62KUU2mSsMDZ/EoTVx4sKBSwHuAbFDstNvVfTqbk5+XTE1EpEpZ2lU
RJJtW8j+ouDcj6rcg4t+BM7cVZrlPauXcf1zP2w0rmR565yf5/p+dMEx1PRVnBD860//7HdvAnE4
J1YNXE1dCTrvmdZlZKBLgp9mnK64dlPxcuirPl4m4qq+FnyUil1B7jGLrixKiPz7mEnYoPw4Cgu8
sIPWqoO79jKNX9kTVcYwXe7q53QFOQPhpq/fXTl1YTvuFwoRK8sVdc7xZItEoRrQr2T2GxJd4egt
rUpFdcphw592eSHqGx9oMuBti0rOIIiGgID2svvjv8m8hewF0TWSy/5P6oVKBJ8Nh9F8eYlncGXc
m2FvRkYXMx+AN+ZaU5K8Tt7Gy6xhd8LjG52yfFo/xgGa0DfyxmBC7ewlV/sCSeCC8nGLzcM7e5HX
AN84tyGxHwhk9VclNzWPsFzGPxgJFH0PIJVeXOFLAbDycBwFlwW1g4mlUv09PiL4T0pqBGPH6s8T
ntfeDdp8yzWWe/xZU+YNLryV+fDCX59ZjBSIkki6SFNFO5ofkDZYJUIk2auKKDwQEPlgdM9uuYHy
jNJP/pZrwuu5XVG0I521umj8jFgX3tskYU5fnl4JBRpxqpCdOT1MocchPZGK14J/gXOfwrXtsO2k
jCEySfnueo4HJtUCThRqwx0DxjswT19IB+MACgu4KwNoId+ZJm9nom89D7yQd4S3H4E9pZw++4zo
ZalLa6QxL6PmgWWnDndacxKfmbmflxirdr7twaS8g36zpA+P82VLnH6PhZ2HrNTw1npF7aGDBgXi
37Hdz+dpySAMePlfCzNywh36GWuS5R+0KYHUCXJK7Lglb1tuJgwWjVuIEF8TdwL6+X+LeMG5AiaG
GwTx+6OQOjgizQf9GGdCxN1eu3KIMro+/bqDB8zUJwZIZgFHP+G3VE0t9Kc6MoMKRvfEV7nzxUFn
CyfbzSvJd2dKUP1V8Yb+he0HDhFNfXOkPKEOuz3dIJ8JX8jCepD7sNdJKwfkTgvKxowi7rt1+Ylg
ZAXrky1xhf4OZJ+TSMZ2k9nIPEfSNfIWAQh0nRnnea8SKKIRmprqrcTjFniKq0wzNMPnSYZTIsZi
F+ehyMcUBapVuqwbRJh5TxUXC/j/xQLkQ90BBCp6m7C6tmZSP8CQMnYUPvphRlNOmn2GsnCeSHdp
dB4y2YDFqwwlXaU94hTsatI6+fIJA4xf7YAyshtbFcro/KnABuG4vTIwqZ12GZYW3BjFOYs0hD93
k6lxv/Ykcs4S5DrSYm1f0X4OIPY34cH+ntu4UU7JQSSRZ0yrAwPg5NFOQPIK7HGGV21MfYZcQ60c
weEezEJskuyQB8Erf5VIds4/oFg9OzWiz3fgjkO3AMFwMlVtZ4ztWkWyssFuW7RBdL6HWfYdhVhv
F8vtsn/WYsFkMPWAUg5VLKkwHkwgMEADeaS5KIyXX0mecvVx+QVKUxD+0KdXvfRR7i5qho6edCH7
caSXDVdH7VsMx5kE1yNcxoEt2yHwMQeg8UREBKHoYVtKevzjhZSZz0XIL09go8zB/CXe+SDeB+sQ
8VoxP01U4KPUhpZbE3wHUB/DWx6goy98OJyCffmBBTucrbk7z1bkVmZ16eZI1GnXGXIzOj9f3y/v
ssfcnAVC5Gmc9GnrCY/nkR70FOiw2oK68VJz/KVbToSA5bMxT7mT5vEJqyoLgqV7THVIZZX3hQUw
HH8mt8Wh+diMvCUqX/4e0E/XvEkAtCjUEVWxA+JPpnQqrKs/w+O+raaG3NsY7RALWvrXSrIB8M1M
2oSkBiA7Ih85M71WoPc8dA320QKlI3hbleoQDM1QenenpSGkvC4//ye0OxwgRKOoi1Bui7J6gTSL
al2Ak+9eKMWkHy7ZGvV9xrzNQ7yQIibMkmKnQ39ToyE7PSZJkIaH5iNNYC1zI14AFe2lruBI7w7L
qCr0vftSG0asV4Np3Ay16BAzOTsaKRBcUow2JyEZEwbJ1FTeCRNxh+034ehibvm3UT65B0/Opg/W
x2+iaIZInPOmbbo7KMhOpz0Tzty8bWXijvp9LEAiMwS1rbF2LOzeyjCV2o1i2C0eUxez53rPKjL7
u1wFCrqC5vtX+asTolLkrKm1NBcUdRBzfidj8itaDSnbmu7yNDb52bb1MiHscKmj7JU5rEa7bMYH
pFvKpJV52jPI/m88YJ+GhA7+OSBqSw2qLszsWogHe1yRgCp2yU5gtzqRth1O/wp7DgLQlB5U8xJN
QFr5CTIxhB7N/gA77tWUgPdZ7J8Q0v2AasL4w5XjztCeQA8nIBVkskKH63py0at+aDyunnpGzpi7
MnPseGEYeu7snSzoOjPut0xybAoipBlxcwzHhdwQLH6sHkNsJwzK/5N0yp3GMJ+x71XtUPuJDsrc
f9lL3bIDxZWKAkN0yH982f54kMPYoN1piIJOh6+R8FomLcq5pKa2SEIrAP8dk2RIXTbPNAq8gsAJ
DuHVsFeodEAOscrHxKVzs+Cq/lH6sLhEavix4e/0jXV66/o5ik/l/3VCK4y99Ur8pLQyxP0gJ542
vkJBBB6OfM8PN/x9npn+pm193GIYvb16oyezcFf38L0HYM5icHpsW1AxvPClt0WM34eY9c1dlp03
8VfA4jUC4Nc1sWOR+NE3GTT//zAN2ywuROFxW/Ru713qvsCtg7ZpkdsJOa4LqNv060zHVixh+i+P
xpS3dweUTYAjLjZY6ho15vtGQfxVg4gwW05EWONKf5G/TnvwCJna3SWU0Ykn7Fe45zp46FlVaX1E
MMK2aSAdrKVVCbFrGRnzAyIfDvJocDeFS3INLdjdVGbjtjRjSgJWsJYGmbp8ai9eriSy6XcbG5GD
p2VuwUENbVmPqeYNsKVeyXhapzPMobOZscokWXL4gzqShGzpCw/L3N90GFL2kqddERbSEpoH/Ajh
HpP8xuoXz7mJoWxLDqYcbCcfhLBVhp2L++7yhQjJG3VJb1bRrxkvVf6NGaGZdw55fn4N6JIFE+B3
jKzZxaRzwrkHU3qtx4/z84T7w8RKHJ+Q+LeD3pyNgQAHQoWBsC2plofWdMzFJe+tU/wuaLcWSsBB
0my7NhhbCXRjOBgAjAbONx7Bx9Flu0jaXtlQn74q90DVxzVeKUbZPbYsNDPb7ZbUHmL8T7BlkuRi
pYIHOMZEMTzgzimgsUGg83vep7/7S2q3DA+8ra8tm6nlfPliezAtMMEBlJKsNv9fP1ZwHuDSf/63
eqKtR0GZt63GcdRAZpgG+Ic9lvwg+ZHaa2H2iu2k5zp3OozlzjFDU49xtckl6VGJ/KqvQh/iAsFK
8qRuWjfAT4aPF8TOfoayg8gMkIIp22x+cWc2AD+vcx8hG0vxboCd3UEtZfgcN50IMYN3PdRaCRhO
4V0fBzdQUwjt4CZhxYvQ4b7FChSTs7gw6wyf5u70jRsE8gH3aUg/gzII0088fLztfWco29Zizvub
HRXTZ24Ee6faCgyd6tpi68q7Dw5OMVAVSzmqodHbHP9oOp03eW+94SzzSZDI9owihiAUBkeSJ1WF
D8gO57Kkj0unspWeEyWCCyLdwSFQw7XZr+eNjBOeH8f32ImXNfUBWCMCckDzz64xiUNhCUFV2eBr
Fbs8o9NFcTfJV5IW0ITQL/LBT5hwoT464qTIk0kcGlJdzMlhbOAjJ67CerJJebXbtaBKBNVFe/E4
sqJW+LvqGlVmPtCg9Mbwtia+VhnAgk0lQQeJC32rehLOV5IJ2go5ImGI0IsSY08+Mdf/QIv/qZ+R
XYXNa2q/Ufj8QGSmegJG5S8yIdhRT0E36iE36Z+7FWa25le2+VCf6251n6p/pUvz4ccTKCcDK89q
sPBtoozoN+NVHdHTiLL0MRfmM4KXSh5IBxrucllTDAMlKOnvwtJNzRkN/Tsf38fiuA7oTZBTWZ/C
3iTdwGVIKfBKxFWtsKwgG2fBRoy+78VC7hykvKNv2ZAu+LFVygIjI5vq42mbVpKdBrSf7GRlX2hu
ZLJko5Xz4urAavLyy4jDLRRZu5E+7sGUY9PnvFAuY6NTdNnUT4hsTn5vUiAzPmooVuDEY5vR39Dp
KjLQy6itZzvoO3n3ybF8qSTn7IOc7KUbHECoYZt72RNJ2EC2hrZJ8Klq+nycZKcUF8Pz+B0+513a
meRN5c1W1GegOaUsnBTLeGbuVBzWVklkv/cP8ayvaBsfxTndge4xn7QkXvvNH0OY8l3osvY+/O72
XvlirxlxVYP3zLykCfuApFVZaS8xGU4DehbnDT8eUNGaXyDHhC3hun+V9uYecdo+MFwsDlzN0q1B
+mHsY9JGPEMRLj53pjiPPmC6nmOcRj+CBfDWUsbDp62GTk5bHyjMQLGv7DI5ogBXiXHFixlr9fCl
nN3PveUm7xVUhB6fW3HvZ/4hm4AT+Sb5/lzFYzwcWNlUvY0l4Ri1BX4LGsy7YKpwzGOWrQ41Lix5
C/D8L2LbYM2PIDBsAR/E7kPxBuSkpGapqpaVycNauiN/QfeRBAERxymkp7sg1pMdZDI0NctjDMh6
/dM7wBR7G7VmP5qsaiy4nrwKpj3Cr4XX8IX2hSYs3KlFBAc08mqoS2CFMhyYUX8OZ+DL42Res287
Kji4aqFDvtbUvZDlV4IQ8FgjlHw6UQidCGpYW3VIYqpHJ+P0lAKY2GESUpngrCdi8IoYp8chAp//
2EOI1NgA1PaJtdI7JvbbgJqP5FhBYrbTjOUklBCb3cuydgHoUWCFLrCZTxu70aVrWo2p4yU+B7jb
oaeojiYucbG0FGH4hmV/1Xd0kbuR5xXVz2FQAWsn5MzbAxR++0/TSnACJCDHAyxSGeT3DbYlhJp0
4hAL/WZAoVVLKVvOkEW0DDJ6GcdjT9y1SKWUMgrhd9qB1zG1OhDUcbFfpUPMFGK0kMcQkjyDdxGP
VkkL3FIBQV1+lg/zu+z18e3SOoo6T+OS0M0ywOXJIUOucm/IbZ4WNfWKhXIS8OmN0oSENRmF3GqE
x1ZjTwwnMr3Q4vbuT6K5dEJYx8YZwWf7JzBXy+MwabIo3qDvdpJj90SRRk7XKqsFAvZRWux4i6IH
y+wQVk7Cr+gL7mbbZbDS5sZNibg/ZAcKMmkvxxv4pBxxUfeC6IQoYVbAwzuTDV4RYgUl7wxTIbTZ
/3vFZtU/VoxMHjTST2K+LzLJBWPUd0vs6FhJwMhhOM2q3j/wGj1LEnDkXe0JiCbWBHOa7Q0Sa0Rm
knjbdCWbjUybswvFPmGuAqXuPKwpoVrZNDRWhfTd1clE+nYsIaT080AwUakF0kiLXxP0uzfFtVdz
SPfo7GHLfSbYQmIJi0GLMQqSbmyNZNcqsVAIrwvR7RErkGX+kVz29mSI7xfa9tQLHjuepCZSbvDN
EqHBKTpg4SRz1yhwhxmig6ciPFrf1wxRi86Q2S1kV+KZB1+kcfFf/ntM/JQIAYLxsxyuD46mJ9k/
DBLLQfNb+WbmK5miUXQxQzeVdyJtYMsKHwLGb44XY1oZ+I7K+aHBJEjmK+pvi3XOnezXaa+8wJol
oPv2+Fu4X0Q7tBm4uradgi+HKeRq5E9loLaewjVtmH4Bm1NZMHO7HO6+SYWNI8E+aK0Uoz/iAVnt
QA53ut+J7ULcpdY6TpfQsxen9PHl+ImXbmLQrwTEu8wC9vBtzJx0a10OS3bPCtwDEFJv4J/8gsUd
Uve9yyZoaUFfJu5NKRuflFOGeukSRiTO8RHIyjFDziRGxd8AsCAqS2gQtbl/Tl/HbZ+4elRZSmST
GKwgHg0tBI9fn3uiGoYo9LHwurG6dp6nmYSmWntPtlBWWLETQYKwnKCPqNyz5U6c17b5uBwVe6fO
J410iuTA7HKxGALKeZJg8ezZbUoRk/+umvIuGYQzmATl6QCJp62c3vNys3V+XDONWJ0sr4D60A3/
G6Tsil8TL7PRYLpRFUe8uwEIRyUi7Hp34nB+yJv1GhtNG0dt+u/iQOg+MvLgoFkDKXpMCLKaxK/Z
wBG3pV/ukgYYWbuKcyHcGX9zBraKl3y55dZyUtR+2+BptLyFbV9UoTu+kiRJI0pU0QEs6FfIKy8b
bxOcGvx0m988kgZm5sk7KlSwEO4fqNj/K8IKWxwxUzc5hjCxQI3VEa4Zpgmef37xkrohj1MGpag7
ImirUjxxgqcOE28IR97YPIENB8Cf6h3g0U9Yj7Yn3Xc+WoqsB1uUdKc8dWaV05xn49MJwOuZu5VO
oS/YZLlOy0doMlIMRYTRwiVm1CnPdRXhmXcaq3XS0N32zKEfkbBE7pVl+vniIEy20UKhCGDUp7aI
wp2Np+8AVoC/bUlFjTYK0ahEu20kPnhhoHb15xcZPpJqWK9Am0FIrLnXU4bV2mWTsY7lBBLe4uVf
BkxeTRYa1y2v2tvbY6GiWpLBuHNvn18nawUBSdNgP1CEu+1XDt61lFUV85gQwTLBxu3XLCYbMX3n
/QV7B+C+bBpxjJTSHSJ4t5AO7vWo4+qApOqulH4xUn62JiSNXRpM2+rsxIHRujOSTABfcgGObKcT
paV6Ip1vPwsktAgCpuOgIbX6TPI3utIEJaCsO132409iXvZWDRRnjbl8dsuGY2QUENgtaoSz8Jr6
WTsvlMLbwBR0qjc6I/rbiIAnh/0ZThbyMNocQ9T86L2y85pG4j+/uce4+7oUSasnEJknC1HHtwVw
kkL3iCQZunMPlas489/VVYOBcxnI9zfZzjCh84hu0GoLYi27HDj+V5GhBtvcr2HMYcRk/wTEGhVb
RYFH8yAY4kq7ZP0d7HpZ/hyz+FcPGoZB6wN8D/gQs1qSFbLVTwUYZ5AsvFvmfHYCqomK6lBUAWeU
cEroNjQyO2wCtU1L+Pp+paTAC+h/3Ok3Vp2Rfub91e1Rx0wwUBLnxKv4OPyraLsSomZ8c1nIrAr1
0ZUnjjEWh33mP+AXaHGYxq+wJQfqV6e27/ju3njv1RHr5zkLKg+GwMkh3W/WlYJ4TO/+ojNItiSK
So777TO5x6iSJ6VTD+KT1UMhXfPJeWdYclNkp4u9p9alon9/rBWH3Jq379rjh6JzLxPebj03wGrD
p+VFZ+MPdv1mztGkW0/Kg3ndDGZE3VABhAoHn7cF/1ixpCvB8r0XbPZFOyMssstyY2B2UwumGQId
qAUC8qF97iEeZwMqZEoePCmb4eRKVCzLiXQ0pu99fAocQcGB7CBcEgR9L2BYUB9Kgvf1FWPEZval
UBRWVYmF0HxOSm1HVmYmy7A0sPMZN2K7+4goc1bkIo4woIqwqOK6PfP40dr/f2Solr3nlFtjsbqj
ZRBWzTYxfCySftTUStWFkVLlyzobOo3Yw70R4LiMVe1lbIUEVmKGWVX+XC7SP0GGvYCIoLMpxwOF
dmdeAXvj22TV09RMad97WLxsQe21JILjPTTl02bpUOZVdCo/z+S+1gwkzVMl8pBJ5hx+faOvAlhO
9SJoywbOhaM8BD5kdkKUJeX9jz+cmsCW8TyGgkGdOY8ITRTwIy3nNf2IkPiVlZR707OwfUNXtVvR
K2E1oZ53GGfYcFatQ+G5WMYyk7qChy5hZk6cuIrYj/RsR3XaPUSV71UvRTx4XcLNIpQ1VbzsMWtj
fTMfgKaCxsLacFMok6wkOirRkIouCM44D6aoVi752IndDKcqS8p0Y20yoyR/W8CU7ixz1RTNEjqU
Mp1qx/DThiQzg2f8fH4vxD0prJ0EnMI/iEncegtEaAd/wafHzkjYWGX198USMt3K2h2xezH9cLf3
P4TRQy3md/xCRIKHJlpTL+nXuxaZvd4/OGfyUu4wI0fvDyItKCEOm94lqOOQ4JW4qqkv6wYJFsTS
mfXeCpZle2iIhkBJnwPcfx2dWMi17eaSw03FaU494BfgTpgwyBR6QC0ltlFI3+wL20quD3uidEMs
y8BuTzdvHMpyyWNnA7rfwTVqQu354B/XF/HfDn6GS66k6Jv8GevOSssWhm22kV2A7e26PbId/0JX
YmGhWTqSPuBcysh9T97RpTsLJjHkuSyiTTxs1OUjHKKC5kxJWY3kMlWxmsqdw1q3CyPvqbXnyWDM
HWrDne/i0Ike/jEZD2WKHL/VFzq/O0pGRX95vczHe4EweUY28Xjfdlo4oaGjBrGD4V9yvHzjKszm
2jx/q53rBb8Q2dzt4k34S9L02uG0u+jiy8ASnbb9QYksmmHBAaUiBevfjAhV3e3Al4Rr3Jb5p3zm
2PuB8eF7Z0lvN+hNuoO0u5IiTwWLtw6jhkARJ+cwLGV2ihkFvmqQgC3J8ASZITs3c8lGsOAUKOTq
tmEG6EOZ8JetEe+sxVhcRGkm8JpytiW0WpXgal/GlsR0ZKR1TgLbSbUM9/89eRTMm53sn6eYD3kb
Zkla/xtTa2QSPpGqGq4PMQbE44cM8RC4R+Aj9g2yQu6bM/kGl7mBfnH44wHTCpl3Gp9vPfltGvk7
nlBN7vEjFN8H/lQUfwSbr1jrCwr10VcNnvCHr1Ti5RZ9GkohgLw29CLatmVTGG8SldPjX+sRh2wj
yBppfAlBkVLpGzxAde4ZKvUHzjYDlwcLk8eH7o0NpMq6Htm1D1JDj4U4u1zIYDNZagLGu2FAOM1C
qW6E8tsf5o9oNq6R6hhNWkJfuSnmQcG4U/bbFjBJUG+bCdVmkJLRvfWiAD7BumCIBgcSo+Wa7/ZO
RjfJWV8X5qS2McQiyIjv84AGnwV5YesDZpQVNHZaTCHxT+ZT5VCb4GS4sNf5JzCLw+fN09/3vIm3
SmNEGy0zNTdYOqIRy4CXXGPp1M87F1j917dU2ij3poNPEVWQgHQtl1BrkKkc8Kijssqiih4vnXGe
lHF9CiLZ7+DOCTvjjLgmlEIU9XZO5fRn1Tzw8WH3z8tDnPvkdwc9T8Q5l4FCT70ECh9FFp/7YltF
sjAZ15oYqBHT0s6/5THt9EOlF/1y4w2577mZUEOlbjc6nsh3fUuK1yVdERCP1NvkiUAKrjEboI22
I5XwXjqqpZ1DI4meE9s5X6CuLXlNFlhx7WTHmhZiN/B68kOCoWIiGhD0Gztjr3jTL1Dd/IQFYQEH
JdDw9UyROGRDyGwq9VnYrJgh6VgARqQQYM94VIFvfd5EmxwjilMuiBHSttzjNYaUpm2yEB5VPEHI
RE1j2YVWWGNzqQMONHOmXppK1UtunYDEIuRSowe8aDVVIVUEHCM8jYIXm4hkmNeO3ijiD3X1nb/q
/A1IVQsHPEO4LPkNRHd9f6reiJbbRoAqmJ6+MetMKVcZp0y8cNw9eYLhXBZF3zIgRD+TaPaiRgZo
6MEQzwJ23w5JAu0ylremgihsLz0himm5GojfJ+fF21MATts5Dvzgu3q1W/0+UmYyA+PYhtvXj0q1
SE8il2iBcFPcIIVcR5fMWmk8qp1S7e5Qf9lGz/N3ycyQNl6N4a729lwA6Xu5W41FqeIqn6E0dbsh
rYC0+UDevA0FBwdUQThbA+IxUjz/QT0rUf5oLRv3GNUH45kZmMjsK2KS2NBTFcfr9TO7QVk3tJcE
GvBnucpvY1FyyIPuLSulpNqpOSych6NTxiZaL3kxTMbAhiaRb7kbkPwz3vJ9S1ZP7Dz9IpBDQjbF
hzVTSIXYNTJqA8ddzZ6Wj7ShE2p2kkqbvz8KdRaaz0N0ZsFK0qFu/7/03OIWZ5DxmcInDl07xU9H
2nKmJ1pFxVP1tah1EFfZR0ECJ0VwBs6TgbFtILnr7x3X+Ox8hm0ILwice0huRROinEhv3EKu2lr5
z1HJdNXaMjg2FWdQ61ANT++kQFqOhFNlhrRSafPFrGc8pXFoRjUXUFwULsg8p/32dP+l2d+nhO4t
Bv5CieUsl1Wve/ncbXeSS3qw/jx6M07qU914r45u09u1C29C0scGC3+YgZGVPJM8gazC9X19Q7Z6
EQ9hwF92xJYeSLFH3ujhGqQsYkpD7RhBu8H2z00kk0v/MLpHR6WOzyAo3oVLJbybas2ncQGiH6CV
zlvwDfzCo1IZT71P7VoLYSIMRnxKXyptZyyN5D9f+9OprJCHY+mSAWE46yLiM8JXWVw3L2hGUx4y
jLFir5UskTg+1JJwOMoo8z7lj+nkmC8r8d3wh9WwmhR9sxGgQOQJauKbjkIwhveY5Y/FrfMGBBqO
TqGVERSz3DeTPF4B7x+yLFpF+OUKMeFhE9fJhQzM27+8DKeTFkVzQla7oIO9vpsohL0Xa/Blg3s6
qbT4opuqSRJhHzxSM9cdjiesDlB7BIoupJHwDHQpuwvn85xDkFV1cpNCFfas1VgRdDQTbaXW3P6Q
R3Sic338wAijFnHrIVqj+60r7ArWBrJB4AYjl+ERzWNfgNV/EWAvmeavuzqgvjuvVAs+9nNqHzoH
Rz9Bivkj//xHveLVh6sbiBa1Y92V3ZqWmCOWykmkeL87NoxlPMUi+2dFfwY6ysJ0k85r7sziYpaa
juSxi4Nu6+krdWmauKvSOam2dBzCvHeLQ8you4Xx6u/NGqZ1x0Y+JPvyz5PZGb4yeympzwe6K4a4
jkTjXMrBQpGXVbE0DNUONvLeB/mL6vK5xbVLlJ1J+Ohv5gbrv2Me3/plgeVTCYD0Pvho5JQ5Powt
jPtZTjuWeDL5G8vPdhRJ2u8i4FfBkZutF9zA8Lw7+IHA/OF7WwOgWXH0ME8xvIRsZUtWdfUK64U9
Hz32IXaMIweQu6zNZm4lKqBQ5Rv35uLuLyDhZpzAxwU2Nz6RIoNNF6nSYCd5AuhZp8ghibZz6yjm
XNIZ89jJMqNHPZgZDs7AsvfFrc0vc2WlDnrLezahTJ2/fU1YATjokHHOlWxrTE4bGxCPfdoaxrzd
p5kjBkxySPXRAllpvzfdwHOPQlU+LWQ8iELg5wXF3vp24EK9pER2eHhb0yjwHAgXLQdvrt/ko2Cr
2wWTtj7LlM8cxSfF8slq8wYfIVDvS5KmLUxU/sJqk8ge9aM9C6tNIP0Iprrysc1ah8PzB5b1Bpd0
rJt5bshbIONfrNNcGpA2DEngTYxeklNIFzOAmeqpGnyBnoaratjqgdNe4LuClgnPrzwCEq+6PPgE
dpry7z62FUHJj1Ozk/GmyNmhiDALXGnpzuO+W0qcuRnCR6BCns2egVrrmNngEQkiPcwOyMn8d++5
trzngt/2uB7XNg3YjdZoO7iy7LtxLmdam2PSfnBIBQNK48eTDWiB42tL08eiYqt2PdWlAPQNQ/zS
mtvw4UUVos2wcDty4hslCrIi1NDD9mvzMbkqcm8KUoRxuaxva2vt9AtUBrBY+mjwBqHPuC3byVCp
/QECqfx9PhI0dzk76xHnQjg82jRu1P6LNmGc94T1Rz8GrIpxkbbxHOkD3dYuu+SvzMUC9UqRUK2c
/4A//CZGtUcpfHYhWcgXCLpkaONWvPuRN+V2HIq2sIIMd4w/MrbCED7+C9PT57ULVtq5IoP6ijjV
uZLJw9KLXRFFkKvSZcd/phsDvIE0Pc0vuCAA8s5XlBOchZJAnts3durm4XEl34W1xv6ypUi9zPGU
syTPSAD9BQjNAmjvHdoif7lS/s7ztD6o+L3LHVOzf9sKGK38l69nqZgCvdXV/1Iy6U+hNQ0r9Cgr
wnG/gOWPnkRtJenCN5Cg+j7pXbircUtGSibSY9SFjYF2Wwiik5wi8dChemqaWA3+GSHCB6TGzzc9
X1nQeqAJGSH42wVe97NECJPJit8nhpln8WXNUDVPOTNaYEZjVb1ZerOrh//j/7U7Lemim7UHvmt5
s2USTQdZU5qJkIHOVVb6ZpNkl3OuOJyJRzTRtoNZuzzeSPdckheLIv2Qepms+Q6fVxmcTp0fHHxb
Vmsxq0H0/1TzRqB8OrLrjbIySh6PqbYw08iZTO8exF1N4rJYxTRC25kMymUFYN0hPp9e/FH6u6D3
5V2Xq1QaMUQz6ucgVOzY/kt/hTizYI7Ed3Z6X76cBgWnZVsOgY4AxiGfl5dGbOK7jun/Jsodx5DN
HVpH8aQTCRy79W5upGOp1xzrqeYI4m++xetlvY8KZmh1Ee3MkWB5aoBrw6+XlpNJxyD7eowTstnv
bmqce0tXA80eXezxxO3Z5I66GUgss6tcXrW/EApa/GjC6sUr/TnYpzlnvQ4NmpyeVGUzY1Cb9oIm
30orc04NZSyvgwiXbEEPqZCZ+BfhsyRKV8OX+7NB944TqSuhkhGgFHgg9Yu+FKvQUszcSXm5B2xN
SoDXHoNaPrDyLGlmznIo7Dn/7rxqv8H44J2wm8/RgzAXiNscNQ/zb5DxlFP+25iLlA2p+GqPtJAW
3QDr5GGyz/6T0zq8NYxdzPG9XrCG9z/pn6r/6IfbTJgWkf1VipEX+FIyzTiu00DLOGVrWkSWLNMb
NiSHF6Z+Wkcd3mJhJRCkbPQ6M+zPm8XkNBQdeBlGh+VXfPSv5T7ftgdJAIOQM9VhkuXklPm3UEzy
ndVO1Lx8s875FGHA8cRIgSjxKO+/2yJfFrf8hxuf3u77GucaQ6mHeiGgIQExJMRJLnUvJEOSo+hx
v5VvfwvLpUT5rZ3FpYP0wUMYrbzuzukd+2YmptCV/1wge2m+DrU1CVipriWFzpL1SnzHOymg+RGm
TufEV4UCd8fRs19ACnfTG0/bZOr912NZOzsUUJGnI4oZVZDbvS95+BN90bQWK1AGe3/RQZVVSGO2
AgjccjphR8RujW0d5aOIA5rL/z3M5rn4L+zMiLDTGoNi71hDpc+QJl4kvfkqppb/flfmuR8/4Du0
6u+ghzammEfFvtAr9jDbgrzdgIiVXZYTIaz7AiMPgxlGVhZ3pgIXGK4i4mdKkYuTVhNIY3/vh1Ob
EQL2IgC1fgXb5ymIK/2i8Pj9DeYdT8UtTf4/MDQZN00m0nCneYQlXwsCawip62eS7ynm8nVw87mi
X19ew4GNhMLMjR4y/BMMBUkRDUt0Lim1UmIL9lmAwqk1O8iJmQ6XPLN0i6frb+pGXE3JbFkv9AbT
cq80TbXloyeYUufEuhSn5SG2IGhA+n8U0wbvKoK0aMe1Ic9j9+qKdpXOWnbL5KFYucinQ4QkcmQE
JT6Gvx51ZinPVSB32/MGton/KMwfBkoM7wzUsu3o7c07Y+vDI60gOZKsjk82vJjAW2WzZvd6H/+n
9fadmI7yH+8JzvTRoL18LhMk2Gupb61+KA+EHMM0+pz+b1Az26gYhnYK7R1N2D1Gee6sbI9YHIuH
7OSms8NSQNnLYwRjiUuY6n6IKlUsPSit8nJEOWRUQwVLK4KqVQo2STEvVBcf60I+KITNhafUynk9
cqAraQ3rzA+F0q57yM3ydjQ5o5G4pBQBrmS++Q2UBQXxP9ykL8i5hEgzD/RUyMCGQz9jWq6TeQt+
JchsQqpCl8DrwtSLf3tVrehXYAaXqNqKvudCBidvoRT7l2ZE8pxB8MIAGnpNMXTdW3B+Nzx0mQRy
ijKVGxN95Sh8WNWTfr6/Guj1f4nC6uXNW3DXVKrm4WNk57DAiRmXGjrPt0QrOwhrZtEsL2QegQ7w
ZrQZLbcZVXi/3xnekL4FLP8AidjuUZNOj+sukKLXAjWjYj+Ksqwd1/hlhRwlLiqs0tpgOE95akqu
lZfy5indeOrIYNbDqQ9KpzVxjH16qth2EYs3BPOA4aVkB1bPPmsfaNsob3omtTdYdAkarjQv0EUW
FTP++cCSllcJ4l37bA3ZzKw2wltIAJhQTg98Cr5w7TwHNwLfIbydD/d19zW25wVjFjl+n8+aaBN9
C9SxfbQVxIEWIcaYsfMl+c6vz1AeUpKBLp+VP4jGPgk1b5v6ei0adJEhOxBv6+ffURaFFYMVohD7
HjIOMdS68BRe37a8oEtTRkAxyA4Rp5qRDjqmKcKWzfg3xZ2MFIreYs/lvo8yOPyXftjQaqED67J8
2oW4cKxOFOSuKzqCGsgXSTOjMmg7fxGlPLTk9opv6NQI+EFCWFq6swyEyhtquZOrX3HE4+M/2VvA
egOWEZ5yL1mDqB8xRophbo/W/I0JibTKxpI4n8HEam4eb3V0qbtpsgjLo0ecUq3Dq3n0IJwX+z0K
tB+JdXLdhTQdg+0H0kKgRhB2UKtpj99stJVmmSlJlfx8mbh4wznDLzHUghSv9vtc4zVAZFG6aOi7
kydhtkEas5KKS34HffUWAVFtVSo5PmrYH0AzGkOyr/qw1mrCgHF7/KWiSPg+2pB+wbZlynWJeCep
VqpMLpndEl2jDP2Y6wz8EBP80a+CF7pwuDN2PE0PTVqKdaH2xf6lb7SRBkOOhA2+aRb6k1UuPrHi
ZKqXk0d89wp41DYLlzgSXoVmc2lEO5ZiWj3AxmacbJ6B09YEQDHZrpDfHrY/7Pg1rw/7SKFWsTaQ
lHgvTHEuuWBlAIIND+2ZmgUJS5hFZK3EEyFxvMXxkwHyy6vKyo4WQ/WrA1M4lvrD6ItJW9BNCUC3
Htnq9pOdY0wvW9QTA54M/h8uIgef6kYfBPlJ+AZH5cY9b3jRqaJviQiYh1pZ3KTEQUoRV0tCqCiE
XYU4JoVkV6CS3iwZPg92mQi6C2EePR2sWF8IcU979KrYry0C1hYmcJxMrLQJ5pzCI+Uqna5uO0g0
jC+fZVqXixyG87V5i3gGnbP5puwgKosO7oEhIRpzABt295TgoMU7OBxRRWcCAa83284RAn1Kt/Mk
sa66jZ9xPs7Vj9+lxqiuxuEzKPpgLyW/n09+A4L1fKuKW19FBULZ+G/NbNAIkBTKpqNldGcGLdLb
NTAISqH2ZHzJ8YVH7Nt/iHhsDGDjJPMCP5Dc097a2Fslg6y2/Y0eIyC18OzyNl/lRIx5XJMYUEbn
/P6GkWM9NyrnWOPIIRQ7Al3wu7XAE0QVlz8R0jFSjQT6k5VQVXx6wIpl09GmKr4g4yiqjMaEnISB
d1rNFWmk8CsMDu/GWV8pf8cIDiksNDHaY9S1jYOLK9MoT2uteL4TR1TAddUIaCJGg4i7GnO5QIdD
DwZO1x4cY8Y4jt0tOqef0Y8b991Mbxv9p+nYqg87JK33Z63J5H7cqbbl+8vwJA/qO95oiw+6BmMn
N3V+iMrt9czHIvx0o+c7N67+u2GfNDt8kQ8QPzG4IVJfdrbNJiI7j+EiJ1hzVXk6Bu6fcsglcGU0
XkY+8pZX09Wg+u/r1078vGMUOZMoW9IMnO8sGwuyQ69vSHRRPghtlU1Nhqth1bB9OO0H5yWm9ye4
42JbNn0gCHt4/bnn6yKynCUGH0mZAKUz6XpcsPD+IJ+XQDNundOp/wA8vhitXAdvjj5Fg3qn1n7x
PIPNLt6sq1Ntx0Xs1pl5J1+Hjzw1CHj+CFZHv/VA5ZjDxQq2iN9fXBfXBJXe/yuy2KefcO+xG1Gk
l+BHJHpczB8ImG2MKInpvDlQrn/Q2CI9Y1MPFAOw5u6scLTxW3HrK6PXkEKhjMcNWKw8XpuBFnzx
l9oyo29tj83Sb+MJ0V0zgG3QAgccOjCexkglg1Qpbfve8Eze8UlxE2KLZccDFeQPrEof3Z88dgPN
OuZPkq32LnPGLuRmOHeHmzyDinwAXcnOV9i7yo2H1IlihpMKCbMvRfzdbkYUZaKlIOGJV08fG3OL
5CBhB77n4/3wuXUSQHiUcsKLmh9vz6w1enmkl8qUlBxkWnjluVj3S1Uf5Pc9QoXkzAvwdoJXE9m1
0QON6nUzxlRfl/VRnOlM1iO/wg9zE9AG6hAAP2nBth0iYxqvHAElwPdS5G/5PSJfIk90Qwtqy56C
oZsfsnBD/pztAaxQy0XY1nAKtsFk0+yVqE2+h63tjLLQyYApbuwiBKqasXOYGqZwnDrxnVi9+M3P
ZvgyQ18QQ+SrvzqYeTEkPVA1PNJKw2AuSo0br2NZ7SRMq1hpPMVbLkx01J2eapMPAKPmisK+bwtm
zqk0pD8cVboy+g9OMxT0dbuEM4EhhMWy6CUtjF5mPdZX27OXtJAuhNLzIVKKR4HGkKocpqVGOW1B
DplG6AyBnUe6K7cpOexh31eRlAEwYOl2du0AY8iT6Amv0TxTAXki0+8S+ll2CbnuKqaeIQxzb5hn
cr/XCNEA7+3ia5u4KNZjD0fWQV7Yxx/tnDw/CxTiDzG3xTXpxwmv4EtD6hfhrWrhhRH9ljXZnTGZ
7K9upQJD75i/a31/Y72u+6Am/gRF5YroMawFD5fdoLhQvnpO3nLOd7EFmsbvrXnoYwlYAAfCRuQq
Tjh8+fprfWgqi/8+BqfELYRzim5I5Dhs6SxxZlFZymrpwu5ZsOQVGMwTm7K9ZYZQ7NF0yzt/xoWy
zbPFPubrd11uAhz0/z5xBzLBJcwYgHSpF5C6nsNOifNB2IZqgpuavdaI50rGGKb5StDLlXtGLJBW
aysmPvJAbLBkgUpuZyMDknEI4CVUnJ6VnbM/55Q+jqLq9aMrGc5aodwaQtVSeZSkA7cpnWFFBSYN
SLijFzo1Suyw9l9/4/aw+Hpo+DXIqBE4kx88uTr3jOcDhASURGaCnAH2thJueOJYK3Mq8HvZ5h3T
sF4L0I0eONqCt93OSl8AjFsryRmRrFerR75ATm4hI+AiGv1ruHunWmgrC7HgvXI8uC96slng8nuR
4ztmLtsoecR4ujZyAizcnWzWpVD6PrJnfolGuXbKcFoHc1ug8aTY8kgiA2Dc98xuR/S5uKKrYi21
MChjmbWVdTGw9L7y5Mg2XazQKemELgcbntU80Y2hgNUjfe1VuzUisQEQrSBkQXY8jsRohZxeNOz1
NoFR6ex42YvZMC4oA7WmLysdsi0vGMB6dSaGbhsDzAhFXkS0m4Yu0VeM3oIhvNdvpQ+WSQQ46RIz
kpFWkxFakwBQH4p2yp8sseIIjhDpRz7SKhavDXhj1e0JcsXtzXk9kyAjj6eT18WHSuMxh8amNO7U
qgVkUe7Jt8ST3JykcexXtZHeRaekX1cCQFE3E44jvUuR8KWkvYgnQzJBkO6ltBAupUW2O6eJKnik
KZORz1cPZjhC67hGuSlbPANz1cdBnXRqDASbvO4lI/QK51WMOucjCqrnV5UUnqExCZBMKB5D223p
vC/6PRABZVEeFARS3T2gWFKeDo852859PG86dJnsWafgeCHauZM/mSRPLgFHbtpjMJMD8GRIMKXV
zVEow1C+UJGK4tvVDFz6A/jjhaJeIMiTbyNSu32rCePXQPIM9g7T5k7sRSZOEyyj8Jd4Pt6ukxuY
OikDkHXqdGj+CLZXoNfYWo60tBztY3o12Bg6X01uKDhaIxH3IrbjtWYkwXLnU5/9ZHulncDaPsP8
x4bPh9sdrYUYkckByJsaIF/ch8ymZgnmSPfbXeCSvU9rGGr0BqlwKdsPs/bm6LO+h5/A24HbRydY
v6kCKMDNyjpFfsxbxmjS18KyRx6+C3h2/9TSsy4hYcuzlJZzW9laN40xt5ua5DQmmjQ/NP9xe0m6
J6QMJQCVfSsKQ34SaqaHOUKVlJXOqdkWpRwx91LLJO9BHL7cd8paxCD3kR2xcMTHsdPtHiO9jkAx
69xKhgD82iz2W2cfUqoa3S4jHtyORSqCPCysv1jlwd2QvcmJ+L/2URbOOmCYuHFDnbCUnC+aXsBh
jXs9U7ryXlzRtN+Btr1e3vhB4M48LkD3UiSQeH+pAwQAtvUaCaTwd6YgSBU6s+rAhyzcrlJN7/It
vm/yUBwtR4C1dib5L7RQ6o+sBv1onuAR71ssuZm3Kr+/yHOJBdCasXLBUepYBNgrWK8cELdU4E+P
uOGZlEfNfRo+KSPZBHjHIRgyeDmNMK4+KEi4R8R/Evc6KteD/yotlYKf/xkwVzBzt6vOLu6/6uKD
jeZEc7Oql4bbtKbVDpCjYhA1mw2j++fQaq/QO+GzzjtmdhXbJAE5BcMMUGjhwjCGSwypFjPoLQpb
8VDOEblX5NwUjERP/nT6TA2Wofx0v5SZEgQ3Q+V15bYz4JEAhkJA95Wloj+R6eaHWCyykif2kM+G
+ucYbBNl7/zBXEHeSotrOakpR8Oz0dzbsLWpwJqA/bYfZLWglQm8WUKrMd75cz2ogSh/JjvI/cf4
o10edzMdgdP5thUcR09pj9UGyCHYQ1y9MxVhrWE6EP1AgNd5ekYAJ9xFhYZA06Z/3GdU4y1aLrRu
DnlHjCeCSIrwTiQx8HR+cDBeHGszk+GgjkstrfHyg5NiWQfR2X+JoIWpT8slhCTxa/jeu3i17SAx
fCUr0XLdV8KkdG7lbVs2Bpp3zUWZv2q6w73VXh3s4aEvfUYIg8fbUZFxlkvZ13r7VYQlZd1qNzrj
2vhGddGOkCc4YioUhw7XdE3bu7145g4bZgTGCiW40NVCuNs0E/LT6cy0+71wvcHXFQklFyIhMG8/
MLToc/JIAcOYOrzWowPP5tXWz+gs/84pYcETSPFowzqw2Uot1duvUEPyYEfKcVJHAlpYbH1xRqPc
omPcJLzn2OGEleEf/VEaVtWW9jZ6109lv8pCq3d2ACK5bhs7RxhOcLdXatJadRgxtLXZthJzFK1O
cC7pdmRohKMiyboaCjAjInEWyoGcUkOCKQqw4Ry+XyzadF8Bu+7xAaYKL8AmxY99KGdkKF3gYMsL
coYu6K8q57fn4vDnBktkMB7MhTrOHI/WJoURwnwZjyzj3qMRh1gu810zHWl5XL3JYpLVyDwCfxLs
M8JOz4623aVnBaz9g/utG8Jy5mVIlKl+VnqIbvghz8kVRRcGwH1i/TZE2TEz0ynGXUCJlkMboalK
jKJ2akBS7f3vPTbuTzCdzRarhEtxG56SvJzksU2vP0OQWeJd9ezwC9qZWtOd5KHjExi8N/o0Oslk
r39f1oDsgs9gkdEGI2L4soEeItUkwlZoznVQ8d+doEj9oAV6btZBhuLRivg7x9nABp4XduLBLPjl
Ny//O0aV4+jekiqfwSjfrQYgyZyT6inNlOzdF6xppodaVo87BNL191txks9fC1fva//rK7YRpgYM
Xkw00ui977JFfOmGnPf4VtHcvDKbLjoQVKBe7B7lYaE9BJoCspRXeQ+tprsLVPrXiuMZ3OJPJr2Q
d0umUeXEiWGZCO7Aad6DB/46nmBF48K4z+yyRCvDlTGlb7g0zYq/mRj+T8RKuNMDZQ5RpdxP1fFU
IaQcPyvCh/ZBAInC16MeynB/+s3nrcN0JvnuBetX97OQbpJM9J+cCY7j81r8y4yeJEJwCOxS/J8G
EI/3nG6dBD4fTs1/xHuMyL891J+7o9DZdLIBpX99ScqyRNmTV4IPR4aqNfmEXcmjke/a8AauoQvu
DhI4zBlhzbUz2TM9nrp/G/nl/Xa/9cfKdWPRpbOHzcu4xhpqBC3Vj8p88ImVZtK+j3L+Bfl6LqjH
n3NF4gacjzCjM3+jECptSo59/STKlCb31FvLhRgffZTEoKqXZNhRohJgkalbtUCGe1pQ0qFsbG8d
ea4dL6s4gObzpr/J6toQ/8F21GdonUSd8JJHLA949QedDRx6WRuH8vlycoY5q9Zm4o+qAgWdAa3P
sFFG8pTAT45CGYoeRISj4XXwRtwV7w581Oy0IPPfnMoBSHgc+kVjhkZFIGvgXVQSdOzRMAd4ZjoM
NL3RBd54ed+X4kaJfYEYcXgLJjzXeH7GbiM+UKO37RzvAiJyv9iuYKbJDkdDaP2Op+FYXe+afbaP
puczokAYudz8RpD9FkzN1iFvdsRsLfwKTbRkBAlH9FiGNGq8YAivzRavNjREV+B5sBc+j12VgB1p
sVBE3AI+Gt6ccg10TRk7rkC8sev8PQu2WJ+qFO9I1ZHRK+tmAKPD4h8+xSW9RGuZ9Xd6t5gnARgo
FhWyDSbeb8vmsSb4A1h7Ws9O6hu5lzbU5uhL7M/4T9/O1J3UuZQFdXl6iM7+PVYeXKvv9XXQN06I
CQjR7fkYFkkwxp77Aqy7NDuc4OVwGU/G1sqVDy57JlaN2HOM8mp+WMEoi6H/84B+ovRgF0vvoP0t
KK6oekboZEysiDZp/isto9egoAU7OEblsmyWYm9+oVDescoZx5ejF7UNwPnN/Di4A7keDwo/KPTC
vpV4dENI+uj+6jIe3TclOfziIfcLpDs/QcCxeefFtAghkCo0xB+x8bD7FLX7+1oqDhrlA99y9EVJ
xL4XpN2FASphYuMP6/PNtEvS2SB8M3+MCtyvZTQmNQ3M+viDG62dvGU7GiZ9xXeQu0JT/rt9PLTB
nVLZVzlBFWjjUUa23hYlAH1xnAaUvBkBt9gfQZJACJOfcBFUOT4HUfdsea1t5dAyZijPW+D048Ax
4DgEX2+5t5FKRUFY0sglNUpkrBmc0ahNNaNqBme45tMxmcv7Vn32wUybUWigzF4b2OpbeZKuAKXF
re6Pb2viRHOMQSxltCEHPi97vCKJEneIp1XS83dEjsyl7emDtLmdCmjhHXVa376Kd43VqxnR9fSr
y6Owo3DI22N4Lhk9VYdzleGgvtVGuWDqzcbmHkQ5HmqYtr6niy/HDl4ZHpZvJyw0YrftFZXYPfIW
m5RIQxRJG6NZ/E0KNCiOvR+KEGHz/sYURlmGJY+PwWVIccfXOzOIrPmXYUvgrtMKPXZTIS5QcYsV
vMY/eq8HEk6g2VLzBG2qtjLOM9iX2scRYYVPtIblRKt6RTiaSuIdpbvMPaGZUedzjNHMTtUscl3t
pAg68VwsQOqyPLH19DNdO7DZZTKvpyJjcmHpOHfJh0OZgujSepmYRjV0iUdZDWyfJ9EfEesyOn1F
s8TRXr+RMU3mYaq87RjziCG/niR+74eTpwNOF4q5gz/suB926t32Wg5lGEp+EYznqbXFAHsSnXST
Qdzfr6PLOgPamUpelbkV8i/33L9huNaw1B7UWmE1s2diPS+1KO2It7QFChdJfw89yhGdtyFkxtfR
7Pi4F0L1lEaDfAECr3rmpgHjhPYbyT9wx6sCyuvz2a0Q7pyt0pab46SzJbyQ5ubbGKgL880fUeON
A4qncA2lAew6445m2RLLU4caKrrLoSolQRuwmaa5USOO83noVUK6NXbE4jTNyaDny2drWN8r9wp1
EzlOOej2ysmL3olifRpyAk6/dIVyvQI9s69ieYfZAm1nLFgaYjyLGY9fqHoE4Zot3WLmJgoSJr1I
iIlePqpZtNknnLrGaH5aqyCQeooRVRopilxdRbXD/0fFPFjVpbdT/SXM9OFWinYQwy+Uv+868ist
BEQSC4nQikKM1FDA+2EnOjek4uCarQHhmIjbv9SFHSEUXPyWr4E9eWWuMVgN/mNzepemlpChdCJQ
rNsGlwBwajy4dj0oNZ10///zD6zjWsIK8uH3PvJrRHTt2u5Jak5TVxAYYoAJhEKujAJC8nynqBLr
O23phbwb/dxaLE8UnBpQWCBFhL05sKGRVKH+nrO1bM9sSAQOW0W2TxMbKAk4ajlfXH0DNEhXVsAG
P6GLyFdBGyXpFvAPDxEJmjc5eSYTFoF8fdvImSnf3WP2NY66IoRKdoJum6D3bW6KKywNx3u8gzq9
sMobQzKAFeLZl8PLmJTID/PyenPfG1da5VKl+WGOcNQI0DKJSohIsC6ODwwz3D8rKfhLxpcBr42/
WxKDkWZ/X7YjWlX8peyOzpfWCUkBTRcGDXOwMJKJDQ6MR1Yn7oSLg/ysPRdG7rnFdAisTb3B8sII
AeSUakqe5/naKl0wiWceCL9AQuqP21pRpijJil6o2r+wmcuG2bVWL9lVCzQxzd5U56Ck9Nn2WFNZ
9ZWWbeT73innTir6yz93z0J3JcUUbKKBVH6ZEb13Jlt2BLFdWnlWb9n0TyrU80NeS1PgszKjMaZH
IPVoMo/xm2rA0wuVRllHCyzOJ5uY3Te2Zxj/J8sdRh7CcKs8Fz2dBLUeuBxpOAedSyundl641HQj
OjCnBr0RQg3DgjAlU1sj2vDGyUlNoKVNPZY83BOvaWPQbw6hGRtD//7r1sA/AnaEwwOFeiE5ZVyy
7TuSShqkF8o0CRA9bB03VLYgvCScGv02ZGJNaxFUiAbPEOcHy79FRHZGvFY+kD3RXfiwj9bcfNxE
6NrIrgOQKLhdhhrNvJV8JzguTjtfZvlYI0szblsVgJCiHPP3gnw+UbTn6YCfSBVpvC6y1p5YJK8t
sXRUdih9IWAJaOPH5cRS1mjJmYQVcLh4lY5gpcXKUa26XjceBFl9xiLzOjTetfTQiJ7EJNi8L//8
1jnjifKdY5dqjNJz9ayCG9cD9nStIT9sgun8n28idtIx7wBOwTq2aGdY/8pwA8Td+bOXpaki/pPU
c4DRfaHfYBv1sRtuZo+A31/xBMvlhUtho88uYU/fvBmus7m8hwfH799HStFHTwfGNq6kT5/STTmg
ERWRnl8oRagt7ZaCEWxNWteO0e4Hf9wqQvRMTM9XGPZwQbS6etvmt8zDtn+eWwo41ltKTy2/1c3k
JeJYEJFthCpXR2InfxKwydivuKbJk3ILNqRLMpVdDdsFtMgYQsPFpdWGN2V57L27ODIB6BrYranx
A579sgq/SktFTdOF9e7OHT7+brHWxxhdg0W8EKHSxGwJlNCB/Tobg9gWTk7eUln+J0mmkHuEHQxN
B3651FbbGVL+Ho4eu3TdTnnv5iVUkZdBJvlE9aw1JOAL2Udwx8hWk5+jYfd+CISEt6VmWYiJuJW0
7HhMYZgF5Ye7+uM5jzTT0ha7egQIw9UWc7qMJ5oBPnf9fMlKZOlH2BBqfUSOVEvpNwQ1eFIjkOzE
F14yA0a3oEff4FUkO3orh1jMSAuWrhmYF/Q49Criqoz9tvSHHZMp1TZ90j6GLhPH7egVRAmlYvPd
oRW1NE9PxRkt+DANdnmJuAjx8rlM5a98FETkuKCbiuUDkaSpT/tvU9PBTSG+hUjyD+k6VPqLi557
pz1979FwwYd9hJjuON0U0aoapXWPIKPTuHFUSqwYwlHhiWaaS7+tMz+rmjQf618Le0Hrm6asGFcL
jFjPf7peChfrJ8lO/HmAnyfhl0s8yMIcuhEQClbcFYGTQFHWlTbFc0mzhS37rmjOKdUO78h3Xx54
dURwIwtxjnP+KEPZm7hhGh+x31zI1ZpBLUaVI79FrdY5ThJ0+lsyC+2XpeWXKDQILmXSiE74MxUI
/qfTeocCtxVpYA1n6+zLop6Uu+BNcbMrxdHeKGJU574qjBGH6qN3aw+N9c6D3v6HSPgDXEiQAyxs
ff5pukpcWLNuEFmGASp/nPLnOD7qpsQqoZ90Bt5gh7ie0owYKGxjPLr5YQLVaHhwvJeTNcgeLnbS
zsdVyvnNT0wInjienTgTaYaEnf99sxp6FLd4S4TW1cyw8YyLzxubqOzHoDMJna7LhKnd33mywZPg
57mhQzs/mGTcg130YVp80+TaSQGjuLmUgIaq5zExdCwEWmQY/kKO+7Jm78W/PO1rVIXbeWTsCUcK
S4iV3PEjx73EV0U42c8abLZl8izQCsrGLMNgv5j+R7XkRBrQcZJ/RbbDDiUcNN+fofBAHDCv8m6V
mknbPIQ6s99ppJ+0mQy9cdnFVzAzueM3Jn9ETMwiJEC7yhk3UqC7pljRZ+KUnHtHsjPAUy7F6tbh
8AQ90wFrDbH2/mPcV+rJmJBQDhwxANnDuKVL2D/KRkxDhu3QeIb9EJwJRWceUCQ0FOJLgopUbjnx
+ZCq09E684GYIsnbbzeRozJF/Qp2qZ7tp8LOEb7fYhrWNqee91uzPfHXt9RWRsPecccdj69q+bsB
q3lybaKL3KAwkBVYyQ7ccmNjzGEMZZVLfEPfRVZqIXCJEUqzQkb9NEklDKVzypgePfwptHIhyMKv
KL9v4QvSEmlg7loO37nUFSK2ATRSSgVlSdnCWJq0M2jV3Yl6Ffpq+x+7hGn41YIuGNB/RosPrjjn
tAFH4HmMfj/eP2ppj5yj4J5Qdxx187WngK9I7//EGELjCc57l/kkq9SD/tAD4I64JVmsrYz9Q/H/
Ta4Q8LQhDYEBlz9c+u9WZdkIKq1jKZPpx4JM52hFuhYPNhR5OaCDBamN01hAeoUtKC2RbRc7j/A7
0cjIqxsOMIA9pxhsVVTyZUWTJAdd8mYgoSJRrNLeaoSDY4kFTdQo32HdENfKkryzgOS2JJUqR+p0
TC0ND9R/msY80vEKqTlXUw5+Y5hhcI8N1Ve/RVcog4jCuMcmM3nugkzfXUO2d+qN6Wa+CYtgdkCd
64Wgcv1HANFZwACGdtZs/RQvUEi8lJOThcZNQH6IcwErP8LjFT22RTtUry2cxONyZZ09YgtP8cQ4
T0kCQAA3VYT2LBNkTfC2xApJV3Wi+Od/Kt3MZrWYDp5mVnuiU4/sOiRwzJx6+cLhuM6CMy0l490A
fow7ZYFIHcDCQ0t/e0su1i1eAYbVwOD9CLocUT3Sk4/jdbxBLth7zAu47nU+UzQS9qupr6zTKdWa
wY+MBbseyHER/9uYSWrjRedFKNpK4zySVy03Osyu6Q+nQDtp6U63EkBOY/Dk7B+d3oscjenSj30M
TdJo0X1y/y2ulTXI2t78P+dB8DtjRPNM8WpM8qY79WDKaZIi5r7oTlAGca6bkvkRR48NLvgrW27b
lWIkvGDkRPdbvYp0V6Jx4eKl3NA/xu9zm+oZVWPEK2DykyVp2Hq/SF1S8TGNdXh6byUYiJ1eK1BM
wsWK59v/BBXop9MsLfXis/qT9+r2krmLuxNtbMnPkSQxXNMe82bOfydGMp3Psf3Yme9bbrPQ853T
7o10XHKwmSBempjgnV+2yDcVE7Y8wB9TvZbEQpi/6yHzGoshz7hnlwbJ6WlNhMDQq751DM9LJ/FW
RM86SEmKAabzpovidtJ+1yQNIclFD213rUrR95eZMR178Avep5ZXUFm5NBywbNqSfY/gJcygTH6F
8Gb10pVyI9741q7OIFPaylkQZFgeOamrf1mAr1peBn016JspcdkWUy1JdROGOC3m6QhlvMWVXzgh
E0WNc7+DHDpWUoKntn8qqLMH8izW2rnsuW2sP9Uz4XSiLS2qTXdAlyb58T8ld05y/Kc+Os0u9U1M
q/yVfvd7d70QqcCnF/SzI5872muZcryVy98R5rmLRr0fPn2Lo/lfyXXpiosfnwDzcXL/yq2x2TPi
ROeVAlPLifPLYxmpEOhT2Z1reYdk96J2xyMjz0dvXL8kbvX3Cnf2Fs2dJwrLJ6M4N7SDjcK0C+8b
1t6/9EZKnsUAx77SbRsoDzNmn/xFGu+k+UDL3vk8GEYQ+u1OjpetEu3D1OPrCVK6KX9NzCePIr3K
jo6Dv+KKlB5Yv6YarX0kzE0yGClMc3aNDNjzlv695ANFq1miP7r0FgQqmPHMHLD64RPMufRN/0KG
vaqPUM/dNw4NJr7m6P0EkAQ+lm8f+8WPx12lKvqp5I2fHp8RoARshH4RLhS5MrA0HTv7GWS8J1kU
vVERs0ziDNdHypkve33kYxm2IKndSVA/cbhSCg3M8ZpWtV2NlgnvFhyPwE3Gy3p0INC2rGEzCG6f
mNCNP28yGalAv2zdgszKVWIKBNVRC9EP0YoHWn9tFoYdLqkGWUr0vh2G7Pe2S4/X1HofVdt6gxgd
3BKQ8mBATpv+52Fopss79ndBW9eF84cYPVzfIWgVPxmQysg+WMEcn6E00axCRquiDoFUfUEnR6O9
hU0xK9op6HQFDWlXX5iLevtaAkoGxE1rZp8aJ/nd8+vPsIHxjSWmgEvSqdVq/VOzEyZSCUH1twsI
Z7llo3Athe7Fj9h/E0mj6MA6OiIk0inYdCENasolpgeI1kJrzcJcIXW+Ho54xnjRR7dT/iJiKS37
laoahX/7zKf3toDufvnBZxxBnW1lMjHnLbbUEdrLV/Jgt7+jRQZZ7+mMCkQyfdZRPFcNLWubpGOF
VuuhDlJpiO/34yYfPMz1GC9MzREUGpXlAFQzliQFtS1CrMerdAARJy3U6wKPAqqa0Zlea1HCBwa1
evR4IfCalzJ0O9k2JMvmssdmmN5Xm+uPfsbt8xRaWCPpNqRL1r5XkcHvd5S1IYdeCro/96He1G8J
hMhWWtrmVNp+0Uqfb3ePUdd6G2FcDA4iQJhowr05pdRFmk9QrgAC/buIS0WxOxbbXwOiZuUtJTZm
k331GIvHxuJBqbdr356SLyjLKFR2UMAlqP0AVlnXMVG0HBwcljDnUefc11tk2OJaFzqb2URzzaLi
L/hPq64KiXUDGIrArp2F+lV8+ntsNOkg0cCEtzaFnXYTj+6IQKG48Gi0WFMxpWtqG3ia1Dt5UDoX
xllFD1SebvhEVyQCXCc1dDW7litdRequtNd28UV/lxXWD2JSMTUxQNo1s1YqkDjswAOS2SMeWKSN
2nC01EnZ7YinE1NVr84Cq+dlgMPMhR1AxTBICk49KZQBTlwxvJCzzKw4oTmIn6sgeCzjBHBvWEof
SIPJXGGOkH6C+FtnPuYtcSCpYTIziTiRapq6y0SL15uDbr6Erdma9G7NM+8sSaQf2xpm1tgMkfYh
Ew47Wq8k+0+1EDT7X0R5t7LWoLRkzRDWnSmhhyQzT1uGOLc8yXxBUJqY0e89l7z8WOYJZV4wAolr
U+vNfSuns1OrMEeI1SK0h1pX+7Sz/S435KGRr88h8C1TZYcGli4rTMJKJlJO/Gg0lQQSv8h4Ybd9
8zsYPIpBKGgf7A1zFypqIvCGXA0INTyKtqRnQulQsrJeQzpbmFo/QCi0z6cGq4RhuhSPDk80a01Z
VtvAB2PUWBkjZ3BQwy5WPHwyB/uf+WtThvByeuhLDh+we5uBuJw9Bl4yqH+n7/eA6ph+kvE8nCkK
PX85kPoSZXfrrlpbWm9KJ7J37JZhxDA8mnsKYgXGDM8kSK0/qZH+IvgPiD4xRigALn1OzEhsvpo9
VWNFG1T17BKQUP0XsKf4VdNAG0EdaIwj2OWwJbi2OykQWwtD8LN1Nt1aKqbmcadakTLKVhXlz8B3
wFMTEPZ/ZnybV3b7cL1owz9BLVXgseVtCYVA27CqYhHGuhg7cSs3963rKgpUZIucLm8MSScrDaTY
E3P5AAxLxwkGHYdZAAITNOKt6kt3lRUj77KXUB6KYLQBgcy1BNDXvHVoRfAt+Kk6v3cXf6JWmrWU
6JC7+8B4PlWc5jS1itBJzZ9hEt0s7SqggkgYwIcoQUh+L+dpGT681L9sS2714hQfT4benR5C9+eK
F7Zz9l8kITnE40znJa6oFADqd8/TlWtIC2b9eHboDv1KthGGzMxq3jLOdH0D3+U8avYApsplIDwj
zysGcb40Ov04vMrjYfuMAzG9HXHEhTgwSn8JUe6QEfmbYZ2Tm6M0bf5D+PhUDjY5Pz3K+Il1WMgC
DzzDZHlOYpIeO8D47vNGX56i/4FkMgCiSaG3Y4LH1Qv4WVNruoXrH2ZNU+Amj+Rwk6dxACv8/kQk
xG7id9jnxXhzdXQQPtS9E+mTsDwBjy+5CLPn2Wro9ikkfF8FZaLm17M3AENE+WWEuDDvn7vZyCzh
4nyQVfvkxl1JgTWCmQGqW5P/qNj4u3HgLR0/N9u90EvbfnL+Gk/9+vl7WtEO6iQvpjekftjK4ai9
1F9rwTahusAkzIxyCuG43tUpiz92wwRZusjW5j/sy+9BZ8gy7WI0ZfpXBYArjvXFSUmo1jhd/0DL
ROEmj74QNoMIIbQhetVnnBIfXzxdQtS8AGTwE+q9hsSw5DVxuBnCJUaRWbdaHSWprpS9eoGUK04E
5jfDvA8tV8LFwQ4xD5ScBQPOzvACM3OZoNTm0ayNb8R2OJGHe6XXiPElQLeNJoiwa7Dw9q7XKBOG
cEiPXUaqI/3JoneSr11Xe5uMwOR+VYNWbskuIbrX6vE9oVFVxKDpc0cgabEGoQlH2LRNcJR5jR8B
ggFFZ4cH6KxbT5kbY7aaOS9MZGEeLHKXYqFLIR9OJgj96QmmxzR+ISH1a+dLxGY3qyjg4y8geJE2
GSptDyfBIien9unJ92rDdIgW3pyr4L4TARc+oheU85xHiTm+r8zUgm7BRoZCYxXwA8z0RpHRE/4i
kVBCH3DWwmPoBlb78QtJeiHCR0uZoC0sirr5SfS8xmxk5WaNkbMl6jQWY2sxARhpWmZq7BIrKTSi
5o/WDBQjSzTGSwGzvyFRIJ0hazv4q0sEa/KwBFAS9Rd4sqeUsujPU6uKAoYcprECiyl6ZPptTIsS
qsoXI2lha8TA4+KcWpZMC5E7aYnv1AXkjxw2jYyFfwwszpu4GXJYOuiVHZ3PqVXNMyvfyRwGyFTW
eM5v/Qe51fIGp0f8Y/Le7bAG9YPYro2lZu/t6vSrBR+AY+eqqrzR+qhMueNBz7yTaCyRiT0c823a
kkaFusW9ee0S1OdTylLf/gsiQpmUBc9S+gjsFkELC3QyOYmM8ic33ucSWcQu5Ra7QxOuW1kV9Amh
onqNhGZWDVLLAOhMBK+VilT9Ye35F2Sw5WCdqdqUds5BLfqToQCC6Cd5YGWtz58/kOxrazH0gDM+
QEIDH8b2SOjsQ1uhhdWqMUbwRePgwTYLBDR0/y0luftr+P0V7pIAEOT6X98K+pvjcQunYQmNAhPc
3leUaOuqKjCNxgwVUriFgYXBaVTaApi2YL9Hba9ZSHoxkFTZmaSFcMi1rdOySzy4cAc5D6DaD5It
s+4KNEfu0P2CuRiQC7iM0g2jQbB0Va2SxnrokV9O4pUMe1mR8PB480lgM1aeQkVM2SfX3jX35Nzd
V5Ab3ZmGAbk79k57+kM6kcjoWcU2v7OVlutR5ITCIaPsAgEoZ8rMG3vPaD2D8YnrOWX/l2zl6Qrc
+PlB5Tszx2MFELqGZc5kcZs6Q4XLSgK9/dWb064ymKnNQfGsu9v3VO6RziB2CIDg0IDgqXh7tL3n
sHUfcOYBhCIHVFIvOovjTMSjga1JcImQU4UF6yiA7eW4qrJ9q6/4kmeUHVtvDQd2hwl1GCSDk/Uj
rRDbvoSDj5E+cbViHg7Mg4NyjQQAK/xp08QoTFGwyrNoYa2V5rrgaynZYOGopeSV0zH8wdDiXuQg
x4EhINnaSk0vOR1oLJ40pwFQZxiNVx8mKyeSm/zSaoj4f+zvudXLh5qWI5B8rdx1lmslV6FyTY0C
jncThlMLYRvnIu9PYwnh0ZdVreVXV78fmK2ew/ojyEgd4j0erTAu0xz2OdiWGfzib2x2H63gCTgI
ptHFiz2cs8bsTg/H74MNbV9898nDfYU6+3t8aAKk3tad45nZlydxfau+XzL0zcDR0uw7Du5Do+WP
47Bd2BqUsAgGh8VFeNmoAeCP8AxNe9/YKsZMBMyOgydcqP5h8byvq1Nt5WM14HI7d38GfESLE5rW
6TlJSWyoVusawGrWSAqTqVM6/Z8dkd3e3/P02Z4WibUQzE1FFP7s+GJYE+WmDV/jFno+wzNyIlrS
VVubL6f6DN+ILkTP2t8ytTbZwpagGvnhEE+B1IHm29JU3ABCXzz0TJF3zXxuQwwf1P5UbkSXBUJk
EmvljlYd3/iQS6444r6d1R1/8bC93AqgFeI0xOS5e/VNEvs3SwCkkVNjwp/xl9W/yKgcwjK0eVp7
V7YI6T/b8Z3m/ON4eSRDR8SfmwFL7/TVPlBoYZSWnJNRm1/cAtJAFlE7WEvypdNzGYCN7q/jxlDE
VGXdJ2tAfNaULBApZodjBzruETdPmq4DJ8uu6A3olWgU4nE15DScZPOkDBarlqMQ7nz3jaTyf3EL
PUZcfKBq8DZu+BxBK9zvDsNKQV2+oyHE29OR+D/3buTWnsVwQtlPv6gYpLhzawtCSwR7GfWdrpVj
d/IoYQm3QH68AOOePUvcnMZZ/ADtsd+ur77vKvBIQ2gI/m3BCMYpKBZTHDtm7PtHo/gA9uEdBYyN
oZvLAf39xCniVDV1jh33HeFRtwMx0VWaKMt7nWiLQ8JVlgbIdWnV8a7v5pyalfcKza6asnlhmDML
gBabWpPMtITkEdHlOWAKrQNNNDmKsovBNQpwmI9vJhSAUmF6uxuRd0RrM1q3MGYqm+ubkmmIQuzc
yzalZzqcKwlnwxmAKeKwnXkN1KAW1VM16M5QSUdScJyFJZdVGMHUPHelqJNNd0AC7A0BQQQS3fi9
jWV5S8sTS/DEnHIZCUrlrA3qk7bsd0fp0kmEvP6octNO7ekdoWl75O41654RTGn3gMLaNJwmBMKK
swcD2CA7OtIGvBOKpoJwBSOPi++SqCPJOxpfZnQsIxNmK46OsTXadfPPPKNX3JlYsELQxfTVVfKL
8H+genYMFjYrdCaX5B0l8D4//nwWamRdcRdKDEMVOfmgHiggzqIHtZmxJz57M2l7fRHo8GVRUjOX
TABerTGhSPAA6SO43ytcYbdcq2YGl7lZmuym3vkWYN0m78JUYi6KF+GiVs2/DmXGyyRlMoWWAB67
y6B3F+2sQURlD+oRDPAReA3P0qn/IQjuz+lskeKEpIaXfYhX/KOL1XjK2tpFQseznkh0IQD3q8eX
00nPhvdUhZ0yc+VGLDyvtVdYt+UQ2t95AM6FOrryJOVS12jaayNNyVDsOsbcP8YpfQ8f3ZKa4zQq
3cSSeiaOM7iy/DrjbQftf816c4vrLeIFk5JmhCtkdzpwtYGTqB4TWANEs0YRY7ZXXdmN87u6hwyJ
kB9aAZ4i1+3Y2QQC23eIL86W4qWTCCxdfpC/dLUhtj8dCZ23Lnp5JMadC56uvz6OSwc4xgtY8Qjd
nuPCbMi+xS+8dS+BOBXqC+XF0QCP+7JaqbsqtkZuxLjxKZYv+TLJd+31J2PDFkmY1WcC2I3u96R4
ePvWE3gN/oCU3x/ConpgX3D5xADgGKYXszRt/MUGwugHgtgm6u7u4umaHyP51mo6rEDmwVNi1bMY
+MWls/E8rS9ZWqJ7k9jzEJJqcW0iviD5Pt5UKcIgvnOwej+dNotWMkW6DKm/G1o4oyGn0HE3YSOl
Tub9X7l8lGYQBCTsngSaUayDscvlMVKhLGlSjojpx3ELsx3ElVVsijD4znWHlDt3vWNSU8hEpRdB
P07AYyxBwnQGll+aTm+/erT3bnrXK//Zsn2G8xMAiZxilNzJSnbgGo3vsRdV38nYVVV0D4wUD/wP
sUOF077ko52Ah66txLRoOTbdAj6DYy82K+83CXeZr3y3lKEZe7Ic6PApRGrhca2o4dmHzV48rUW2
JQG1GRPDafE72oAnuUx6vOsV3nNqREyckO38FTAsCHUdFX5UErIZ2nY/cspL7cUpkriDZczXOlba
7A9js6ICthRbEw46uioiVeLncKgbSsJ6X4Xd0pNtJ8lZLJkgzoUQIa3AGs4ooDTUMXUXDLuP8TfV
wfLxwxf2PlISMS6Hifx9UTApVSzefqjedIFb3XmOnVdTnflM3RIRGS6mMQPLp89Jm8VIQor3EfGp
19eqcXaepTYmNhWaOnEEN/ZibZ98iaBoVuo5Mt1PiUEhhLkJsMYNxQ5whwnv6Yo7ej0VYmJR9h3q
T9m4BDnVLZBh23CSvx3dJpN2EXV8TjyGgiLDE/AlCaLKqFGlKbU2WW44it4T4VksJcMw+Qn0V67r
pwIPjnYIvxmZeNBEqqGcVrq1foAx528Zq1UF1MdZJdlRlbGUqLrQJZjzlwQkvIZDJkUbaoBRfgdO
PjAi1pKZrzIOovL6vkx+JyEp/tOn9MIq6adjRmAMPiWmb9xq1lfkyf+BdgvkH42KVkox80spP2An
3RkW+1s0zZ//Pd7wQFLaio4TSqNEov7izqiau9nwPfaONC/lVQZ0AZ/UDgK/2N1E8MB9/s5/UNXO
OzQFoiG7g5jSv1v0NdevX3S3SgtmHmy+/AA4f7757OUGpxM1l54Me67ZSPZ+PToptkbbGWE1N4kD
S/8PlI3wZyCmvJhVX5ov4ebW+ZgHs1n1YtQGZlaOAYgp2nw/IDVlZRU9F6rcmKQxy7lI2Te2acqj
THpg4gASNYkCNHE/stIP0grxCsTlt+R4X0iq9IHFf3hZ3HUvPxgePFhP1vvLqa1OdWmN1vftOxiS
SXIGbtXmxK77VAA0j9U2ehrPUpJNY3FXtZ6Z9CtA42IkyUcGwcXlWmwKW8bb0j6HP8u+GZt4old1
r1JI0YTIEUST8ZL8asggf8WCjtY2Eu1WKuYnX2s9kJLUqrhvpUGlCu9GiGQNNIIdvlunQ1XhG1HJ
UXqiqbhEKw7Kw6QxYUCqJ0H2KGMCYTWCwlApafuDgISub10mYIaiE4UdZETZXDRTEhKMC3yAEOzt
0PxTZabsek4UMJVALDO5lNNrCffkIkoueRUvHs8trhQFww3wQcIbTJhgd83tfKjj5Q2t3J0atunr
vX9V/9xChV+w0aqfLnArgR9z3N0r2XvCs77Epu0x5vc7hS6DcfqpnuswoaA5fgQRQ8/Xe/WNiOZ/
jBdKwq7P0V5ORmb1VgD3jP/RE02Tkfc6aIeOED+63slUSjiOnqwo7thr2zNEzV8+91N/FZL1XUw0
iRTZjZHcMLdtQF3cwgl4sTtaQpofsk79Di3W2bVXLrdjp1LTlxhBLKgqKjMkFhjCsgG8RfFGiB9I
zyt8dfXQlp75iPTehLjsI8BLRsjGzVjqf9Xf7ceLlN1FbNHM8q7tjUKXqFHHw7t2WPV3gsAYPJco
n8M4puxpblmFVO/Hrp3PvjgxWJnrZ5nzHv2qqALoiuWcnwjrOwPiTl4RBrjlH/DBp7yem+S8NDTL
bXgnFDDreqO3hPB8Zg4qeuRZrOd2lMw0kIKM42wcuAcj4FUkcS0b/JXNPMh5TUUX/6MTpUPTEPT7
VRgsqsdqjLb044lyMRA49GByoImRpfHz1ctncr5/+Cp2u4LrOqcAijfXr1jRpyayPgjmRFqoEpEc
RRQzzpejGIttuAcORcWTjq5Ku/rYN0AsQOTLjWFwRYyXNUgXOMLgrdkbBAEc/8iV0eEB6f4XHQpQ
UUTc8qwsMS10n4+Wa9fPH5gzfMZb7sjqxyfL9FSY23zb+TNYSdEZatzme0cqn4etD/+9XppkwPSs
kbQ4LCezLi6Eb6nM16zS6wi/L1RgnPQNLZXB2kIOekWz6ccOyw/Tf1k9Y6PF+c9GwzBo40d0mHtr
IJgLfu+Ii+0Af6vVuWxHB0qtq9AARgbH7VIndCV1kWSmIuFSpz6n3cqua1QCZ5ly2oW3e8DKQKAi
phoHxWH6uGmUVYa9GDbC0WfBVC21vfpMYJKln+1/03dHR2pdthgJmWoEfGRB1Am7nYbjh09O9JSo
cdHSUcZMAtWbfgV5jkVfID1RKItEtQjuvWXVqzaomvu3Nnd0N/xIVKRpxXZ2yV9gV0CrPT1C9ICB
qAzPvHfzyjwvoekYrOyi52sViNK+FeykY104UhJhmFXTwfmBwH5LzJ/Lrh0NkVdMOcAFJQK1r98A
6e5ulAtydBrMaVYvi256p6d9mIrefJpRuhEI7jYYnEQBGqP2P9w9lVSCrRXnVULqYTqaROLKKjrx
B8hrKrH5Pu6Wej7S3ozXwMD2u1oO3Kd4E5NBEJKeEZOWy4nPISB6EAIAnY+Vd7p+GEkqjwUQALOW
RtkjJpBNv6qIQp2bDY7jOC1GkFdmbMBcdgWluBQTLvkjKS5yGxgf2AQe7wMSefOLrQjArDZ6OCgf
rx+OlCTHm/X9yZl7ZVOrv6kAlQFXDK2Aie4eRxd8fO7Ui9K/ULIkLqK/WgjLJxXgztDdOGbF16F0
4Hs9xGNgZrhlczJqtU+AqzfS6MaZ5QTPKk1FW88KJ3HIQL+hOUHOvfCHcDlt+RiYsedCQ5M2PoST
DBPh76S4A3U8iILPIS5Kg0vZLm30GVev6LIzq11VEp/GJsYAdc8QwCUIRSadgnRhOFNR/+WnPv9B
EeXIQllIDTTZDCzC3D5EZOxaq5R2mUB4ki39493rLNq4hxoOTTGRIrs1cusmgeqiG+lhDO7UcJyc
bbfsszpVLeFWAtCcKx7Aefgn+kWDBtImT02LaOsQaddtmIsLbaB62jv0cmtAdnjHZokVJHPhnBeb
QZg3ctr2Nd8kERB+f+kf6vNkXQPrvdAbCusdSmOBboEHe2ykq1PPFfk1Pw1asWSEqEUetBAQpWls
4IHgGIiGnZzt55/jJfAotPdfFJMMC48kEt0fjsDFtn4vJeuRH2bO+WAKY3SaclpKthBef7e4EX+n
OZyE3Z/hpOjCTGX1rXa2Oz1sNabKLukkY3yqVs7Pg1l+MIQZuUEirSkFnyps/zni0cwzc891TXHs
sRa87YRlT0r4aBsZZUASHGD0GZhxfVbjf6kOvK5TjF8mMo3ERN4hEBKrr/LGDzROh40Qee1dPhVC
Ajuss8yVKFMQK+dCupFvALSjtiUbTgZFFEgU+lWN1Lcg1zyVDyZHhF1taiLzamZfaCtQQxBHogS8
LN+73DpvsHjCpSqc5SfcXZm6uoqo5gGbkso688+d1H5xE22TDI8llnfC80qU3/DvaLQQZ2IGeiqe
qbZ/qwXzhKcZRch6dfr6Bymu1n2ys9yQtnLjYF/rpbEF+mhc4vuMjrn9S5ChlPmNlE1t4NDkzrcW
6nPr5nP+aVA4a36ov9Uy++rX9BY+oXl2gtTEsj53VholddlQ+yWc51OqXhyOot9MTa8gJkEHUIp/
OXonKZD65dEmMkOsUeADLDSu3Y4Rg58aoc3Q/qOJqMyKgtYGC9auLAtl7KBZdJJg9OlPUjVWlY0Q
ukSk8i5LrHMrBAoj+JQEfsCurPB5uF4HscDJAHNPzVS54BQNrvlE7tWmeNZ7rtHwyScYvWHQLs/V
p8XoM8Gu0y4YtaIkSnn9BROiu/9QNE85Zo7SxWHX6S/lDu7OABiSJG2jccRbeBNjtoSM/VXMkvJJ
4n35ygsXVGZM9Ap0QT5pJu92vQnDffJKGtW1UtDZx0ew1OOR4cg/KXXW6qCh5swVNnoGdLAKXH+X
7OdfoOd7sTrPaCHDm1ySR75TpL01L1M+7vgXHy3uiBd5Jg8IdQMZq/7NoFedBRMVCs6/DWBHVvkA
+YTOZ4lJgz/Vz4tx9wGVpmyvSRKZTQRQN6OhAo5yXGWyxoHPb1q3a6oly/jIF2Aky3HObpGZZahc
ZUHrqHWzzYfKG8uhQKpB5NJZ0TsrMhj1TEtZ7RlNC7JcaF4rOFvOB0pQrK1y5khAKvGfI7R8VK00
OzrVe+v5sqNRCMmGjIKHfcBOQwxWxUoKZITQ8vv6Ei3+kxY6E6+0kwUENKbLbNGzevx9TT5sFyIP
mtqdPCJvYO7bpyepQSvNwpov2HPKwaC//+ZxYX+I16EKNAxUpnG77URkygiof9G7yBOJ/WYWiGCr
ecybT+ODiEKdTf10Y/jFvHsEWk3wVNNs+f+hb0VBnmmfh4h1oqWap4iqamd939uLmDr0csPfah+O
Tzz2PgSatynMA3N2Ivet/fovpl4HYrDnduzMniSF2+8wRooOqLOkndUBbjOw9GQUXY6jGptfnbbK
5Vk4x9ljxbyx7+1Gua7EQmnk0pUklhgldWcE2mmolHQ5vMp3YXYv1Xq35XxhEu6W3OXR0PP8VrJH
2d9KKfQYvNRYLa91Qb2LpoFQ+OqE2zwQVklKNq2cvMPWXefx3e1ZJnLGId29FsbWMwhXCF8AqkFL
wD4pPvGAouJtHlE9qYvwnxzAwg8QU9u4cqts23eoYeTQUe8msHCe2zn5igyv7gc7jO77vJcorPET
B3HaAPV4HqZfG0wORBp4JwP5A0cnW3Ri0YNN683qULQOgJUnIM1uRdSStKrWE3c1JKTHuXWt2CdV
eW5AEedll8Lu34AfMQ1wzqtfVWNCSb31OQYOTatohCMgHItajkoM6mPZzFDkO6BeygoXlOM7O3eV
q/fKE2ThBzPxrW0LL7q52SWNlZqzUZ5x5oh+nDhFnO5HM4cJXCu7yUOLptGZLHiszTnJBT7qzqU7
qs6iqZ69NxRpKPZQ9AdKbV9EUzUIkmhds6S0OJUbzdeWhPL0bz++PEWfXVrBNq5yYD73gRSsDZIk
IsIe0TvOEJQWoTM8xSYg/WJfzWubf7uV5kLsb4Y4d5xVetIPg1SDaottiYmhMYDeUysUB9Xd0l8Q
0AseQ8OW3LDaeB70H8+Eb+fe/Qpi/6Tsn+f380cWJ60GSgEf10JsdXha46dD/tj9aNVm4l1xb50O
Lctn3vRK3YrtNbNx1m7F0yFYxwDD4Sisfq3EV9CTM0yaXf/ZB0+rkGJk+EJvHbxacS5qvAqDrcTN
bx8vrZTWEBoW52xtipmMVNtUuKU0jkMs4XkWNFeP85C7/eS805rUtHyIbLd+nM5N0pQIebtxWdzk
/lKTvIveUETYLxg3FfRo6iXconwcq/9QuTXrLqnjCYlm0Ka/sdMWhbDDn1E/ZUZQx7E227XJUG7M
njd/FK+pp1JEKrhDE7EJfqeII2Knms3Egl6S2MQYYqMA9WaRnTzi9QrejnNX6Mo4fxPjk6X6dxzp
4IVBvmdcQAMewQCQdYWUOkUyuc7TwEc20XWJD1jo5Wz2WgNl7wCCkX5wNqdvxGtXzB/zU1nvTRQh
kxODciHQQujcEcGLO0/E5M09oC7eEyjpKrzIL81c9EApZOmVrNevZzJ1eNRMQYHU3IQpGD1idCpA
Q1nJIJGU7EFkRnvKPJ2KIs2HTyJ+GcEeYUvEfCQLwxT7xDQsOpPPFh8YncZ4z4cD4mpvpVizATqL
/cuB3n6fQeHIyraZwb9sE+dLJLDouYbIUi99whBt9Uw2muN+Ofj1lABmZlDtORH/XzMInIq+4Cw0
fMX3Ijtcb+majARFA2ZWdmaJE6a3kxqIrv17L8tt0Xji9lQLcxA9ig5o54bkLD6WtZM/yccMA86H
wCr2Up16r4RtASBQ64jP/9KpaNqs0NLPO+0ttUA8ltyM8hOyj5TjkwAeckl0c23WOtHNQ0zRZbIQ
YJok0PppyHoytKPI/bMxU9loYlOmb+ppScSnYzjLe6f8n0FMy+Or3YUJRyR2HKwbH8lnkb8eB/M7
GrrMVFkxPx11OMUAGeH8uUvZq/uf3Qwhwnk8JD0lPg+mUMVA6tUoB5Mx0+/eCCCkC322TWnhIoN/
zOXTIMIVx7X+iP8u3KWMsOzzv3BNHfpe+3ShcNyBpASWOfFqytNCw4Kj6Tg+LjieVX3YRvphndS6
wzfmf3NNWc58j3mtcFIB2Jh7u+sRu6n/mScli2EZfeIX7SJ9MTk3+M+eBX5/Ck9ZGv/tix3MK3AF
oaNtr2eKVzQX8FuquSBbRaHWQHxBLcVEtUd8HrR4lMereV7gHKnuoWtndWwNB3ihfLOE0USNifs3
46fYwtGeFGzg3ZqxBvNWgdy61huAN4wi6QWaih3en/DwjV7H281ae9nf5iEeb3uuemKK0crvevf2
Q3/FjJD/6/nsRcpwPPiKRAnMJV8ODEYyhiP9/JH+h+8ww5bEEQFkUALuMmr8v+OrMmTbgmwupNpf
BBbR5UAuVrYQsuGX30gOC6IlRTdnzpxL27qrZ+d/0S4gX0t0h26HpSholCULHJqaAmLSokix97z4
WZX6YwkGyGMlm5xv+Yx+L7Dhizlj3R/oSL9f8+sDSoPRyZqIANqwSb6d1+IP7swRROnrnOsp2pk3
DUbYPaY6LE5ONTbsCkQzN8PvCD0CsWSnOzLI7d7cTI2jicbWzX02BxM0GPW47PBU3iUJLflR8LCj
kI85b8zJKfYsZUWGL6OXz+gsEkbP0y+oPBJ1MkkEHt8zBINRZFhmJEaRx5GYgMy5l4MbzTsauwX+
NBq6zTxXKRXYhLTkqTCoKbtcQkp4+wbmsyfqEYNLIP/wrb62c5xYrNvhubOflbwRTj63xTYjz3/b
MH0gtKVYa+9OrUqqXU3XzQuqvz0GWAYbygHiWyzOgNCHWvrZ8+MALkwwSbKHZxUiSvZ9MvBJsL+o
qSABVDvPTEBcv29FQSOghYsNh2q8L9L9dtxIvDtiIy9/YDLKBRj74z5Ha75C/DpFTSELUpWO9wBk
IRISMcO9v6D91kn0by4WqM4/H80fNU6wCUC9iCKe8jJZ1eKmiT9jT3c94DIDDvS3G5oCyiD11xj8
VlKnPhsBEvBH05YuZggwZlwo+NsWGXe2SsvZ9C9yP89GyCVBNMFoodkg4/USVIQjBeWaRdSEqSQP
My+xifSwn3WDiT6BzaHnr136Beou/JJuJ+2MtcrzbwKiwwq1Mma6eHvxW3yU7bFGwgErUhKNJiY/
rRGg1ZZzWeoAkCsjHsegxUY3Du1A64IyGu43n4T77vFLM+yzNDotosM31rVeeiYk38ofG3dC17Ah
GjCSRNca854uI6HJYXvcrtkQO/EIeBnYu7gdnJ7aV+c/qJDe2tI2B62twWc2xV+U9OgSKv5ScdbU
6WhEfLxT/OBwcDw0gSyjZbmB3WD0J3h2KDzJ+/XLCvgxW8Aca2DDSd+wHUrLPlrJJAsV9ou60X1C
GwlTExmNvaRwazZMDIQEp+XhuBuqoAmbFw4xEIMrlfnQGrPZc3NkoB0Xw6kaI1LUmpfYXTnzZlQ7
iXC2iM29V8LdzZ7Heea/olrEKxIJ9fjUrncmegpFW3bEArDDlnZjT/ci6MtyRR5bz8aamthta4n5
AZGaZd2cHh/7+uwClKPDhXC4K18l7TsW+NSKwbJDgdXX0h5qRMcqRM9bSC8z81iziR/Svu0HYh/+
rdRkswFrO3rpJA3JI7AILBo5HCVxYbYylbKnwuREyQA926jAXMubKx7kKFQdKLXTPTUx7Fzjen12
cC18chCKgZEMVvmXhzlsYX/xBNG9d2SWGGbjitQoW2X/iYcqRo1JPvxN3dbFUb1+vezOhvatUzKa
BPpwKfZHbkF4GvXaMSG98GVqdAtpAQ3eigMt91AY6cZw38pzSk6NlN/vDxKG2vG8B0/KoAcALRD/
x+4XYT5mg0xJDwrWPb645C10mceFa3d1BhVfESQkof7BTtt9tW7oNCLyMIuicLOG2RX5UQF6t7dB
ZRNj1/Xx4ocZShm2FtT7vx6YihWGWGSacdg0rbV+UqJq2gf9jPS6PXRYA6v3eI9kxk6iAriatVt7
ImZCmX+0CzjpTzOKYRoew+vsV9OUSFS4xeaCTd+4fAfxtaqJCy+iGienHUzvX6/elk9LaqyROs3W
Gu9F+uqkHNBsEPOjb/czy0Ss3E9XpUipAXLw/HYNoDcJ/KEoiVNiTqxHIlWzWiGe6bx7xTbnKOmV
8piRDXybB2QU3TSLEV+zwL3tfmh2ISgKlbrwHJsa0wn5webpvTGk0igMCiCTUfw4BAbYBOHPtEUu
rzEJE93Fe8FESRdx06gL/SSkpJn8lYdIWOI3C+ASQcuNu7LzmWeUJBwJ962vd95vpa5q6gKY2dVt
rRQdf2B96dlVOz8R1uzSYik6zcoDuGb1Nql1E4JzZ4B8pyjV0H3TvGKx+wecbz89BAVk3wIDDmR4
AAL3aD9ru5uYCS2L0ajWXzfuD71BvD7i7XxD9Q0gK3UEYxS5ajLWa6UDSR0GdkIsR+FQOAxZo4a3
f7ZE6KFdh59e72jUFHPWLy6yxOwuN0K2pN4/rGb8Tt7ZkM56WVr+7E/hdWtxdXKBuDgyPNY7cEe0
BKqkrXTjCxKfIXnyWfR0kX62+PT6XrC7bc3zu1Vbp5MvWmHQhKrngYHbqnq/kCjAfywFpGg6CP6c
b3KEYyoMVOFadPUm+SH1K3n6kj7h2stxTZQZ6wcQWM4u3lsgwfA+pgDfnHyx/cCpi+aahBZPH6yH
WflNjbuOtY4iQO62NcGE3pqTSYyJ/dwt3pRGFvZG/yoCwPNSpkDw7X+1EsRZYCYsPQHnr83fu6Dq
9M6G01ysYi7IjN7o0lbCBUT3kDsj19bDLKDdkkjMc/0uUML+XYydE10csth60ZAaO1DWfPdSMgiq
JcWTbZNuFK+fEA0Yk90gMok3d/acYzPedrico3xP25luTgXzJ/sYBmiwP5XKKQHfbQyO+fuPpqvk
vBvQ9MSHx7ADivBC4KsvkY2AFeFC7hsWhxtSZUKM8tmY5o3+yhv98nVStG0MexJedSk3Zo/EPdNv
HaieGyNkoCdZ/26Nf2kE9mnf8WMKJ8LuXai4f0GjcSxPxYj+YMY7qa3dgFrU9vIuZSmwV3Gj4CND
oMpYp9jOmyP1NZISqed16t89vHlN2tZAC7yQNe6axTavLnjhbOLES9X1kCK2PGjvQtDuDXeWxH6O
K+i5Fq7WnZz1oJ3y98TOdiHzUOatnc1ozQwZaGm58wjbcH6/IUAnTZCtx2sVlZmB106foesQyCaR
GqSElCxeF7Df/QucmrJ6nMvziLXNGt8YgSAvcP0xb7UQWgzS2cHE9cGC+AVarwXjI67Vz1++TBI8
uKOICQYyrrJniWaUGx0Lgm8ICnFrfOrUeWhgPs9hOpp46+7h6PdBQ6wS62nPwKF+fzPEMyPRfTTA
NvXdlKgwUB3Gr5FQ8rsU+Z/4oM0pBQCLot+4naxo+SwKBs0O14ty86R8Y37htkxJO9yEFOmPIU3V
xn3HrWrWCUf0zNOqxuJRmViht9SyHxSMBKmLHJjpuIC4zY2p0aPR0D9UT4y7C7+T/UNftTknp0Im
5iMJFYG+ud9CdHSKRv7UPVmgYPGYOjNqVpDU3ybmWIWD/idolNlyh7ArbgHDoHzqlfLdl3SLn/EW
pE1GxKQNfTVpLass3KJi2GLPWfZ8aCjnd5LEvnjndCQjbvhXHAOqffUyR+hMOfKG3kcsPLNwFIiS
ainkHAsSZOmIic2UhagmZcXLPZZ5OqZk+ru63rSnyyHWw1b1VHDPO+LnrItHNkFF4u8KZ83Lh2/Y
5+0gBrBLohiHRTrzN8NgIoIkAt6rxXai2iSSl+mvkfer/1aTw9slkISpuxlp52ySXUywlC/NoNIL
bl5vft0WakXk2DxL/kRAmOgZSFiW9ogKfoUEaCPoasU1t4EAhXmU+ya0r7mDqUGhwCOVwLFsutS9
TzA0ftdo9yywoxYWyU0ug2nCAvuMNC2EKjqpEke+ifcoMiwnSkpFoSELSeBLVzbU8utqZqsA1Je9
eIT7Y0UpY7za5ybF2mV8iGidVem2zzlzBCU3aC+MjD3YieGsHdb9FNXsadGmWG5JXM2mDg/t8Ii1
4OWcRxNmxv4L+OLb9TOxgZ/KiLzrdWGMJyeDF9fIuvfY3sMlbdpsX12838P/yiK+n/mnE3D8p3rM
p/7A+anYeIOPhUCwSUPZiVYIvAibubvJqLMB1AtStlHEHW/GZcrcV8wuuwVMSqMdKnJdF5caGthw
2GgodYpqaCVS/PhJDcZBLAhv4RmxWK8UhZpMPw36n0r/ZAqPhUHNf3rvjgePGZKf/a0XMGSFnNPr
yTs2lNe25qJlFFZEU4v+y/lO236a7y/DNz4Sqsl0ihsAbjC9VrDoxCicqJW0ebYcbwhtRimdSn+c
sEfHDssZ04AveEdZ+6XzhVNZbwyP827COCCPBZZ7Sh3QiexGzKnltJD9YwyJtIj60pMzSiQC44fI
1njIhLy/UTKhH9abwhDGUNo/3u0devaNgsewQmZNJ5KcWnFJFGCCidJIGmdDQLjI+QJT9o64c2DA
u5UxM5z/yOn8tC3aKtlWHX4cAzxQQQ6hik6usjqSB3SHuObW1+B/jmymL5Sa2q8aWExFMMGXkOys
CCDmhVjemwFVdvzaD0x1Tl29kr5SXahiFPiOlV+SY3pPl/qciGbtZ1Kr3vwuqEMeh4D0dXRYrtt2
8GAnwBDuSy4fb9isHIYfQ4RHo6/4JNCQoW6ORkcHubK2GSm2KssdV8Z2SHBolVuNDUQqoq3hjRBl
Aw4HzLwkWC7DZLGaYR0Jtjys3obH+bX6yyIKDW5+dPErqbbuOwxeLwmOL1XBVmQEkd1fCmG7/b7q
sAwXHeYqxNdbP6YQgpVUQyUGG8uZN4Hgxtxl18vQlKkFRTO6XfW/xidX7owWp+HsR2fZlE4S4E1f
AEA+fQaTptPqljf7+C5VF4MIVItCn9FVBlx/0D7Q3wIazQqyXWaUtYxPJ7GC1kVPtGEUBZXJLdfh
valw3n+oG2/b87nc57ZL8YAOYieoEb8SH6Jn/F+C0D8Er5oduBH9IEjHcB7d4lk0t63K9syOh+2h
tgPhVaaMWAsS8xC/Eyn+iIt63C67Iyz36Vdh1bZLmzyxNmBkBIjQeiA2nPxBGMwsBAPCBTCyrRB7
IetpcuPzRU08mSElnFf7ldesXqrY+9r06hHUU1+W/fNJ2Kerl1Do1nUhbrF7BNOkWjVY7RjHybgd
RimBoUrmNMFwhRGsX1i0sIXcH6MFzKBILViwBLYMvdknIbX6aasRMVQ5/ByTefKfEzN6kuLLP66V
bH2tSBQX7hfquuImOIZMikwuBAhuG/jYOJvd6OD9xwI55IS81O0MMU5+SkfFLO+iQNBE2d+dlBKa
L+LPZwq7K/0MI12BkP0H5ym6ZXy/YSa1RXzgA2fOW9+IzzZJxllAlrOYziWfM5xvY1Ek6MfzHiXQ
hcAzE5tV+iPLDHNI8MxTTPEJdXKEbOm23XZqhuPJd1AGJOLjCILPrgVGm6W7xOfssBcQ+lQlcg2Y
Sb6nJ494nldsB0j2nhAB8uC4/AIMqoignmLsO13bLsRiwaZhS6DxrGgNA8kKJlo5No8vUG7DlGPl
verhQwIAJWOfAhwJNk3QVNDwT7KqySIe4H4EZJUWy68Vo7QJjDWfHDaLr/A/Qnegafr1vaPv53Lv
p95r1KSpUslKw07E4Erue5Lppixv9g0EwmUKMljEAHr+sdxbzilN83yTjSLoGojEL795tap8vL9R
ZpMJuVhz3TNX0ehA/fMfDCXa6vSsGkSenr2ZovHhDlRSi1XuWAEkxldY/ThTgmI2QdrJxKOPOApV
e5PAfN9tYvjXga3Ybjt2Z0ReXaELIRgRxLjSohbSCB0rOA9luXEPMlTCeRjKp5hDvEVPYs8Rewrp
Nz0Gqj7x1nMFcyc/C+/GFSNZeIqQ+wRRnkjkz+ewt5qX3XplkpklreiqMk5B8I07EYhPhiK1/C0z
BxqEcaz1fYelLmHBaeH+8cE+JLX8LrwiN7x01hWtRKXALPyk/5vcjYVbsGEaF31zI/+NpwBdp4pB
CPe2KbjyCL0I/qrEpYVLsmV2TWlFze5t+uuTrVolVEq4q0a5noxzwRDIZBtPCNEIwMAI5/PF+4/v
Uz5vo8UbFN2mNQwoMVeTkHlzXDrqlS3uFT1x6OM4KvsfBmHspWXc7GxiZBC54OxlJslpdCbW5H0n
M09tHx+lJpvz8/j7vVeK/g4dGleZ5QI8/QZK/i3dnMzYWlBIV0arFemQFr3U7ogbwGoeKK3MhEDM
nlrm8RvuM7jXE+i01K1+yL4ExJtTZDbHNBvMD4no9STcsZm74gn+o54ONtdtFArRh2a5scJpZNu3
TfSBTu+7rjrJdqOZ+7whQHt/iTXO2D26B97kAc+KhroyU5y0qqCrc1QKPPXrFzRLKl0rzyDQDBMA
9myAGW0h+ElGLBWLuUCSkLiENp5x/1lMjefY7kL2IYwEaDtQx/liiKiYg9ltdHEg/yHbFfr1ixRE
k1ZxR543CEA49ga6U3SjZiPSr9N9aI4ea/ofA7FE9MWzG3U5LvAVqAzLl8NrQAq6mv5w6yScBgUq
iixjSAs4QK4czSJ9FRsIMtOOPXV/rJYCn94+k2DrujRMybeid6vd+VAbVk70NDMCNAitA9TzWv+J
thJuzu+NP4MK4YOFXMeZSxJoTSrNLQG4bhIl/sa5v98Dnv6OO1SVp7RXX499Nex7j3HWJa0Y0i0W
nVbJ2mgCGS9c8NqU+W8B+DmDJyN5OLAugBMPBztqSewZFdqJPLFNHbFK8116NfiD/2KdoSq5OfJf
P47pvzvtUi06UiuHEh/mF8/0+99xFb4bDxopf+8ZgolpClPnDo5yNj1C0m0pzXbX0uIPN+M7cpxO
nCa/CZSk+tsARTsY9RQHz9hVVN09qugMcerTCxXmMPFEGRKkYV3mNZK68nzdE1RaOMBu7b+stzuo
u4VR0hT6C0U9+s1kNZ+0NIIjUUfSaOTscugmYXBZ49DO1wahCgtf/KlaF9HHhMFlztt7dwpp0Erb
ksm6r/pVRcAqgzxxeJtpXiXI1cHeyDq9GWOqOr+UfguhNoaVnGSSCqgfaoEXOZbeqduhT3cPw7md
ZEQ1uS7+23azW/MgV5nO5NMHP9HQ8uCoBoLw/ccOvTWXXXK+l5Um1J0HncBIC6ip3zfGIWWMoR9f
pKP7+a8Z8MTOjs8gP8ijLhnFbD7YMLKAPAvLsZb9eMGpEpWTki19UdTNcJtMOziYsOGTogFpggGj
9QFvtnkBnpT22jZ7JO/osXLQ70utBfq7sqvc3Y51JzspF2kKso8mB4ceOmqeLV9qGY2813MMxI1u
FWKfJ0gYKHTGhoFT6a9mcINsyZ9TzGxvrQcUs2lEW42dlU5+YhRyF3YQXKaVz/OaLPm+Vwk97upY
XMYTUGPKdKM8mk9y0XqQIGQJLUZVAsvjyv+rtD7S0UHmx8SZbdqj/Pmx75CF1x5+gVxbZ/Adtwsh
b+Vu1V73E1csmOYEYZ9eL1kBQdboj9Q/ZaMK/booWIDjA+aNxU2QQj/jTcGADl8pOgs0vJHssyck
VMIQJIUeo7go1PRuqV40GX3EcXbBGCIxTP5xpRrGikTl1sJi7tJeRv+AjGf1lPWxHrzPy9ojMLTj
39Vh20XHz7NwgFNx/MpqeBW2neXXBk6fChYOYKgv4v79lfU78xHeuTnsqxcEpzLHd45O7kjv30lU
y9/EXJbTMR5RCWhm2DDBxMrl/TqS0kv32a8GGCm839uSXpwoKb0vYwxtT4BB9X/jXAxwq5OTZ9s+
cQsafPJ6nJSaUo3j/r+1TJ+XV0lq2paTbCoJ8UOLgdsk8Y25nO4Fxc0wrG8oZzl6WDMYfFZ6HJmB
6ZsdUb4VwqHcaYz7wvkAicPmcdoXZqfwi4kXXFgeKJpUicmJXDUa5Nfjuj81FvXASKTnP7Eqz4tK
cQuhWfjrzdLDy0wItgtIXWvOFpSBrRw2g8nQVWj1YperBvbaw6s1R8isbG5gcclOQZYbJ9IM2831
8hdy3TpWeGzeyuDuCeFudYU1elfd9faKhWl0NEar+US8BsJkP49hZTNN8+190SxyX16xOaluXKtV
hE+ALngzZb5ECq8SsbCcuke3BO5yhcqjOPCJHXiwXK/t8OtEaPEFaiCpjaL/8sYYyLdsJm56XFDq
Ldptp3smoDKguWlKSGZt+BUf9JWhWwNNuFD2tfRg8zzcDbF+DLSPtAGKpp+jVVlxSer+hnK2X0q8
EgcaWZicpvpZGQbNg0WI/d+fsbiw1N1hGVXD6Di/DQHq6OmxYCA3pG5NwC04OB44NoBciksBsVWj
cb5L8ti/VbLKRbeGnuWDvJgbZmg8eUbIZqRPkPcf13iFZVRwiKbMyN8EU2mQKDLjodjx07i/CkSp
uEaLCZWbuy6b5dTi/1wN4HuSrntpm2qdU/pV8G5SD/rWDXDn6mI0ZjKrWpYlZO+d1r9ZF/VAG6/J
ysoX0jLk+6N3YpA83JR2JxFp5QILkGFY25LHf128fHC/jdZGez/NWnjsfC+v5jIw9V8CghcGJuys
6dJYvco7fD6oavNaPwKAqHEKIWnzLFMW059dil6/kCc8n2PKidw7qJLst7SPIEX4hgi7g65i19wT
4SkSWvYd+08I5zPmWgV+nZF/Cn1OlgOcTnQSpQkI5ydf6meDXZQXyWKUfT8m93z9mfmGW8a3ulF4
+IxKiaTjDfAZG7Jxf4PYht3ddPAq0bUzh2RohNPxSuVVzz58zMPU8dKZ3RTBeTT5RFmj4s0Qb1u+
vDEE2Y1RYNP+xZ0/EvuYFHRGUOQgzVvueo1dR010pYTxQKZNU2o+rWPTAaLnfopm/Eos5r4G6n3X
Avh4sZDmpsS7EW61oEylmZKjptm6uY0cCN7H4jOenTUKC+Mdgp2OsijN19v4ykfaCFPKzD0tZGsD
1xyQFDBBNq1RLwTDPv4ZMtdZANdnrFPN+RujF5Vg8LRpnLlmCzIBULV/Un2wYd8P0pBG16Ajkreb
eV5G/mpqYKaViI4siVrWtzT4c2hzpIekry7JiKdg3+ag7OloP8dtHCBozNo6Spb5JJV8C4NclnC6
wI1+v6kGR3ECoUcKAOmuR5W9y7/1iSHV/MPKKQOnmsjxUsWcNBYnecxemWfPTpQnIk6ovqvEHuXI
6mSuV5IHNuIHEorqwqAfR/xWd14s80Izv++ff/DQmWDTHKTTRrcUYvLqqT56W7IRbSOAOR6DLDbK
nFe2/rXj8cf8iSjigTiQYGOcKmDyTUL1YmSdqaTbmno0FobkHpLW97sNaXS8ehCjlc6PcKHtcwJx
07PcSOygugvs4r5CTm90RPE7bsudPS/iaTMjDxxow3YRa5pTQUBu8FPQPFogaR6nfKRG4puXnSe6
lQknW6tah1JdcmRHxVZFX7A3qd+6vaDq0pyljJladTqLVW5kF0FsNI5LRh2brx9L0ZdxTxJMjS4b
ckYhmnpiMMdgzM/Dxl8N5YnRQfJP9ZK83S6n38R1ky1RN2Ix+PcYg5kiCUCiG4C9kV2j3CTTQ/eV
RQDUQ8JeZgcgsXe/MdUkRwe+o+jmJvhEJRLYXNR3+iUgRi9EXfv9ilhU2j0fgCpInlzKSS++CEBo
Bb8wfngIz/B2bgqjKqre48wEtgAFaVowNa8ibBWa1eFrPJ35U1tAjSiym1tAph/QirbxDRHcgZOq
49QECiPJPLsuXi9k+CJ8jgX5T6wfPq+GhpnERmCMphkJ6q5jDFb1scPaMX+VGk/jNWegEJO1aZ6p
pTnyV5qH4SMEQVD3+iY43vzuFlO3BWOvLwemWoyhVaIpKj3ya2QPnLFCPgZ8fnykm5cNCTkFPTAg
wHUgYxhwEwaifn6/bSOeQnToBNVaTVitxsZifEt2GUwlOLtwTsUaZUZ6hsUDLcvEptFcz/0aZEou
jpAZAITZUX4Z0ruiIJqUPH75IYmDkcGdRn2pNgKWMqiZCyypKrYulYSOG47C2LcGJQeyJIvqH2VD
O+h7/WFlWSA430xLj6ulr++NIqmnMD2wH/WsGB46Ka02wh58rRbsd5owaryq2G4zhSSePgj2fGSJ
MZbntbhCeqGVdO9wyg0XDlt6NkxVLG4FzKHOScb1vV8worUVZm0nU/O4wmfEiwM7GZ+GQV7IdlUl
XF7EzzfI0osiXY4NMIvmBasbPDXvIY6LZZ25cFg1oGP9DyS788k3GOu+968n5PTARNssbJjwqOLH
y7ChzGbYhKnKiUbJs9+ovWUvB05/whVXGRdQj1c5Kt1gdKmY4XOv7BkhPIa6eIC4oYpXpMh0+FHy
WbJqgduLailaiExCKKfTbz2Jsam7InjQ+s/JM19j5ZtKHCHEyvs5O2jegaHg7U9c0/aERSwaaG0u
7V2o6l7lAN/aNTC7lXWI96ZvftVWuRRdeSNRUd0BZQ5oenKk7R7Dq8cM9iahINGKPdfxVvIFfu9/
UJ/MPweZjafebLj85B/01WLaXi+j4bru7jzvYMwtnBEACgdYu6+J3Hn3QoaZepKDDawhoHbhH/yb
r17GuT65ZqP7k4eR/X2BcZGVcWJjwkKkvHkFx7xpVpIV9Oi1aAill9T911sL+eVMQy8dNkGfVMaO
19XYL7Ml9O60aJ4KLTbtGwPUjy4zSSCeygnHOrKTv66yFabUJm1yLbpMb06r4a1IJB+vGE3xOyjk
z9by7ARN0owInnuOEklrpVI/H+8rNZjQKEQTEY8PZqtXVKi81LWtGHQCArXsxA54z9s82g809NEr
hRTPvogVLIojXDEQzvcNcfV7+FResOETkW5zIBC4edWrSJcZ7k29uRNnHMqcGHCm+3zc3ImjLkxF
aXcQAMorlUOG6HyWZW0LrARVSZaDe/BnE357JHAVNyyQc6VDlzGeOMVHwMvpOPPsS3QXC3ekiC9z
bJQTRebY8X5xopat8fsiyhSb6l8dg4a9SvWtIKaN1K9UkwRwld1IF9Gv2eUmus9pgvWnngaDP8EB
dXiI5aIWGqqlepAx1DrXwBo+JGJyJcBxLTYEIjGCvCtLLaMhI1nwcFjCIui1bQ6s904LFn99VkGZ
vHcr5Ns26jqVAAod+AE7e+kN00Rv2Kpbby5S7wzy8zjW0ERV+rfJJYMBK+8FCI4Hi++EapuJoHOJ
W5NG94cso0uNtAU5wB4AouGEC2ajKarM65yAlA+7vq19o1dacxvVE3eedutA3u9qdRwFc8G7HzB3
QpiA1IP6IovTBw/9zU/vTaRFkicJf2oz+KvWKt683HZrmkbHyQYZVuhjeCVcDua4wlnLwHk9CSRv
a7TqRH6rPmWWL2D1EalaZzcOg/C45/mmr/XytwM7cZyc8W6/GpFD5YjZWRbpo5g6SNBGtGq31qWs
nEzdp7UCPb5MCOETzimYsrO6sVaYDq4kyAWOsKMuCib5Ii1yZ0NQr8N4/bZ47z77ueS/fYR5YASl
sV116MUPweZjXf5P4eUQxZHRbcRxsGhkvTU4VKI+SQ/wH8ijbyspZdZmWAANZ2Nl4cY/DGAHo/82
t9dlz8u0ewitzmADdgcZ+j5aPSau034/0Y8AG2O6LaWN86XfLdvBGZoDvs9Dfnraf8LqXlsR4Gct
3eAWrJcz9CJriUjS/lYEaf5cnedXgsrCUO3Xp+/tyE/QKGeBHzBmBkUpCZI9ycHol0na0c10t05Q
jeZ0yeHNJhNgY0MfdgFquE9JO8Xg54IAJ296FtsTSZ9C89BMCwlUa5eyJaMtUfuI2yWsF21liArt
K+rDO/XazzreBhJKFN5+9DWmrKka1B2/6pbwrqpBOyLYpJXNngT2v21HBUnHQ1Zwqz379RH1zuo7
NMB+/fQEtFjRCb61F4JQ6ZpnMV4jP31j6ZImvvaYcN7gfRqbHYPBEBCBWVHj1lUW76vvZYFO7aTx
pVZYfTdauZw2LrterZMR8h9EV4PnrhGZ4mx33bW43jUgsJAwP36xJlDBkZgfAKIOvpkuag9s6Q6j
4ejV6fI5vYuMtKVajAHzQVwAnXYg21BARoc3imaDrjC1SVmt4yBvxjaoQgpQRx96JmrR8kPqK5dE
ulF1xztgQ0Idct2SdpWQIdPcyf5/9ZsEvWLgtpRnQiEnlDjSoK/9lGhpd1STbKtKqlnzP1K0dzZK
AICESHjnWMjMUkxtXmTT1msHqUkjGL8naNEaX8J23klvZDrcX5ipCRhBmZ/zCeB4hXffeD/QI0qO
ETCDiRhdGN45MOkkRGm6tX2H9taw0qBgBQhhuf00vfuyqaWsY4FPI5P0EkkZJSh2cibnwvnqDRCY
yO/oRaN5/aBLkwAJ6GjcQQtpyJnjDgAx42AAXwbwI0a/iZFC3vJA3ZesFT0ZKtMKz5/zPnTdoKrm
v/Lbo8jSJImHcBJwKu6dUeNJ2lSEW/g0VN/GxAjnfLElKbsgFt+XXWhR/ddgi3tnuRkg/OzhE57Z
nqLqoK8p8ZDVpJ/EGnorPh9F/GfH/8m87hZhwfAwp50IKIdetT5eouPplhS8rgO0+5fVFZKc7WNa
4xPdVjml2NLj6ZTjvHNj+BztDQkjR5ygd3P8S+xOd/zHou+oO+qQrwepJilh4nhduFQYv+GkJKLf
9nMT+U1VeqU/YouD2bnJIsWWc5KBJ9fm3Q2PNrDl8IiGjMgqtQ9x8jwZ25oSNSf1yGUSnw1l9sEI
WOxFHS3QG2pQ8Eu59cplloHeqMWPx1J+mH/kJRCb9gwRLlIS22y8VD7OpwdVMJTb/eUIHkYjY2kb
oor1pA0bYrjCv80EFuc4WKuvpwNCM8Brg+AnuihcTISL1gPtvae8JJBwUPye8nFj2brbgc509qPY
AUsDOUgShSIMT2zUSZR+kuKc3PpkezG6TqmSV4N5RLrJCstmKkx08lhsBrGYcvdPL97Fx3qFjtqQ
EsLfTUEerStolUzcIlprz7gbo/kzFxU8OoARX9h1dkE6h4sMnS7Ag0OEDCqPOZ+1DxJk2JhYXWrz
NfdgRDaItgr0KOQ59ObjP5UEhu+PMhm0MEgAxLjH2ClX/ipyEdQOthA/6Zhf/NEpaR4ckNquUwrA
AmtSzNIphh3vpKgWgue3/PMkM7G+QYGg1BMUykhrcmtFiIbXvBdmpqDje8M3FQLPoqojlyjT/0gb
6hFlIK+PP4jh+YlAE2O+YPbGeYtciRamBRsv9lNvHeNjpKclCxHGkL99/q+fnvG+HLfcJOlkYl7W
cx4DFhIOmZjLkahmsRZ6/2/ATK14OZAnH3beenmLy/0KEMmTvgwQHZ8d7951pI9W/znG8vtiP+w/
/01WsxxTt7onRdyJDEc0wb11NYKBMyDsXNELhehxv0xcBomHRedBFu+ipXRwGMPLgHH/zrkW9P83
AseCBqYeMUJJPIpoGTckd3oBCuMO/pyuNwxX5/3M48c7xYb+DbhqSo/5cqv0kAmZDX8Ek9RH3SE7
kGy8fJPVErhpdgF5qTqv72hT54nrMQTPiT0+0niANllvyNKaONvrEkOiFaQXhq+PItoqb1F1Pq6o
MK8ZHodK9qBh1wUWYN6XO38Y3lPZHnR9HRKIULCDPXPgsTY4TSOrGsvYwEFZevSE9vO73K5WxRnO
Zk7cFdEbyY/6u8RTmEir7uIuTSD3P+FWW7b6ZANshD1H7eqq/umveiOqDDifK1rXBlpl/hsl/x/T
exYotCkhGr1Vuqpr9rTky1y2Xizgobddns9kzgOhSQcWOHhQAvGGNoFhoZLf+mJ5dl/x5EUanRGs
TdCbOtOWtnYb3kcD7hxDYvUdGrdiTxuCDx2eZTiiPPbL3Anpyf4eOIVHeq8HX1r7vxzEpS4ssiZ9
KdPL4lp9WaUyz8EYegZJVaY9JW3JxpHFGLRxwSJpLuYo7tkaPKvjjid2z9mmVamyQ9zvKRMG3Spr
Qn66fDqLkjRj12hH73KZRlUHHoGYMOcFkYw8kP00+vpBddnmDSvUACvtsf3IyN5k7gFUB389AvhW
SLOVE8qYv+N6Vp4B9CCagRm5AWyOLiaINyvxZs7BwIgc8QrzgjM3KRb+dumSPkb0iS2J/HGqHV/2
1JJ21tTbX6AxEcyeHFuVApieQAgqX9+K4QjUVE7BfZbPjzH+oStyMOB/Ez8VFwx/jcVIRSPiLRCN
TUUQUKTDb51DIxNDNdTROdrGIQ84T/KGIBgm2BFWBjqGkWE2XnpyY8snXWmDWUGal51gW37dcLk0
76egqmiF3LYd5kAU2/N65EpcmRVQODFzXZdXTvlGAi3j9e6U+KiBfwXbqNnM0ooqHKlQkgU7PfWW
Qe6pO8XopPFTkqDWmxZZJWkVqCMXGoOoRM0lgoyHnkKMjw2uuwX9p3j/QDXNsZDk4Sq4Z7IrrQwM
vlL09KEh7f1RIgZUfEc6bgALgYN297iry09QxdwMgoVf56xH++Dr/sxTqEiTczDwxWBj0s9/3/KJ
uQ54+lCwSxq+NgwGQZW9TZzC7gBzgiAxYzaRRAdyA9VWU8tNZi/9IBbU6YH9z0vXe/mNbYQkxxOP
RJaLFVMLRceOO+epP8j+Jo3xYolZdg/Y8iEiv7Cy0RZ+XEYomU3HEvGq0Wg0z6CbZgYbNQWMeOVQ
F8uMXz3VfYt0417s+FHDY7Fz/+8ckreMujU7khpq0PCJAg+2CFjIstSXJcnQAUYpYX2/z6Kq2rim
NmHEzsi02yoIjwUSaf6235dIQgtl17H72aMXZTJ9hJPD+a0JfFyQqNS2gRqlCc9Yz0KVpREe+70K
xCSS4LrItT3U452eyW6qpi26UjobchHRmvyHdoOJHBL/B0AygTCymZjJ5uNQfGicAgAixmmYLWvC
xH6YJ4vk++cX2v+UU+BH107Q/747mwCXrfPpTEKyMso9i5wtkVu8h4GWpKeLxjlI3baRFOiGiy2H
FWJ6ZWZqle/W2XKyZz6EgjHE6cWovcTQeatoEP4Sk7BsCBObihEnOI+4xfViUtw1lMtt9K261168
3wcitXqg8LuS/Gfl4E5eNFq7/S3XuEoARNHNXoSHQ8TDS428nNYGHCYqweumfK87VZIPqtkatKmE
Ikl4yf7rhctZmZG3R6cEPVJLnBGUYNMHWt0tluOrzjYwBzb3jEXmiogsVoE6qo9IlCTaN+kYhJb3
AMGUQ3NgB4q1ohDPmNlNkCxcLybsaJwztFtXXMdF6C+8D2ndLrmeLurtmp75ua7eKBan1Vk9xr5E
LVJxR2WD1wE0xoIe/u5LiR+VnZlA22fh8e/iTD8l1bCKr2g9vV1Wxc6WpQOm6Ey9mVIqrfaSA5aQ
NJ5lrGW/RUywrKI1xZTN5wc6UlacMihUAjbom61FZvptZupGKCi5TuOD+rhkKfx9YgIhtydRS+UK
6ptdQfnym+EJmIJrq3R+hp2Rvt3CeyofRrEpXoV/9vUwgKenHKM7WZPsZ963ChOAOof3vYpgabxm
yHJWAiqP+9z8KCmoLq2VNRc4TbTcdwHiu6I7WAC31QTy8Y1iwFPYlpVMdhrfSGewe0qjUDMEVV+I
FLYvLre2gMgODesFD6VFkQGamWdDX/8bj3HlcJ628wVNNBZ46aJhgRFs3KRW3aR0nZU7SV9ICfs+
zI6/uDFn6tU7GWQe7pqTlUQl4eVQyRf4grSKkzBD5buFOMowoe8YD3u3MO/YFq8Bfj5BZ4Q6JAJN
3IW3c2q1aPqysB2mFF+M6Tu71LPW/wOEotWTMEDV0Mas7BoQal8M5EBXWKQbzRkq6g6R2pN/2ps8
gyvEHnsNLQcJWf0McEILrwps3nIQbD6b9sqm0HCCCAUKK0MZY2upGMWiec5ZDP025hqciNaIC5pI
EIWCpIAaoLtmDTbTHYf0A/SVUtulpxbXE4lTk/OXViG2iZYC0jeMiX7SfuqpJsPW8X4jdPkMcB/l
Dh72iiIy7WcyY/gBCpmvWqEA8i1E6vVlJqfoybUF5BsV0yhcU7SL7W12yWep/Z3j1pEQaK7HfTgK
28qL9cVAcXrVTNnAgDHUd+k0clqQSU4PNY5LcOQKrZsUVtsBEJhKRdN4IyAwtRdvD93zGwNfNsVd
pXmCDj/nf4snenhU1RrZVa342/Vjj/H/clivkNv6DM8iCtdTxAY5gbDa+Oz1U8m/ddQ0zlJCiz3c
aMGtviSooTIZvxEpczk7NmeFADibrr2ahFb0b5Yl/p13MzR2xK2+H/K1SPBtAAQexA8+PheIG3ng
yJtrU295qAKWV9eNhDzjXWJw8xMMwhihD8zPqBzbvcRl/lff5HZfr8oxL/hPSJACHEm2gMeVdzAF
VmIE1IEbqq4lxqReu1B7hy6fHdll6WilJf0DIIivLlrFAx+HnSAP8hfIaNAIGVo+bVH7YCXBFBtF
WXri6no75Ac1O1udoTYHZbA+blQ3NPlijEdX/IkrVJAF/fEcs5DECNBzSORieFAosxK5dtve/nl5
TxCdziRDk7Oze+YrbYQUVaT7RcAOMmk1W4gir6p+AyObTmwKzMhyVinsB2F82qWDpm7Osr071sSb
x6Auv2CS+mDLjlcsoj/FRCGlfD+fACEOuwFSMsfISXbQhVvU9E1IAOwLHdJwdHexF5YYqLm/68kA
aJa/nfIi8+qwvNTwxdyJB+ZRUH7xh9vCyynGASJR/XqLnD8u6YolqyzLHagukcJhu/Za4QsgK3zk
jA7NwQXKHPllLuSqQlwEzCSOc3OMNeWsPZIZ/HWnbyMQnt4mfV8KKee4fLdO58F1wwRZgqi/oETL
rt2m2hqUwPQEeUjclcl+LLEu68fZwjL21vvBWEq079zyMQzRZFoIfUgF0xuUboXYdDc6lGZWqUv2
sdXXvRqfO5X4pITRZmhHY8uhS2QtIhv43qhN2znuo+OBUOMIr4NbdYOC1mOKXduQynHNpMKpc4E5
fagXIUz81kYBP2CzTvgshngkLHrzykrZbF+jdVbZvXNSXA2KdxAukq7siIMpGDSS+B5GRB1tfZlA
hy4dHV5v5x8bZkPFJCwdGZIYXKXGnipp9qYO5zGP27HxTQj7sTu9pDsy6tZlkG20k6oU+QmBS11u
we+U5TBmY4neejf11eWHKayKHndedPzMNZGMIePYEzAVm9MlYXWMUSBU6L0vdOeFoI+6dKgN6WER
Td4sXaLOxj1O3TudoGsPCFum4OXGOvmWA/3iz+AjPAiAbU4B+Ds7Bj64d3QBhFzr8oD1wmw2YBPs
HTajgnhwXoVRoNCb3y7kAVCVCmSlKGrYLFaYB+X5f/QUeD8iMhx4vYrJr6QaK0SJ5IoKeO4ibLpk
08Pq9E3evkqQyOfuRq9hvOsh91tm0/Gk+8IJc8W5WVk2bS3g1WAWyl7rJHUOdCEOunwAR1l7r0G0
YSZZPr7Vw6tN3yPcBWmJkoFRHiXBQ6rOnw6f5bbXjJpC5U6vMpvYA22CBZ08MV7R4DrrTw464agf
/Cl8zKLlxbRePhMCA8OPzbi+9sSv0vsEpvQJBsX3Elnxz71O8TPwEu2D3+MMdgeD8FzmNr2A7AgZ
F6HwWp60ZtaOVjheZ3Tl9a47DHpftHTV1NBR0ADTKPorD26il6ivKoiLfYvH8Cu3Vvb6iS6//5Ak
K5HunMq0c5heIfXdEFI2s2j1Pr6qtko2u2SkOVhXuavaCI04KXQ/TOFmlL/74+5UxZoEIdXa8eVg
p6NI9YlLYTQAaD7WSQ61MUXIo6BX1danno0YU7snIMbU7vaKXGLmSE3JUaesEzMOol02BlH3c5UE
I+xY7NL30ox+PXrqfLiUo5D4fqhCZpVdh0gUqaVmn5/zutRe5ZkeAMTzz1gWfxHBU1wWTJyUGkI3
oqLps+ucAD+5SYVj7bPZdCGUx/ahWxA9XWRMYRfaNWhCdiSF9jOA94MVhPOxs6FYlfT6IjiYZPW8
E5XlI0OuopULZ6bX0FXLHM7fv6/w6aUmFfH1EOAwweDADICMB3FcjvmwzBS/0kdLVmBLU4/vBAkf
33rzuwR6iClzAwHRASP+cNTOTiyKP7ZaFUbx+xXgZ1TwJ6PxlOsvucJhqdCYvks8Rjjra18/ko1b
qdM3CaI05VDotnKwI5ncejejAmXtUDrcPH4/2mDyfRJ9kqRuh7bLDhwgcsaI2Y5ITFbbupd/37nw
pZRFFo/55kpiIPOSgcP5JVEvnT4w9TQldm0cUtjDodvHJvZQRx0Q1k9B7CyiXh1/dPyZInACNNRu
3eeGrD59BMRfgh4c4PBXIJhQb8TZcOTkXFserIMINKhxJ1zgl/MTgZj5Ofgiqzp/096h9EIAdqkJ
7m3thguZrDJLbI6ke2AAQXXUpWy9c5tnJMsoqa0el6YCyc2woUl7xU0EykjcBRIaW6bit/N4LMix
WnK8sS0B5FLsvMA7jre4/1+g/7UGe8//LsC9gHJbFe02ttlG4v/n8Ar8a9NepNgLHhUjt2ANU8sg
tiQkSzqjFiy5Bxo7SiMhMIUX/8ilSfEL+WWnvd+61d4Rc718+D0y5FE+MMlXaLd4ASwlc6prnyN/
JhJfYkXso4KaLa1YQSbYIobKefrpfeYTEAH8YHlr1xM0Ky2sJMCcn4BiAcNKSFy1QNV7Y8T7fnwg
N1q8Oyltj2sPRbfKLOqjQt1YINB1dhBL3de4YalCTCzakB4e2U0JikVpEHjNM0Rfau5y85clpz4L
WbP8c9EiZ1+QFRM6Cifp6qhrFkDZ8c+gfgJFNkmFBSl7554eIStAMP3YfxfTZieNiuG+sZshs0jB
GeL79YU1Tu+Vhxx2XGsZE9qOXdLz1G7DqOdRWKicG9rJNG70yPCfuJEgFi3I25SzaBOp2l0HBLHK
e0UC2IbMJ4cQCBxCz9Gp7FjU/GQyCj4g9Y0qOF8d4YaRNb7hf1fR3dOh7Gw81Dmavga2d4+JXDHt
bQ99q3D7TOSxKzT0/oc5DnZ8N5MNeIdBiSZC0TSOQHK/yDXUKjBuFJAMzwqO8PzGnMCNdWNVnBdE
V71TW+2RRrWPavTljAdbALWjw0X/4Wg/vHNlE3zxVR2tS4okpyFya6tPnWCwX9f40BIA+mnQ0HaR
1En4Gbg7vK24qHMqLMsSxC2637zc/gzT1NFoKsdH0X5UptZWdgjdhLxbHwxMgvocGoxYJEncqIR6
LulRLGqxdBqzQaUHPcGKYR+1EMSdNAMlq6CgJ3KRHdQYycklK7zNQu1A2471oT57Xm6UDm5UxAm6
io6uUXeTjqWslK332X8XM4eybAPfBHHHs5lvyGAT38nS4bBmxW4DR/T2gcpFNNMkc779CnvqfT7U
lGIo9mhTZ8GeU9stsuJQFqazCdZRNnCdfjTAwWbedhI1HT2vvi6GH3WCNp4541eiHXApH+G0lRLL
/H3nWKceV4UnC0ACC2M+WLk8sAn9nGT8fOpf5svXMRPZXsngaMeR06Q3IvKs/zFZIWYhYgl5wj4i
7xUIfyrUcJMT0RsCS0Z3sY6vAMxGL9ldP/L3m6qezqPH9WZaTPACoGxVZKxlFMp0bzkupX/m6afN
75+upCkUOtMWBLYHut2xZqpTlIxR48+lVTXKqpDbGEXe3wuA3nYITdkII5kZDBL6jxb83ff55Tli
04Y3/qRhF+5Mf2i9uYQgGgoWdDUJHtO7z8fxY9fYTegH4jeSoUA5hAZ3xn6rZTqOVEIWKPMvOgAy
F3iLniPkdVnBvFfdAo93e8G4JlziksbxZfL3JUUNukPYBe1EnG5ihmpiByQuTEy55hyXlCvGWqsg
5myuLbYaEcWnPlLd9XV/6FfvqAXqzDCcCy5YT2sktrZZxgcNe043A486lR33CARttk/rXL+9p+kh
mGsAKJeBc86ShN8Oz9EnLolHIdE3O/87QXrIj+FbxzSPQT10BpqS84o5Xqv50efgREtSdRn7BBC3
4w7SN+iySdipKCApbcNUoM94VQIj0Wj68iJMnCS7yi9QgocmeJKRRXZeSO6nr1vcMt5gNZtVQqYj
8SgNZFxSmYxgqldR0Ds73xAffdyO+SW9or3Ugl7tCqizDp8TviKT2iqn19ylUCxbiB9q+RW+PcR9
4nQOzvxwMIAtqPs0SpQibbq7cTNUqKpX/4UGDyv53MtQPfIVdoqbZzVpgCePgEZoghsyFSgN6jLm
7XTaJ54DQRDwEpw3uPkmZ3tmamehpRCjhoElT+FqbpHE+X11DEGGt1DkpLnnNQwO4zwdLxkpg7RP
lTzhAreoyyjZJiNEKoE6zaY+7Ut26UHTGbwoqmlm2QW1J+2L1tPpB7JhAOHAZiUa8LuVTN2Ogt5X
BLe23KPM5hHBaqxP+MhCgeaUc6eUB97HgKvfz0wXHmFBYlZ+uCtG/2A/anjEdLtPsRp0oiWAcLUE
9FZwy/ps0fUgmlgtxQuJEJx1PcWfrb84v4HitWAjdrp84SxG7v9s8xqv55Rk1nud8H1uAbswsL/L
NHJpTjTCZdkk4p0zr3QpGC7LoAVtGYxqitHuP9QOxUb7cKGegH72ZD9E/L3KZkbbn0FwdXsxQP+s
JtyBL/5oK3MeysDi+8h1pZnPIn7zvrbVNJW30QRjwBZGq0oeW/0M4wmeccaGdI45mc6qAGigtedq
IUfpbDnD5WytAlV3ubjlOvDI8o+WOOk431fXzoru9VHpKxzuocBck1YX4NSx7wjzj5uOMejP7DYL
LCpjn4Pblqq3ivzOMy4l4GV36L35ZgLjxhIIHvV/+bUN5G2jdOeDY+FmPCMdwV+hmb7jE10xrbvo
zOE2iGluXUL9FxEQNllOfbrYSzs7FgLGA8jc/OzuPiW7zL6cIyXEJBi90M99mbOdZtn6hkuOSHfa
UatHgYRbEKlEomV+AXSxqwd8OZ44W4+SRVx8XT/V5ROts8sf0Q/styo9aln48uiAvxm67oFvjahl
0JrzYSTpoPkDhHWyhv/nQOOVqzvUtW4ek0o1dodcCrzXp9VaO7FXqxq7N1z3ewRd0NMv6xTGH4Rh
fehqRPTBrUg403dMqLcwjAHbHKNhDxkrlunWm4UGfxm+fXVQrl3wNXOdJInBs1TcRsogQ/M2AeTu
oCH66mqDDr6HvqXitzD69RgR8VPNchBv6mpXuBhJY3b1HgsQINBnabJVAE5B73xjbL85PZEbQkqr
UFNkCUU1myo/5N2qBqxjtWNNALT+lZsEHfOJa+lcGzfEM8GWqJDQ2tkvCv9lQF+K49jRCZId/dB5
73oPV5HrXUXnXvsIP84tBmv4zWvDxmxDP+AJkLSjl9jh0FufA/6sAVUbd5L4ag4987lgRn+CzRT8
GWmze739jLUvcAxl2cukeuL88jitu3rFsjZXVknIfWhbNKVpuQ0o0SN47GRyH6uuxAt5VibBzfsS
hzLMgB6g2olD6D9ijV0PUidStYSctQPsRssPGlx36I98tD69NnZyPJBiSDFurLZl+8q28ciGGYmx
EQvbrt27cESqF7EY7AmufN/vyQ1BherRjlaxiU3qanOYHPSl+BrOkBf9VghS6N8TSlpTkS3pJr/o
Ma34gUTO2HiQ4KfkWwmSOAkf9WyTCBh/afU8tPS2LLbH2eHhFjlThrHkStTjZS951M2YWIbE8IU+
t1ARAvXhDi0cfG+7szEug79St70IQOg7Cv0RkcRgFhoC+6d10J7y5Pkjn1WjUB24DAtRwIQQ10f7
zZdbIOXR5QaaQ2CX8VlW5dxcpPhHA336gChvvPZaewEAsEmkGZJ3omkjngXmZVdQzI4aTcCHwsUi
PIyNRa4+K9fn0vagvUTLkG0F2zs3wGF1ubXw0zbzd5nU8zcjbTNmWwhUTdS5mkEBngoMx+bxNUaF
1bqsx6QgOzaDkmmlBIwr05SXWmVIKcyFM1RaJKSgsnhQW2ICjt/APrFDeUqAjHhwjy9O3xHshxRd
7KXHgetUfy7S1y1Et+4RAvXmHe3jyBtWHIILZWm2UqPDTZhRo82UJr4xPr5ZuOOjavEqIOffHSR4
r6GkPZIZ/tcPkozZlGfP2ImyjXi9P5GWPV0YDpKtzh+MsqAAXChZXldzzLv+InOs+fBzHhcV6BTC
fsH4XWlEtAX8uedtH1i+T6m6NMdeJYJ1OBlRVzDNNQshIRKyIz2jMVbFYbPRs2bM+9tlMA/UwAB4
+ujibHbFJZy4ULBfW3uhIa88Ymztn+JSn+z9JGjB31mf4sLiJirOKj8Zih8V1SsmgIwFSnFCDr4A
pt0jTjWBwKfA8HFl861fIz73R7faWM8ulweEXGe91wbF0Ta2Cgc4ocQ9vAJ0CXvXWYwPhkhowdLn
c8VEskO0MboEYTMkz2cXNEGfcE9CpDB7LDAcpXfmUm+Iyh0dIH+OxdRveu6vTK3dyRu/B22bLmk+
/io08CrKsKOGCkzcltBmmkRiPAf6k+LqS+bqaiSpgRPmCrokUNwSiY6zT/78lDxIJOb97E1cyom5
5AbSR31k1FhQ/Bb4tLA/VMmQIoU7GzJt2GpcUTLSft7pGNa0Cbc52CQoCug5UfJ3HrBGNAdF2061
chvpElyljooZ+Iofjh28696HwwZ5WB6cUfWViIJ+Rkz7eoOJSgaGBkK/BMOHFwTgngMwW9MA/4uK
e0I+y8KVFl1Mbr/5MWNrnw55OARjLONAH4Rma/rkY6WMtSElL0dtrC8ATZEhgd48uyw0B2+aiiHs
mcVsPdH6YY48/igkGGzEeCWbfAGv5tKinj0dYbTCbeGhO9Q61DS4AkbZiuT6khTZRNM7m5T6CKRH
lRmAhUv+SwCsGoDgn4WkxUPLpDuv1FL7MTnTuXLTqvx1GsHLI9kAkmzxoEDNXfGmXG/ODCj9QNRE
aaHJjpsYvmAgfVUJeVznYdj4nKOHI75/0B6lqkmzKPXICTfj/HadFvVrZp5P4ZJ2DIEXDlgxlZzx
Ow5W27DyeN7akh0LAxI9dPggS7vZCJfBC0HMPLEEc76VD+fwNH0Yr/vd0vwg2w1JLZ3LnLZjM3ap
WMSZaF5J0/9uUQJLeFTW7qAk4Zc5tQBwwog9CqWOYnomTYww1FURco69vfTq35PhQ37TlSRZhr1V
Xjik12oKwchUCgYAzNIh9Bz5NMLOG8MTgcWlXZhkDilGe3DyJODbFVHTiNvkjonP7/LJIfR9H2Z8
A0qGnjs1ZeOvKv7tvTKDt5vEHLtIH1n4ryVh/n3XWM+Lpi0ys0iQhOTSl0jtt4i54nCDISjGzovx
2JvKEw84ghPKeAGY6oAR8ZfF9m+B/yqIkfsC3WY7LNpCYUWPpCih4G0vKxV7J4fRrX9R3VNQk/Er
RJjfy+2lCyqtt1IAP6exPFU2ZLRV1LFe+4M68NLBCwXMPKstSQQqpFCIqjILOgjAOZfTZFVgFKKO
5Eg4YKGqDh9NCTJOfGc2SAiypHlUErrpps0eR8XX5eShjyEEb2pQ6RAaSf4haguPW5Y3bvHxHhKR
skpRsuMtAL5epoRxdQiB8bBZDEi8JGOaKSH8twN6Yr3TQ40Ajc02FsHPjCe5kdkup3MITezCF/W4
iGv+NfRfJJPtnnY9q8xFctYQ1hYOnuy6i2cIXmEPTdtNZMK1KTDqg5v+TAkD3aqj1itSz20G3Opm
TwB+WqoDnxh2hX4jK6N4ybv6qHAWQbqIX7CQaZzV+HiiUizIPTvrtstVOQncZqIoHNtqrZ+4f/Xt
zDZ8xpAfaTfj5yaYezW+Fl3+YvPJ8eba9XoWhLwz8sMZNQf1WEU3cDB0N+AbGm6qauVOEStuT6g/
aJ3bx20u+etYn2OggipGGK9GPj3ytdIaF1u12o3kYAS+9GGoFlzSahNSFK/8YR3LYvdJfiiWOUp0
4hRIXY6qCRyaG8MuDIn79xi42L5Vp9Qp0l/iPJ8lTHCiqZOFrsl7C2lVp4smbIsWQVfqNsQBHBZO
tkegS+4iF0JZ+ryhkMcfLsKjArhtksaWiaKe7vN0H7o8EWmWlENaVk4urHSWMdx03AkNcoPm0+Tx
aMuIqFSBd1Z9SptCdWTfENMLyoJim+wwpOeVvPITNHE4AhkfinBI0AXiY1WFONlPRpV045Hql3bR
83PnsCCHn30WaQUwHthaX8XTF0GjjM51zJqz+l5NG9ROBshbY0G+Ga1QkZ/wjTjiLhZjutBQkNEy
z0nKesD6dN5c11X5vIyR3mPef8HXYqsExh2q+H0BNFwXwubQc1bJLhsS40UA6qid4p8ZJxqoG2R/
aqW724Ucq4QkiF42aQTHkj7VhWVNMd68EXAD+KuoysL5OGGfaZkpEUdYJ7AkdWi6z3cuMn6Rvr7q
JIYCFqHmzy75Mtb/J7NXCUZoCfJRlF3KIdq86meeRkNVWl1f4iAgv4e04Bs8vKJFIDjZVjysBRkK
gb3+oHmhITkJa95O2XqJsRVmZXUkwamC5nJ4pGagfJKBOCjsM2Nzw3fKepz5KeD2KbovL48GcvGI
vtOaEOBIT8o0v8QpDAFGxVeX8x9lRrujRGRpfUSKmKMURvrMk1B8HsuTS2PYAFYhcplCLz5sQR+F
kcC3GVu/JXQk0u1bwGaCUwRPsdWGgoxrA3EscIMhtejIPYJgAU8qHxiWEBRFT0dzlqLhki7avij2
Xq4ZS87vPz2E8jHOFjr3LQmcQ16za6KIaNjNRDaeEsBaIhUOyy956P/OIQS7iyqtlZsUw1OWS6TV
24aMw6raAkrNmkxAKoDYvT8luC0UAM55sPaA43JRF5nApWgG+8TH9u0eurU/w1C+Hb+/GSOkO5Yp
6KcYKHAKwSPnUFPqvLK5BvPURz66gCYnNhBy6IMcdLAFCIDWi3LrWXpQYssHuBogrhbzYISg97Mw
WqEzgttvGji3ZR9t/zqXQh+HMYgg6r8gwG/EoixZc8PLxyTtqTzNRsacQmsLYsc89jboyPOqnt/y
ZAgHxmwJcC1gQCLgqHnVu4VknCwQnH0iI4+OiLrfFjABdwhSYYpj1+a60u3bLIqkaenNzEAKCf2W
POC5PaGwydz6EsDX8RA/jmNMIL/GWdTTxQC8CqVpVozZcOM6YAah7/C3N97jmGSnXwB91Av/we48
Td2Y9Znd4BRZ68/1fZao0wd/TewJP+49dXvAVrMbrbRQ2/2o6JpAtv5K93I6CViPwuFJuX/b9rPt
d8339BohVB7n5FnHAgWjcSDgF5t7WWgU7IujdcKjeIteUptTzVgrZc+ybusB+eNbC5J30AuWVIgm
OdKcyK/igsEUd44d5NXqxuIZ04SYi/8hbzrkAUlG0jnc9lzXM2C/9XOIZzsatiC96XaN66oXEOrV
Ljvj9i0zqNhg8bUithri3NdEgJh1EXRunxB8CuMMQiORYmykwMIlu4d9mil7LIctS8IDHRgF+USo
NnSuHF11n8llWkIpnyF8TJvI0Tb8aks2uIt5sdQUGbAhOZx+xDPalnSezs7LFoXnF9tXX9MJRzQS
5ktyi6DL7MJm+vqkmX6k1n8mRNCqSMzO79XCdj5fkxvnZyrmIITbFjR0+FP5lV3mnFVRuwuqHSgO
SsvFDamz+ECAFBG8lU3wyA3dwDkHmci7U60nkLlZJOL6NFTEmqGcK27sEcfsoXYHrUi4/kcvbhvV
wjoP0FpdCoAwk73j6WolUBMvzcB2SgE8l/+wpuW1zwKXaqnZpPPZp3+gsntiI5Zzjz6s0WbNf/UC
Z7GpZgWXhvp/29OKqWBXUSGaRl2Zrsy9FxpyuEUVHHk9JV9G9IPdGVHTr/WeX35KoanMy4+fwTZ8
tBissnmpRexFEpyhKMd2LVuBP5ScVI56f4FVIkOrxDzcwJeqjlJRDDeTC5he+6AXR5yCplHwUcsH
KlOJY0zQZFGgv77HKY+SdfswQKoUnqiOTf58XFN5MuHF/aSF3jPgcGBk6KLJCjpkxH6x0x8hNYLt
yFMgaGp8swcMiJ4nQoIcE/8lu1VvISAsKuVqkgkqLVZRnscs0zFHltf2ZIQL6THkNeqp9sQoKAZX
PpE7guPDvQwGl1SKOWnA3594WeogubQUIYZoRHrNd8wghMuRm/P7JvfgU3UwninJZnm1Lp+vMirX
Ny32dmIVxRoMUBfsW4WZaYIIfei73CGNO5/K4W+SdXVhg74MvOnrxXkJKsKZc8bDt3735FzSIisu
stgfukTqtPIBZjHDofZz4vNAct6Q5ZPiRDfAdPdL3yBg0Gyk55uOBK90yc+dCdrdaLmliCtyrjLI
NJbok/56Y8kkfIAFs9kJGbs2+SHDV+xo4zyIe3WyS6yoZVGozaflcKA3nqbRc8s40P5uw3d9rjMI
zjuglagZWF4R+FUBXDvvEeZpxmmfDWJ2bqsmAiyugKxPFgfrLsdJ3PH4LNkQHfXFltXVI3sPHhjj
PdH/QUBg1YjBleqjU8gyt3IL7N4Wr0EUTFlbDKBFyx7nb5oPde36Doz47WBJ+tJTYVHIX0cXId52
OPrfHtP6TY5J5Rv4nOltsa/K5gsyNxGj2B0O6TtqklGmQrSsNim8HU9S61f+d8VIubZSE2J7Nvpa
xMgh5JwGBboHStG1LpLAAYAqLpaNYTrjNoaRUG5Qos9r0opGw2/gqeOrlcQ4G+tg4pMEgApSBQqv
09WgcKog6nYNPGmRUTv7WUOv4aSpWrJJYse5OflBWA3nZnyYMdtLagaTvfQj/zXHXNU/0AYa0Gw1
QgyAQ88krOLE+d79oZsIarRxHKPWTd13WQIacPhofYGH2oLnzT407kyn4zrX59b/yYA/krX/Kgvs
q5wX1Gcx056KauMRRIRXuzP1Y6io9cf6Uq61A0LbwzLKsLf9GG/m+EDND9xiz2gU8gvPSfv6joUi
wGyyKhS+bvKVySo4vPejebYGIdwfSG9tH3DNrh+fH6G9BqmbNyUvXoTnLM92h8WSUyyIN5iYdmpF
ZETnyvWb+4q7YhaOioQTKZE7XrxNkOa+LhjdtDJ2k6MoJGPhu85rwu7nTYzIiY4WR9freUAKeZ1z
ZriV7k/4YZOE5qT1PexsIo6uci6Tmvfn7qqgsVo0WPXxV0Sd1aN9SBBxZzUs1j795nlMr/YxYIRi
1U4fhzO7Y4Me7P4924YigsKOuyguKBkVo5MRgcWoy2gAFXGbwktt4bYrhU/K5/zusmPpiYJgD3fj
Keicx4CKXsRWPS0Wlct3W5KKZ5y7TciSLXvy3wBELpxnwStvH9cAIN69UzNdjY4tIuGJOFsD1TEb
PTbVp03OKo9LoptfMmFlB60hSjdsMr9khvJ2dmGpTcRs0er9MjxJZyMODvwVVq1gMifkFUVImMMB
CZNILV5PXTO6HfqByuaTBXVIEP9Q41xHynJpwfkcMgXHMyeRotZ8mkeDeOZ2Lg3qIO15hKbwKUYt
mqOaERo9XrleN7BLRXFX8LFk73drrbZyEbrHvU0JtSO5EZpFnJ4QOhyeNk6bFN84ZPG0/xLM8yL2
MQqAFNRl8wO7gZfqjNshU3mU0wOUMsTFy45Zf8mf89ZLagYhpR/32MlopWz9nob9k5/VMiQDhGVu
9ZTje6xd83pWQb6su4IDfUywkbYLKtEElmAqS+9k2yg7+JJJry6IpifCTvTTvaZ8AP0dz/mavRli
q4WxPPum3OXITkPVmSy7BcGHW5W4qM6230Sn45nbnSF3+h5a2pV9kDHW8raIYNMwSu0zJACl554O
lcN5+zQewjKS6fmHEx0iN/QgVolam9E4i/b1Ff8Kz8BCT/X/xmC8d7TTJSY3Bq5+SeBQId+XO+sd
DvzkPORgdFnrxCSYG1lBEag5eIb05vFmQbFZ0EW1vK6SkfJN6f8CReRUtjfzMQYOJcI4eOuykuzv
q7LS+IBiVQqVd0WepdHprpcU2CuQ80evC+DwHc8hDJ5qYiK8ehJGfHUxATm4fH5GmJgN6l+fvVK1
wfmikJKEpUk9aqTW6WVKrPL7hX8r7ugZ4kTb3S4bfLhv+modjrKZOvvZOHwcPlWhBag5kNKFo4kt
OoGutcRr10CF6OqdPc28TiKO7RIUKSFppAiCbvcle7JQTiy/3eSlctuX7a+rWznZxHC352KDzrC4
GWcjaSdvry4lyI4rBfLc/j+IqmwA9O06GGrdmqu+dtRezp56Pi9fFmZFSvxsIXeFvo7XvzT20WIP
haM2Q21Yfyrk+LaGRZzxflLmAVLfiNEc3XhW58emCtnbOLJwzBjINHiqmfleTp0uz+1cGR8orZ8z
EMAEJ8d8DadZ8Vp7PcLvWFGxVk/DDnGHZuzsSbJzxf+n/XWPHRnI/5w/272VtbywiZznxLW0v2P1
hWsX8elTev7/PjBIhhO5T5jE34o8w7ShMikogoppKVpbCjRQNE3n+wc9/rCWX7ZAwsDH59C9tM9/
yc8NFdDYlhhaXDujn1ihe7tso3426DakU2djNMgg3GQj7P6hTJhtfe+I2zQMnsAfOOO2u4Nwfytl
lwKbj+YvzcYbF6vyxL0yWJ9xSuJIoq7XoAk/JxRURRCkjOkc7rAzAdbu6UBCffYlLzboM3PVkDoC
EezopC1jaysluGQLZOEoOZsCAE62rOhRicXsM/ghyTnLXjLrbttCqFauqPoaF/yr9MNGzPgImCl+
9KSJVCtIRRRF6R7oezbMif9V4WN15gitLEuNnHhN+Mg4ruXWf5twL18F8sao0DXqD4pM8SrnNWnq
to+YfDCT3aMMcjatSwDVwNtBCmz3ZHcrFjUIiZXbj3HiZRsI0bcwneYqqTnTcxNO/Zuk8opRtjJP
ie2W9gibetBBvsSSsS3Uywgka4YuD1w4IHbfKqy2mvJcVNaPbZt43zMufOTfYv/nZYBKTYI/6ga1
rXVg1UBxq8h63UvfuS0D2a/C5gp6HpxSwhMqoQUqPrg0ASZpTBfpiD+2Bg9QrkTE3msueFxQqxUA
1ZxtDVZijDnTqubB5Oa0ELXeKLWmnGkPzopWZeDZKyA+5GaUSLZvEcB6mH104LBKpJJrHK9ovnVF
eRD2MLIuK1pZkycaJ4MfqauhT/IG2PMP0ZDVpCLoKdTruDcdcsu6lSij5WjVRIl8aDMdXkIFUSdB
0JR+d14+/MKjN5yYEmxZmAHAv+26AZEgMwnj0Q6bhFYgkAHsLsTf375N+xYX1ZcUNG60lrq/aiF1
XWR0LIsWX9gp/MLWnixoSPiD40m6NNwr/PpRxrcswWqPaDU5dX/LhqPO8qI8Eo/pv/HCAGWvkQ5V
XkGl5BIrQEi1be0Ojt1DYFMeqtpZ1uVyXxnMHcD1i0NJP+sUlrkhtci6A3UXgfYeozr64LTVh/iy
KAUT/PeWTm8NUqIDUZHqPulLThH1tZDgRjSSaU1YQZE3JXds0LSULmh0NfRsaFPsh3WwCQ03iLvG
CbYAfB+HkMhmuvMpPVBb90gvRlxJ4u7ZlyyJhZH/v6+GSy2p9uNZQNxRfvv1tWcfUtXLAInHQjYO
r2xjUtUx2fdqZyRLTqOdA64AjeBewxmDqVYQpw6ynoaaxF15G8Heutntu7ldq5cl94z2ysCMvXBr
RXvkR7a64QQbhBQnpRmwjuWyNwzs8aO7CQLUQnqA3CCxTLyoEs4QrAtdFJNyty2yHEoqNlEONNgn
r+7DrSjnnF0LhrY/DYPWfXY9e85qmZIr/Ibhkip2NJ5JZV38Ll7ZKl9ufcjCOJUvdtF/vpJYbdTu
b/U/ztUkAvOeN5P+PvpwZNWcVugAXTD1V+3lYkuIlSjxuDwX46B1nSRgU7xlmeOdsUoktuJQp7Q0
FbipTH/kEMfWdBL/tJ4izQSRXX/+xY7Iwjfx5WRFull86Anse2Wk1xQQA4EyGSz91axg1CQlmpfk
lWqi9B38DXiWU7MVDcOiAjYRJyQbF9CnY8oBdgLJxR5uAa4H/NjOoEKy20/0mvO74bz3YEfesIbs
u1Vob+IkTd3ey4xvDE9iG5H5Pna0VjmfwyRBYvReYLUaZ5njtdLo86IQR6YvENVcwvhtMypYWpco
+fytr2uBGee7oKP/7fB+gPgeTt4SFcBghEMFUcv8WY+xQWUiA0d76TGKHQsm0GtQT+ZadF4yME07
OA4ImmEBSpVSspUnyjSZ9XekBrmGPHZjDiyExLhTBs/mXXvTtgBqlyTOuxkN9dg2WxnyPc1xKq3B
mw7dkHvHYqiyfSGNlJb+PlSMEsLE45pDCXpVPYwn2+i8LfjXDzR2i9oa0DnGU99KSS1CcVUwqLpY
c++DCJQALrKtzD1rg2JTXHPdNJIZxoo0jESQKXmbOwqSsEVv+n2udddJEliaL7BvzsywJncr0zbF
BwzCoLe1uLTpObOaJgVsppEDnl6Eo3MiOC5CiqAGOsq8xFtohp9Q/UZJZy/nucsMLJ+44SajZnyS
V2WwJEaYjopIvool5Uc8kCWEVy90cm1Xup/hzJWdCg6DXMEdB1tBWwbvROAa+oBPaeaR05XyaJWb
a9BZOBtPddf8QFryvAc/KgwioRP7vuNMr5Nfkw820+V/IVMcIG1DraF0nVY9A97OU4KAfY2LthuW
tVtx7PowNPmcYt53RSv8szLMAbttozIwYL4Uy5DomXBTBP4WHNl9EhbTuEHmfSCXO1nR9nGGc3XJ
8+uR6dzVD7HVAn7BcMXLg7+0D+4YJvBIroKYyRs2xfSYj1FLmoxzPg1siffEHHKCjGo4TiZu1cFg
qL0AkjsgmSuL9NSNJmdG/T2Hz/cRY5xB43jeaLMXfCyi9QKqZR3ZQOaBZdzMOM51mtTd8VmnrK8G
6P+iTsNGR9YgTnKihEB6UPxjhRknw/4PVIrqkqvxNP7R5kntcxa3eWCSW/gtViaIzgUFRYA39ZOm
pvhhMWj4zl6U5vhc8j/q+d0P1NrYYatNzAKfF+ehe6LZLmFyekrmnjMaiM8xFr4egZvn0FWcy+Xu
k/Jmz1LL+TknAMWg8dxwj6jE9ZeWOfBED7Cm3bIS0P7xi9gVGtTXz0vv1DDeQ2VkMBeWE6hlbYD+
AtCKc/kRPVF8Ra/xQR5wwMaTXQZiW4O5+F23IgUMzR89I0Lnv0nEUcVBF6eCFZhfA/odrfeUA9fC
dNGmcO4OHBxW6kkDrLHaqsjYwhVqZghlMBWrYa0wiyjiR2LXxq39y4HbbdcHLEFmoabLiqdtetmC
LTnbUgoM8jaC2zCb6psHt1IOB0qLujPNufV+DS+kkv8TIZMduh9debMD/y7UvUeJBEtM9s0UvduP
iaWSPyFdictSGA3JUiB0YNyPw5hLKfoOXBQn1QmbZAn63hKy8X7ZlMKA+QsSsW20yT/X8SuuwoDa
lnESaTQWe5+UIrucAwTcSEP2MLB8V237rWF2jonZG5d9KmATrDGRQIRdqh6M3ZSHOz1qSV/o58wm
7gbgMMXBtyq9l7IoG53CGxAtxCCECJIkUf0OfSSQcvUcD1O1BGTe4ieY6oqjn4c7JXdhE2UYavip
yllZRQiKwS++DLuRG0v2CNDxm6g62cKDkbstfaocPuxoHd6C+9wpvXIfFd3fGT8NrtNUp+L9v4/j
MMsUV9xSDKH3RL74gYlGgjEzptuqdJwKhuAjG6ePaMkxoGOycNeW+lr1p/3e+oVKmt95X6fTheZH
VedExL5r48cp1PHY3RHE8qEF/EWK0VxaP+1O3F68xz7Tneyd2Doq2idG8TJshkOH6upxo/AJGoth
Ftgzp4U4/BuSxT/LpkZQi03qlxlzyw1/TyEF6u4xcKZBCqOkUYZFlWRq/vKkYXUeJRd8ZZwmHPYK
kBii5jjkrcBP6oCd0kxmN83nglY2lkIib35mzPn7HFtUkUAyLSyeilqYpIp0FL2JaxuiwisQ/Mm1
wawqLxWNRy4Aqn2WPZCwtwcWd0Nr37YmvIQakzgGQ/FfyV0dXWpGqqslF3KqDTbWbEh0yepE6N0h
oIFUyTi+bEBkExRK4P1Au2VGANtfmgVIwjeW4rLHdR/EmAGeEU9c7tLKJf16U7lO5o2UO3g3ZFjE
TUJo5ewK7Fq1m+9XEaI81gFaNMliNvTqhZu6j9l8zNQiZ8mkyfEw4LtxAglsOAw3ZlGEmJ39q/pf
fRmkfoFTRDYXfkWYffPZbvLyxzVQMLBk53JbZRrD6YFwMZhobk/GBx7odv3amJNhz9odSVvm4jyC
rkM5HeYnmWU1wdEwzMHim1k8E/jzOaksZfJmEjo8igcTAJtp1WxJNK7RwcGr+0LDsBLBX4rn0QAd
o1S0Cs4Ou9zwtwzCGclW35J42SOa4bMOeWmFEfcbRUqQYfo1pSiS3O4bPDiFoR1hWDlqkUKevNg6
u8D+cCLrFqWH/dHiVP5khIK35ccMHv/ys12pLmH+UzYb0JxsSEG3Z2jYeiI+KRNvIrXGeoKhCWsK
VBTO/DOX/tpREGCPZKKqn+xiUYBCfz/cIojPevADDb0RfzscfaaFTxEKhwFbTkgo4as9Lp5sOIeB
l3a3jAI+UHogku6vlRuKKBK6nU8p26SAIL9OLNMmfA5mLQbmJxDkYSrOGBYhmcAT8AMHiKpA6mKF
GXVDdRRqoCjbYGnbLz6SkKWy67v8H3TQanKGTe3Ieuolax0dFiwcFYTMtAIrUvIeSWpPrpn+AU8a
gfhyumMMvJTernaaiZXkOowsDDgecizw3Aw92mY+5cTNxXIWTrFOdbo+8/8I10B1zaLcTkAQLRsc
l7KjAIdFIMQba2qa4KfC/Ptn35yvBylTwgk5QidMJS5i2CDr1+62GGI8JMbW1nUyWwgVWAe2SdIH
f3wEIQ8sOGkZ05N/H4h5DSVzEZrcu4rq8M33lJve2kTS0VhLbxpXyi+Mwiag+13mSOOE984G5Wku
zsQIJEhodo3FnhRmbW2UzZaPrx7tA/yb1FcyK00IPfLRCWkbUfWTC1HOjQDVRH7fufvepj/O3um8
cEs0E7wZCRI8vZrcubg1SceZmIuld6KV3UHomJjxsk+FxrawQk+MHuAo72sWWpBrlAoxWnBXpl2G
d0iEYA+sl2jYkas1dYz9vMtMH6AU/JsfgLn1QZ7AZPYO0vt4HpUODQoGGrnvkv7E6jORPMUKP6mA
Ps2SaRQ/BgZwFkXB4LJFvtb1BX7ftSQ6t0ASEgTAtE9g5Kmh3kL/SQFxONN2IVfDO0KCBBQVpW1X
9w35l2ebVNq5R111ynZZVaOgXNjk7Yvz6vA1muMstJBE33SCyabpP9fSizVfubEB8Kj1AkAdREYo
vSj69qOwl6M2gYeH4scm22mwwgZnYim1BXlRzMzEL/JAqK6LIutDw8vHl2MGnF5WT4/N/rPmXt0C
/vMa/FoFv14AgKJJXT4RLf6OjVgxuVzzA8HEu7rcvEs2h4PzrqkuPmkOnxIUkkmmV8DJnsXYNOf6
GcqjS6zlBAnYQEkDN8TYLA+2A3p4SV0eo0GyD+ydiLxV7jT2Qwyt1JycrAjxIPaFqgDgG2dhRdPo
Cv05S5ai7f8ptGSCEfOYxBlU2U5qcjR992SPhA4yAleKpadh6PBcvyMdGNMqWhP6lE+K9bvQf85F
KZ0AZGJ9qT/fmVpg29whSu8RKvRd4weJ3MuiAHlU6mmRT0OXm+T36skncPjKmYdCzAeW0H31eEmk
0Ot56KpyyUYMq6/aO/71AUffuAttc4WfWvJHHz+NzUPbsfZ7j3AkPrcp5UHNuBcfRHS9MBVQvOsK
PuhzMJV2/Hq8KpMX/1KEmw/UCVJiG1lG+/wyfcFyTM0ROlx3g1dbuVK03szMyrnzUdoSvZ2E1pmC
zF6obt8uAHrPoOTroLaJAwLFrwdUdG/1yCPw0mAXoPq2JJgRZyMA+RnIonsi/6od1yqfjb2j/qoP
scQIoKIHw6v1cyCcxdGqv8R51cOX620uiFPdTiJytQCkn2Kfv2QAIiSEpuSEWkiJGWfW4eUMdT2U
QFeoe0oXQzH7dASgCJJUIjvHCY95CM88ROiKMrams80ver6ut1swWs5+fcBIiuQ4FvBbbcjgrqyM
9R1VUFcczG6OTYacZpjJ5JRHESNA0F2TgvRHhfwFGP55wxfDt8dBHRAQdeEnQK+UbBOGpBOp8aJd
hEquSol82LCD8uiuPppPzaOOPtKCmXRflh/PfXgcoRP7lMQHk2sJjceiQEtjc/jw61w7xhhbYqDf
NI2LzSjMDEZTNHb1gmlJLmE2Y1mQobLslajl4v8W5YhSc2HW12xN2caAT2qKws//M3hvbkQBnMyw
RTCCGrDzCah9Ruj4hGHX2y0+OGtyUDRGctWOVkmK/jqO0J02E1WRxYFIkebbZgAPUqsa6JMCuVnN
32FJpySUgbbFR2XZcZwcCgee0O0GwQtlVji2b0YbjG7b9AaS7zlaz1961rFFoH+x8GgdTlwbOtXy
F/r2rxL3FBPuvkL30sO+DG32TYaQb2X1ROkdWm3Fpd4+XQFLlZfxvOHkvjHur/clIX6YwRx75TDs
12n5PXrbS60uS6P5ZnW9t/V9Lj2WFfYK7jPbtaGp53dqy8Lmfvx7RKUE9lsXgBEi6t2Xyvd0DlAe
4pzBu2uKhSLeo8rQFZv1Bi3I65mu7/IRTlj05xq5OJceECcuAp0A9qjnw2eLDFrPBRjHMInZWHSP
Va2YShKZi1Y1fagM2OpQE1p4sa6/SrrB2iBrfRKxpwPq8+7jggjWrN0Rrl0RcCGN09UT2F5WLTKr
rpZ+7XyG4m01qTpdXLaGeCj0A1vVCS6cCZY0rJWz5O5IZ+Iw7DS7fsJ1Z63ODd04XBvOfJiqh8v6
1jq8ghYnU9h7xc34KS4/1Il9VwZS1lcZ/NC1Q7f5oExtyI7dgxCl2AoTUQXPncXg0lJpcQHnBtAW
6dmpoNq/b1DX4omuiiVx1mPT986VrKpqwAkqorDJsxrYXig4wdi8AGbNz+iV51RCQP9phM330g0p
R/QDQZEjhz5lCPtTGf4EGgAzi4ptpSTXWKMxFxvqhfZq509lMcrXGkChwaTvy5s/nWZyuWrjyk6F
vf36Tf9c1MpdHC7cT5w4H79gmmjGG2Xtorn5Z5ln8IduSUK+/hVnK5gcZH3oqva1YrhJJQrg4wg8
crU7WXQPNWM7R5Ey60kCToXyOx7VFPFSAa2WWzuFpiBDm5V2nEBR3m9SF/7xvNYIl2MGMERQMcCF
DJBTVRzIoWBBj+GeAkDkizjGM9KJYjTkaBzL19nbhRXRrTfxCYoEdlqlc0ZmmeM4VbDqubKZI419
5QF8csNYpcc1qgRGFIes0rv86HaaB+Gyh54iriRicngZQrrCrqlG6qkJZ3BHAJqMfR0CXRVft4Y+
GaiQnQzXVCOux+UvRQIGVlMonipP4pD4lQTq2o7OySuPisc5q/BkGveleijef4MJoRimOS8jVy7Z
A4dJVylCQHUOMooStw5TCfe+HSFiLYuJvyMPsIt9Tw30akgamBjDHDDxgcV3LV5ycod5q0Gz/g1q
wX/OtQ8/DdvBP+JBtpUxmeTAd+1A0CNpWgfEd/9+RhTFR2bS/ZMg/5rObVqp0S9cYGeYwUoDKyxQ
OW8xUDaWVf6BpDwfUNSWMI+rfasRi41vZXs0AZmCq+vj453a6nhCxXRZLGRehZ1mGQetBooHY22N
5RUfeM5P48MurOnOIm3eWCl/LASQwbi9f/SBvXQrY2g+yjMAEpQPOCpsRnnI+0Kuwe0b5uv5UunW
YRox3y1tbZwyB56wIThZzSYnjTXaQUPogGQWwqq2oKJEJTvAHjVDVmwMTfYeU3BZu1HpNULgNhq8
GhPF3IoFeBZGqiSsdDfTK51SMQjeUskycqDbiAQL0JxdriwIUq8CCoNKQ0PmOcmKOrGUGRQs3y/P
bfbKOHjdcuaCDU5klMfBMhLN936hWfC5z8Ki25fdRUZtObpPaAHnHDwUStnsFF3ZutjPFWIrtjQq
C8d9QPvheppshft5SJGX8WgoaBQZsrdNGfCDFLBDhpYaRvuhvzVCtKv3SOgdZbijv78Pk6UoY6DG
0/GIdpNwK66lhagIMccLcqGJArHFzSm3xPXFnGpYpyJU/fASHuEUlFc7mOCRdUPugagEhf3izAf7
WbgNaDeWqa5vnLlFEBW9lWe0ELjGbITJBbGBu1qnjeA5ELQRBnzFtc3BBhGqDFUJT/H3koGDI7cg
4m1qkQwyabe9Y6+YHchH/oXQky6Egn7J9a1/kFm9pDltMaGPlOfang+C8/ttgz1LyLqb1sbc5FLf
RztrBdGytjvk4BGdTZD8oBn1PzEoUpZsVR0zADI0zDATexeJzAQjwde2lvjhwgz4L8azf7RAeHiI
PBjYNOl9b8ioUzVP6L+oAaiRQpNdRRTIgVeav/vLNXiP0VJ6Ww7s0Ld8M3VJbuE0Z7tTtmSnsFZD
kn2uW80ny2FDFztxQaGtJaV8bf1as+ookMHZRRoQPSRR6yiZTAibRI0JWrookxSGq120ICmGe5U7
1MM7dGIs3o83runnTRtzQu76KwmhM53igH0js5z1DlOKeW2rUM8SAsqpyWWM67KzcfQt77t8lebm
HREwdNCFrX4fx608Arc1qZCz7vIGPKsF358wfLdtxApr6BeBujJtkiKlBfj7M32U3AqmYEmVjcgy
OTwDJrsLJyb1hRucfDBKpGhIrB+4PX/5hrLGo3OkLOuuvqkUfb4wYkOMBd21689a/qYERnT9dga2
EivJrvNZRHCORVQC2449sb46EwbknhPOvvv4XlADDfXyeLBXbnUbp7foqpPGO3YlTCAH7fdlQ59r
6r6cE91GXmIWJaBF8QgF3V3LfhO04Ev53EptItFWtcG1+TsCs8XqCWA49jqLqK9Ca4RNrXpyHG1N
/QKfy4o2J5D3oaRz3OLQK8+WQWk9FDsZyX9hf5I9irLeQOmxmOr6XJfsYGBE4RehNHhp37NPuu6N
03PoD0RO544qjrwhVFyJwvapUBR3Vw8vgeRfs3kOUqOA9c6RzLIgsOyn2sNpVC3/rOcSwHSeFujY
NVK4Ktu0+NGvbz1GEyrJOFC8lpwgYXadQMMcvbLAg7y214h4xd4y6DWeKwYCg1eH0OJZZ63/+6I3
qgeBAFdN5LRvg1nEFXRViIJ3ithXEEQQGyyNdKB0ns9bZFCic0DCzf4igpUv2eFa3GBSZb1wiupE
+uRCJ8z9aU3XE9sKxqr31GMs8enpLZ7BwW5gsz2ew++tKqFTyyJ9BxMY1n1CSUS99bww74N4AJ80
idQSWqXvy6zfOzoyeOGO6s6NznXjVVgYvJfpQx5c4kH/T+RIVqV+qIwH2cAfZUxsEiohIGgCEIPl
nsd+E1YBzrv++yOyNA5q3kh8G/ik1owrQouGojP5hXFeaSE8utBURy4H08bjpejTR11BToMuzfKn
iAN0NUH/yc0GPs0K+4uKB+potREk0vjXtTH2qEDosPuBdnfs+EHiT8+76TCCTTUmITWwGwOo15t+
0XOP+p8PVbTk7tDQp56LbQmW/wOdnAtfcs7gHkeRZHCzwcniSUB+X7nIPCwquxiNwa3+YGlQPmOA
v6PRhyWndjoxZbrMvkYiGVDTczhWaoCElj1+9ya8C8ScAAG2oPmG3iCuuZEAp6dl/M7fCMVnPEgT
k/KJQmxwLsNLDgco1jKE8HtUbTSdJK0VWLk5Auui/KVokqY1Dfq4lrk4l9rn+jeiE5pXb4Nx0x78
czmDqM5BWjEuXE975ikuUZSQGbb5w5g9wYGm8RYj38HLu00XxtqUO8J+ED1PuXGsdXlJVmulg1os
LOJpbxEasaw/eYvXYCKV9yEbN2CEC7vtkf3yKc/SvqaQi+MQrnlkWemiMmCJoHyRRNkLX6RfTmRi
CNovTcSMGYPx5Qcj0UPIhVba1vDFEOOTzqlBakpsXFCcJBPt6dopDlc1MVY78+XbeZAlD9Q1rAnc
yizqAA3Q9zqFr+iVkP3OrNUSKAbcvheTp9lWu87vC21duo7PbR2AarygSbFYVpknUA78OKUlOSTQ
MFlfac9qUkF88EZkUlCNllX0DXRbNsB8RhoG9uzOzKkktHl6YQWw1KC/zWL3kB3zzgwDucL1f9Zj
YtfOaDr3t1INZceny+wWH6egRvYVAcj3t0XzXIASF0ylw93t1EFPeBUwjERxyZhLx5oOGbwlrvg1
G7lcZkD4vPAtRHMSGE3boUIYgdUaNLF3E7xNnYqOA5Fpxy3S7ZuXf7zM+1S9do4Xe9NoR8HlaupP
jyc4ZXj0A2eZ7X3qM5u5FQze50ZMUZFJCIiPU+kM1aUuMN3wpSo4jdzWRmNcGU4QfQGn2Y+C07ET
0sIwh+ZUfIGggdQfD5UqJ8vOFOM42UmVwGGt36FDko4qWXfa3B96E+6pJROtlOcumraJfQZnVvAK
cUC9twivRPA0FW7/2kfcKalzDZ7lEwB8fU3MpNB3RAgYXz7Xm5o0wn8V2YBruR62NpPJpiAht4gq
hKXI1Y8Iui+W4E1O0ZzpTx2OGc4gOZEaRXEEuTUsxnipyDTexZQnl8BMi/t5FLsczVb/K2X6QZJZ
CnEj2T9tCSk8IdId/a/Mr7MqhNbNw8OuvWa3cDg8IoXwAKOh53/nPiFvdp315lCMyVLfjHq2/xlY
PxGq+vuMwWvgy5n/MAnev1/SmrNsgAakJaGuqzuiMqWrP2ItNvZGghI7ZcXGi0bgW56hbHsNZrVk
Q/sIK1DlisDshcx+2It0cQizovbX0FqPSt8NyyA2puLyx+XXT0S3rr56378/c0ec5H1abwSJOW7H
8QDn0AYtHoiuwT4FTDhpQRQJlpL1FIawIHR1wOgAYNgw6msornVmsZnAREbjdbvkya/FUARJg8/p
dzRgdWj47P29cYzq7CVhuvJwMNNJvehFBBdrxQTG79U1vqU0YmznfNR8B/HctzjncqcLmt2r4BYO
ZiYZI3qMSumilyeEGbQTnaGFRbFbUzoC+BE/ITGQqct5KCTFdBJqgFjtE4hqd0KxqEqhwkcL7nnf
rQK+tAota8qxznKRtrxVRDX7pFW3H8Ot96gCVeSKKzc2rxksEPzoKJVcYfa9t+yGTVHBJLhsYQed
qbBcDy993kPetHjImCSdPkj838l0WfeaumPQZwXnWielNuCJ6OjF+hqcEdiH+iIlQszWkQe5CqPb
YzoCzelsGz/PMOtBR4Xi8oH5Jz1zof4tiJyCJtx/beInttOUggDj9EoADoQcCb9xBoGB0z5fZ/nO
pIrtRVKEyKu25drrx0mFIBgsGanXSG5wYkbp2CAY7v1auHE5Ldhp63XAJ+ODplLzQLs4WWaSKu0Y
3uua8m+AToVLkap7MoK3HBOdfUec2Aac50kQCPsg0k5/NcS+ArNJi41wHglmxvjusDKC13ye4lTB
E3dJBvVxoNGmX+0Mav9+0EMa589FfCibUKYLAY5FPXeGZrL+AcSbnwjqXTp4tXDb5mUYuysUjSG7
lgeG6fSnSfHvLM04xcNVMH6xl3CvVWud2ZVoE1QHvJq2b3tgAKsp/H2LVhO80M2tlkzblOE/PTky
Z7FqG/YmBWp4Upn0X1jWMks4HrceFCIK/H8MOelEBu69b0DcmkCrA9LLvcorSrPnji+b/ZWyBDxQ
m1ere+j2AmzIN4BF/fv/Jrn//WGvz0ibSqE9eU3AfI68oFb5beJKUvwNQXb1pvzN9VfEq2LtMDSX
at7nl0pAoajg7TzCHqp6ETTuyUywJuhot772MDwI8me7JkPwY2KfEqV7tRKCz8Eu+OLg4mXBQukd
QiuW6b7uT8mrxxXKSVOayFqYRRC4vkhwgit5+PgD3zMDaQQqyNT8P8E8vMl8PSVrrctxygiu+wVC
Ukx/619HBit+j9qxMBpxx7osVLmbIZNN6yJco9QVpc9E9JxXppemqF7puS2LHwyOVV/fIa6v2x8n
7oxpkRPwmNwzZvsSDkr/oCCUHFyYydWY6luiZu0hUkH9GwYnty9//FvIcN5BjbiH26FIjkOmtNdZ
noeLlL8qr/HuY7b0ddE5dFV3S4my2tc2I6FjWXuzY6TwAbpeAYBtVts7vHGIq7TZAe0tckW3Uh2B
qgI5DJbXMtuS3PcBMtdU28F9WYLqFomFN/UjwqHuqkXRR7eUS9+lb5tqbvmql1Hu5vC82Q0G6kKX
hDkxtr4U+48IX1WKwDHM8YjDgTbQoPO7ABRClpF8q/c4TzQ7IzUXvCGpxsXmmx1pbQYusgX2vYxV
iQD1V10P6CwPeupW+74UtjwHM1cOsckHFsQNKs/XZbpIl82JihsdYvEk8DokSx+eLsKUDtZ1inB7
VASfSz5h1paArnYzI0FwzXWFGVZiaE8zEu8I905VK3lzCBsjJbMdoi+XvTFMOBaj35efsPS0iajf
dd+IkOokI9+ShSrUf1xbVVSjYjPecfrEzcdZHXMKdnuki8MB/8Ga+gVELCCBukQvC/UlPeBNKz5x
Efj3Ti4K66u6djZRY7V8aAYMMscn/MfZa3GP3yW68k0xIm8oGuVTLTH0k9SvadAzMDbvGiy3NZ09
vamdTpw8xMfwQxw6QhYG5l+AodQLTmpld1E8xP4zemcYpezwxDZJ4B2WJpFEtvdVszyZuL/2O3Ki
VwDG8MzpO7b3Q8WGO6HuXSijk+7omC1Pa0tnLjLsNPOMrEiMndeb2YzRQV5hzPv8nvJL3QPNyTQG
g1FnoNMvcWDbiBiB2oaSt8Tb37GB1ZkfOKKmZW4Mj7u+9SjFfsRZg8AY0RC2H6i5ASqN8YXwwgNm
b34FhlPOTL1aV8gAlztjrxMOz1KZeKGcbL7k5EPh0M8zWKyPdcuPu7smbYbb6rMdpLRuaePvkcdR
+21/uky5g7TnXsx3FY7Xcd5LTA3SighAvv9Ging2bBZXAJsVj3B+hg1z2ifUmjJeItjHDqpLx32t
kj1wF0BlIqtCmrAJjJnhE6kX4PVbTku4iK/6CYiqKGUThOsRL0oPNrT8JlmRZc13t2IhKWXrDdJV
jpim861AZi4hx7fVY+mcesVlfgirA7N36XHEsEq2kjktpBy7gl1xmYR4+iQS1KLCOvYJLOwm0/su
8B103BiHcxcNQrMqmBR7MPNBkMitlUYkEhHLSgWmAMAFLS4HOyPvoLjnyijdKrIBF9EUZQ4y36xY
7vtLyzcKmTNgP+A828y77RgYTqdhjWpJhrJG1/Mk/XkRsQeN/SOvFSVkAIQ19lDKc3L7Zb1MqOQR
MGgrWAIvduwhQaIMLjwwfN3yugkcefUoN0YnFedQs47EhCYNeym9gxPa+meoQ1TAK465DE31hwhP
iQAF3LIqC3weTm00VE9aLtph/VRJx6305UubhqC54u4IJhSmO3wOgzdBwv+/vWzsTr+xZjFAytAG
1JLaMsvqP1eG/ilgYNBBZseouD0p0YzAs6bNM7a6F9YC8hfo8atjDICS/bvKSclnsyF8SkegnB7N
KS+VdDhxTWv/xWf51ybOcwwYux4Lgxljg4Gt4NuVrwMy1UKx48/APo8aDi5BzoOhSjNd55XW1H2Q
FLhd8Jm/lGqaK5zE6r6Nsrn7i++daxEsfzWREfzq+PSE//jcf12L2MtW+4AbtfV7+lgqgC82KDt3
RtcSLbQrieIwG0Y1MT9J2/cRJ5BPaOV90ZrHEvlqQYiCcBhzuQOYWOp+UrMWR+klNPSNaOVFSbl2
5HjTbGOv4JYPZoLq5XrDa6Imdeuc8PwD8jWGnfLp7rKe3QY+ckYW4hQoTFCxH+5RcBFTjVY4m1Es
V0CXEQUgSS52Av9A/MNSdPxnskU4KsU/0u7LQAUxkdsHDpTHIx9XBxMbShfd7ZsENwYXsFsM8tA0
W9Eztp/NMZClOMmwlAXXc/b9csy/EkV+OAvMUPJtegliNqTEeGwOT2EDsLI4mZohiRO/2/5rlT2J
avBPUzPnB0o65GSTvBll7KFDVsbceQdtpr51CvXuuW3//Ud/1WxrOzJbx0JgIvxul9cfLolunG9d
pKEUbZm1DJsabHVxlZsPqhGooh9UDoabAUZKXlahAiC+REHaV6pcXOaptvWzIZGdfCVJrt21FlsI
x6SS+yDJxt3Z4bTo/yimOxEC02y9z7pYCet4L2aDcUoZ/Y+JPabt+rRt7jZjfMbpSNrtGSXjtgZZ
IyMj967l7IPJeBuxySaSKSDte2KI/lJP9RDttNbh03D06f+3knM23rCismq19A58Cn+wxm+wefhV
BwsLhCPqIrv49ykAgB713iF+VqJoqSp3febytdQPblCLl9oLVJrV2J5j5Mgybsr+4NEynFQMZ4V5
aWLXZ4uEg4Pt9YgZaqCMlXQFlX1qTON0kmoXDZBE5Peeq28pqkfhiJyhIVc268rdGyMI8vkWDRRa
w5J9sxbQf64+71xRoOpFujRt1V2qwd/yOv443Y/NUX+iWfR+vUtugFQ7qoG4ifTvgyta0Hx38nEY
+aqlXxW1thjuLR6JPliAG+mUvBWKznWZw0xUfui5fAwQav17Pz37YlNRqNfEvDiMWHmZnzim1VwC
qxpcHo2YsrIGT6zBRrLGEea3LpmKhNM88evVT5uXdfUOPKjb6TrB/qNFTyvtjlhfGe3dYyPs10u2
5UmWBoNosUeJ3AxO0el5/wsyTTs+/IfMgvGpZq7L7ttI4U5XrEYlMJeV5PbHXda4VVMsNW4HzLTD
R68K/TUgYZIkLzPyl4AVfzP3D2k6p0V9dCJtd4yPWlUDIQPcOrGcNb/a8EE7uazK4/PgviRuvHEW
1k/g6qsVbo6pj8FHjtKxqXo8tyx+D/APGxPq9pP/MROU8e9o0QjThdwrs8fpriSxjFZnLH0USMP+
VEFXUEhme7nXCpAEYnIz7ZqL60mSn/CQilOI5wF9Q1Hv2SvXXrv0SOmKMFwqZxcaoNzbPapxUZbk
jkPxfpWNmT5xaDZqS01nlQYFmxi6aqv8f0668qUk/KxnHd4GnL8MIKdYc4r6n8CroPTsaEAbQQdQ
F3Z64gj3gNq7qpzlBP1KQ8ugVH7226VxOm/OqHaYgGEzfw/aeU49AELFM9unhhbCpJin9NJY5CtE
PDHGGeDY/nrU3OOI544mjDeTfaka8IU1UflkQOmSSV3nYXvl33Suq1aE/uRvWev181J6aAId1+YW
1U/nut/cH9rqzNLLTojOdeAgaBFeD1lYjG5Cxi406lkUvc7bHr3pfGkSAf6wkk76otv8jnjdH4Hp
pdfc2LBFE/QcdvXMuljnc2Q9nzdmkgYqtzf8oUjH+c8tzODwDaR4E5Hdrd10nDD+WKoFu1ehIatZ
Rb4PRspOJPffNRTINQJAoPQy2gpzmwRlctgRe7nF9KRXeQVGks4OW/yHmZSwILS5Hws++lVJnYKA
FOiKfSGOJ4KJ+ZBgxsa4/Hzcc94GYVkduAILzFtRDs6jEiu/IC0czsLKVHHF9G5X5QYOQ3e9FKml
redoJFnRZLuKyYqODAJl+AF0cvElAJCCB5fDMTBzBpc5DRovEEMve7gBrSDr9DLgf4he2Vl94yKV
/tUE4XWwwiCnVxaUaEdLTbO14nDLo8wraI+VTKEmGqAXvKwvas109qaQSygOI/K72VjDKFkhoOrX
PwgfAi/9AIzEdsu3wpnSm72C5OcAMIhmKbIw/43fI6tdU4v58O0urhpMsU8G8qg1vcN8Fx9IJFxI
UeKtZBVrN50G27mdamoJTbTgSRVx2niMIuU5HxgLNaK2IShG1jkZLSskrMc4SkhCtQ6YNNqHSteA
KX9RybhqxXP7tK47D+SBX3GjyO5Vb15huSh91W194rj9w9NECtGudd0pCqBpNOn73EK0uu4QpTMP
LeilPYJcImTViVCsbVuNTdOCpVrty0qAjeoxYY0GI4VS8y7vKrCKX14YMr4GvgS/ZyCg/6YltcyP
wNbHvHlHWkb0ufqEjNBGKlLuB6m6A9VwKc2xZP9x5AdAtKC6EQssKZmqZnVvu3i4HcEvJC2oVBVM
J6aMm4Q56W5XF9sk9PMZS6xWXC+QDYJU8ZS4OJqILr1b9+6Zc8/Zys2tSnJ+2mC3CuKSsyrFYWh/
Luwe2s9xRn5E7VCC85//VJi5dQUHAE2WQ1T+o/ePY5dPPh/BRU2s5VAT3RwsoR8t/RizVqGHJyaz
H+xt+SboWHlyFuqSHjMjZjwiWOfKAsQtxFC0LpfU+7YPtiF+dONOAkkQKOf4YZHZoEVPtP3SYQnA
nro6XCDPGGpP2z8v1Mnkdg5t/4/doYEh+JC6Z0nbZUrhOfXB3MSQjrPJG+a7iv9rQVj7EfK6A+Uz
HuRD9DBDxatQDk9IgLBt4JqdDpP/Fv3v+kK2mkDIIF9TPYFjK5gi7cJn23sS8T2R4ssknGEau0M/
X/eEBKB3usYv+Z9NJmZMKvzo//gQs9KcZSQE2bFZJj1QT+mn4MBynSfp2TG/TdhrxJMg6IR+EEZC
cVfMA6z9jth1flefZtb/piTBF2gvpQnl3zTTjJWS0e43vTR573J8DLPoIesuA18karOu4l6Zf4Dg
FE8Vlo8u7A/QdxudIkSA0xJHODpmI3gVhKs2JBUnTEOqeR/f9x4JrQfgYe3yxZu2kCqGSj9u41qq
iTILQOYI6u3GcKINgTkIyEFfJrgxFnYPj0EULu9teBirSgXXqfsqAIsvv89B1/faI5/vUZ1GR46l
emFx8o9T5CxTlZ1QtSAhDBk7tw/G1wWLXNVJQxApEjaBLDBmD7C3BI9stLja6oDhDP/HxEd93P28
E+8yUHTQ+S01Ou+oeazRkO7EXdPrdNUqpJkF7KJFHlMUptnkwSUFX5VhnUswhZ/lR7Cx0Ugtmef6
DABRSL+HqfGku3FCHMpDijzLhIhQveNvJyhsCAuQ4dhOhRNg0DZDChd7fsPXz5qz+b+0cb06HtUC
rGaj9Q52a4Q4I6UOEG0jFouBntepJMV8h7HGMKmu3OKYiDLKATu+8K0G/jYBaz1R2yCyh4G4iwAW
ahU1mC7IabmWhkHIAOf4nsYI4TdxfcloLzNE+1PH8lszUYGb6hGj1XgBuU7ND27G0nnt5+jLWB6B
G1x7G6qI9bH917vntLAtM7mINwdsWP+mrUxz6tm5xq2104ZbeKOTRs3A7B3uguRTuy0OjPzr2nWV
KgsrHx8OQ6akyOc6VFgOjC3I8Nj5ts8PrXNCT22gz0QAzlUiPtBmFdKvk2B8QqqI/mz3Kb1of/DO
jVzLY+Cs6AKifyedbQQbjB6ESHZ89/JZ7evW5OmCV61wpovnm7/19YuNlZ8TXk6Pg21nHGOk80m/
fHnBlLldC7OV0CYxmLugYCUk2sO2Fcf08eD78mbe1fG1tZF1qhsoBLY9svB+kb+tLCc8uRpwrZVk
B5B9JaNgjMooWCprHL7c57s4wROeo0zuHYEooomLnS92p1pkG+WEqiUZSTelaN9ROemRDwDlHzIS
PasypYkdRNZ78xnk+PWwSm0ZsZ/hhjb6msWXF33PRW41VV/23Djc///+519RRFS6+IbTEaPmIvHr
G5RLt7AMKxm1jgqAq7zjVYrDP8xI3/APjqXUnWY8DneqfI8M72cQHjG1tXIYqpcsEBaddBxzUW1w
xWit2hW3SChvWbfSMpg4YKqRpxN6iPIR4NFwxhqCwZd4a9piqEx96etgykLoWKHxlgQpkOU8X5Eq
giCwwz+r+04cfGsWHYUSU59X/qnwdap4R0L7YuC0DS9jICGbjtFjFbUizBQhnTU3IgEpU/KX+bCa
GALa/jTZTG0XEa77SpY934Td0blNWZPqzeStn+/fcPP4Dn/8wwImxjQ7nehad45Lz5ba3u1ztFUb
hwePQ94gIjvxS2pRLlSfhlmS2QETwIP3TqdoYBYHqgU4Mg6ndqa4RobaRv6twg9gNxwWB/wqgTbo
lsjFyaqVNh00E4T1knsAo+oFnvo31US+bAeFTQoYj/L6YblS88nQxI3ukf5G6Wk149gXVu0w8aXt
a6/xya5P2O/XfcgSE3o/rCQLXd5WHbH2jBbUWdHUUJ3NBwNdhszplCOBOnAtQ5ae7APH709+F2Dx
k+oSe9qsqU6lQyLjwbapjDISP9gOsyUvoIAB8UaUWWdPTEqkX9LOh/F5bg7YQY9KS1CQ0rxdwpPt
AYnEV5QmxxUWdFzoNDW/ivSdq9O1FA+9EnLLIuJXTRe2ysFWLeNyQLP0Vw+6nERnqkQO9c08vFGY
qkhJLWKtfGWdw6pDakHWuMFRnKmObfc5tARtd09bDfebfnyA/9k0rFrT7SzAYQDW4M0Kow/SCDJ6
f39bNakMg1/R6U5eAMM0KfZh8D8cyBvVmHsvz7I/WNvop6fKTTRauEk4zGRrrPDGXYJj2zlV1ZsB
3qDgzdQr9Ev4//zROQD6r8oFKWIP+9gCQ079IuTz8D1HDg1ZNMflBaetbJcXytdObX7is+Muwrgk
fK3u5V0ekoDxtK+m2OIhfSWG7za5WUVWSoXloOoJ8OvZvd8Wdmc66B0C/QXEy3+IwwF4e+Gg6Fkc
TZ3RScs+5mVDjWU8o0dldGuPDpV24h1lAOUPIwTp1Epc3YDjM4MLGQTmx8K3xezNxmdxfOKQ5d5x
wIsFgtvqeoORYB56yjZldZwEvGTpuQTuyoyXWukwb5SlNKpFRMemVOQbdzAkd2LMaNxnQnuHs/pG
4CiLP4nbaUYBxyTQRzuOIb0EsPqnoDxi49Cq12SXTalLB19fuFvF3NHxS9dsySuwhPgXim4tX25j
THJ6fBQCNWeg0WB7Ib1HqU6pVyFCh1Nl1rP9KLQgWopyNrRiOAsx7SjkHPWxJn6kTyyqIR7O3auO
ePQSWt6fxleL2FHcYrUSV+zCEoNiAK6XHrNh6J1S+wOUARK/znW+QblNR4RBs2qUJB56KaupkF0f
HT1iRmtCpvaBFAzFbfPlHMZh56yHAStGQJ5CdOKuU5ZUXM8XgLKPT+WgEP2/rN/srkeGeBIdrZ+7
vN6GwtIi1QY/lI5H5fuV5SmpeAuR0hF26xu1JYQ7xFCYOJ7IL3M+ISjI1hilPo1lF2Ph8NbEhEp7
YDLop6L7UQzqxIYjh4KTkbOc9LfDygwikC3DBJLmJmfGTpzLM8MBE6KwkCaiJWeXmzMo/kggHrf/
4WVWJtE65w8efl8iMijzef0rnfACwNVczTgamNMRAh1FZgb8mVP6T4vJa5zjPZfVGu3vQiv4x0O4
tdX4owpMBBdHgbSmocuxY7sUnGiyMuvPnvwyIiDv/On+3irCt/EQr63mVdl+tgjuGsVqKEmtaRaW
4AVAali6+HBkfGIJCl4zZyjieTfU9L85F1JPH01Y2poTe9jsbF8i0KXOPalaSVfEvUF/UbiCtkS8
ltwoXT4TbZFYYjg4f4+c11eDAmAzw0dSpQxcJu9CpCt/Kz33cCkLF5W2WCywN3owlvZ0wnlpzXD9
ZRAxTsplFmfPzrOj6Y1WvQKkgL5sWjzn9VrbaUdrzQ1aP4cY0ksttKVWaCS1q68IpA3aLdqlEp83
N4EposFH+9MX17FrIrxBRE/r2kHpMTGNIvgFFDJpWV2wfSiadlQnVa3mkZzIpjU/RR180VCXceF7
6E8p+kqoXS3kwzEnLGg58GL1BhSZxS9n13FqiixT07Gjb0bosmMKw7JlapU/21xi9azA781Zdyxs
jZbK2nqlTOlNox0sIoT2S9i7WsSUJ5vjfCgPyVpC5G1DLl1BMh+Q0BaRxVADQyVRbpQZ3IOOcVmZ
kuyfFILsL6IhVFBJU44r37cMaqPFQWHu2ywOssT+8uGP+8wnNROxYeLqAZ3ifv7LAsLZq8Sr5oox
vMyF6NK01SBjHh1SdcoL5++uVTOg5ycHwUVb/x6xvCcL8eVwXX2dzkuHo+qhkTuNLK5pwTgGrHJR
qwoV9kYs8lKzGtf2xAmt3JW843REknz0EQmzd5OVYWhbzbkMm5duV+GMY2zdy+q7FmixHI1n+jM/
l/9RXjsSnViHDh4D6cUtAi3EZnErPwQdSXTx7j5g43ggOjQ1kN4qm7SVvlvahe/0wmHhxiQ14Aui
CqPuZpzi5B0hde9AQ/7Xu83ppc1A6o6KW0M5phcZClK8Qpw56uxNOQiRgk5FuRG5hB74dy8dlMtf
lfFO+waiOIhCo1ATKv3EtlyfQaqTu9qEHwpBaXW+EasKyt5i0pAl+gKDyOt14oRJkLZccE6Wpoj9
2goC1jySwvJa7X/+9ZXucXxZZIY48wLzSFIrYgfYNFGHmc2R7u/pG8qV1qtckaN0W0FiKAvuJbpr
eMQJ0nvr0YuO33nGUMYXzGYPqeI24SJcsI/CTCkUMone7hlhMGm06Icdgc/xi8sMUe4QL/NaKs3S
KEoq4+Zb38+XQHL1D0w6aeys665Nl+yTSBUHbRrpOUf+8FXpsIXkWzYnlqCh8ROIdMYVzW5FBgJQ
IggONLbC6B+U3vi3yKYoujUsUz8k3IDpwdsJhiYqZ9lyWBQnVZnhr2dbUlzOFQjCKvMHtDxEPj8v
OuTIHWLyOE2Y+VqvUuY/HTQqPUMHGprx1RP9PstvKhPeKNy6VF1HqJASU3YhzZFSLR9QAlzEPzdQ
0hM1KktEXRyKe7mu8XBTHOMQQQfOtuC4XigiL10y9APVQq6HOIIdLudd9XSoA3HqIHSenwoRkcvq
oAzafD0JC/jzAYZrvqSF9eSe/DlVOB6txnF3N+JHi1/dqfZt7BLFMg1E/gNLEbqXfhiYptCtBhsO
PZ6iUUOQtolgWHPnUbLxOiALacsz8o3QRN+MZBDTw6wc2ae8AotlhJBNySQKwEWmM6iHCQoq8bgK
aplM35O9LCWU3LzTwabykxz1Q3akAvpqWaADHnmBd+8DckWYBvWYDyI6PL5RpzxKuGARvE8JMsbl
nuuRFgTafMpj3tf3ukQuvcGQjWgOIY1HdmiDqBN46GUxLgvAF8sqXm9oonl4AG0+vbrxsHSUiDI7
jRSaot0LuUCoVPEEoXqDx8amP04GypRjMtLLiooqPjScUxwUHuu5WUSjraFpYGlPQ443dgDKsE0W
Ho9Y6vz6ODcbs4Wjyh0CU3cxUNB+WirEW2rWzbKs2yCVLjeBRqrkiD/LR2WkSlTZINyvxrTzMI3/
QCOrL2+ulT+saM99U7r56eO02xQ9LAChDwrU9yNt37UDv4JEgKNT7X9OWh8nWhAW5p4gOlw5xMDY
6kZT/k4/tbyNEtzFxzNgatWmNR4Wu5Sf0TdxSHojGEw1MnaxzHskyoYta00ltIRybkZKDdjzFnSw
rgUq1JSdyc+DiOkqWvqWYBw3pozJGCeGvN9024bqOzQ+DjsxXbbVcsCINABCafAW+3KTl5xs1YsG
kdHHyIU5ftWzD/4mXR4jkqC74sra+xjyWN606LXHDLtnQ/2BFPkQm2ECsrDVlJlL0TDfT5E9prXT
9LqIgGR4aTIS63uK9xci2UETfxyK3ShP/eedOp+QeJF6YdctdzCHD5IX2UQIBu6M7c42F+TfFEeF
Dm0MYKGFJrLbub7SzspFpAnWmM3YprWWPrPQdDZk1eXbsaWqvGPIfwYD8QYcyQc0XaN4JwfVLaDC
WJ0PtWHk+kI/mP3Ld/Hq4+AaO2EEaLCPAXGCPxYpMc9aQT6PbjcI8DtF3HkKRXjiIiOLeytZZHAc
unKn4BuWYnMjzMskdEAjyOZS/ut8fftUnc0xmZa4+I4Ru8ZKjPvhwjuPFE55WpkxDHLYIOT1cSIb
m2vh/2igAahF1VWN8GelnzxhkXOdC83Ik6HPcw/JCYh6nk62mj5GFv0fRA8hVG34Fdqps+nKlFoJ
Jh4nQu2accCC2psqkvCdRvRRflr0tMGhNoFk15QSs1wsfj4cSNgXPCvtadtHYXiDcrSILdfMquP2
rB1sVQqJ7u6nE7DgFg896aRoQQiFkMgVd57BMzOA+I5SDXt2EV1IyrQcQs5NLcSAuS/sfTRZYL0l
q5Kd+JJ7B5CRuB+/++WnUwUBRnB6oOFdOxQzZ6SM7DISqHWQo0LaMtlprmFTyeNFCgwJ/GRmpS8I
0f+7GyxYmiB+RhsSYGrYPjSNgGsR42a1+L2NhY8Sujurxr6Xt6xtDAY1g/4Y6ZnaeLn1OA4crWuv
a7AZaTZhpDH8ERk5rJXy5K0ATbYNoKkLq/zD9vFRMqPOa54nk2sfBRJtGoXLFfCLjFeC01XL/uMs
o95mv3xCJ9CyNnHAjMohvp+lz/2Sj2ZKW6Qn688M/a9eYUimaoTnZSQu0L/9ygR8cmS2a+xRe8nV
7TkR4XivLGVWxSWar92EB3sv+h2lXtpWS8lZofWGUx/kTE0kQIuugUzwpEc0dvvsIsZirNq+Q3Yp
t72Vj7oTVynvvx8OD2X+Yt0IUNOVdrTE4oLGozU0qoGQA/FSI+30BC91TnSpifKN1UF8H9k+fsF2
DWIa3cTj6399gwbLhBaBClxh1+p4YKeiA+N+cNz05FNrQY+hzdp7h6eJjy6vy48MnrokUCXie+lE
mPF7niuDtiTUHUewarJdP+0x/Ih+ZUyQos9zDnsLF3nx3l6IRvKAxIvleRv4s2ffD7s9YFQSR6aQ
lsn0Ki9MhhTLvR+B2tsW++gEoAySL2B7hId1ZPXf3mLxXNcCRFXO/Uzf9GsP3gLTZVeXzJGrEcDv
N/m8zEHwP6VtwN7hP7mi6WJ5s6Q7Vdne/+h8wIsKZpzaDAKmHTXya6tx2iAtEVhbO+sgoiuXamII
SsCozRinYh1LtAqcKFWPIS53hPDNjjLR0A3uy1kcfI/Rk3kZLgS+xMRe/4UflHgeKAu8vabm3nRv
zjv8XLfdEdNekBup1B0330tN6gl/FrtFhpSm3Wxw64cpuxQUP+nXhTYNoKTxR53bAbDB4iD1uak+
YnAZQ7/5/m8+KAvapWgi4Jn8z7rOYGzqLmmYgeLVzOpI7TfvmL3RAW1T0OQeTtbQW7pDgG2itMVa
NX3X1h1QH7wCP79o8gt4Db7uIah2/tnz8qZgy2b0eO5DWWRXe9xsnfCuQgv58WX+C/TLuj/K0dxj
4QUAdpZlyPdTQLA2RFVhnoBTOVn+VB85V1uNc1rLljBdbQYt4SEWIeSP0U+adP1uHWfXTDwdgn3T
AVQxKigUXObeSGMwKoHIg6T+kuBjVY8dyklUd7CacKw39FTsOUVRJmvonfMvt8Qb9AP2IVr7lteV
4Pz3YBRdp5LrbFG246p6oqTtxsrXS28wrmZF21gyF+JNzsjg24H2OirDpgAxn51ztlVKKWNEBD/h
IuH6OsZyay+t8rijKqlXepykSXZ0dbFgRki48wkHd+b6DAdmogOmZ5iELb5BdfjqFXficPkyVhtU
BKy4nvGXMA974/e1Cmm/DRnGiUZ7ehsWLbXDVIgKOj2XZ/fB6BNkr3xENjGI5HVWXpST3j/NtT6u
t3UFX730403D8rZVjFoLboH7NXIrdivtPt/blnieanLps8+UOFPI3KlUcSpEgdXqQ8WI7x1KJdLB
0jsdnfteKDq/mulGRq0RVVo/2f3lnBrj9CzKKVy56wIEzGpWJ+8EOsdREaDWySntUzGxoNFyuKKt
GcO9Z8UCOCqR6TvYYhNYqNL2RU8P++YY5tSHB4pf5KIKO/21K0iuF48rvkznzJJleISY16Mjigm3
VmXioI/MUZcrPZ3VAmcwvhAOIgtp2G8LrGh5G3hxreR7T7wv81wSt1YvScdrG8MgWDsARF1YsIdn
Mu/oYpx4ESp3jhSMh9rxKMACrfMj4n6yV5mprGfMDx1Gm++nxpYVnOCgXBl471MuB7bMHZLEg/CS
iNA2og6xMOdOI/kBtWN1dyjNFbdliL8PzuPI+V32vYXmkNU9PZ5SwdrWwyXSKGBFEbEAip23yeaM
w+vOsEjXSR/3kwuk2XUIxIVrKSY21AH73F8lGu+6X5Tms62vWbj+8g4vnVr6VUlh52t0hMlGwas3
S0xFwrxwlsCtrIZ92bTIiUyubZUHgjNWl/ICTJMv6npaE2PUQLXuweqggwAD09ucYrMUPdiklRXL
yf6IekjhBSbL8mcpJ2x5p5mTapBTdg6jrPqSkb9nIGrkE16W+vIWBZQem6w0WDcWqdneT/60OoUr
pbycO4/MCCmWi8VM4SEHtSXr7e0TM0hkl2bZLv7f307oQWl0T3yIghajNf5XUhhY7C2GvmPJaa68
iMd9TpXTM951XA6QTqXg0fJjl6AiijRBiHSngrKEXVEaVUM4C45gx1mpFOnjmAXKhyziUe2PVOYw
Nq8j6YxWjg/EZbBWM/SrQkUBMTETAFJA+/Kmk/ORE+UPf3SJP60dvqTxfZa6Yb8BONssP9l5jkXI
oG/nwfBg7Ps0ejCfEEuamRfwFzY3kv0bqFQLCoAXw8fUKj6I3wDKjXxj8QSuXVvyXjyRrdTRnbdp
lt0q9k+fDVi+xU+ioCbPe4QJHlytrMD+rVL56nCQthFUpPLtvR1UcZq2GOvnMfW99LbTrOCf1dAk
4GUXXA9b2lRyJX/BV4Rt4EOtJFLrM4PRlLgpwKy/RGeQUyshYu8zdGXGLiNzNcR9aKz8OmNWb4Ab
VWKLXB0GLcOCMhlef7HMdMxHf2+0fQREhjedgJLDrbu7IsCdnk4CGccog7BYe0mAcbI/+fr9pwiR
dF6EbIsa/IJUAOJquRV01yrfuonXPx7DF3LdIITkTKUHqU9O6pXMvlur0KJ4/cjtWpEAOVU8a6YC
KAZdecQpg/ehNPZ3DWMHckdj08NHEimtGxEPd80xlFMyB+i0kSK6myTDBHr1nJfzIMJoR/wkGc4w
MyY+7rGD+JPbfWKjdyFprqwHLEOSIAisVISWzf88aOInOrhJ6vXklSvdfwc6/bdKE0AgDVOlrJMd
rBgRsFqb056iL/TZ3XS+N9PwZjz+leYtz2TsGLX35nJIb/3SOwDKo/HkDUOTxjR1nExSzJ/wU5yT
VbDOe1S/ZFm9EB5DRNiHlfYfNopMbBLCs2490G4JFNwKWI6dm6enMcXTy5pN/kRO1ss0/nXYUoaf
JLAmM42WxaAVei25D7j5ApOJeeNPaq+4xLswiY3dh81TTfTqsjrA2mBIoLzb1L44sw95t30eqVaI
zSV4KZbztj7ap6YGkdaKCTJkWX5YzTFJ8o7lowDgZyRdIHq/QelgwpxmY5Fo+6z8UqxFh3qcqTw/
2qRqyagyLM5T7+xVuDp37ceRvdTcrifMz4I/f3p1fm04vpMRea76TDC7CSnx3N0sCfXvT2Osdv6x
/C1kXr+5/BZDZdligZyUEBBSmn45cDXbDuAPItPLg3BYweYTCJDxNLdq3IZX7jno1MJlVjuV4yB2
J1IxghOCrDh9rZhZ9s+/l1P6zC1LY3rsh7q1FMlrUEQlr/cIYfq3yoEEezNoodpAKamEIxlv5AJE
cao8uEz0fTx+Jdx3WcnQAHfCfy22z33nJ+eA4ShEIUzhk2rRO21V7BzHoystfjpfZN3Dbzwo4nr8
YSZ595rrogfioMlzYZ572oWOg+V/FnOrWxvxsuoHD28g7UDiB63MXc5Jo4XOOsKHsheUjxTzlqMT
Ge1BDxeSlRkNatzQKnvbKLXWcfV3WbuCDGxKVlBUHnw1STZJCH5o5OYhNr7/+CxU64Y04mzB+zLu
wi9ZZ8JSY8/SzI7Y0x9ewxUNQ+nV3jF/R2lupVIO+jL9NHpo0qudGTIa4khcG44eQwqZycvfwU5S
2JcrCWP9pWY5c0BCm5+nC/3sUrHfR3268neOPNB0ZABhhzsmu1jqk0WUpVt+VQEqp15emRMKJbgU
WIINOJpprrDFuZIrJRlUuOzOSdG3LYdeq0aaUCIGut/SKl+H7/I48caZCS8GXOl/c6ciBV1897So
l4wF8MXn96Oj047es8USwLaimtdihzgrhvvcwaEMKWZnUoTeYNpGQLD9QO5v6Y3MiFxLkifGY9A5
lwPeUuoEzzJ4LRUC3oEYkHjLW85sRT/TCBMah4M8He9Pr5AWvjj9sRQFTqXsJdjeiH0dLZJgENoi
PEF3KK55GP4XhCBn/+ZG9UNFmK45OxyzPJ3f2n6FKcxZHKJ5WwD4a6GC7S1sKOy1a/jv9n+0KkFj
C75SHCaC8CTAH3bd1T1kuqwicO+fXQJjzMtcz949tJxPVByImAQjpzCaMrqoCrT+VX/hwgNuy4Oo
sQwT7axHhtOlPN6pXB0xD3/Nc9R14NUaqriUVMS9FcT/GdywKuTcdt/JXOkSCI5Rm6oKvtdkIP1+
lCyBAmhVhFg0prT0TGSkNdvwKMRQDDdFF/vv1oA1eajeJ8zJgXcwNCPlUV1r82H767/G1avpgof3
fchsp1H2oRqF2+SedZgv2mMYXWnp7c+Fw0XvRg6jwtsP9DxhGCcSwP80glUQ6JwYs3SpeJP77l9T
zCesqsQs31sAWmMvCs8LpaQGa5XggQLHHZ27QDJ4CxA0n+ghV4f876gn9iHCCWWny3sYomo6nNgN
ca5wjC93nVXyQ97s6+ZImFDEL5wmmnMgKjfb6Ht4aBKnuLOJvQTZ5ruMpF8uMe5ZvMQZBT+xcxTm
F4BU2wSpgHaqAO5pgrC1cWTRiQOrvOMhSfCpyKGL6VT5pjthcV5QtXwXdIBb4JIqR1GIjJtTRdzY
9qm7KTqS0TGB+/NnK1wy1iUZ8MtAqYHdi8xpsHq2lu9CA9NayRKnzD6GDs2lJd0q9UZgrkeIUkFN
83nJBM/y1qV4LH/N5I3051RTDtqrnvj3xASB7grY/VwD1Xxju9FMQxong0WsbaavZsfjLpQXIRNj
4owzwSI+MRNNon9nhyocqaihNVLI9wxlFWAWlwlaN7nKGSxfvPDJAN9KH8Ezlq3pJfTbVxKuExnY
kMT8kpUphqjOOaMljpid7p/9d08jW0Il25QD91foglld9JGAIRLqMNLghc97o/6vHAmcXA7LfHtK
IxB7ZHqGc/NsKkJJ/p47C5oNZQzz9znKZlINatyH0Fn+OBjDogxxSx7dHftFEdcd0ZN4PKHYNmK4
sXS5/JzwPlmA5eSD7Ppf7qPgyxxGvVt+lYxbxQFtthLmVX/EPTRbz6Yc5H3wiJzhgpagSTt1A9hU
Uv2hfriTk80S9ybAS9Bk20e651RWPVbmxJzkI6BlLsfC+Q0JA4ClXSXmNUCSdEKdSS6qBoWTlJJu
kcIgqhlX+ICGtx4WnPOVf2kO6lMUYkbKoHLvDNDnijU8S1n0XsiDsMKd0FgpDDhlyYI458gPrRkN
qXMurUjvRFMOyHUjjUUGx/7e+v6M0lhDN/WtfwIKf0ZvI31KhYZ0vf9eHE4ur+3alWopkeC6CM+A
s3gmYjkxActGixXrdJ2SwIMBxXZPoDnQ2VmLMG1iO/0rLpL2pKWtgEDXALFNb7sw13JmPoMhpIBH
G49Y89PkLm4U9lL20m1l8WAev9BjCPmqt5mMXmUJY2Ilb2dCiLS8V/ZYO1oN718yN5oWiz8hPGnY
DL3dvsWjMHEhVEEvdPNbYFxM0yf1aWxQm8s+L00DMQnL5va5nG4pKJDbSznu6Fhw9/6UqBIpF26P
ZdvSCnjNCf4jy6vocKIYj0y7DQpycPM+OX8o8aQg0goH1Rcz4ZWpqN4GguEcGBoiddfXlAnr0OAX
q4LwbljJG7358oYuoQ3g0LYUbrw1hsyKWZyEpWoGhh2klhgS6wAIPlf2ijEufJpTchP9V9/ET6mx
n2xUDounxO4S42N4RgCsoamc59LKEIlS6ap7H10zmE6aFY6Di1rqHq+9U3ymSSJKrKqRroZFraOd
FhQ+eiV/adZTquROPxTRYB5hBr5DfrfmL53Rux3yNP2P4+9/Cc07GWH+nLtH3c9tdX/qPXKnx5Qj
LxEOhV8uXY8tt9F7AJ48oSJtTsMt9RwtorVc47sfI4+O3WXzTgvnj7jyrgu+8rmdQ24NX42EKzbu
p6EC+LZH0W0EGwekcwN5raGCRmUJg7liqkNGnR0fK/u+UQYN0IK/5168ffIkNbaWjsFNP61CqrzB
CpB3IhSWgrxfCALci/XzeNHBKA2FFgBRyPYoVMUJU4/1S7OYGJd1kl1OCaENfqNfPw4CVLCErTn3
fx8EYIwlXhY8KcfbFs2bahghO4xOVFFMwxIpQReXVc10kmWP90WzJJOX16UpBvASKFR/VL6f556V
z/6IyxKB3Am109K36+p/UXCWgzWK3aBIKDDlaiTK9K8Y7SSlmYbCB8f8xrXzNhdxHEPh+UZGQk+6
PpOW+pj21+P0T2XMX1sn/3SgyrDOGv6Weu5UGZKzvyZbAkAJzTKgPN8vmfGi1u1E7MwPgcP77yL1
zKG5oo5/XWi03qqBf5ie4WfTe0txfE5KzfbhampAjAj991/bqbiEkwQHxDSi9A92fbZRZokBpkof
oFssNJLCiQNTT4RgdMt4jYy9Yai2QxvnSZO9QhHSUP1KprvI5dyu3CvPE1uPqT3WQSgUASu1+9T1
etuELEkdWTaO+3cpwuFBSofTVQK/JzAETRoZi1sLJHGSJDZThyhLT7jIAxQPEkiKR8g0oD96rjVh
ZIbnD5Lx0Y9gBpajV6p3JWqdRNGfrqbSK2SFOfoBCSqXmOEX33TteCUqe9eoX21ByKNk/EE0i3LC
G3vEaxpuayhIHc2moFzwUev4gdTk4GOnb1YRXOg2sNl4zblxoxdfqYDUz/RbaRMJOP7Dqvgev20S
AV54HqTVp2GArrRXm99XJtrrX0QgV7HXrbubmAFxMmi+kv5bhxAkHJiB+/uLmXOiSfPjrhVm+oL2
kw0NbwVHbRWnQ5ljE9pNzSn+hEklqTqp0CtSBMKtu2Q3FoNuxOT8PQUBksypTIiEf6Abfs19UpZY
s0H1zv5Xf2MsmapD41Hm5bgjEcslxUP10yqUyj8VU+KHLlVAtOtMiDhAA42jFAOVN7plMc2EVWo5
iIUSEjGX++vcbAiOmRvdyToM8rbyIXOwLE+YqUePkjFOIPOzPOnnAgZhEf6fd6Lj+YFjhSGVNQYH
G6oonpZwFksA4/QDESCoPPy/idIAIs7d6tIzU3GwMwCdTwu9Tref1qfJ90dT4N1GRIyVnYUCS2tP
QxiuEMwy7xJklA2kmOTQ+XI7BL3/kibsHyWmzDQWEQpmJ9sKYxAN3wMkOtQQMb5/3Q729kSXDp0F
8SXtHd+IL7HNZvDkrAb781jr6SYQK8v0mwW3XT9jMRh+fmzu6n55yQC+R1o+J1D0kvbZ6KkkeFzF
lPcwfg4akaF0mNLd8qyAxdXNm7eImkJYa+Ok3mKE64kyGTZVbQNjeHjtWzOLy/v4zfwzyLni/3i+
LSvcTX2RYkhRXK7rCqmM1tH2rlAsmrAdo5kQxQpjMClILMs1LT9dSPRmhVcouklLnJP+Mn3P915q
YEh9nVkCdEYBC69k1di3AU+5e238C5SMbJNIVx+D21AYJcrXHuzQkSzSoetCr6rBKD1pycYpH9we
vLOlmifNEUcXwdDoX5V1w3FxNQOSIa3XCvbti095rSgiHDgDL3JExvxKvCcmK9Bg0cFTKwfzmksA
jJpYC4z7e27M0ROExamnq7R2/PWZDLRyT+NFutvhX4ior9nUwp2qUNWoPFD+XStdNq2cunuDi8VU
YJtsf7t11W/kffgoYOYFrTUU+9tbqt21msVpgeOQFDpu9E74ymbgPjtOUX4B8knG9Ot/H/4gbDOT
G4YQPkqpJTQ/7xfgm/NxU4lrXsRA3n7cEtf4scQng/7gd2R5B4uuVAqUH8xlIbNPs+63yIhYozuh
pAb6ZaC8Gu19fF1DdiUJ2PXdSkhlXk5s9SmVOerp+8Qao5SGFs853PvTfzvm9GWw5zQB65U6hnSi
uXOACkn2sI+6qSc7OsFiKkgpqZxn8TD9F+cP0bsD4SEh0wRPBkiANbkDFj7w9armfux/Cl9WKH+u
IitTBNkGVgX8l0r6KO64Vo7UKcpoTgiNSqlfjChM2oNFCMG0ezRpNxieGjWO4YJSiRmLBePYkkJp
u2VB9uKYcnaxxBsekndGZPdgTahil0QzIkwLEvOQ63scVhxatFFM81rz7Ap3o7649o0Zf/PNalZ3
HUJ2yzbFWM9JNa8ngJ8xa+jBffKua7089pqmVbUYdSMBs58wsrR/ARLWxVtS0/YRUE5vsJvZuSOW
aruIQUzv+rjsQPakKNtYyJ9f2wU2Mng55zpAdWYeuJBp80elomw1zz0NGWHSytAIzXFcf1EP5R+C
CtKTk9qxOR0mVHbhhWh4WZ5raPX1l5Fg/8VbhQHmxZYel/DJ5RR2077wjwjdGejqTRurDQLkkdpM
SIkoS+ggKXX5jmA3DN/wle+jzI9MSMWo6bPFixa1Nch8Us36Xjo7/MrUIz8JjaaBvlE91nWTRNcw
ZJDTs+4noRKIWQYgUxr5iwq6dHw9h8spdvOCbkMKYp/w52OLrOEFbm8Nxa0S85feGlb58wUo87c4
7BMF6IiS96Mr4mXilzBCBlwKi2DB50cbIGehp8kNP2TrpbeST2Pp4xFSqMZ308HbhGiFiMwLyw01
cOi1ojwHA6wtNYbgsG/lmW5AeW0rRnE4aZgsSjQPszf5ZbiPFZJApAe0d32+Wu2AVqcoRcRwz9jk
+aImXXLlg/Ah7ZAwV1miDkjRHYRvDPnJ90yNTahku/sgfcan0LFmfUpgjGYkKNw+tQZwAjdRY7VO
GEKK5XC+HTccTvtOX2Y+ul3vEO7jP35WQ0b55GztcQDPIXfJghndWU2sAnqfZsfyob7O72DGOahH
HBOrB346lEeDHIZusphCrUGz66lT0fwMhrFfQnYp1s1j86n4jPkMTRCqbsDx3rZwPcaegyLWeFqw
9I1oJQlJeGqGnMitGTVvVBlqDc6362yHHhkqeMDGuSLoUqpfarh6/QWrklbyh8X4lH/Z7jBP3mS1
SpBV1jo+SiWDDwjQPWYXMMMMXyvOkESRXqbWu7mPBr5p5NvyARVVVVlXWWpVWKkuOAZEHmaes12k
LNbYzC913R3xPmGuPGGkX4AFbybLCapEiZd/LxBqoi6SMX6GKbXgv0kF7hs+uGWhsJ7RMm64ZrMw
xbL1mRAr1MtTETB53dy8yZlPC0hxAiRRHioySBKJKvyvDt+v9QXUevikQVbith0Kczg0pRs2GGtG
8VRgpq5eh2/Jx9QIZoKQGzJCUFejk0qxRBuw/78p4Ht678bo9kqvLwEkd0qqkApe6ImBDBtqjg5N
x3MU7d3GPr960K6fFfqgJ3c2fb/7nFGg6Sgh4297XTjBno3zLHNZl35QAeEekjzr1FIH0nYtASmm
CNkHreSvk4o57bf2rAmnfsYHLz7i+9MRvr4PAsurTxNbM8n7WtLPvp/CGyx8jjlQh8qjCmQqcNKh
pWMW4l1X/wF0k38x2fpz6kW8Ff2QbLwCBEHDcR6zgB3SZ5ZSm03C55i26rH5a3P6eocJqoxn32Sz
kViUdAVmXGxesoLkdkdbImosBOQ7pajFdxM19yfp7sW8ffiKsxFuAvKb6kjgR7EIQ70ARkXFiuXR
QDYMtkoT2duXfX51+POxv16Bne2MA011S3nlypPjnhvzPNLRR5D9Seu4U0/5nXAJKD34S1IOtDby
oNZrcpaSoRfcmWidUSAqb5ZcP14NOCjuUe5eE//ZyVf/FplSz71tX66XuhuK9aR4XegmipWoQVJ5
G4O2pqU89ktit1pc04AHH+5DOVA5glgPxnUK3Yw6+zjWyQpJH8qhVm8p22kKMPFgBdvtzPwMlKn3
h6knWH0s1wpCFizwH8apcrQCzpRxeBAPFha/NCMjQ0ZmN8JFTdgIosCIalEToZGEENkL57QunSDD
tEfawZp2miNfIO5rEzhp1N16gEhn63setRMV+4h4v1qUVehSFek40txbdwSk5wHO0ihkp5CrMkxQ
OGdcopp29szYJAMC4csl7etvahQo8pqmrDSYqH2xcBWZHzmFJLMEoziUDntSWXJEnNTptaMdMLiB
hH7oMImeD2jH/xBHpl6zOXVUW4Vj5RNE3NnFMpdfeSMy5DUedliHd9lN4vHqE5+owAZHca5suFhY
GSOIBURyNFJS2FSGOzCzzApgFEe+OJiO8qoW/tdGKPetUFaU37YN/cThSqjrdQ02fCPISsZwlDji
+B960zjDz+C0+ZAAITr6q0Ut1NqbvTpjbphBpRV96FldiwvOfJVosCE9mgkIL5uqojiOITXy9Onq
U2WnxPwL2tPzqnozssGVxu7tWwBov4as5+VkXTKJ3BY0wcZTpo1ihrhUl2/KVlgoccSVAJ7pNQgL
x0E/mW8weULVpY90TutTQxO9YUrcyg7FKafR+4lYiADNoKYbCEcLEvuczQlVP7umjgRI/Ajz3lMg
7MioYt7oY9/akf/LwfYVD4pvMjr9sy0Zo3HHyQ5E3Qt88yQgnwtWzyrSaK8AsgZ85TQ/EQyd/ZHm
lFQ2w0grnluGTUlT6UToEs3GbcSl2GRwkWXiiR3R9BZ1Nq4XVLe/JtTU2jTCOYMO43TrvW1HYN7K
8lEshfQyGyjImW1Tm7Zh7PMOz3nNfdeWHIoduHIgcjf0TqW2hDHfq6yK+KODXnTvVIGAd7QTIMsZ
1YK7zLCPBNg0J1hP9o9452r8xObMOd6MUIMVvgao0kpe+DuVNiTLXdduYR4/Sk3OYHW/6Z3Qgt/W
PlhcTCYCIjyJ5c5g+sZeGjM7lnhYIHiJMBbHT8cmNUBLzZr+BUAO2lJJiXYYx1KFk4oOeUOzb7h6
zUo6j8hM5/nRhITKYPjIyl9ydpG2vTPNHXwx996HclwZa0J3ug4ZLwUuRmrlGeIzRyNKLfyr0LoZ
V3vbWr+mwrmh+jv3TfsBmpLwYuVx3N536drldLYd2Y5bAvfk/iWUAYVDtGCe/aV65eohgoTgKWBw
PwbXlXdYC/LacQ6kfwGRoKl+TAlhbcF9qe7dk+AQOz6FSJnJuSeFAg8533BFL3/OZTTzv5qwdDqn
W550JZXcQcw2iG/UXYCN2Ky7U8ZrTAEORMdYZ5Gqi8ZEqS5eNVkdjSgABoBk7vLP58qOB73lAhPQ
7GaivtlMdn4ZZpkwYxEbN7i1RVIxRSGeU/4YoSJOk9b3iPT5ymdUcQKUmwJD9y9sdiIX0TkdyI/3
uyN8TbvhcYc1I4yGOgGNDQK+yJEBCUDQ8p7rYtJLYHaOYcjduvqGSApIDVZ49aBpafiaJAQVSNKM
DBXAILCVOefshX0pMgyfR5Z66CIliCqJl1S94U4hVYqLR8d8uf1hOfFbQUTbTy+SN+/55GspXzrW
8NSwwiRH3STVdmM1i6ZgG/G+N2A1rxJO/ohUALMA/WOArlsFDbx7QocOYhlFKCpzsDRGulQwuGDI
+1frqsg0dK4jTl16GP3eTJt6U9tmo+7XjtYv14eTChMvS3x+lqybCuw5GvZZBSnxDYoGVCGb1bC4
ePqNgUQqw8bZag022fNbRBX60r5H4cHxcuZ0utek0L50p+qmCkn9Sc/Kt14hLNYuFXr0p9sS//dG
lHVtdhajtmyRBWPNHzQyrp0ay+Qz16qdPXgWlAKKshuv7ibkHZKjJslKbAzO51My2IUwGcv00ITP
yUX0HaAmowXiEn3ZbkYLiJngT+GwzsGlVt+2qOXeAFu4CVOM6VWipkxoC4xk613oLBXPmaIP70MP
lz6w5j2LWv1yD9ilD0PpU+wwuCY8dZvsvp4sqP1mqlWGmJMncLecNw+9nP8IFm5W1yz46iSU4MjK
m/GFBa0rTanQldqPAcgJV5iPMmb/f9ihB0I0OierbQYTWgyz2/Xu0dm8cc6/CRFRq9ZTSJer3Afn
/LRG40pP46o6dmAQXZVBR3Qr1fuu+9BSlAtXjMOhCTLVnvmHiUXgEErD5qSub5fMzcaSqht9aQsd
ifvSlknjrwVFriB0WaSaOResIyg6WKdSIuajGYc2pI9O6CMagu6Ez+1Cq0k9SKcE1078rj1pbbmq
GtOVgANt1QXwBU/gt3XH+ngxAs01TP/r3ZPOe1jA+K6GWIu8VTAXexzgDpPPVWHm3cxe7xchbxaN
r/xcYNwf1Ebzaif+h+dRj+YSJIqpiQj677MnJEh7lcEnXrm0SFwZHv3Dp8cnr2KgytjK/HmfnSLe
B4m1UVnDL7XrbrFWluAABx4Drns0kan6BaXpDRixl7ewekFzEYKMzI4qba7pNo+mpJI18R3OF/5n
Oudgy2Y1oQIrZxXTA2nhhM6mGaQ8JLhT3zQl4FY1fEJ0nWUWh2wprc7bOAY5tRBptyC1VCLylwAQ
6jwVUwx+mSMImcLfbc4ba1olBVfdbDkK7hMJgvbINFYjDjQHt4WyhY/f1KrYZ3bM1c6Kcg14tWFr
iq6DOdrhnTL+63alcNUCpThUh+aLOy6Kt8psfp17n88hq7mOxT3iThpBSb77Zf2OmGw26RDroW75
MV0WBRFN2J1edrg7VZzabiFF6H7YsbmLMgfKwHLQ1wcsnafOl9pCg8seXIc4meEZqpbKGpt8Ispm
+IEOmAunGq/Zl6xbbzGDfw8starKQ1Vhc0dio8CQg9bPl2sfwdT4dCxjEQzzD0eTKN/3Dotds/hA
Bb4pr+nr7RMnxc/dviprttEOB1KgyoKRALInpBd2fSMk2W1qzwGsy6hZ9lrg7PqqQy2yPFe2BzxT
oLIrWVVvQQauhLxhM2/Ia7M/E/sspzfkjd6mcjybNJSxbNzIPL3nQ3Ay5CSWUfIh7EyCl1bIiiOM
jKpxR8OYfBQ8h2pmlDK3pTJVHpNTywBRcv8Etej8ZuD/pg5ZC+C8qgw0y9EgNEz5fjbsnS/hfXGZ
Y+1aj3nb0LDYFvF/43qb9O0LSU2RvhzN86SJtPBsbYEp3LaadK2whaUpNjP4vH7rj35AIspkHgcI
keTyeoIewqVZy7/ar/97iKgZjrlR7fxX2jokNxQ824sbFFe/Vy/Y3ExhqtcecB34qFLMSPZpMlCB
g2/DC0zLfa9pHwPtcUKt/MikvKE4W5l4QwiNMNplIPk/disCtRC6rAi4H91TSgFsLFFJI5cacNsZ
gMMjbCBrF3i+hvr0l/eT1W3HwtRRqWR3qNnAbr2PZQVda3xvr/muY+4zH2plpjskZDqbgzBXoJp9
q4lsw9sCqDRBB2wZl+iFEd7bn5JRgP/tk9D6nH4UvDl0HIaP/SylNwdr+FuMBVwc+DfgJ805td0u
ZkDMYViqvipmN14Y+CoHUWyevNIQF8SfdISw3GpSTZmPdVghvK4CNEgkIx/bqXrqqcm8ltNzZqAj
32H3CxhSQq04Jy4S6OjCaNy987q0j81kAafcrCZmRJVGQDn8YlhQ0hNlXaLNyTPNBeoKInO8k4E4
uAzu1O33blnQ9M9B0y8NbTMmziS38Zke0nzrYSm3hnP3hO3hMtRjLAvjjoBdQuzgapQHym7A7FUR
9dsbE5Z/bzqu5qIdE0N9yfzqtXjMpWjXrmbGCdLEdd/bLG8fkR66XIjuILc2ZREA27oEjpJ2sSSu
zHxn1rbWHqILegBAEU5N9CbwTwNjoCD3qqUuf3d34mI7MRobmMu2F+6Wp9+sYpajYhfaXPRHtmTA
6phq47dArQTTB3Z8paRl5djf1iN41465lA0ojk9HV4zoWPAQbAhkRLZ59HFfqwtRs2Os9JWPLQ1o
zvW5NcQsF08GJunweBpT37k/twS37h0rU7kP0BlO4KCYNd8ZMRvUNrmHQwRMQGWv+Ge1v5yPeeVm
XK96UjpgVXJWM/HY9aeMDbpmH5QRENS4GmbJYz/ybQkiBJBTp2f8Jqtirn1GMlkRiKvxxfLYwJTi
bpLrTIotc6qbB5RwHIwHJX4XZZfJZHjAeGg3I3EnDXSYmjxmtbmAZmzZQAsS9ytI9GVxt/cyaUEI
+mA7ltVNEy3DwkLAs027H4KZDJ6EKk1TU84ne5Q/j0tT1SsTC419yq7SNt5yL15JXE4Fo9bTQnuM
35PbHnPLJOvuo6auDk2l+ywgbSLfO9daonA7O+0QtUWjlY6ddEbujJEGrC9TLs2JQNPQtWsdvS+F
rtcTK6czzIi5fktIW9GPPSgTQ2N1T77zg6uL/ruzJRv5j9OVae2kcaZlOxgUdakKcl2MsHd9d1WE
P8klWophjgUtJ6ocENhZbxBulbKiDERAthYbQhIS5z0VgqXlV9yGAygDsoCGDkZhg9+KfNKZl2DE
oNYDsa+V9yASRZtfS+xTHnyxsdJtbgm8IANNGK2VBHSRAUVCOrKmoH+flw00pBE+x94TMTuaaIbd
UAv3fmCqvc00Hppgt4vcJC2KPSFwF40DLacL2ri51dk4mwa8RsCFATkgIIwYDsuoiw0LaYKDjbyb
YNlsblde2niQxVysF7TbFN7Wrbc2eDh68bUeEk/HjdHrcwGL4M8eNnzqKQstDk7RHKvxwhbrENkL
c6a9DgvWqJV6/4zy/2P4nfTdjEHi8iIo7SKTluIq2R/w7wC+Kj2iMEQFN8Hqm8Iqc3S5+7WwXq7V
bFAiiMsq4oIwZSIsfwdxdzIh1xWkjH21Q6NmfbNF0zTVsd2dhPFPelFhfGRN9xpunam9mP9CDufD
1qjPA6QDJgZRBuzr9pvAF3VrNxGefjQg3ixPSpO48eQfZ9Kk0CELMwk5qdF/Lcexg8NdV39TlqRu
4Y/ztZigoOQZQDB+lAV52PPLdx6UEtKucVIn6BVP90yxhrE9yUAu/YW/YHodwpYM4jmrc61e84Fu
XxY+RM1Kh2aPSjHf7fFRVUj6e5Se6m1Ypd6Wxj0+41H/c3krJ5U1siinHiCOAN6JUSU9j6kcRs8Y
llDlYk+clPfPXJNrOWZCx19w5a0CXsvL88f8DfWFHlVnIrY7XB/avMAmpOF4lQ7VDKcXUIZSOyG/
Jalm4GA9iUQ/XhTbKy9ixyQBtULnxeF96ycXmvU4NNKPLBlwl26vUy29CUu/FierG3z9a5ZdLv6r
c99Ow1Xgpzzps8E1eox0zMDkhD+vlNDCZGrrkhlYBRBB1mx0Swu1RowpZila8ERnqfIC3DEQK31N
7dL9CyKcIeClMaFgKvmlYF0x/MnW5OCa+wNHAWRRtFEwZunwFs4egvVo2G/BZxMpM0iQ6ZmzeIBO
fJQLoMZw9QZFPv+/q5megS5eAZK7VuuovHYqM9RR8kQTGJmoOllOH7v12HzU4yD+xgUEth+on0FT
8bq7YudgZWukZck8p4VwvQW+sreLk28WfJuJ6UFfSb/pNE91dDrsFIIFdoNoGkfGzQdazeW3oa29
ezfwPs8UrBAeU3J9whxr9o3e1gVaqd8Je/Ic9cCXyW06Iv32ayF+ve+owJZagnZStBX5NIkAbZlM
LJ+hT8pwGO23IbfHsSciMDD9Te6249e89nHEdoj0p+osNe8B1vs/IpFGBp8/MiAPfxGccC1OwtVD
amJDUhl6VAEWHKCfQGdjRQAlI+OVZTvwxkIL1hmuyQkFy49NyYxQOiZzUJ8krgPplA9F+KJ7+GRb
IfZGdXXXRicBQV7JEW29/awW6eBo9x14lLO6t2vyKQ/mgpFlIzBnV0XoOolK1DRjTpUjWY//2uMy
G/EpOoPwBgSeG01IuBrBVdKsaRHVsh9oDpepDBIQeR4iyiv6d7JU38T8wsh/wHUzCUrEBBYhu7Mn
F3ZRC9DhBZusYnjKrqmM3LSY9MSXHlp5D2SgCunmYJM0HKtC1ptd1jIl1CxXiervqNXvbFGJJYnG
ZAv3DlhfLit9ZoxuptpE5vyWGUtKb3jv4q4CKecHvlrFlLYj9WPhixzsAJaGHo/IqgF9V17MhBzv
O1Erg896Mxzs+3GXVvPUnjKXl/pdIrf/HqESmlYzicU3C7KhpnOspgBVWTbbTq4myrwtbg+wNtLs
XdbBOfQ4vOM7wQX1tCGbR6i0/U590DFX1Fww1dldeSFrh3tMm4j+TF24QDUtaDugFytQcUyVYmf9
QY3/PW2MEg12pn9qG15eS9HM8yhIx1kA9+Qu9gyjre/E9oZhVC4YWs2HIrPPyWpOGXCO7YavTVKE
1NecQnkE/GkEE/HHzVo+2RtjrvqxSLV2sSozHNZ1LiJ1E6Vwrwa5xzQ0uL9t4d760/8LY/GkwDAx
HcqrA8FlryaJbWTXYDJIc7gLRFaaZw4UhWMcO7VmZuQdSg98xsGvwBc9IFjUl5HYxgxzUZGrcXiu
yHvbg4RLuV0CxcnlXDqChqgzHs5l7T46sPg7cOck5GdRsfc8Tg/5gs0a3bcnFhs3/SV1liAd/cMl
Iu43v3ytYiWi+UgrGzjTS1JsgIP+mrmE+0K39uo0CNIaDQ/njvSDh65bMsYjGlPc+qLaM0jDkr66
bbDfikZi0cYuk0Mh7BBeFh4ORat+ROAnYaaUvql/zuI6stNmnVy6RIq07kLGcti4udDBmBrd/IKQ
2hHdIizyR2LEdWkG2OSPsrChFvQ1MdaXKvSvwAEIcjOmpC7WuDAXdiB6QHvAr/eHD+0r+dnGh14s
uBuzDvB/KGKZUk/Bk9UrkcR7FSMIPRWr+/pgPZHvTZqCs9FKgO4oM2gC9Uo4qAsWqYd+PUUSVppR
bXJKWZJw6w1HPx2yjNX7qYdUdqDb59MLHGCHZIdjIkL359xGqzTOqtb40YRAVz1VJvQKnsmmYctO
nuSeGDF7KfbW4CEU2/ZATDmy5V9e4J3YtVQElH5k1hQyqvJqomEflvV0AOaboEiIhVuiWec+TPPF
YCBHquCvjAfWXDzXGGKubBXKMLt/04llfLwaqG2FX6e2u7thMt4UEADWHScXKmV3EvyzjVgXhVzP
BZggZ+bkkcRAhWSzOO21NrfOYiqIQVN2/6DfOs1yywHMrxKE+JH/9Qhy0Dw7SJZfSGjobv/1Xmcz
uYaIs8DND5p1iYhKlchG3y2pmKtxz9hEMJY3D3gdYHttqktp+F8usHaJF67w3xH2f2KAvsv/Oanu
wkhM/oAd/+FwxLPw0jTq4DmzfkZKMgNJ6izFfyoihLoqzUWZgDtdMMLaPYahOYiodIBatZ0xiujb
ov/XFmjUVpB01jdnVf/+uMaW79bsUdzBZP6wCms44dGaB7jOdymThQWS+BamkWerUgBIViqh7K+5
G2g2Q14Vg2BQb8eqT6GPsNDoolvr2uA5lo6KswTypbFMLa7EF0Pbe/OCBZTaUQfUta2+dg45NvNq
DnCP6nu2Uzsi6yVGObQQA4TQ8Esd91PNurn6DBfzy+q7cxWNeqHu8uaOKDrjc9tRJfRPkbrmPYLr
IyMKPuIZzaRgkxF4rsGw8T2zk3qwHYX8tB9zDRx5hgjjx50X1SWI9K8RGaCC6juxQSp3qKeTm5hJ
Vntme3gSA7jwmHElDiyiIBOjFadcFMdgaBpdbqyEKXVjyQQJFN2si84lZ+ixgaZsI2Dg+O/Ce10u
Wb2m+i0u9nAsPodtzLz/QepK6ezjbW5yyvquSeC2s5KtHIy/F74wMCEPPYidg9Gw2OZ7yhvIQd0U
TChb8duKagUXUPra4iqcvMi9YPsMZFk8qu95VLs5u5mBEqzQnT9ragEUW0dj3oe+nmOZJyAor7DR
AH1Hx6s1KsUsszZutPfId4sLJ/nsJ1+lXw2OHvhatv9j+KjojoeCINLXQRlw7hP0wGBOgpzqFTEl
cjnSXeUK1MP5KQeeu/wUfKxBak/JhdGV50ymtDSEqdI4JHw3ADHj9K3TEBqlqCq9d5dOTFMB/D7s
kjIaJCEzaRoOeNkzaAV6bLbsmCTLZFE5oK69cJga6Bg1ceYdGRoI6KPHthN82641gp8A+bY6YoYS
tBr6Rh/YIOas4r3y+RbkFDdzKAx82wxbPnrVa8Li9N/G+1qJ4OgFVM656hDABV92cI9ER3oDzgZO
04bdH4mIA8u7jJdzmBfQvqP/JSdy4SxwubCxpC3iCjUtK+o+RqxIz7pzQz5XH2O7yDDFlaJAE4jb
49+6u1cTb8E8Ebe4Nz5e5yGHZNT1fMyLc+XvpoCG1h+/dg2U2RJfZrEzu1G2cXzOEN7e06CDek0Z
cGka0hfI2sRn/r/qYBXM1RkVsaQx/UAvrsVcaUoY5rhbznD+2Il6tfUsFdE86I8A/XB808XDBFe9
d+L0/7/jmiIEfRMfUL6vrhgvtl1KVXal74FdQt9bWnAtCa4rnXQLQWKiL7WurtfNS0h1zbNKvCBn
WZUomUb+MNICoDZ9c9Pk7Z1xdiY97EvSIH5gl+M7+mjDk49BEx/GyDZAw6MOX8PU4Qe28/xgAB/z
KmDQirmwxSIzeE2C7hPVOza+7ooKjZtTEN4maqNVJ9efppmjQvoJmPtmZEWCIujokbRh0Wljk+7b
SsyKZOR4SL6JxPtDf+u+j2l8sbEJzbOserB4gz2ySSXUdzhIo9BW2pUj59RwLbejqJCyUZI3Wey/
eSRKKZepzpWjNv8Jc/6RIwMJxnKyqve5GEAm15SEeG9qYV4puOTf9UcBoSd8jXJckLL29U5MeCWW
EEs44mMUEHiRKVEQSTTGUZUIJ1dgaB7GPVconFA98m4b934ukARhyqUnY+isozdAhtbV98Bf5E5B
d6S5NEpuJa1/esF/RSZuxnQ+27SFkf1/7/vd71c6nUTOoN212/kFqIxWrbBKBhlyaN9r8z2PX/Pi
uDIYfFgjK0rchKAjDuXgJfibV8lmi1LEg2LIMlrZmGANZdR0p6ZBk2rEEO/a2PmabsF8Sjltn4qL
nponAgKEAU8ByEeofNrS8AEMmOgmXR2bHEMQAmMO519kh3nhpXIUXS7D3RUO+N3ey+3hSyD836oN
M9RYEgm38zemwLBAXo45d4k0qxYyT0sG9cyyw9STvQkCIm65dgPOq+Hv/YAn+DnmE+/vwWtnbXxo
CFxPm53Xy7v3lwY32Geg5JZuZfHbE4TpMvZEuIhNRYG4e851wjuRfAUhyxPKF4iKHxnAKawrkrQY
IWHnFY6A1KC8cN2eam52cpVn3Rrh6HPV4p97TM/vFp/wez0vRGKLEwvFBwhduuTZnBNk9SFTTyiG
atHCm5nVh18vHClVHVMjNWCljd8xsX7yfeFfnmRWEwqO9ZrTEv4Lm47zr4FmogR90YURY+MYb/za
4RN0W3M0huelTrP++yC3ufTeNdk+QUqFPt4H7qTZX4Xsn3TeythCDY13gZQm1//PzgiBh0J2M4nB
/OP8tmw4Fs1RPlwOe+jalnXuU4D6utkuty554spxfsL/FQI1YtrTJQWUBvx6BkMxCxTJpuU02vwI
BTihSAAzEIBRGPYLZ/61ZfR/C7CPOd4E8Uvi3+ALMSHwDxBV+z01+KyVNMJla5Le/JWdCim/0tvl
9XrMgX9yI+haqlwWSFZRYFTayFH1/TRQMq+8rupcWD1uTzuphN2fkCs6pSy9Lb28MxWveJPfeLoE
oEY6F2ogrdw9xV+PQMB3dbU032dWvcFCz7H1TmhOry3dhEEufIrHmTVIxp+7rdiKsQToMl4ZaY1R
IHypo70FtAEXd05/HNxqcDCqZEZni6GBnj7kSvq47XXdliu1U2QiRcMl35KiNBF0oq4/3Kj0IrLg
1585o2ECu+sj5kVMuiDzPg+YasFTAMoK+pPw2eH6/Yor/8mog1VahJR6Zv0Egpf8AFTkj2B/BjpR
sqMIXczAolWOMvVG6dZUQQGH9BNFoCHA2OQR1XyXK6s53hUWec8fxeHslNiMRnYqsMI2NYzU617z
pip76LR/WMUmKbuzfB9/ISVRc1Kkb/9SqL9+yn84e6ZOeDfPbfq70mxqoU/boQTv9Y2cZ77R1aA0
/PHVqbvSmmSfmx5ShJTgmrfx6z7ZopnqZJAgv4jK0qvmDjgoJkV0T6r5C02017eba/zWnvBjCrO5
u5QtMtRi61O/l3vRdr/g/BsQ6HqFAkcVCRnNS6W8DzmwG1ay+MpWLBO8QtyN7JRLFi06BN3H+CZn
OP5o6168YJNdtrS3hb8cEbNU33t4yCK4y3nbm0vkKy3Cpoln9VESiRn20AYDhNjKn14nPoBv6UYr
Dxd+Hxgmr62hIT4EeeY/C8jUA38b3ioyM+8Z5xgUIHFAs+Fg1D/SM06+SLB/v66vZQQhqa/ff/3z
ld5N4HFEQ29TIDKqn7BGcUfLzmgWXVG/ft5wNKe3JpvB4h5jdIRH5JR9tCHCD1uodErJkw5vKVrJ
1l8IcxXu7GMYoEFq0wfkUx1cbDb7KrgtAbI18za2wiaCGFhuYVydREWrT9blQ/2sHay2YAJ2vuwW
bnTPxXcTYolNz5GDcOJemeXFlXZ354O18HbMCSOr5LlajoY3nxsBek6AP40OuOCbKWK5GZTriFRc
Jq7+d/jFKwOaP8wjx7ony3EHqJ+sEvV4ARnRDMJP+IO1ONGEnmtpzAv7LL051PfaO+w4wK4/YL4r
NDtqYmJFKryDUA2hSV4aWknl05XrNUmXObz2Cb5wT0Er242QFlLRf7ABpcAOFYfGBs9GBeJKfq5h
l8GIZKi/eXvkHYOBgXo/e8xt2GDODPQRkwf36/7IztFmsP5XDYgGexoUFwqsjsOTmhJd3Bd/pqaD
OnALBacJB8VKRcU4ZbHDz6jvHVpW+MMCmzyZnZjZqw6E4Hmb1seAYbBwuK6dG35hDQ+Jf+p4OHmQ
8Lk2xhtcbJKua7B9uUY2W3LnoTSDLmG0LQzMTiALyjvQumLaSp/fPxa/hwHOor/1VsHvHPsmXmjm
OOZBqilRW0rB27MTT15IKvgNwtk70WDsPtTRwe2bx2lTrgmb/uLxfQWnTrY8/M7WnA2Nv1AlxDHZ
k/DTVsCfPkAeo4VNBv0bHi/rctzhQBoRp4+OutOuc+bWHzbrEfoiyojaKSNzIQp7N+kSRuzJxV2/
L3AjKRlOaq3lhDiqjt2PUQJdk8AWq+aPkezZEyhT2Un2J+nuoyb3rKJA/OFdbcf5r4kZBWohc2zl
GBYWiV9GPk6cblme/U5TQtCCp4Vgwy8TI3WQ9ph2s6+fM2WZB47l9Gh07x0sPCO8fci/uX20b1p7
2HIBWT2w0fzY4DXk+FJ5d0heGcBqb/uin1k/CkRq8rxAUPcpE974SuJvQDtfcavKf1ncX+Yk8aTd
yicWt2fiWUhrNCH4sjkzasQuAWcmhf+eTm0sGoRLj2OwJYRCM3byl48oP0Cx5aplHQyAd+PY+v4E
wGR9ehmcekm3hRJc8uf1WyTwU+TxArvIp876j4dqVpWVkqR0uORvLJT33XVghjSucBq0txh0eOVB
ATMKJfFiq2r1nHPb2c1adhMirXjDZ/yATfr19uXFaLcIBuedPxO5VZG/+/wZSc46DehuAskwjTbz
l7/ZxfzLG1iTVvSeCZuGnNgJr8ERtaYEUJziUluVrsnLWmR1Mdo9LqC07z767zEycF/xtj21LqEO
mWyq5jz3dtg8bQoJ5N7pDBih7Di8rYYPupBhDNmnl23IwVhiYM5mKOwTKwQRXNUhrUx7y19yPM2W
FqbM+G7GVG9E8IIYFlBWjpo4+be7qjA9Dsm5m2FZQIzsXtolWojCokL9NMwBZoFqskXNwkYDq7GP
HirwHKNWINBObdCS3merEBJ0ueH5fUvSxkQywVLpjfRLiAgrF+sIKiHx6B6aDpyyvmkm05XEkYfD
TBFnOSrUOOdZhgC5qxDEao7Jjj1qscMRSXQDoalIHgBIo4cTb7x/ZmEha4OTwKvFbipn9aH/vtUB
sBznwdx7oUmzYEHV7CVWu8sJaBDMnXGNgf4858G4HIVokWLQ7/qCZbZaxNA2v7L6SLnQ9C+TgV/j
U1x3Him5rhd7LLskjWRGjjd+mmfdFTpcXbj1UwT5e7n8HKCwdl9tYB8P9AbE9UNO/QGRqAeHayGa
0WkTrPbt0M5qH9Pnn5sN8AVjU3N9mPltyb79cuaI3MKk0aWZYkM2wZdM68z+Ypi/SqiN2EdFPt5j
hUwKhkyq02+In8e+RIX+JycD8NzNoQesqz01EYM/Md1QF92Tt3UMQ7o9ctj/1Y001nJY/LEmIRgi
mFha3Gp3aHXpcJyhfA/3/Z64qnqMEexOJosatxVfOAXrGCk5eIifvjIwBSR7Wgf3AXA2CsAl2Jfj
qQsqUCErBdetm8R+S9Eu7+mXzVdhGEmCB8MCVjM3/IyBRiUpLL+kZjpsToxu5B3uU78Liht8llSl
fPXuGAgF1UemHxNQ05QylafcBnv1cIm504OE8ZFsddOfw1tWqzzDLrD5q+PqQwNiReJ/4nLF8vDn
70OyxPvSLU2uOV+MvgXBIwd9uKhrkwsWzWAaazYCyLkangK0+P897ELqMqyzFzbbxnx0AC1EUhSC
Ql/a0S8qVqA4ykKZgC8oZuZwNAne8LWDx3ew7uNIAcAN46pfTgmbAfbIankiwhXSKOznwL49WVZo
AFJubrG1sM4JeriOMahHQdZf4eX2fXGWRzCk9oJRfaRk6QCqiTnByUIeaRfp5nGcPBCpweinWl9R
8FerSerEYf+572v6kkSCZjF5p8noCdmLrVbgSrrdBX7RwxrVqn5ojumAGXyrBIjeBaU7+37Jr01E
W/7fmUL+JtyD8RiExrPpCdlWCLCdKDee24CDKNc29DftgCg5PyWgpGffFoNZ52HuaWHYnjG0PImp
a8D+2UmAO5BxlxuenRFbp3WKFm58+peU/ACoXgKmjRL39fl57Fp8h6bwy2LVdTqmyNmjG4sjBCfT
U77L5+zLxJd8ssyWeugtTDr4reQ2OYKFa47F9uXDflohKp4gOSZQTiqHD4a8Gdw+dscP3OFLsT+U
6edvxXT1V0853xHjpAVTc2xdfYiXUtg/5HwUI7WpLgBCsxifLYnK0vSpFHapsRfGEyXag8hO1wUe
0k7krjEA+x6T7pF1awhQ2u4/UlCmnQH8fQG6QO1IxHdhnzwzZdyuaA6NXfdPVQQFA8vwhLwMaETG
ZrezgJWpwmpXoOehz9fwiQfFYKBd1XSyGPWxF2rbD490XjbnfhjUbrmHwikdnWfM0eKvm+QfNupL
y7Ynv1xoumdE22peH+z6wWjq9ilTXjjkMx1D9717k3+Ft9z+iU66Tua0gyZO66W+6IqzkelrE9LO
2hW3C3uh/tlxvvSH0bCuAr3AkBUuHGFLM/EIEtySek0zYmpLJ7bhp8w42PohPit1MadCUsIgrsDP
XGwp88EoybUzHHNb/gf60zTULMweFTvJvy38+i/FMpoThAMPpz71vzHj7YoBoe5Ija3yuLU76kVV
AnV6gjQaD1Yn42xNDrZ/1jZ5r5ABIW73pdP5oNpRwh/uX0JqTfVQZyitN/LzUcAFGAEANFdCRNR5
YfcdvuJvlbTKzYSW5/1j45tWb1XVsAIlghFwdOpcT6P3KPVM4Jgfz+KxChUQ2HrpkVqEJjTXIPti
YA/9S5MnrOKRcF7M39BlZnXOUouchkRAQ4gb/CyQrBpjec22paSNXYrexxeNFbuB4iuC2YyP1IPt
+yPobHBBP6oDobmt77Ytl+aE98uYxaZqlq4gA835dnX8bNL1bjwf9XW12i1zu2gmol6madUPPp9h
9wR9/BjLRXoGM/o+N6lQ/cIKaOnVnHYEnGV4NRxN0Q7ttNf9btemUoyhsDlXmGB39+osjYhKXRHx
WBqoWKWqMsM0zCXwMPoaOzszkBsDPItkuqwuimF4POBWqJC+/BZZ9hc6gsRAGLHjNHWP77EzqKze
waE8lt6NsXO6/aPI+Y3BNIbJDvB7Z5ax2kBy9lpdXLdQX5X4OnFenZeh+ijxr9D5IruDB99IDW70
+GJAewT6WhaAF9G9SNvF9rSJJ2NxI9/5tONjnlupI2AGFQxHI22Z12KRms/IjYeRqP9kBmOU6S/C
7bAMjYE6wuGwkPlQcGHtpX7cUQzJcIzN/4rmsZVZs2470AX1tPbOAkJ33qv+vUF/s3Ccpzk2wfFV
4dwm8iZGzTZc0gVgJQh6Vz8HELi3hYV49Hstlms0I0BCCd4kAgRjdeJWKp31f2hSnhS6gDLnJJV6
QyJ4W/0pU4QfrosA0LdZihOORx8KOVIIGyWhgMDp1pJOWajIbM0Oei9kDNjiKYPQDydcFDLTuN1r
CqZh1lB1hR4gXcag8qlSmLWfxkYM1+z73eVpq5caHxC+yCa1ZoQZ9lSyUumFDzOxyJO82JFg3I8M
NSoZWGEy44x3YMmu10OWUSkZHNy6dwU/23GDII6VIBxupJh54qgq0fDQjeMKULSFNUaq6/il//tk
KCq2Z3ckbk6+UXbKAfDwwkCLyuKffb3bn34gNyh1mQD6DHONOTnsKORpwsG8ep2D4J0xttZtet7J
QJmPviq+lu1uFaQe1PGp0zRsetgQHCIQiSqqqsRVQnxH7WlJ252hJSqya1zwEWZsbuesBcam/W+W
bePORBt5wjirGZTgvCO3gNYfNgzQoRxvMSD1lr6bL2Q7Q9SLioPm2imydTNgtpPwgSkiZ/INNq0n
nW8DRjELIDYHsjdjLF2uMb0+PngnUTgrgoMtjJKFLKjXpegpvki/wImyR0OHmfL5l6gvz9eEeXm6
SptFe7F+j7ViE2FUxgZLUcjFh24GXtpMXcSq3/rGRHKLljwb+j3Wds0n4ukzfepiCQkNaL6/0aQ6
sc76JcisYDTlg0vk1Nwg/WSNgBZkhHGyGjBTKbk381HRgwfOjr0voGFBkfMdLJNvU5X6gcgfjVLc
1wCXEPLB//EamytLIeVPkP+FSKxICYsjy0rxXBTR85kFnRmRyD+DEWMEN3FWsHJbXE6McJcjFrjx
UOnxp7xUTvub0WxhNtAW3sGc4p0ijD+G7Ti95J8pSZG+e+NYvC/bpl5sUKjEcNJt9I/cdcCWLo9+
AFFmrm76C2lV5M+9YmIi5yHalTgDwHqPf6NXzxDfTunF1qwfdVrt1TMNWxG4yXdcWEEk++dZA5T0
A33iiM7FxZRE4MUgeNVqIKeGI7tlaucAvn3D1fsFPSj+pIfMOaY/sCjSWggoKQdT3LflLHh1CLys
DkqamSTXnaSmyBJrYI59HrywzDIBs+EUGd2MiDfr6epNn4lJqdkM4Nl0LO1Z9eqaux3LdXQyDlpl
8xIOUKZioN5AiD0Wd9mQ+EViOvuReOEOPbLVQzFnB51TmxyUItLhb/MMJjGXpXOC5GuVfj6rBt8L
GBd+bRhu5PFNxcFUetfwCKhc4S/C/xqlAcbnfRxuN9Afe2On7VB3+MBLz+CAQts3myOziMsN0Uht
U4GwFg2uhoDHo3LGHU7+UDFSnKZQdqbUdWhhb0yavuhouKCnTRCMGXChUJhjyOwi2hp8E0YbBtLB
Kgi5Z224yWlOdLgQv0kwCAe0KUEcryFpiXzeo+UN/xLGvjKp1dW0NGdmKn6Oh0XYga2bfNO9OfRb
YJe1GHph15eahMYpRJlxq5OXES4HXOTQ+PX6cR1sjLg+WYDrECSgs6hSTa6fxsnnGvFQcMmAu9fb
rkFUmX6jDrT8nbReKC/kROQM2ow1Yp4vuWWnHqxu+w6bePtwsU8qTnWZsgUWTxljtnqstUWfzctV
kgZiRncL6pgU+spDdW+++dlVy1XJbuQkHAx3f28PCKD7gM4rAiITIrf+z9IY/8FmtfH6+EGG+9PJ
xC0rSi/LYGPs7t3NSIKLeTfU83ZkJMV3o7nDmYXCcrGAtlBy4WRVEyvmbletizKeyTwgi0j2f6zL
rSx281CIj2KZB2T6uYCRH1p3kfLZzmFc0ToKFcvDKeJAHa6zyVRyeoKn9cRqh4DEEGzADxKqPDx6
YoSVNW4AKToVfcaNmZtWvKC53CvCDjzMG4d96VykoaZezoTZvudKoioy5wiVY8HA55GlKDw453ab
RJ52zEfqBDnv+UvxFc5j2ibKEcvSu3o17JcDEswQSuxQk2WD3hUe43W8DbGLD5hb+h8U+cfg1QbH
aLg46ka1pb4QMXoqQYws+tN6sZGl05tnd6yeoe2X9qA0yYUGlI/JdYpOMzX1DgRDfY/BLyYiFvwO
BQnD/Rb554m+tRDL1Oh3Jq2pE7l8P43bUGIsVwCPeNtis2jf7paf4DKGpUOdAXF26ox4qAOSceDU
FtYY7JOR0kPqC0rg8lMleG2LIY1Fi8Nn8v632Z/os5fTjZxg4c0VcikcRBjZX4AIzvfuaYklcWw3
0oYI/TQDIlGSML34Sg+FpwVB99lFBlzocL0tjmz4d2mChxaPnWI03zWKWcYJDXVbHXNsezFW91I6
5yxgh3+Pjd2lC+okgnxnltASgt6/V6A/41vLO3CLoYnVTVTLrPCqv5wntogHry4T8ga6E5V85Ww6
TZ1Qe8SSrWPV+6mpigNQOB85gnJWLG9ZQ5YH6WX71ukKkmEDNSF6uryInFaBQjPIrUwer3b+rBiI
Y78jjDDxutvg5NEgmOsW1t/u2jtEg3bCnfRm1/+epMwm95VJZa/i5Gq7JU0iLL69RixueOamzr6F
mhVt+RjJIofOfCRS0hdJ0PZxLiIEIp1rR4YEWd5fYZnj08R5BtF7r/RsWuufcRnTeyGHiotCk80z
4XHH3IoC9vaVtJSwQ0YpQy4Wzk3gyYXxXbirnUc65nghV/N0kFUdA3RtrYgB9+SK1vh8Fg34VXZa
m58EsHbqhQOMB+tGx8MRVtV7Q8v4IroxIAKwrZG/vqaTzEon99+zVbDko062Vho6LalViPnYgKhr
VV4OHc9AVXqKe5RiMhVx4Y20T22ESfadwKWqRhZUewJgzXz+EvIWHmIk5sVHAg5zjGisOPd9SiXl
AeEwNCuGvUS9wusd7t/9lEXvjns1s8JvL0YEAMkG+Aq3ARHBr97QanIZW+VLAUz+QyyNh/IQJTKW
k+BUu4JQIuV3e3eynfQjquE0xI5uBR+CV3ngHLXcRcSYPnJ//aRX8blmflwH2CjE4lDCaGJdbC3Y
Q1rcKx2PSfMQA6jTNYm6NRdoKKz684LW9Rzq3P38OTiU52DGLh1F4PJurIudIC0mVLn+R684/Okl
V3HSyQhSod/rtzDMwloeq+HHA668pH74HSrwtkfwUKzmpTwaWyqSJWYmcuYLaUNMcpCkOFvlC0mZ
oE30yr/RyiAJEd8JHtC0k7N8fFXR3vtl8/oQPhs73asEZPUH7cmM5Aw4Qz5tv+TsGl6ocoqaXLJL
QL53OHv77BqAWRcqXX/BYwBLnjzffAPhBGODrx6qbs7qLgimxxYTLcqGPhSCW6zOSu1mVTx7l6qx
XHL5kwSiY67S4qRRJfZYzImqlhpv6/ZO7kbVarWg6iTChIuz5wAM/cmmVnf1jxTdyKNbTjaL6CXZ
XDUodB59JPyxHpb7sFvzZh3823d1rlwTOKGF36gxXppVJiWWf8jflKyDyHGQCv0c8jtnj9Dm2MRR
0fgfTuchHWhhBgA3221+ecpyVcWMSAJu1MxztKkl0n+r3f7PHsIafCxusHhq4Gw2DXjatSubBZ8J
RZIj+X8B4kGkkMz6JdG8hz0aL2WPfcuPW8xP4m2De8doMl81SAYpTAvN7T2iVB0bQVsYcHTCb6Cr
eUC3mrjODFdzEI+QEpoFX2mjJcQDj10V5QohrVfB5siiUx8yHUnH8fWhn6We1RJdULYRe7Oz6Q+r
Cg7gMnNpaPe6aJFDIGEpKY/r6zLHGOVybm6S/GpD4CXOiC5aNxTfpQ49IkHzaXDfeShud+OR2OLK
uqkz0n3a+GgviUaejvbn8KzwLb1oxQaVw2/mLenlOWtBoxEkWdc4apGjtmOLdSBD2SqEZO+cbKGc
amsUMCzwrVIxnbXh+7BqEclWazzZUJOS81+hrj0/jyz4/U7Cd1h882k/z5VFteC15c+62QzzqdQk
LDpKkrUdyEcK7G6wfG8zE4d5i255OgK7X+cUF86AnxAGFoWFiWB8+VWoWRH6TOo+13rx0ECdLE0w
7y5rqzW45jtFKIZj7gUAATgQqdiwQy3t6ulSynDZdHKlCTuiCTCw7BYhrzxrSEWsw9vNkhfQ+xVo
C1fmkXB6c2xlGOOwBaXu1KyTBH5PoqPS4vOgDB2z1+LOzT2p4x+7ztN7VG6GLPaavqM1kJBWfKWy
xmodmdiSx1ksu4ZZI9g1g2noRzvuI/hPNgRC0Bbe6Pz+Pyf0EwVQ1ozBSjqivcccHwa5u3hCxwhl
hbmze0izIW97H5TKsCyDKIVUWyWWL95UxVbivmsQ/I3Ia/Qy/dlzsGrbHFMKiUmug43bJx4dXbD8
q/TVuaTY+Fx1L6suqLoV4fmS4Egrveqsoq9gfPHgRmpPLkNEWCO9tinX2y157yPoase1PjRMg7jB
gju6gmzSzp+DaF4sn+IFyCUferzd3Kgb7vq5WHZy7CXai/3r2X8J7RaxBJdc8nCAS5R1bz6NPoiT
ZLqLAMSDN64OMCBalGymobqduj0POA0CgqRa5YPw2zbTU3/YYEob1DRpHedGnV5vUiQspmKHLpbN
VlfI5i414rHWm0h6HpGVi1wv622EnbkERtNUsr3zQGudu4NnHVt8mNqOC99TcphjA/KNaY9BdBXI
fOMZIagnP2cpSg9e8LdBdEFfkvJNgapD8cLQvvnMGWeSBrNQ3/Qjn2NC8MvAIQl8gfC7FA64vzu+
bF1Izw5OJELhHtCk4lkGLlfpKw10jCh4DYDsbYgoXeL0Gf0wxQ9XnaSBOPEX6cMR29KkzkeParlt
pQkkzM9gDrzoNpA24zDU7S9zHpOvKUkIxDHghqdIZASBRF4BviiGmOIqKBNFGdEG2KKXUpIqgzRs
cY7IY27Ix7T71TylVQI8FtnUgPGxSG9fHWbXy2Hv9maQwl0OAp7Y0fZ1FA8i9dbFM2P3XP6vpb2L
+3+9d7v2YAmNjdJie1Xcq5SHQ1sZVSQmM3YUM0dVBoiuXVWnoiDfefB2iWiop+DiBSCVNObrNaFO
ukYioMNh98EYh1tWTLA7tlcBh3NXekugn2RpLY3iV4QGj/VmsEYBCVDqoPSQ5LASF8qkjEu6S5+n
IHGZTsBt6fzG2Sm1WjV6XecOCaak2Hk8KwYkTQrAX1mnYRyxe7uJQc+uvIPz7P8kt/ARIzINk2hG
rWwZEWQWuRFO1gi6bHoE6GyFkMKkczDl7kRWV87S/2BsJPBp7Wu1x5rVPagyEjO2GNJ1MqoOe5jW
ZJfcYa8xir7ZOQn3LcycJCzee3mv8sMKErSd7suSMnZ0zo6/x5oMo7UIe8JJ+pVRfDbJoYXTOI9t
Cq4YP6oILAQfAoXmM60uaPqCu+hxCAJ0pCsa9KtitNSxAsrAHhSdXeZK0loY209FCCdN56H+cJeN
YzP6pulk5ncyBliBXkXYtkrgwjT+0glDimidKy/FZfUoAeb5LybGOOmKzEFYvzkdR+W3U/td/sji
MWyISV5x7ymWSTbfAhe+qoy0LmxpuGCGYpPapKoEkj81LAiLEEkb7g4R9OWEVuZ/XXvU0D0eaqW1
C7nwOdVzaWO/3JKTlUgZyqXMGRtfed12pqNsWg9btREswEU7suAZle8DWBrS7ilsldwDsY6nhCrP
qo4zDJzLwrGrBo+zFxPFf6O8QAcH/MOzgBAiBr0cT0gZiwMWHxIIs9eJPdHjQ3v+oS7k1CU8bG2q
GiEqygDybR/Y02+eWkaOS8HjaZc1uNe7DcxS399q8Lmq9MFLYKA/3X+dV62KmA7sC3SNDYb6EhSd
a8SgfB9P06HJPNsLuNQwZmjMFpbHNlhfh8BuW0P4Y5YYgHSzqpAAwY/+W0pTWMp7bvpl+yyHRqF9
3kga7NVh6RNK3hAgnVoQT2Hcjp5+6SZDEI2wr/ac3nBoMSoQGr6I5EI3q6/m+3Yvz+W8OHnZrzj2
AgxASleneNpgEuVf2aKZWvF+uOa3VIgBQhTS4Jet3nDsoyGehVaEFgPE6JuovifgKACZ7ubqY70Z
Nsto6smeK7f8DEliY9ne3ssyp2BSW/liFsGogDFhsZ2g4HKx3vVHHtF23/Ed4QIFwGUtw4e1Kvy7
uJri/1by8WdfBd5UTxYXU1tXgLrtNzAKpZL3jmVBoGieN56CNDNa/12ostGGkqszYVPv9yCJWUBk
20w77FuRpWVQqOt75It15V37st5zngInJp5YzpB2uPNRPuH/1V4FRatN2xa6F/nHsBivjDfIuGYu
15PejLneQtA57TdyoW4fc7+SPp9BvlqjLspdPe+ZJWK52Qe0SBYwL0BPTVqpsXaoQUCja9ynZsL9
YtnkX4WjxuRKKnH/JvgTh/DcgyyJjS0HSb4aS2Hps6UY7qQv8amLzilwRAKBFySIiyS9NR1wXbS/
0F3Ie4S86ZMxt0t1tFF+TBJAJVCjEbRKiugv1o/lMzo21bACS0nJaiaOOKBJa/RKtAz/cbic35sG
ETqfi6iPQoYg4eXgNamGPGldbHFnCjt+m/HVIbSgP5C6I5EWHkPo9dYxgzJp3Z+1DX1CugTG0mQ/
t1kuhpWmEBRDYHFR7qCfUtJtryCIU3vhAdN0nSlYPrh32rqFsYwoNJ5521VDP0gESGY9g9CAfQme
A9cb7+rKqrfk1+HbnW8bzfx7deaoRS9blM3cZ1UBEH+Et6VHlWZoRI/H9mnBf5hDjsrjnWC9G8W5
4Qy8mMRt1eQiRip/qEt+ufVZVwsfIWkdcrBRHXtQ4zS0ciejZHVbfhIY+b5U73DItNBQG9f5C+rv
9DP4QcmZlb42YxW6bTWsTco7CSp1toePlpjzjP3iAACyB5P6zei1OyLeUopxGLVxpw7aZcCN7HSp
eXF5QxzBjPK1FWD7q3HopxyC1m5ILAnYz0bgk0cei50821BBZk9LguSX6S6yXlaAwMbSe4hexzm/
kBQKvbVDuGj8H9+wJNVOitbA7ee6pMU7Z+3zOrYdf4DtY9kl3QNadlFf7XxoHPvVoI7nSOxHkd6i
2oGXjkeVwh995r6MgZHLwvuaSMIlNXCvILK+bCu0ICtQqaqSOOlZEqgvTq/DXrMnUVQ+d9XH1ATL
n87j1pEUC9ZmZN0bYfld7mjN01HKCIbGAwe5XBls/PRRT6X+uR1Lkz47RC4pAjZMHXaONaAzPQzh
HIJi+czcpp9Xj3KCDjc/59jwBji9wTgoyA7QrekSRWpusBgyJmNccnKubBdKIjn1T9xgdTbuCZe/
U4pqeBSN2zPdiq24Ft7PvJCk9Q2wIxQPRdP1awY/GI4Oabakt5ezLCGMBtB7uV9EWKD16SRLS6GR
Vj3cOEk5IgzJpl90x3ksV86x4f42Gikedy8NX7/J2BhdsmKjr5qyMQbl10DxUbbon3U6MRNYFkWL
fenfq1q9+qAkEnRuOuswEigWGKLEru+uCuRFYU9A65HcYaZjrkeBLqJpOgrl1QpOIL3qzZbG715z
OTvhyF0pWtQbmHo00LmREwxaNQVEs18DNiDDSz+itdgb3e7Aoj9yUHbfJbI4LOPN7FXdIqzruAcd
953MOefyaAyYMCg4ZbK25i54gdvJHBpvQCqFsxq/DENtKQABeAdRE8Tutnu6mB5R+qBqmvxyIXNz
/PlPDZLXCOd5nsgsRA0hxGYNX1Y2bVuFiHLyJEEoSTVB7Z9DBiJJheVdDGON2bmsP9IsY5yao9ru
Lj9TecQYEQMA2kLVGxI//hayj1NWV59xydKwSAyWmKJEJvWiP9KO6AEJTFTvR3AwWAMHA+598XXQ
HVCYwYvtdOYiqLoAw/FWqnJ8n59hmDx1Cy6Sct32lASpEpJJIbXhcXeRfAxte4LXFd0gl7EPHa0y
+RYlmY7/3xbYSlxvAtCMWIxv0zC2YMjpT+SQ45FHeuambX4VG8WKeZcU50crravocd1s7oGS8jHG
dPsbQ2fi06jo9rwa3mWBgBc8cWVyMLkC17G8Fo3hJzkIL041Z3s3L/Ai1RvljZrUmZ0A4woselJO
5F4IMUqRRz+blL1xo3OhsBFW/WyDh5ZGF9yBH8Luli4vpaMXyu+ANSxHSbHrQePwkbmB7Sf6mZMb
m8mfzmGZYS5CxIqUdCNjjBwV2T9iQ//S/LfScvjAlYake/d5uT7JBQVgoE/bkCCjfXoqmDgL+msO
7ID1WKuGWQisa13IZASRqlakIAtCP/iqOvdv5w4tQD4bxpWz2h6grEfIW3RCX9X9FXfgo3hQSHVY
I+RZVlgBuFkBG3oV+yDdrIs25ciHjAZ+6bwx+apLs6/whuzAOABOCLCaKmf55jNuwZ4/B3LumrtS
uBqJy6eFHfi4AzzuGdzqOoJ1qSscEFcVKG6JRtGsWmWpL0Chy24eLL4/akSz1YRR5T4Y3cGAeMS6
OcXdrkjIBDbkiMBXH7Lzqu/CGoBhzigQ38/J88jug25F+ChBmPE5HZ557+2xrYz0CiVrS9i43wav
4byYJt3BEQ9L/gyxaHC7wpYfGNMrw+HXXeh1t8UTxENRfMz3d6aWjUVu/zKdCC/bsF2hcmm0m8DB
gjyTJXsRmm38VnrTrGfP2YbKxLw1W29z7iHNq/FQPwRNXWTB2xzgtEgaxufkNIPwUkUXrc8olpvr
QAGl+klpUP1PTvNAALlCk41UA3NylFFqip10AwS0F6d0P8OHm0Q6BD7eIgqcKfge4LEMmpmewTba
IKaeVdQLRzdKXjdEf3rmjmRw9mju8RbeCvltup8tfv9CI1/uAt2v4ZKhxkNMpwiRpKe1TrSlkkl3
1KiPsRGXhnV7WTbxU4ZUDMLaxZ1sx5PeFe3DbNzOyBrayvXjUk3+fMcM1/DvxZv/izV1OA5cUD0D
lD28Sx8/WbVgwrJcpNk3CE3jLzqY4Ro3rDNHfdtT34Xkh5vfFBOZrqIU6mraUg+JULrng94neQZv
ZWkxbGrRNGolrXPonBfQvc4vrLgVQ4nJbg+N9Zd5uljOrE5Nd1rkqgaSJFR3gyBMnIIJ3AL+GDEO
munrFzxwqzbGCrTlYJyBTWvvE/X7fYRwcnOIwCTv5Tahcf/F5NVE4jk9WIgFdFjqdQQd9vqNBuDK
18Xl617jSFQLcAm3zyBmq70ItTepZzTHr26+hqoFZqhdnC8SGESdqP5BiJ+kDg7UhWM8A67M2EYm
3u5sssKHtKuMRVstMxUhXPmbv3BLoY5q3tKaWvYXIrQYl5Mc2Ll9xs9ubUL+/2DaMDf66FNAAWdX
/Ub2WKAZCyLlEQzZ09mxSYYHF97AsKHVU122xRmWGqEF620MmCUWL+oMdD2YuqUcLqYaNhcw8Mab
mQGniTDLAGj0MI5vPX2DnM4BlQRcKSV8CcJoXs+MToJxosp+LDW0cFxkL8d0+kuS+LTyAImGyVAG
r2qdl4GBTiSRyQ/3HtC2sp/+BU/y8WSKNxI0A/o/UUHajQv+3isfmAZpkhEi1nww/312QPZ53eVk
PW3ddg3zYleEEemqJYGS7rk+9aIaM03LU4rCBKFuPx8XifLyX5U5pCJGNeBdc+n6Nk+YyaTtypvl
EspQxqWm3cHJyIkYkCdTEU/T1vR/1TToeYdY5tULD1DKgmzm5qX9aLF7Lc2QQCUlqpIwjUDzCeI1
IU+HV/nVSFGmH022eZj9R+twBqvijvQHUOSsYn7f4q/QAd57DaL2bLCFw3I7TyeF7fKD4wAD08XB
cZRWKeqOfu0jHDmQIikvEGR3UDx5WDHRChzdIqE6uqaoL7WvK8yiBDNfs+4mFlHGKo8MWHYrSnhz
1Z0Ob8ZfbZfMxdyARGSDAYUv96H7u4zh6meOYygGTUyOmxy9ci4AtlU1Kn14JjmxSc+P0RWt1ZIM
LeSbgnoxVSGwuyJsmDzk4V+ZkH4NrMdhUq4zB8dDWIjg0aQ0x4RSYcOovh/O+sspgfKX8HVLkV1p
Ylei2WP8NqdxIiMh1mhJPsvudyj1OZL04+5Xt9hBbqzORdHtbWONyDG5ACx1rQnCIW9yAuDYAN7f
07FylAdf48Nxm3rE3qLsj6nQZz657nfVU2lkHSs5Bwscs6/aZBqaXo3jZ7kOKrdGka6aXM3t2AD7
Rdt1bNl+2gP/PiYSrGcm3VqsVU1t2D07ZpRC5ljnBKLUbtmRLA0Wm4Cl8B53TYfaGFs2Rbu8t/GS
80IDwZUGuggy1iTXL8qQF7KfLnJGU2BqAC2KH+kIW+uF2VIaiVRYcg8jvcU3WoxY+fEJqQCv2avz
8VGt2uJV07wadStl3Qr8bmuDONPCpfM2JPcEwNJZ17S9Kipo9zZolTD83rK0jtcYWdo03TPfeeMk
C65pdjSdNe38BBALjcHBcH+fzgxZi2cKB1SrwQRDyn37gIQM4Evr8fEgNKCbz1FgrjYSO7PIkn+e
Y5PyPWo7+i4dDZ9DbzoXSf1u1B9uxv7WLW8SkwNetIY+B2Pe4lb4+QFwNH37J+d91odjygzK9jOz
WAbq1ND2vyNGxUulf08OaDhBk4CBueECDkVnzMVGko+IedCHkmPN1sAUH9tNTjITeREt8sRgjO+C
QZgC48O4OmlG3UX5ANjTf04Fvf9wDIclpjAWkhEV/l//INhgMttdRANEX1e1M6FSrxtRWJsaCgXG
bcEso2uqB4SSyRE0Z6/yUsbPhjU62Pf0AOKAEh/1+9gwahXvQ8+wxRAlx5e9sZF+T2smOtFlMnld
YybEh0b2IZNUrRBe6N8OaqRtPBJ8tdao9OOaE7xf0fV69OYYFMls2y8hSfJnuvS5v8tusD72C0J+
j3JaSLwjMrngy0aRMdiixdtDgu74p+Nfe8EOl2o01z0iayqE5S1+IV2J2F/rVipWZYjoszbpfsNf
hDmXFw/unzYh8GOD6OLWwKSW+MOmaXvP+O0fzy+WAjsXYHN3Bg8sihxyIwRWRhpRLM9HZyIchGDV
YlFtFrc5V+gGq0QrNH3qMqbN+nu2VMkK9W73JyvVCWU9DRLQ/ocwbRwrKOwNRqhllQ8p7h3B3a68
kE0ibtjw7Jnh2qNrceRVr8rhPfr05taB080yVPvPRED0kpEv5PLPePV/3LK0OR2U+sO77kazuWfw
Y5HwhhFVHaxJFcp5MIA0k8gfJ69iQdWdCv2mqsFK1GJn5V0ha7h13Qo998DwdzfXNqQlJdGaUha7
1TXO8OFc6XFUU5wB+2pD/VHOktWFMJFDoYhypOpLqbwJ0DHEgXSE2HX2IKGXQ/phO1u0HRHMo08S
VgB2320kwXmv4KvBXcDy0uWs9ElzeK+qJ+0PvWLvvp57x19fW8M34k5C0mJjw9vlZ/78lr0VdbR6
Ph9pJO2ffNNpAlViHKFxDyMY02wqm6tRkNCdNj65V1w0rYK7S1j2SBEK3DfcSsJnaA+HgoO/Wwz5
knxrllRCv0aI+duRHWfkQdoGQ1Y42yupH9zKI6KiJ5y1i2ThN+Yed4xdWQ4KBW/yev10Kp8OSXh9
m0jyQ0ApeHmZTSoMbRzJg48O/wDDFga4HtIyDM+HvEwJyS3v7P3Ir2UzStC6GYrQK6l/VlJMeXYR
WP9UxLL5EgPhfijiY8Ln4fqLmUFj/jS8IWqvuwZHi3NnD/NqB3nrv04snTTM0/PIoCrGgrXC5c4E
LM7Vz2uHK4ACBr3OeO2Ax8bZR2ztbdeEM8s2As2ptwPulR5tDz+jvcKUniiriP3g4+jHW+trEOwX
Qlc4dBdHX115AObzQ3Bmwj9eGAumeoQYQoSLs7jzpCmMg4OHFZDzn8xtnmj71+pM/NOoNPGiXz/K
etkviCZqZ3bKAWvdbrx0k2gXCDqvUsK7TTM6RZByW67bzmiQ7f1ekMWX2XdKHWeAyEWtURRy56Ak
GDu2mzKECnmmbKgQ7HFl2b/aDwPa9HFwQal292E4KmiLBMLJVOr/ooWwbcNTVgC3kZn22JNXp9lL
kfsdRG5+PL5B/rAsatXGwCeXcdGPu4+uCNeAGvP6ZhKu0uqt11CFrDii0JN6KSi6La3fLrv1CFA1
5PGn5JRWBQKS9QIeWLEWqjuIGZyFs7g6vnfZ2Kb/hkolWYbLDzOGRLLknEe5uRybfO8UowzKAuW6
xCZAJ8HtBoXSiCKvy1t23ZPOROiuqsyl4lQCxUKMK7DvUFyj2ihNS2XWOAmC+YlnfsbVQPjdN9Vc
O9IJeCEOQlT/Hlu/zhW5f+eY/W8hALOt9e0/nzjLokac2Nq+/XWLskRFZWsK/wUMz+n0jr8enR0f
jZTN0vm0xUttZxdy6VtkcUiMM1rHU+qhQF5ygkGHfGWhhw8zzD5e65C+0Nr8HaUJ2rixIP2/FOB1
gtxDDTwSy0Jwtr/vj6nhYq2Xtg5Horh7pp/lmY3gY7SHNXARPK+xFBF8tQj6Lo0GRLzjxvUIDL+g
t+LCIa+ECN561agcgHtFGk4hf46R6dxl2ci84TiQZU43mI2CgzR7Pffv7q6C/VeIN4W1CWESdBe1
o7vF/pvFkVzFMbpjGmcC2/buaNfgb1Hfn8OvM67sjGrYbFBoNE5Ho1fVtCjxrYOMKjGgIA7qEH3r
d/zxyrkWnZWL18zbsJZPu1zV4mTKCGGIr0M+Kwld6baoqPdZI2SRPvl5pzjBelm360kyjt8U+9Gz
Hf12ZLVkofyuEN5o8tWx1ILC9rATWC42cOjYmOZdlTHBj0dHLXw4Tf1hT6WimK00OhICZyi5P3k7
dUsgDZYFpcj/xqwQXeD6B19mygEypXwn1jLg4qZnKY/c+iVtJSOsCP0+dMYIiHK/4ChHFdBNtmz3
f6dtKlbjAicnPqGm08PEH3eJ4OSVkROe8bpEx+Z2AGC1VxqPE+4w+Lz1pqHjr28BhMVwDI91GdVr
TCAVKWcN1CitG240lEPc8TDzq2IhAkrU6HH3tOEGQxUHhA5Fm8gefeNT4jj7DvgIWv4if0G5qadF
6xWIHtndWqH9z1Km3p2+wHNiM59EBkZx9tZzvoOb9FbCpdWD7zgdOAjm5aaQ8qFeF3PCg9kWpVnC
HQmf2Pd+VZqbtYA+kvgDKh0cEb87ghFjnBYEv1sHGMC56nzV3dLJdZCCdDQkCeE57OmXLqMjfg3H
aoUPy2NCEnCIgj+NbsSgWOZ9seq71uKeAda3VNf20yl3ax3zQ88+N7Vw1VY4BlDoRR9l0Rc4/HKi
qh/HOiTa8+5/kqok76ms9y8tY5SZ5/C4o6EzCQotR7ecb3pta31AfKmZGmB9bAZ0LOgZa1CUYFKE
MoUueb7wok0ngTMVEDkvoJzqP+OiWvsWgMQB3EDVvla2TiZltSZomzIOpyWBSkyOcvdOowc93WU/
LFR0N7+gJPzwzivrIHEBQPQsy7dg3ti2pS18E8MMXOhfawdiwU3SL7ketWqpfRyYi+m1jhl70bGD
PTiw9VOXqyBJWm3dIGs42ZmSazlf1NONo8yOuNHt4oGs8rP/ru7mDDmgGnuliDAaGf5eCGctN7zU
tG6Fk8tZRTUMjJS379Du5JPwWpSeJMXGdhdAtRd1i2YFEIkYtgYjN3ypXT5UFIsjEvkiaryRjaAx
dOtGlyUkAXSRSay4XjuGF49NCBsSAxXFuUHXqHMxG3KLNUw88mEoHeWD/+Q+fjGsljNQ6cUOxkUE
Pf5eGXb8a2pZtdK9a5Q+8L8GUqCI7jAsSU3zAZzI26IM5nBd+4Z9E+YP6HU1LzFKMi/Hz7Mg4rYP
IrurSuLwOORSgKJkPlEFefOz0sTvD6B16dCOerAuxq0ANgQJSQIeWqlU8Cdxesz9U6N9lqmiFc7Q
P73cJCfESF59bGc3s+qtRBJG3/LZSGdBhSZsOGp9q684N03HT6+vywk0A+SJ1Ae9LHcOq8GmUgHm
znok94giZY8bkDwTeVK95mioJxjQmzwlIQ/aO79duZoxlLQol/7i2pnTJCoinz5GwLNV7a8pphWh
HcZNtTyXf5mY4EZ27Vh9Cr4FmedwxKoMS8i0QP9wb4vUA1vPjduiRTtgUewvJfuBHRrugv8P7o2E
1IGNOwmKENrSg6VwDYu9kWIeqdznhKaX5ccUxY4C6SQ5TgUrrPwzOCCvGv0YN+YbUKi0FQNpqLco
5MtPkf/JmjpIBsVYSCvdy30TK+x8u4kJvW7VGYvtoNwOdVZ+yXHlUKolAEkTJwAaEoqPXWwcASMm
uB1dLVQ5C8pJUzgyjAjz/lAjtvWvgHLkAX0ao0l00sT8u5ws8FctMoQu6c+789XeBaNvw54OETik
Vs7Vqy+KDQSiVni76c4tlRz7R7ksaKGhP7H922PiZYKD0lQ3++dXgZBKn9SbrF6q1ReomS9VF8xH
GU6sPad2Lho3ug5BB8EGMrWouwQ91UC+H/VSGH/ze5YagXrBXDljDhMuTYX9W7EqTW5f7vhGQt5j
8NdLGFb0HA6ro8Kn92sWyFINFJnXGlEJ71xJSV5Nbiug7cH4vRP22qoVEZ5AEZ6go4y9DCh8wzVS
HaOocSsJtRPyWB+LLbECliG+sOZuTBhUSVggMNZz5/lLRpVVeXKSNRwisSum4g30WlveAJ1oxbiW
WwFXcujPRXLfiEUlFKh+MNwpjVzbC4/QxXhJj+vaqngFJJKFkqnU46Wim3HtJDjND9WY9Atq1JJo
yaNOKfbnJXubYomZhuT/FhQ1Xqd7hQo1Rw8RfG9QbrmPEn//kBr8YJvps9UsVvrioLVK+c09Zao9
iCbQ5qPqF0RRldwJrEtb/fW2KDc6uoORqDF6N7fdNFc6DiFYg0o02JDIqwkyT1f5Bf3tFv2U07I4
S6GQjOv5Y1rKNaG+N4xTWeVB4oaGfgrMolIabcLzOyK37l9r81xeOOTYp8GyY9DFy41VNsgDayMv
UxXTD++DT+G+9jTg2jeXbJpTbZXUGLzh/XurcAJ5EfhERgxpvLa5xxOv1P1Io0yEOuR55lhejQfW
+UpgBKsFtZbFM7LfhFLHyjdjt2eViXcIv2ce4jcqYikbqDgWlgvLoHXxnZ5+nfvDmxVh1bqHGWl4
uQSaGdJiZG1QKHxV/V5IsiV4JO71ta3/lRQQA1bpVUsmbYQ4OxanmPbfFXdVMRSYC1wiUxf5iOfp
080lXjTcoKmwOmUOz0r0+6EuXgp8IhSVI9x4NR4AmXQsv3/pVS/lP2jFqP47p5gNbQiii3GHtnsy
oUxDZcYSPXEU555+xfw/HXt7vibbEmWqJBe/7nRvCuK2ZMfIlhi3Yx3UqdulK9SDivuAuAfOLcoh
gqqto1YPLGFbniQ0ZXjaMb2M1O20+nDdHzewiTJ1sG0KcB/DkUxL9OZU38eM5X+ZEk48YOD7Np3E
deGXZcwTiUJgrjxJsH3PYqNXQzFkj+cAAMC9aNXw9q7YJ4sOqVLxqBan0U5aKtSd45DnCFt4KDpO
pwvpZPifrabxRraDtO6gxKaM7LOMB8f7rvq+OVjtIA2ZQPE4rSvIFchTN8+scUi6ubJ2OjLgac9A
/Hk5wGu27X8ZwDnijgnwkzjG87eh48csvPYKtIcGgh78CG43bx1Isv5++TLu1I6I7N7ca4x1peDK
S0U/zgBJIyG02QClliDRWu2O67z/pN5Xvj7+j5jYBlJrKEE4/j7wPHIM23o841kIobx2SbM+v1od
wr7KefuXDIOZlgyLbTVR0R7zpEik61AG8Hv0/wfVfWCyS+zSYerpSN9KuYRwMorauZy4/fl+VUHI
2do4tQww5nReaCW/lCHoudPWu662plLD22ykNwtyr4YxVlmcDPNx+M0cqej2vnDSBN2XuZuCR2NH
jkBu5SbqQvAouydnEKoVnC8EfIzJVR7Fec7bymu0MGTGZqnKe2l80ocI5zyqBrPtEVdN5ezvvy1G
l7jQ38DE9y1NPs0pL+myy+fNsz/FQiAma/34i9JtrmlNZxW3/0L2zGjQRfJBHdq0V7ejMjWxJkPP
HRFh0QWc9Yfordnuoa3PIzIbK30sGE2jWxLn9VBafmc/BuyD8aoR1IdUf3zowz3uNwUxPIGMtU+c
7sz24vMOFcJViTp1S9WTBcvrPUbUSVaGD+2FDJKZXywNe39i+UgCBlgWWZHkQumMiFVjUmAPtjd5
V4Wwy4kFp3CudZhr+BEBpbORz1Gdcee2xtfaOQpdbdyRf3L/vGq9Lmq6Ta8wVQYo8yPEB5Y4WJAG
R+z1HkP4nFLIwm8SuBtdzK1T3Jsqj7KuZ3DEyzRTgOPJiivzA4EZiPsu7VS5UW26ewB8qYfqWfB+
HLCyh/4Gn8SPYB444Z1XaEqixavv362cWvstZf2xZlg4Y9gAmGUzNEH8TSeuIl92j966F46LcULP
6kfI2mMAmzALoy7hALx0HWTm8i38smb1uPjBp66lJyuLyrQSc1hWFnbHdowFFvdKP2xksvW8FsuO
f97/CxA2XGb1pQbz49/N7ADChsHbxBZamQMu8vJ6XuPo8w3S8rDRXF895wjeKg88hT2xZrq65HyX
dxsyM3oTTKZ4Cwc3T/wIKBmyIG3Cn+p3o0n95gfIcMOrm1QrXhGXXNURst2QnOwveBs94k8QMdNi
OjnZQWvKCMGNjNMhJeoNn6t8MYb/5ELKMR1db2ezB37Let8xqVKiA3k9TamFh7SW+Di3jqFrdu5F
x7yeygErF2i6+nWkFHaUuK2K4AXhh2NZXSHDEu+GOmKACKUDAyj6bIrVo4JCl6rn4LY4T6x4na6y
hTWuOMdXz5a7ESKfjbJP31XcEVxS2+caqRhm5ep0QHyDthU/6qtleqZgl2MJh4TdVA9DqAii32BM
J9syZQRrfH6PPa/KlNP52sqvGbNUJ1Nw2nFU+bc3ebAvhUFj8F/D+5Z8ECvWVvcoi0ZOIi/maYdS
G5cyk/V+XByD8CcU+pCjvEAF4j4C3IUp7LeG/bbo4uJuQgcwazDyhhF1ns9lTuFTSJxbOfDrnY8O
USGMMLkHXPCYIS7f8EzKkrhMyFTX5s/28el1I4BUAxwr9t0swIiDCmtaEJjmOM5COWYHegs3QcCv
97p3gJsL6iejLzfVdX3+C/vPiEdcr3yBRhFrzs9S6KogTPSMETL5RtRowE4QQ83kAHUoeD50/6YN
3xNj6x9aKED7KgjmqhB126kFcL7Rl6pQ54gSm0dPkfPsbhcAYTNFgmeaoMYzAtwTKmQ56qMMcU+S
QelPdlODcPstYzkR9oPSD0PhcZfLehxAMR7/w7s4GHjozcC3zkbqDapX8PYx8UCKj9lr1cm78UqO
925rcB+gFHKJL2BYUHMFC/ssf8Cm0486/67FQ83kZdNWIB9bt1LIsPLfoDDl0mk6W6dyp25L4So5
EPnnmjmqmLI3VWfcAiSoeGYQdz7P8hxbvwZUeLC/d++hXdlPKO6sWdHDmQJPe/tz2OQ1QBKYOIIt
eT1jF7riol4CdPPF+YZ3oP8t5mgsyMTJdLZjHP3D8ofY2fyxwqfdyUuTsAX+mHIxI8kXHny93uqp
pKKVl40LemBOitwTew4a00S8eG82c5UuI83KcFwS5KaQ9ppR/Ptzp75E2dRB4XTeR2IIqM2RvnOr
4M03+aTY6hOXcqqwNXoWWj1n09jTai6iah1dK7amV+xM+DyfzwPGr4n45ntt0b4KjASCeMEIv7pp
FqXfGj9VN2GrIfktMZ2zrYTemxl7vFl19JpMrWSB+/Wyb197TilKzbZy4BI7f3lCXvt0cbZ92HFQ
9EcjqX5U46XvbXQK51UgzsJdYPKENlEjYrU/3w92cht0rV5TKKyRhnwHMfCj48q2vASObVEHpKT8
gqZVaXk2fNg8TXAPpdpNCK2+Pv7gOn6l8UkbffFeqSrbZ4BAJse8/yOYJie7vFM8Qwjl6hNtRFqY
C5DsTK6Xjc2Ls18/ufHbLJ2LuhS3cP3zP05yYvOCv+5VnEUfbkEKgLj92bwjvAhFPCFW3LbcEnnW
pgCXW+XKxBi37zaiG4+1fKfYza6vSKzX7uWXk5KaDQtQJDNg1aaWwztR0ixQTwCTIz/CNzL9M88A
iDsa3SZ7t1StU7Wj7uBxZVcmorBHAKS5sq8nwxnyK6hsRI4Y+awuwmEUvig4PokGfDYjyu2N2tnd
l5cZ6R29ycaVUzTh7WjkyPj8KVmAgKNZCCmAJAMsxf/1sgzglKdP1VSZuw0gRoVY6170jzoUjDND
T3LWx2RquDDGIfVZPcU3DjWH0kGXQyp3/qzsgDlXnU4HHQC5ke3D9Ed2hRJ6Xc5XtxsUGAMnaNqi
Htg5aqolhVY64Q3YfVjuI+lDT+7YwDcqnk+pIVGDU9mUFW3jVoOOody1S9GvN/r3Jm7QbYzGSIR1
6bbb9r1MLm1iE9VWI0ZXYllJM8//7a21PtmbHPF7HUfMED1opSvUHdqYIXq/R8hIm6JYF84CbfXP
2n0Q+vwg0xJPTbMp2gMEGTl79kzFDLGTUZfHhiTSLs2ekRLH9dw8BHYH4xS/FRys2mrIJtELVUGj
l/UtS3+9vUH0ZbfoY1UTH5PE36vLiHSKJtNtPKdPgYj6yF0R8CYRV8sXwMQBpXYwZzgwsn+dCQRT
ke/SXUSsjntJya/Phfj5dKl/4gXnDhEC9CCxU3WGs2x2Qxuggv5s9qx2/OdseRiF2aP6qn3ew6ne
dDefXWI1AT+9N5Yn0dpIsec6qtsJCHoeOMG8RysVnYsrWKTDbaTBSjvk5loAKkStdJxwvVwYxJzw
rKEzfPOaIkfZdpN8z/ybUSeXzJhuYrTLCVm9OZir1H2gH1Adnh88bCcnrQcC65V6AxhqAqj7Fmzr
7cnwplnLnH68+utGtg87d67120MVG1lujM17BkzA+v067bbQIp3flZaD7NDRqFFwjEW/yMep2e53
Vlfk3c1lntLoDHNrOI1lKlR+5jj2lvt/CyrIcrA6moZIo8eLpLmKK8CTjqFObT6eX+l+ePcLla2c
yVLB7NPdwmSO8OEcOSRkHev/89sIB2CNob8Nm5j+/cy4Gc0J7X6qF2R/oml9x3rPDTyGyr1ORr3G
Rc7uY5v7RFK5CFxsUpa9TjF7fUCmOWyzcHYzmWFiBkcyjQO7DnbhnlgTpSjDCYP61fXCpijAT3tY
xpn+KMkw9VWZrlVN88MU5DC2+xYv6Caz9fbDnLGw2MEuph/mp5wml0KLJ1zT1vm9sf2m5uuNXw9T
3DLIu4APNoKubJ9FQE6g0B1xCk9UIwDMkWdH3+7fCCzb9qKLBYcRITAXG3QKhL5eGRk0mdWkL7oo
5ecqdfeqcC2uK3pYIuk6Dw/sk3Tpskk8nggKP3wrLV3ZwzEVbhYQrbs853BE2WUuYnWOcFcwg3I0
8ZhjETTYHy9kqjIy4muX6eLhs9liNCP5HDoHIPAoj0NgNlHVx4hw7i+DWZ23OKIV4Lplfc6bgA99
jKTOIo40qgq0Ik7aH97TekUbbQiYvcv+84V1z24wTE+hATD9Mu34W2FmdIMt8//lVewbq3s2Z38S
FP/tIV1MV+bspVeEz5o9oN8quLtOSo6hu7u9GaWYpVsvqurWTupRjMT/PrrJqyZFzYcOnQKoW6GX
k1oHbAfSQTtCDC43KGjXK839oZLQlvi+05NxQ5llxedPGP6UEEl9nHjpkLlZjVP55XTcMkTu3ZbI
Eaya6Um09e7SXLoMtLW+X//h3Z9J5cGkCheqs07LvMu56c3PH8TPM3kauVKXVq8HuNkwxX2Ru4pK
px0xFy8x+gE9MwpIvJRiHMTenmw6IZfgGL32CmmI208hwPgVZk4DdXoRN22wvFtWp6cXEdOClZ6H
/3366xoCz3Gt6Vjw/wZ6+oSuXYnoH2qjWbibXx929rk7HhRK91Hy3+FGJv8w2qxMchFd3MJyvese
Zu56TFN57M56E2L/ZG8ehVZZCRMRzt6TZIukJjyO3llBhpO4RMLSKY7FwvMEbeDDaxuXwrnB72MY
Ow39wGkA5PJ5JPGaN/Lh00TLHgH2YiUHD0OEeqoVaWowzB1rDSoCEfU5VqgzfhsTUxfvlTmso/Na
dJVmvmIMVWJ53Yq9v5lBeS1jqvvGoxzLkW+cgJAfftULfJDRqT363VFsxxxB8GPvw7G4nTZUp3K5
gXYf18AV9tTWJJRH5Vm+RdrDiUMk2XsXSqyAyqta14asfRxuxrfmECypYBX642Q47axjNQZMJly/
W3+ingyH+XZqQ6YZMCFy2Oe1hvjfirU/l2h2+zeYPuSkzanC6EyQpG3wBRGuLkiB6+rFfYWZVxHr
8FnNOUeT2ctrgeKqX6+u7/UPfATxrwYOEfa1RSYYV1FCo6n+1VM0B12kQlKgtaktsSKchQptUbUO
r2hj4/mb6ZpOZHSAHrzP/c6BdfK7BWnhXbFQVoeLBz41hfR1034eSkk48u2qIIMfNpd35dPmSFAT
05zu7WGyMVay/0CMTCBVS2kAgEn04A7gPGCyzQQG3DwQqCHUs7ZStVzSinB4PVsyNlscsFubwxy5
LX18gBYFpGs/dFYtFI0ucYB+xg7UaCpDDe0QsFN6zPT2P5UCxE3ckKb5xP0jD/ixiwSgDG/tw6xQ
aR1KsCINhiERqPvePUEgQ9nyu5u9cqijKrdOS++iDN+MTvTBsuQllRh/YtiTtL1EUTVHtJSGoUHB
BCWUk+zukm95mz1QxYsEVLwrLGWzqhFxfswzPAMiXdCvCjAmhaCb0hAh0+srQZ1o2NE+UdfwnmWh
YXCWfd5gv96iftYX2kUuRP4Caq4rljMk1Te8MPJ9y1Fthh/eJL34NDgcipleT2f5O6PbxdfOgSxW
pSyCPm9j5zbBX5TX3eKbe+w/GX5pUHIO3adsHX/8/RvZe1cUzTr9u+L0CSvzh7KXZQjEwtdswXQA
5hvAkj5LOUSD1F3Nfhu+1YZGEWjRwLfYQmTiZ+uPV3MQr7O9RouBdrNXhd2pCbJWP0eYEEehJ780
HM8BRYEhjupVo5rT2oWVwE/kNG/4B2SXWSfUonk7yx5oqsVmU2RZlXb2bm0MUr3N//wLXDj9AO3t
GvsAm66GDlTI7I1BF7IQKtrBUy2wB8pxmBlx+ZP67g+2jvlVpV9Q8AhJNKvCjZTkFo92jrAGV+La
g/wwcfL09L6HHk7tthvOFeZZNCeGtV6EMd25EcI7MiPM2c5lFXbBLSSfwIdoDkNtGv2Q56wZ4Bqs
HqqIZqToWwA0Kf/rACSwSAeXehV0Q1BoHHPuuQgBhd4F/CZfTmS6RT2bQG8+i+osQqPMPfx2GVgd
DoCVPoswghQ8ix1Uxvu3tIZONVyUlA5S366KJVZNjKEdhj274bm0dVb9+nFuIMpo337gdPOWhKrH
P39RIWXCxX/B22PpImYZq6pGBFu/PvjSo/7YArLrN//z2pbVcVL2m56HpzSc3eybHOf2u/5cO+QN
V4FoTJ3K0DQgFqkqFEetaqPtgK7rZ+8aX+W0PNn68dqo2EJXVliOPMAOgOMWijBgZFZcTGnqYNU9
SHJuFavS8XtEIun8ePAmYAhsWfmEL5KUivcALklS3YmRQj3p4A90Mpxv56GxMBPHq8dLDGwKa4FT
q7DfdwDOzPBt3PVY51JNFyoUJWrfj24wuCBzz9DkxZzr2JL5tYJ0ofYNltHf7S7nr04VVmNorDZn
77Mg+hqpJWxT5m7JrvB23eNpdmeeO52M2xfFhzB3HJWOgjx9qeltuHYKZf310zswdWVFg5GuWYWx
hTwj71Pi6exOcD6M8DsMjVI9907KfLDvOFZ5JCQSQSzAMsN2pRf4kgenM1aD0uxwQjO6i+SbcHcN
h4PDbiceylrrmKb7ufcT03y3t8RESdPCMWapPe+/ZzjtyNnnXkkGtUFis9QeVg6B5AhUqWXQ7D+0
dWlHAtLZ5wkEqL6ySIMxTBU9bj6QagH0msjdqQfKtUFQlw/S5ka0x5GdRQjSgYgKStCRxj3+rXlj
MVaHY9c9ijBSh3quLbvpFIkr6zOMgrp5cUkGqZBjv9OYalsGceIWRXHALVl6/baMlFUhnNe69rOn
e1EJMiUfMD0EFAR/KpwTqHgeW8vemAA4lBAMvLWvB8Ixjkn1rKPasyWOR+JrTORtA79GhEH46QP5
xLzqHAeB33THvQDymV3az+XRl7v/MFZHjMQZGx7WjLlqDjkWOasVuZagMqQ00NwXG72mbhJK4+4r
teqtaClyTxbTOBWmEBYCXRFvGG53CUV2LfIWglYqZkLOmfsyVVo9/iTARCAha8dYlwLYyF5jj2FE
N85fJWkNslEijVBL2dEe/wMw3uUF2P6tI+bns1zLrj6RMxG/t96qKWQPpM4QXZJHJFS9aYRuTYsF
15zgCW+as569hUJtlpK83rafA7JIAOxmsnXIyg1XIWYvQZjssATDIBxITo5XyCk2EvKYpTU64Ar9
yMzVGYu7/m6ZNTC9Ju+OLW9uNSB0c1W07D54rSGkVwefQCabgnUEc86sziP8eCee3pAW+41h12oO
IZMXEx8Lk6qQviNgYmrAac0bX1Lcb2lQCnebUxqOExPf/9pY6KV0ghZ2DE1Wj4USAgRqDU/yJduZ
QUhY8XyqFQ/TRpVapJ9OQnDw4DkG9nNNT/G6VfkpOknB5hYpLIiGEIniw3PONcQjdn5Wfo9jfgOw
Ih3SDwPKu+im9RRWN0N3Xt7Xx1MH3Om8fIqgZ5aL/i9B6w6B4c+oLX/mY6vehmYdIVRpbaks6vm+
KcigilJaeb01TQcObmp6ZSZv7i2/1hN0uNBhjm9Xu4hmmmc9w5y4e4vBv5eTE7+kQk+wQDMgIIqp
5ex09oyEVp1AAVFJoQAynaUo0+L5M8a2gzOeSUvMsuWN+wRLQa1afn+93495HG1Oxp2/CW61jARa
NOxjm78gI89CxQ/HQ13uQXLJ67MF07Ibjo+spbOKyfuI4azS1d/G/CMhUH/bQ8AwOxkYlb3CFwd0
JDjwM4a5EQBKTsWg5OXvYoJqmaPj+E1PgcDhdpJD/6CMQjdpc9yk49tLfA1Ni2ZJmU1EZhdD6/8x
k/eo28avBl1t/jVFQpsxQ/sBf0r45U1EWvXFIxq8l424h1KpejhKr0o3UF+aNMLAzNfnf4N3+XR1
4B6CKY6kMcx+xlG9gsNpHRH1/vaWQXS8FMK5pVK8FxlXn4vZLAf9bf3nXmbiLrowPc6T9dTYNEt3
TcHibt89qtFJXTNmB99zS9moY9o9e0jGnrK1fswMfqecQ7BwJzZ9aBuhUw/bJ/E4CzGFwtClMVBI
D/GVkmDd0kKboTiqnD6cPWXLCHiTRcr5+C/w6UvyGbs9t6kLlveGgxu+7Fp0dv71D2/jOzYhgdja
GWfB5mKzuA/d9h+xK65sMJWCsIf5o0OVI5nEeg2hC34uOfYBPaHm9VrmvafJivr1RZJwF7PLTNTJ
lEbGF43+lA3BG0a8mYdhcT0YypzhTUEyXjrNmWI8CUKOg1NTwjwLjRDpK7610KeYyvDHejZwhL53
NsXQH5n+c/NmoS1yNbadtVPzEyE3Agk3hsLISwDOZAn/rNjWj4nu+PYfqyVtowy+2cabeUUVu9NM
OwpXF0qLSZ+5L5JmI2JKyDe0K+862rr/xT2sqv/Ff4mxhgGYpAfPGKzOWVMMaiDeDm8gyNautpQ7
ojbbTd+r8jb0qMg+PEyMCvqNJvg2rTFActfzuLs1HtbC3kjVcyNCnmf9YMqtq/6R74RwvASiOvBI
AGR9ojCi5J67FR8gWQTm1ROcEEBObQuARRvFQ2zhpPkJqkvdHskemcv96kXtvlaCkZYEBiAeQZVU
JiUCF7b9pUf9MHR3qusxBI6ujr+dngAAimtHuA5bkIs4cGdnlksulmp3NWA+4dJQWwwBRN02AlCy
9wf5MgPAIXc/uBT1DWpm7RxfQQa3An1LLrwrNGWJMYLzHmEahdxwuSo1w4g8AzEREIjJSrz7kTcT
rD7DsJX4+TczIrZZIU9S2GDEh3fOiG9v5XyW0AAKu537b2iBqOizZu2iLa9zs1fXxiraL5BHiey+
oGfMOOi8CZnhVceI1dwaOqIVy5G12v+Y/FnN8rnsMP9TgwWOUcc4e5SIN+1oW3ESlw9sYTPrN3eo
5RYnGI38g24HEKuu2ll92vctxWCD0lTAkOAHu9yPzOZXUcGROiNH96326hooRXdwLv30OybdC2Za
nkE5mJu9YhMUBl9AXsXEJ/sBm6errkQum3j3XIfy6l/58TYGJSDAuPyh/3zU/FJdV9Iy4ppqIY/O
a8Qw1P03oaMUvXZOMTKwl+025z1QCXKFBtDR+okAjBfZYLsKgcwZEwCa0haqdSWehQlVVDEKG2Ht
qqda+AH8ig357spqBUI3ZojfF+f9L5l3BBF1y0iEV3WTUJa5UFPCkG527D+kUj938fQs0Qm9iHr6
nBYYeYSNiSyreOotBtfyZOc8J2IyK2pLEg29Ll6aaV82sibTmdemRbRtHpXp5TMnuWBpIcpy2HyB
vLX9c5gfJK6mJOt0spSXlsuB5aTwIOAFaZGw05h7fHomq+uqjcavSP5zd+TBfPYY9ZcU51Sty1Bs
sy8N/v7jRZ8dVvlSj1BDmY8Wukg0l+509p2vHh7sdX++g5WGlMYJP5j+WEqqeGJZbQPLLLtgP34E
1tmV0Hanqk4GO4y5Kutc+xD2MfbJmRjYrqd9/kG7h8Fkv1syxsY/g5gG9vDRGuRVDvszCY8w+4un
RMdMl2YQfdE3qpJPpv14ZZnMi4t7aQSB4cV79zNgjF8JE6yk+wC/3ci6S9prX/rHEMJeGziJa+mz
642dFfkOM7ENLdzQ/wOcvJktiBwA/9JVtkxKt7s6UFAefYHVAGejnYARKauj8f6uAmzwhh8AXCAB
sUWOawU4cW3tEn8G6gnE1n7uHeJVLov+OxQAM/T5m+83E8payWh1XTVibDPf+CDEaEnh1VfCg5b3
qlQF8NvacHBNxITAGnpO9R1724+xjIKbV97UcSlDffx9OY77PspZ/S99xtu5MxPKGMTChhFOF8KL
PH4Mu/OI5wRz/Jrbx94yBoosCvnUhB/vg3rrcDSE7MXxmBEVAG34hl77IbgdiZEcj0nrvgeAOExk
z9Gw6jtYuJECTDkAQWoCw9H6eiB/qs0kkrJ8m+SKu+E5M2skKMAY7egbesnGSEpKPsT2UiVq04WL
cddhgyZ1cuYA75h8nzc5ipIvfLjPCsXsDK1NCm1VLr8F92hgmyZtrVarXE2twcVvSJtJxfwpMGn5
D10NzrhHKBVvN5sJ/oJndWtUgkpKfHkei+ICxkMWo2I0/d9FLApkxNe6BOn6LIzNSz2JUUmnYfdl
JK4hdwynvGuSBX6myk7uLReIAOsnnrPYZ1TKLo/aXCK6nk6ocCmCKvukqN4cr+tO1A6pShArw6yr
4kBRXnYonLiX9SmdNGG1yk+ztJr/lh2HKVqb88H033T4m5hY1tyPXdsw8PLsUYPtF+mMp0C4TSaQ
fAOIBZZl8C0PtFughncVJ46a/n/FNBr4F4m7EDNB4LA8Ra6nsoh3sIEcpuDttkXfce4vImRg1kQE
3+ihelyHxHHa41fpmQ6kN1OIkNZn0ohesPK8FIZu4Hjk9CR30qb2L5a0U3MlaGLQM8cjgXjJr0Ie
zZnXqky5Bytaq4okJyKjNN88fQ6LVR7Z7jSo98G8JMbHC0zGgK6ZBL1GqKCbiTLYIPpVR29PDaM6
qiMdzjudP9tf+/Cc3lzZ2puWG1x1TgLb6tKbDfTFxoXjP6U6dxhbynK8Pt/kJClv0ognIZQkKxaE
wWFTGkNYtTjDjeOmYrcuypgA4VfmsYOLijNUYrn9kqurR+IPuTuRibx4O0A5W+qOKNy8vBfa/wbZ
lqzaVzTBj15sQnfwAOe5D3dOZzmsVq7Q2W5kGnWAADQawajhrtqRzDucn6+tDHUEZz3/xoTjebO1
Ov3jixM1vC5HJ+WTlDydEJ80zl/SmCGOQg7Mpbaurv8ygQvHetWpp+o1H0pc752db0VWR8YjYCw5
H6z6Jynp80wpCEET7CyqFMCu4De3MKxca+G7FnalFMZyYWnoVegwVst9zds8pn+oSWfYlXt9lRW7
K3FT7Ps0hm88EySljn/Ni423MOWgCBz7GKlDxvajpOOmv2tSHsgLZ0rOklw6KmE5CSD3h6PqOf/Z
JcRzcC3V49BmlaPRMWkZwseMphyZQZMUAQrMasU+QGWKYW5QKsH4pVto/zrdEU6FbNwO/Ub5zBXn
tG4RUVA9JCUk5vFE/oMLLZxg0nKxmKAz66VtQykgCvufY+XWH5UPhGPBkIirptpIdJnnGjdOxx5/
3jPYQ316jDAgC3WawqIagRkjr95vkChs8fAl06d1++7SFWWVXHrU7Wji1bZ7DSDoe7P4fXinFzxs
HDGNTRvhf3z2yZ7u+guG2sJxmB796QdNeI2yzNTcnC/pSMo9oAFoOIaH3/9HZlb0E2ndmboKlB9i
Y7wDG5xJBazpgyErfBdx9d7bgDVk9v6GQA7qBQelMRIKzUWLOQXibDmfcsRjdtLhj7T7vCaOarRW
LcAoCFXbSKuPp6laafP2/10Vb132pBtZlTmoVn0ezmmzlg1mRlsb1YSiW86DLB69JSRBUeoh4xrH
OuheQq5LpV4PnjDw36q+SCJGfXQjgA8vPTx61bazHr4PdNi5UVKYce8gZxh7FTeoxsy0/RuqhoS4
zCg6a+4dHTOKKJLes3CsSAeAvzyzE8cmVylEONXARlJy6l5OJf+9kWtcAOH7f24Yr2676y++BgAK
ikFeAB1CrJr1JoKvHS/IM8l1CtmxZiAXU35fvv/yyhnJKITNU13yfknwkhO5ERwelLDzp5aI+ju/
lVwjjmgH83PPrpkArJwWc1+sln0yJ7B1g15VXSq4dMGsJxuSjUBkCkySrC03GBLlDo7Qj3BAZh5Z
sky/0/8bsPX4ZgL6y9vCz5zOiIhxmI3yfG7EkHwO3Dw7ihdn5wDZbWit2GO/yO+w5jNM8x3+07q8
2KT9rvR2uHGhh60my+1JnnRdTJmWybksGvd2DPjBVPU5YGvS3q5WsD7oPL3puoQPBBvnGW/smggg
k/Lm40Xly+6yAH2/l9G/0UChlfwgcQVT59DceTGcDOXTfzMJvzB5NSg0OGaG5fV4omPZ4+DInW/s
pJvVu2J2t7cbGJrDAQsfTRgKggWDuzncs4wYGuMDnmUkgRJnDJxNOSAFYT5v/lq/qa/pDO/JTBhE
0w62TJhswHKaCEogaU2ol0OjuF0R1UBF8iJ3tab2Z05xN424Z1nrWKp+eiG0g90uDnG6+aseZ2Xb
A5qJWaxoH7EL1Q8UiI4Mh0vKjN0fBGs2zjIUQnEiOrwuc/YT5OpCfxXJmMGlArPkzlANddR2XNBs
vgJxJiq3vwBKtrjp8ij0eUlmQh0s7TdDJT2nry/+lvtnUwnGvMLcO3F+fvVP4ZFUS8/W4mVWYnTG
XSTbsl6abiEScFV51nlM+8u7yw4Iple6v7HsVP9lsqMG9q/OTHJxdoaJfKGVc+KyoJoFvfN3SfG3
UZmUEpdlehGMbtfK0hOkqAerpRj4EjWAxG/vGlJ564Xb2Xs+pmJf6HtRCvCK4IeyR3bmyC/Di0tz
jdugfcXg6uXQLMOy2BK1+HIsklXyfWkjlQfoJWB/ynOvI49l860p31D6n15TX4gk67mlfptLoCRM
soGcBxczrZlPeXvGN8IIgvfL/6UEu7DQOgd7QEXsUkN90GImltslD4OPDrhwnJCZBZcv7++C1DFJ
7mBKXLiCsAC7T++l+UH/ZBd0ZFruW2yZ6RLp7QGQJks8ZqKW0yO7OWDFe0QO6rsrb5pp0VEi/3Nj
YIO++qHkzJSCQVeXa29Q/FAtmN2hE5W3IGBwWHknmS7b7W20rsaZPbK6PHe7yR2xM3cmEM/bk1B/
O5Q2PyK8VrMNv70Xl/wt9A6vJzpSNLJV6cewulQ8viqQwJDzrC7KPuan4dt5nT//OHItbarKqYbu
SrbO1IfzZj+pGO5AaK1154gF8baafIwGxT5Cy0KuayJaJPV6CwKlzIvgqk806E7zy4BrMNGU9drN
fqcjl2PL+QlaC3bCqOftTyARKq9Q0AzUZ08LA40fizYmEoUIXjG/UsC7Qye6h6BRoMJu8kfl4qOK
qTjIULyl9mXbvICBXedjh0z0E8LxDKit0XNVXSoR4QK0+nKKxLLzptJwjM5yoOE1NBModaWtimrT
yDEhhNMWWB5U0G/wd33WgpTAgvOP8WEt883PTTO3PYnMX2LkS0eI8Xbu2NWO2AyiB5PPv4+60qNh
tIIs0885zOSrfIUFD0XhZ6MXF+kuSmWUwAQ8nH7yNi9v/hC3x3gjMSAEvYKNwxga7sEiI/ncMGM1
UGWMGIoBRrZjC++BYFmUHMhidTkGRluFq2PhJ4mXXMr/WO5XPjcUkEv1k5fxJZMFXMn/R5a6PliK
ugUBhklJEpe3V/7p+j4zMUzs9GlqjX17SlhN74nJ7C2oTl96lL2uSFHsloJCeJXgkUW+YcRGTSNU
iERmbQ/mScn2JHS+xTzN7UMdp+Jj6nEYKK9c6xr9agkks82KjjTIr+mfdueh/xExo6YTsSUJ23Te
m3O+Wuo2espspFoKfcGI3RsLhQ5yrleYKgrlDhfsHcUx/dNs3hbO9n9lfrJDwOC9i+eIrNzAfb9c
N4we+AjBhamevnDD1BRFAg3mIrXEsn5E+SPauuWT2F4N3ZhrwxaftJBxLTfaRgsM9ZLJxwLJa4sz
xalm3EpYmp3MSjrgyT8YQwlziNzqFeLM/N6mhSpPgQYjce9dXgfK0UwEP71IIHXQGVqTNgucjZVu
Bs0he+EyIORrXvm+w24vVnwGXuES+5aGS96KOmHc8BWjR6cNqYTVJjXP4Yx5xUYq2p8/E4fz3d7J
fO0IOMfhWQ25X9uwU09K+EezU3s3yU1RF2+YwS3g+jfqiFRR3DdGwYb2WT1zpMmV3wrTWUaQj6dI
9vq4VwZ+x+cStljP1HmiqBVrsdKrVd7Ut0oQ3k5154BEyAc+87RYsfje9jUcZ/3vY5FY5UoETbPx
c+VFbc+vDn8cabhf3sxLAZ5De66UQcGKmK1qZAoFYbXgIsRz2jN+UJZXp290tgVWnYJWs1Ym1Psb
a5Gkizy39PuLCdDPxKNI/Ut/Skxc5XYWyo/KSQKa9ICOne/fQ/pB2xB6nzoIEHkWVKlc/mgXIANm
j/Cs9al9Fw7YW4r9T7sdce+dCO2T80XkxYDB38YLRR7rVpHifdjNG4W9US1dOad93b3RHfEWSCQt
38DDXBmo6mv3edsUUx+Ke1rHCocAfPEtR+tmhgegEh3ScoozKE0Ld/iqIP5VXno2+qt0NlgV04sb
aUC7Iyzgxxd4cYkbA53BOTJgO9FanG9kKVlV7aXCOZCcRhotVW6i+onPXiY/NR6EzkYdtAGhqw5G
q3xH4l6ySqN9DAnczwhiVoPJwZSoe+E8xxF5ONN+3rf+Af8d3YuGwU7AbAImblXIQdKwLRyTw9/q
R/CQfy2Z3fg/VCNUzvx/P7/udP0kdveXhYrdZBHFjy2DT4l/HEfVQGP6VgavqjPtP8OPencaptUL
ZyBl9D1jDaemXRXX06vR5hObHVlybbZ5KBperrMyabfCcLOJKXwrGLT98ATTph2y93VmCmc+U7J+
f8Q+eVOvXDZIjl2hMegfVA6Ol08x5vbv6adnuEXf/cwvydop8GqtfyP435GyB0O2Jsez8olQH9m7
Fc544NH/7jhZcSUU9QnZG123d6zuD3uAWOiYHdS7SBm/0kln9Y6AJam7P6M8U4TrstofunGfxvt1
I2Z1ypARJ3QFevS7QZ45IswN1ILx1CHH9rtR+PZcIEoHggGF7TIqIrYEyvKVLZV7Pbc2mp5MnjuK
wgOHiRvZzWAM2FHkUSd+PqJuAb1nKTRFjND6FlIjG/grFcnsuu8/wzQO9wQZqugDX38hr3McUPCY
mFE4tsbKNsPZ5oFgkGB9stTnkXSQQGROaD57RvhildorTEEULBckFQIfx9V60RXxkYNGNsjz5Ym2
Db7I507R6KGwvuws8Ul+Oxule7CSQKz+UPW4sqTQg1YMmknGELNhO4OERKiNDgZQakRRwADdODBD
HUG/7BlSRcP1rmVEHlvfebirY3bN0f2OUyLd32ZQqAg6otUev8ATPWPUsHzeCNPwC9xjGsmv2Jcw
1dPXJ+qa16xqPxIRYDbUFb6moDCCD2d0MPR4DaZqhkoKJcQIbny2e+6Md7tx1UAZRJi69DXiXBkF
3wcARAHHPMraPACz/C5rAJYijlf2/NrjvA6eeQ+DQPhE1Hqeczv3N+MiS6ADr5B7RusIViVRapun
GVMoUJEJ/N1N6eIgnCkBLyYQwrHVNShCYdhNHKEJytGkVFB+mj99gqGJGiprn6i8oQGm0ZlMI2b9
RUO3unkxSA3FDTmduoyHHHHc2vBZAgTJ52poS1oaBgN3OOiqbCtDNBomksOyfDuxH9IXLR2R0JLt
0An603IHHvrb43LX61yr5UE/9LMGxWvNYv4FFIRE2u2KXIXttRg+FClo5D463tq5oEh/Rot7vx4H
Lod5NjcRnunZ/IzbATr3obD9i3bAw0MNvIARvKIvqr3X582l8vyDjyTvoVuhJDivs+UQDi0ZRJHh
1cL90ddVtBTdMfeNFDHEj/8pkpMzbmN4gFdSL/paetUn3eus4JPtTHXtCmKQVgMGs5MbBf2/MFLS
nIZW/m68LAhiPX3j41I7hPQp6IxC7lNTORpnbePiAgFeJiRtMZ9R4ilcB73PnXrAEt//VKmesC7A
U3DpMrjBDFw4hGrZ8glKPRNfSR/v3MdB1As5m3wSElZxHeSCxSMC2wFe5G/LQitsW0vRW0vjWLMZ
H/MNe9toftvzJiPcbHw+T868Z9PqOF3UE7DIZMzhsit9Y3E5dgemg/Vt/Ci8h+xGnIp0ZSIn3azJ
FOmc7nuL/jDeueEpRmgc4I7yIbBIwpCK0g+H2y5GSZ83jxuEyx1UCUx5hIQbkSEBmUZCRibjMVfc
SgMqnKt8nR5H3dwgi3U+j6t3dpycgeSd/5RiJ/LygRwf7xqzb7kG+WgPUOMNI+2R3fd4tU8LctSt
7IkA5rPBd0aH4kD6MvXlwDIrNW6F9usE7tqAJrW1Pt64u10A+Lzah/1ULkfJ0UsHt/99j3AB3CtD
gd14vu2QQTPDyE1iLsS6StQGjeDDOXodWue6JdrvKD7Sk0/rTKydPzhVnhEL29nu3ALy5lYuRHKR
7Gwl7CQMifqjeQAlvyPjPuZAIC3Gln0jCQmMLM9m4AgNNdhzv5V0k9yj8Zbaw6WuMVrTTnE9+TJZ
wARbjGpj4DqXlxs4AMxm4irkOQpp1udSh6efrP/UdsHpxvDI3sy65YEwdTy5P+FDdoRWQHoVmKSX
KNun0YLXnEwJgNb+xJ/6GesjUMypK2cdPInAifZMqxMK2+Q1AdEbI8Y1xc+VQBx8FwYs0gRqeMlv
uhd+LtV5M1hDmUcsXzYTsDWTeouxGct1ZkDS9CVogAimctfytGZ9xL0DZK6yyGT0rPVRHusmLdT2
douXUP0lfjsYBbdAro4EjqUp5tBrfQ0tFFPHsv+/qLxmsYZSLwczJvDiVosl09FhBnR5eJu8EBn3
jGaakVXM28iM9eXW+9SOy4gr2w2C+vxnKm9AdjpqdOjWsF1O0zuwUmeH11Eaa61sdhbAGBdcARDj
UofZbmvnnbT9/2TM9+7OjJ1vdKcLPIuYXncI3mbr9lrsylYWBkUY475OKHEOMsNgn6hmt9hwbjj7
UIDONSST5OeuUs2h1JDC0Pn5gY5XlCpwqRK6Ms4I4WkEnRXJmyGPfp909ZjQfbmsFly8q3q3piaH
Ebt/OOl811xNUgGqBlV/eHr5b+YwMEOh5DOcXxDzaUlN4I1wLHYuZjqnPIReI+REJMcmqOImTDp2
hnR4wH3OmqfHmOuyedbBJqc+TRrvywMaal7PBKGJbC867g792DSgOYuRN3h/DKII0XF/ueKTkrx+
vN/q8zqC+d9ExTUB1kb7el31dqWLyqnt3Ccl1xvo6PsqwdmwQV9K59fj7ftrBEtxWln0frfV4tJU
IWxJizauq3o/2oa4XEB0Hf40jXCBf2ZUnu3D6Ug+s22F3q+0HKLWQ/dTE7h3mdesW53vVUJFeBCI
2xRZCyaFQfZKI/DhTAl3xpydbE1hWKtzaJzcjGd+sPr4nrYGG3NAPYZy76IO5ZOTlBQ17NM+6+YU
r16IkteQEg169oDvQHB+FXYJ67XEs5S+CnTZFTjAI/qBmUrXLhUaJSzzHbmb6SuziMpeRaTOHIW3
Llqd5M3XIXSxw70DrGwd1SF4IkGTuWwtgNqCUi6Jrp4tfxNiNkVgGelANH7ixTOABsUJE+tA5+YQ
jsW8p8VAfyBC3wH8IhtoOyQufIojAHfdRfiRSeup45baTsW3TTPLUHkEdADhET7WKb1ZMwqRiDka
9t+hJXcnt5mk+/qfcGTDCUmF/mmNjvNRWibAZJC4EHfdv2e5ZQwxK34d+l7UA9FRyxAMbBWameXN
tZ0Sa7WiKGzlgWdqdhBNbuUtYJYH7uSqtBzqNWQ/8tBq3aoX+v0b+rarixp3AXNQPRQJhzgFT2RW
/EQQMCA+K01JGlrm5Nr6lNMi214EICw8zw2kjSq+NOFe3PZDW3CRDTU2/RsKpDenKZxelLkxeSPt
9kQRKiRRJ7CzVzSzEO/FtPMyaU/2Fste1X8cmewJv42YtYfUr+28j3XTYEiu7KR/LkT9drpqctET
P2NSKwVo7H6okHPWagSIHkAIjwzhIxeB3KYIahtGNnLSA4BXAMDsqbvQK2t0FU6uJVcRIZ2mQN2p
LLDIeuQqOkquyTOBJGC2on3IJUwI8HqtGytC1r2zI6co4x5pRi+RbA04bv3LPoUEgCleu7DmKwdf
vlKmEx8ZkNhubc+HMpJ8uiMDkWNqELyh7eLAC0lnn8Bj2Vp5j2xw82vMkAe1irGSMqo0UUCnOdA3
nK40qHQudwJyYnTERJunuoCynhwBiBPI6FUPfJspuwMRijTpCaR+NKX14Bk5BV7oVE3iu9dYzlbw
7+6dLmu/YznL3k3u7LnNyn3RaKRWNPEXK2ZTasqlKJC8q1Y3yMWhYqkFs8QJYOOW/ouS8EBnooPX
iq2l7gDfux1ZYgKJ0t/PZifB1Me5SzJQ6vRuCwkx5m3uYmpzAk/O6tgx58bXsbaFiVm7PRbjZ8aq
9WYASwFiSZOuHKcuLz000SBADRo9LiW9WM/cHEjit0P9v07hWP5GW42ldAJy6Nlwo1kRDJZBZ98M
vyGsW/AgAYIcBM3r6YbIzthoDGXnMT1+fewTYdR9xR7ydvYTniJitcip2SPePjIhP0aZvcD4plI9
2WPq3PCetPagspGOtDJ//XldLKYjkjZGc6sXwp5btHTdK8uZ52Rxlj9DvAwn0qdVNl5xoCQNHd8r
2QsywJzi0kpUGDAxRDjK8E3rxGn9DMRliNbPV1T0W7PzmyZfQLdDKT+b/jJp5n6roES9myBZridA
cBpWyu4uTazdk0rV3vOkAXW4ThvdjpfqNOQGjF4PHRCyOkOOJg5+MitufK7LjXfw8sJbnEMTCBf5
VbqdX+S6G9tdnHc7swWlFfXOALtDSU6b8ExdFHMvYESGZBNrXlpNb5KhLSZdabmXgE2aDxprSEUb
N6mokjdQ1kYazbTK9DwGy8tl4NIGbUthnLtYLrovPrevLLyIB4MMt7plqwI3kYZhThQmGz1ccqMx
e1F5qPBBr1n4vMeynyOTJ2wOOxhDE1I2XCo6Gz1v8KsSr9FcfW3qreunhNz5khIqR1vKGUux+6Cg
Vg7SBSFEA+0zfcYb1c/rPZoznS95zlzbCJP8ieMEdR3BcVG4UmFFbtPYTP44/odjUI10j6hhFeVi
AZE6xsvfLWPil48pUtj7q9zDyiwnzQjR3y5SqTtmPciPOfHhqfYba5XfTwO2t8ZMR+PuYzmu4Xpv
Ih15pL/88X0cpngBk67iPPbrgbPET5Ljgg+ifRdlQsNgxSr63aGJCaHLl5fJpQoxB5Huuuuvs7mP
wv7j8U2/84dfmLufgnCfvsEtY/np9jc8GfTUClZV1TIeCeu8YOP3fCVSpFg8UXcxe1A3TRg0snoW
EOwT2vC+TtQLqBcik9y84otjmpitDurYJj4swZY0pCKJB9mDMjbiaSMMHp5R275PE5tfCH4ed3U9
Froqp3nGkMK7kUoBjySCKAs7WESuSibJjAi9yUEKhxoJ67HXEG2BIJFPyNzE/e2teigA7kORTyni
h54PqI22jvDHelVwXChuOZKPlOow1H4Zh0XPLpmNQxk7FQLbRfMlPn8F7dsFsxJP8/teV70Iv3mV
aHhd7BMPttj+1NUyvTT8AB3IXEymp3smg9iRSLvgkmfBZGWoO5ZiFO7gjoMd2tG+cLueroavmcRU
9Jm+ni9a9xUrbiEaNx8iRkRJsF+Y61y2g00l/uVs2cKQOKM2373wp6kBIDcWtBMyEwRPZdUHF4NI
lXhjQZvk4VrCsMszJ9pzTimF+R7jWkT2XvULeEmYeLu+aY9EZ+2T8Th0iYtvPe+TmcAfbdwFmlWo
Ox07/gOJGg9rkVMdmOoj0P8ZcE54522B/CInfsCHM7gmDbmaRHxpiMVY/wEJdrihpZOywLyP6Jie
TrLgiKGo1cr7FxjNPuvgstUS8LeR0Rzg7GKC86dvvCDV3ibZaiytwHTHuyUMefnJCz0ULCNxsydC
bAxAO6Dza7wZ+Bu/sbdU9OXjEJfw+Eil+vCSeiGrmUXDDBTKKnGRdsndW9FWY2g0uKbb+KKLW7eh
ua4gkjvLf/CQt7lnAF4MBE3eP/kQDabwM0ooHludSjKjmQN0c344TuR/P2kvWU2SdQJflOCAPE/k
he8bGyjpLdZRHA8q95Tir6XV2poOxMh+Ucy3b36lWemzFo/9nXA+VlPOuzHc7M9rsKXztz2JcVXD
AZb2Z8lallZK1WAIcKR62fTEKhoSNwsmljkPy8k0bpScnEVB0CZe4+KZr4vT7Oo3kyu1zg+j/xxU
0SnDXul5fHEVxIF2MIbRwKIwDMoQ+CbIHWsB01UbZsjto8+MbSXUl5pSCUbrCfi2+XewsuY7Jcmq
swfRulznTda7Q7E6tgZ0zrzp+n6zYLRm1okh1a1x+U005TbeK7HcRRF7WuE05bcrndhTI6d3NO40
82e+HtSoJqZeyzvJcuIycC+R0Ak+7rxY6IgIH+YZyv480me7ulGQiUAl3xDtO65KEz5/64zdU9J6
dqdxhToppTSB5/6zt7neaKShV00BzZoLR5TCPbhTWV9RW1VVrqTwCVb/lR9lmIo0INPsh9kt4iv/
WtP8YOFyqBFiZW7ql2baSvjYwHwazNpsArqCqbxXlwWMy+F0iIcNHIyUowhHNcVpV2M+ANmBKvjq
1cReoBy8RbLfyVYVnPpipRl9WqG1qLudwCNm5Dtcs8HMF/eu5WTX17kLoEYn7nw56ijWsdDBpW8e
5uxCTMidZ3c9AOpp8GXOWVNLgYtrwkthxcveFfyBLhziLWyhrEKu60PubYQG45Tl9BrBCpJfhOpU
gMcY23SbdYHOLUWzBTuwzIoK9YUiTd5qpH7ljAtiulH98kdLL08kvy1XMGwdaHt8Izr/jtEz2Zcu
yIpvqu4GJgMbyV/dZiRLcyrjZmpv4116/XOat5cAQKJKGccuVfHLA7QoRGMv1C8KJ/+1YJw6Y7ys
PzjPT/Mg/o8gLT32XRU5oLtQ1b7Y0A5R3D1SztUmxEum2A3u477jRk4S8G5B8B48oNPTq8ldclzJ
Nf7APLEfFPtAbPIVLPHQXZFi/LXIRJ6Ea430jjdK0fn2csJpeLCTt5WS7kfg6EHNeGOgGCYta6tR
M+w9IrQms6aIT4HOr55L9WPsy1fwXEHpmVPtefvDUQpKaZGkFTYAzv//6Q8XlcG+5MkZ4NIk71Ot
UUPocljS4hMFMUeqLLsCHdrXaIm07HALQ8FBSmgZMnDkfi6foef0pHcBhhP6k16VtJ9qvnQdPKtR
6Il391Rb90rROM8Sk5gi/8A7zDzzyakp4yNmSmaDbtqvTnQMvze9+Ceg012EGTZ8OLCiDVEBz+33
uItcm/RJts/egMQgnbP3VcmrlBBbgRbzUgRGdy3BRuifalJMJyFjR2oMWqn8I3BSx1iCqoF3z6nW
i/bsMDRWPt2rdXnzyGlERTDNm+wLAGa4bupuJCKVAd5XQTKEEhA7RTcokLcFjPh2RyWiniy+Sf9N
womgP00pyESqGeOEW+mpnk1i2A1ksX9d9M32wvWX5A+QhnIMU8jdYkrXepei7zUyE4Z2hX1fAEa3
fN7UqdvaI6oL+9OfvzsFliBCJ7epIScj3/ZiBGIRcQ7cgetoIhgIbuFCF5F4iPSUmY/UFUt3WWBc
amWQfbH45x15HC0SE44LKXH/n0iozefCHGYIIBCknNjYy7n1+VQTlXbPEHghkpYgQsL1pOmFr5d/
Maw9Vr2rqTmcgaqy1BswtRkCCMK+1pNM4N5lAiXMCTFd+AdvlgEUiz9uV5fBHxrmXVV8oxCB7WK3
k2jgdWDsvReFh7pcc7m1+a11Gl7IjxT4nRcDoFDVJSAJIzmjuUDp4f7oInihfHWAitDmvTQS4bDX
rvp9IZ8I3tn2UHjtZkMQctZ1zWdlGNzdzTgPvIcHLFFJVwgdEzvtuF9g+S0pWcq/pNfx/xQ55Zol
SjXZpwYJ2tsiSMtrxe2AgbGVRwK5buFhhPqx8KBRZWbTw+gzIALDlhplrz3FWBnHlJDTFy6pfMAV
y/XMKA1wwU3EYJV790VvMNyFg5e2jMAO++tHx9NjpDcUoBkfdq0U/qD5VZdc2AIMmGsbCMQDiCtn
lyi6mUi+4fgqhfQJg1SBd8wsLsirLIn8paClQyUwIQgmIu6BWqzlolzlba9/k/0G6Ub8WhOTJtvz
/bRW5Iesbs/OnbDOSKpL9OviYeNyty3kAGyziARbvPuuLSdgrm6Ox7fC//w4gTighdisVT/1qSjA
AjI5B33Urz5uJhPeWU0ZcwlVm0e1ayLMnGnKLZnMgN6bI6aMvrEymlUAj5NUywwoEH3ChBSgJuej
Xh6EL3053hCyvJ57HwDyeCPrOZC+P+xmKUlRQjiTnb4AsecLdjCz+/mWnZrL0gY1e2B74O/xTFIX
d/bU8YySQNFayQJ/fOMUm8fldPdRuAbWpL6vvn694+W1ejTrPq3kmgLJLVrM3ObtrxcQHSrudLSU
AcRyneab2IKHc44hqTq41p+51NsJ9d0fqSz8zcwWJ8JeYA+4EHH/8IMyQqYk2DhLvIQTljqOxVLu
5pXswoZ4CNqUktH9ao8S5R9IA+AgefZ8SDQvDmBqC68RBeCfkTQ0H/24kdKvRzetnhUuNSzIQCDl
FEaSRHHyGaV1uV/pp7O8OIUugxPcGbs3b6R6mEY91BChrK48Um6r8wWfhUW9NidUJ0pEfBovj7Ot
q/Jta8Jdvpvi7WM5712JRx1vVWkLrihqQ/iKkIQ6IvF+ZAhDzAO5Rr+ITdwwCqySyux2yDuyyBy1
bwXvZbxOcEOdCARWG0gfGiMINYaYC/jISR4V15Ezu/Yr57Lszm4p7eRBW2pr6idon//E/P96KWk7
5NdxG8//lOP5vgC6DorakaeiumanKcJps64/47ye7CJ857HV0+0dLuKRJFdt/gfZUr/TdMBhJDl4
6fV8/M0sR/4uhgO+jYOn74iLp1AM6tO2ySanr3qfxzXbRKaffYCpySY5sGiBDINGaegBXAjDeN59
RJ20QNti2Qd8zAa27BlW8E3ZFCY4brBa0UbGUQZp1S64N9sJJGsDdNktej12XA0uaXMIVQI040Up
XD2T8zh1WPA9b3Oe3si1r2bMd3IguAeGdpRtASZDRKw2oqgZJsN4Usl+JMb/gVV38KFYtFFMcqyS
ndIx0tUq5S8kGFbC6npT1MCx4okpqM5iKyLp7+FTH/jA1N57QO6u1v/HEv/eALLRW48mHyO89U37
XlH03pTcS5APG+neok9oCkmgErgE0K/aASWvJ39zadBVHl5FoLVjv1CY3cGS1JKnejXStf4SJlQN
FsGOSl7I77L73d19LSGI4p0E13gVMK1oBHG/Jrdj86c5hN/C5sFoMu6Mx8NYI7PPpLZrQXkk8XJk
dD5sRmUHNOcQVGYnAfQYnBJGIlO1tfHGyk7kSBQ38M3naNeT15l928s4AWyekO/TTm8sYOMFc38K
9obBy6vwcLZVotfZVN8vCOYjpy/C/1ESgoKzXdWvL4F1dwbLRIR/YGLiwVucvpWfFaOGwNzAJ+MT
X+V6tEqqDyfa7Xg7NeCJuKkr+51oIAPMuV9Iq11Y5f2cwG5zQtEXoU0RWxM39arGaw2BLWsTmlvG
35LjX1+R+jU5zhwixpUM6bkijTyFaFzQK+adbFpZm4DdxCAQ1oLpIIsupdpWTfsaRjFscErxPbEd
qTrw+otpYuannYS6/6qQJy0Juu/wqhEa0lRKvJA3W+Rweg4Ov9ibvDGxQ76xaP4wqLLf43LapuPi
sdtrR9D+524td9ReWK9+v3lCjmhasGz1LHYP8FAO8Iw0BWrTMJieIOIh+fumvNOioSu/WhVKFKbE
DErbMcNe5gxYHONv4Ij7fpF+ROL5WTgNlSCWaVSu+rv2zZ9UR0bZEIhP5KxThv5Q7e59LRk9MAtc
AM/Iu9IPkOCLMXDjFMKvc4HRW0Txea8k8QSvhJwFQ8UrMjMZ6u3oZVgBneOT949FuGeW0/4WUXUW
egYfdg1diJYCsjt19wOiBSzbQ+UM2bsSYvb+VD06AJr2TM43dcPepm3RfQcbVulNWsU9p38pm6C5
HEKAGUhmUCQDIzfjxyirgReu2S2ZIssBvo6oDcl3Rf/bifqL1hlzJhDzokb8/pjc7uBF9JvaaNod
qE/H6hRwS8bjXqTdBG5cpq38AEcFhHq0qLRMg2mkdjklPYv6z+5GhuUWjjLmgonNbPkaVkMoZvPL
rEiHk4yyXaH21QCJ3cTW6BHbmqvXYDDTrVxPcJfjjfDc8yWzSwYH3Bkz0VnO2QeITmiH3JVB4ke/
WnFQxbEKMhCjDaO94GdxKb7tyJB8Op2hXJCZD3t44nP8V19WuwGkd7mKmthfKZ5RBfg4H2DFlWnq
8uJZ7ruTWlftEPHhtkjiMDMsigbfnVI+IUVb4hWl0p5ewGsHfheYC1f3LJR6htx/DQKJrhpVeFOk
0Rzc/1UKZoY+02gXzKjJ8M3Xb5vrNO5Mt+Z32NB3moK/z5c1DEMNFbP//6DghRYguJQPoLlG6dTg
ekBXvN1AIebYVBEhiSaxg5YlZ9Dr0Wy8cjUojYuw/+0VDv5SpQ/n+9GY7LB/EEo2g3QDfNhBNqsH
DEpIAifD9vqTF0A/AChfRbb9ViqFjbyIydUv7Ahs61eAciaZCdi8xiVVUS6NHLm6y6KV6rrtFacv
GmcVd3It/IFcO2ZPO5/mRXFRfDe0DacRXz8fDYBqSfVC/JJH0OAzlfCNmN2Fb4QA6K1+H3pSFykS
IsHUGS3hQGD3uyEr4LPY8CQXEbmyMO06AX/WaqztJkRY4aFUJNDNz3He0yImdvKIX0J2A5fkZMxH
VzcjnfM+ARQ6GUMpjswwtVbXWqpfEd5QLSOds5Ba2PmQYqMvC+rwuYLXfzccsGAVz1JwDI8z5TNU
Ww/7TjxShmJe/PdkzwY0SdpvYDxwBTc4SjdzhOdlRKDOO17khBWN1jdxYLHgTN4i+P3orL47fM2W
qgjkx5VTRRkS0bmuVV6WymARU+25nPFv2oCxU9Y5/F9Fr1lX45ck8r6l2IpC/RzkKn53LMMuCHyr
mUXEde2j1W7iDpc/yjNTZUL6Fy6BQpxe8h0+wFnAzR4ZXdC1/M1Wy1sknNLy7VbE//DOL2GFbhhq
ju5WNQuF3Eop4YEOjFoz+YQhAcItW+F/cxaP5SB7xHsLOkNrYTzBA+dkGLBcHsGZW5CWlP3U5Zup
RVDpGpBdtuNxy4UibPVU3rsqc7jXTkBXJ5yfoQvjkOnKwB9cO+5h85geXefKxHY2dHzTgaTd73RK
Ez3Q4QLln68ub/djRI21mn9oehGjSWbdRk3PjqqOP61uFgCrBqFRvzD+W+gFPQ3ZjyRnvHXet+r5
uomHCU+zfozfyniz18GVMHFLc4EgtjHDkA2Y1qH137xN5TTrnapvH7jz1fhE0KE4D44OCyjlo3wq
VywPimV9bbfMfbssaTSFecFnbfoH8E3UaFfCzMftzFX1rccmiHWU/9vbbcaWeT2Q3dFK9Co/Me5i
j3Qb2TJl20stPg0YLyKpOeuA63PrJLMBh1NscTdCoizSOM/uSDfViZB/N0rWi/K7I9GArOnDo92U
yxxhI+YXXtw4x75/ryij2e9Ckk7nky9AyC44c4/QIgYvEOXcYe90TxWL2nLDH2eoGVAydGBKMB/y
1SQ6o1uK1oiZ4BVL3YBzjf43YGWNnVj9oxxJnB5uyMmdcBgh/AxOWXn4Doq4XWSMVORAC8LfvBS/
apW5xxGwTXwqeoROpFLiQnkhrH4gnCEw8Vw4cH62Gp0oc9cPVuRJKsU3zn5JaYVLuuJWtqtOLcsq
4bapoAyXygktH4Qgkjbk17oI4YTzR0Hzg4Y/8a1LWl6A6oj+g3fBmfRNij2+bKkLK2yPJak7kXL/
Jh9L1rijbQhOVxteuGyQeDEygdR461R/awHnjNVfa5dgS/VIvct4hUrLjloUv+GBSOnRJBBXrhp4
ugTQu0elnaLFOHU7wPD7cWIVubmbpZU3VTsPSLtiNJ7Nf6ME9Xyom1HpcxbDKaS6BLYUbB6Umjyv
B6MmlbhPAEygmaKWBI1EP6Ul5AKdvXAX3dV5gDW1eUIzb0A5OnDlVeYT0pZ4pkEqsvN90AGdud1X
VToA1bkKdugR+r19j21IW9VbCDHPx7ZEMuemrQ7/hbiPVugDoxL81rShpSt3Lexwq66dtHyVz4u0
G7ygbketKlX+ptUaKKQP9JZKYNdYh3E3vun0jrHWkPmus5e23x25LKHMKr7iZ4D5XM1CYswvciob
ucbrvw9XBI0JQ/dO5mYuIMuA3na1pQD82IPT3sB5jAuHH1QJpNrhCSb/eKImEk51Bkbzv1ihg+Vy
GH2mNxNZLPlz4qBGhu8NXmuNT1JiPjw7kSi5q4hxkSUjhv64bCOsJm9m9g604s2uynCLEldPbx1v
Fwd24hBPyrOpqE+zjpBnCDZlm1zfGnwMiPFHRZkpp9ZnKPWfbqqA79Vki7bB1XeYFclXRzt79ZL3
W5Ry6YDCaXaSTFmta8XdoovN9MrYsDceAE/hpuEcMRYTb8+peWSbzoUHvmsrHAk1JFw5app8LYPL
sf9cqdic6voPElK5wrXxAqzdPQZ2cSjpnnSCO6MZkknCU1z2vAqzO/vFTuKR7T30CNt0/DlMn2Sx
qvEOQpFY7T4gbR3iTsLzedSTlmCL5R1rouiXuQaljQ9g81bpAeQJbKusIMLcCw9ONcV70AHPrIEQ
u5N0Xp9hJqihtC+PM/0RHuSTvSMlNRdOxicgFax7kpkMVpMSkkMx/kS40ChAG44AQZ0yyBaJpHEx
EdigeXH1RaXlZCt5bJbvZ9+Z0kawEMswRCVngruZgT0mJwwZi1EU8TLVyTYd5cKxKy3ab9As79OR
hxO/qvZrF2LA2li0AQYNBtCNz2ul1sEZNs5ijmBNXcw0sVdREYIlRRbwPlbboSi+8KlzyxzKvENQ
5dA5JOvifgGXsWF5OugNhnSBegveFNLySqiZoUVBf7W+LdRlH70tetignXINByXWX3b2dXIuHQ76
WRcJo3X2p+lA0W0areC4JtiL8NGQX0wjHLp7xFIppAWtd/kyY5uJ+ShS2Psy0KPGcG0i/btddq2h
5FNhsi5Hx1WLO0/7ILjSV4J4SNxzFaUBXG52G+yuly83afzmvnZR84kMILRg5kd/P73480+46UIa
tYMftv61+haxKJN3iBz7CvkkoDdR1Pmifr3sQLE/k84Ewu5KHKj2A5fTpKd6WiCdE0z51LkKL3U4
BkLpxoSV4LFVWcuAz22t8aLj6MykL2g9o4ONOJ7YK2/cQPtRsRc1pQy5w/dn9ZHsMMWG4oHNb5WR
zjsD4pVIIIxh8vkdPRyjM4753EwwJDJHgOx57H9ELsPE16cDSI9JjrOmT0WQBa+ZfhH+tmv5xvos
j194Gy56/n4ShVvtiPnG09J8LfYQiuZhiSEHPCgWKBguWaTOEHAw20RqF3n+TJGIV/0qgUF8rine
fBGZ/lslzvTHEuWnzeW8cQgSKWwEiBK1YOv65W10EG4Ga6iiod+hxbu+85A7w2BT7DL2evcrsUJG
hu8cToUBVgtoyAGMFVNUwCGuXd0/7NHMTb4LULnYb7Y6vHgvViVy5yB31xb3Gd+anj1EZBmSE6ub
q5/gJA4SFhOB1e4UTYVvIM9cDaH5kGZ1A5xb93oQE/ilL3PAKfJmswrFAq0PTLDSApLqwywjPvUh
icr21HznUi9AuAehkZnqMmRHEHLRHxnSiaWgSahBPduLkNqe8hd4S+xRHA7dcll4o+lF8lTrd9op
3JfV7HuA44zuSmVRBc1TPq6TetIApjaezuuft4AzV7zP4oWqu9ad5wT37NCfYnOx/hv+lh8Mw0Y7
HgzVDkXp9TqnicS9yBsTlE4G4lW5C5w7ZKFVy9TWoJ+O+j+ymBg+PF/FRWdZ89ih9upiXgXXuhTc
nEl+rtfo4KUgGBD9EQLydc0hDFXrp68Mty82BfWtETKDRJpd0yFSHX8MbdDYBMri5fwfSK+BuKnB
AXdxGGnnA0f068PuLoA2Du+aDpbGXKUUqcTVULZ0OdlXn6R+sRJ6cXxfDIu8eQ5zNjNrh0EFXE3x
uJLqw9RcD6sV1qxsysWHxgelJlMOZ7/epbki76lxqLLU4/4/qjOjeUW/Q76XeDNUJmrlP9l/HJFX
Oa1XpKcMDVPwICMf2+6A7aBGsn5QVF3q6P6kMyN8kqSjm9cwzPpUisyO5SFlfE7bIrBeDZvQT/mV
ealMt6oMvw0qJSzTfljjhEzkjbnks23/HKbhAFBv6Iy6S4MpjtZFAuCALgY0byOxElIMBWZsrqI2
ob3ek5n3QxIasbAlLNnqQkSmyJxfS6aLNbTaujBpN0rr/4zA6lZMUsylR376yyS04oS01e9lmsai
ucnMjV3Y8ROftg0dds7suHcgwu2Fll25dDTxxAgGdRFJpofpSxMgOb9593y/+tMQ+WLpRvgqN3UF
tDq0mSN5/VUamGNxor1gGNGU/Sf6fX98bgS8N2rI7qoJrC89UGgSSPIjeaUNnrm8pOT3R8S+W7+k
w1IIcqKSyn6Uxoay8Y+F0PTnH804C2ucfJoE2I7u8yirnyK1HRkSK0y1yDIBce/iFLt1CDmR3ApC
St4wqOduiSeq7LhN3dhPLNtUW6IIScAGcDSR1Q5MthPGaIf98q3D8QUMYp4JT1AEAAFi5eZKL5F7
GoGkvzMyujgGMAV/lxOR90iVO4DOOyq9LXvitOw7MvvNJxeeZYdsO2SCYaltySPD0A4ikxO/USg0
9KAL8P5cuA+Y44ZunHqY2+edx2dMhme8+cD7CcP79rxiya11N5TsEfiLonEfxol5eFP2zCaSMfWF
hxLqRTWMP1l82qTja9Z1muMfrv+lpL1toLcKI9riaspLOH0DDgLO0VSH1YgbiUoSmye2NshYkDD+
TG1ByKWfUJnSzjrktwlHd4VHEvxO5l3kAxML4aM9VLfow91wgLT0MKJrgyn0UyCH+q5E7x+Lz33o
XzZnT+bZze1ngXfOLnJpzDGdeIzkPvCHNfbROpjV4uUvjvrapGshOA+yGaZl1YUm9/wcD9XiwfXK
whOtBr5KHb6rjXwiRsyBX5jt6E+dDDeXHSCKvY5TbavdID9jCySq+17ZSabDkE02Sn/sSBfCRwQc
5IaE1R1aL8yis+wELHkqZET0Cyx9xgDTqQ27oTkOK93lSppDg7n6I+U4RiY1uaBWnWVUQz7aI9Mo
wcZ6zvRNinnaNlnuPahzYSmK23JwK0XbhHTx6wH+4frGbjJG00Od17dtLK+FYCSuiZz4fdpkzcBC
D30gdsJfOyWDvvEeoi2aDQW+V9QmYoi6QOWItAXYTiNyQYFQ8DaGmrNc8iuDlgy51BqYVzRWDZW7
vtmps6R1shVil146pHXXn8L69D79Nmk2Do/1BRu3NpMRwS0Kl74nrVbgduPDF7AmOqMpiDQCERbR
CWWMC9JxGbJIguic5pvuX160OtkQZmRHLNfJrGX6XBNjIJMjYaSGbteDCDwuSw+KNaGepievNAic
LY7yMEYxBiwiG4LDlsQ4GqTutNzrlJwubMObdTpDdT7/S4j9y84dBMId+12wozd6K/NjRdBcCWd7
GtYXna2/YCFGshmpAHDQvECAGJ0tYQtmacf3LKecpdxukTuAIoJaVt4lqgaB+TWtVInauly1A3G6
o99jTEOOxxpkIWMr9/EfKg6LHQO+ZfaHFLONVidC3Y6rUPzTCf+aU9wXTcAKDyS/lF17r8WIl41d
kSUbYApTeGz4fP4CkXuz4Ey/hTDREkez2vj9THXT/iynvdc4zI43/4pOM7fwI8ZDGnN1tUL2uX0+
TI+wQ+8acyJMdBAIxprye/bbiW/9gLTjpZ9SuV++EHU4TSXupscn/mSvjBECBDmyfF8b99wOkeT4
CPsicmXz15jZj5DJs3q15wPiT8EO6A7xE1MVre9sCeAwiN7u7ZAuMAoGz69eWN0q+b1bO1QVK4/O
Mj8xCu9MkipgPkz5g0eryAzQrybtqFFKZAibMNVOwVum7NNS91xuq3AXgAJxMaRjfvH6nlG0iG39
PxAzpsNHrjMTQ4yzpt1zrco6fuBWSzGP4ZFGGJVyzVrN0tcSR8+ZhIdzkRcHTngjb5bex0t2ZE7P
QhlbY9sDqSEHzBSC3c6AL/5iD4JorE3nSNU8NJ3Or13Y7rUI6C51QuoiuR4rQ3v/gD3mpGLD5FKq
LMjOUJyaIm4SUFHIoB0FMsRdz4sNl8QVjfN3CbNgoS0dQamHSz3n2MmrrdC4Yuq8VSlDlZf2IAgK
SF1SUoATzUqMubl2U/4cuDf0Ya+Lsg8QoFAK5GVnaJXGJchtYiVYzOWaGnObI0StxVwSD5jmfftW
n3pjnsFl0eftdJX7fuwiHbB8NAxB1i3UeeQFfSTsdViow8phsQ+jipKzcJheQeh3NxX/MXxpzQUI
fmFLcvahHcRMzH7klfUDTIV22UIaTRmViyCEqrwlYI8Y4x7v6uSBOpl6CsoQXN7yJpDjowmFoya6
RLrE9WjyRd1uSJlhMYIzbkQSnERYgbmMgjYzN9PXhABmLMdCJemlaZP3kodJM9gDslijksgbL9ZD
SN/kJ0cbD72yUo/VZTGdu4ClCXmIX0GblFgbE3XgJPiE4hgyxZ4xP0krB9a7Ev91RUmRbDjokjke
UUEurieGxWc6Ox99VK2DYKG8qRnWafv8jCdJ3m+J76FxMbzZQw4FrzML8uUT9NJLwWigDT1J0QS4
B+SyzfvA7PjSSqpuOxVY4BN7WSLaiy6ebpYQHFpB20GaZoE+HpkvYCzm6L6U1t6b5bXJftDI/EgM
1MjC0046DFbJWdIplyRdriQTl/EtpSuBaHyN8ZMFArvKtI0Eh5chyNVgRZXO74nS37C+GEkeTV6K
DQDWQMw7lHaBFjWOef3rtbBeZVqGXzWbCeaK3z+JXEq9qgNAqWgmlQ92rUZYfT2NGLjW25DdTIK0
CrRFQVVCCQAEnu2P2/zgYYZ6V4KIi2m/03ZW/GrI5LZ8yFyAqravSJLumGKGC+62+RnVS1/f0qAA
oY0ufQJ9+jYEiIN+8Lif4atCDCoMlzJaJbm2lybC/IW06lLoXOaFeNxAlX4ve/EBn6LD2bl7Plc/
HzI5KBn1af0uKfhfkRbpOY+uBWjJ8kTYAj7KSoCAd+64njOprBkqOb0E82XdPVRFdnlQ2/gbZmNH
VB+j/3hOlNpyoyL4ecQkgyR3UwEI0i1cNmplIFrJ6MQu1z8MaXkiwEPdK254V9tWus/YF3MqTR+y
BosKrANtQqnGBQEmub7SIH79u15ge0EsW3oMjqA20Vmlws6J7cF8Gwf5vEYS3gv8pCioYPAyGYOv
MGb9FBHGgkC3gVcXQDv3+0eQFOECv8xS1sV81gIMNuZcoPM6Hybmv4IpTg1X3RY05Iz/eCLb2dWV
hwiPHByYnaTXufyT0DzXhaaBEswIX8174SjskwUMHyI12zyVmnqBK1nGfYqbgxPm0Baf74dwBSnL
fh2foMT7P3NBfPfC5FNfrIXmyqBN3IQbsNLdQKOIfg2pE4vM2dffH9zGqCE3QqMYrpMClEPNz0Sc
yWLjQleh84uegl+m7LVSD2BTFF8aDFWfomD4lvaqw8vb5oPFIqc8w0onh9RrLR3iCIxrGi0rqVch
dDQJ4lZJKJBi+AGVtuQNXlcZ1TCnuJOvScpRHskw41GeULBWy8+CRNoh6gdhDjs5xK8ZePpou0JK
oeZ/F4V2OmU3SYreqCT4c5GIzjSwipGDW7GA1K+VtravuX8DnYz3HNxXWtMyibjSrYVvydTJJdTo
AIUgYp8Hcd4ABfyeyfhOeqdnPvPtX8XYW6+YVDTkgJCkJcIkUq6xJXgvqMvlYrsaGtkvCuRfA8tV
8C17yunu0ECdrE1p4aTQQUx5VhxbDN4e6JwLm4Y9SveipU1B5QuQYqVux0j0TbfNMCHShkYfMbW+
fNmgxSylKnhShAdHctZIJ5ySgeS4RZstQHCwtxUZoTAO6tXUnIilsRMXkIrpFlooujvyEWYi711c
NUQRUP3i7M2d7mzvB+U4gsWXeWHeCFsWTxJAb/hQn1TiIxNHCMKGszep10O0SrLcYxCBdGUc/sV3
CClqIs//YjilvUc/t8U2q2UwZhdDdKBtbNy35XHMGfb0wfEKgMBodvAGsvcYCzFGpA/mxM570Oe6
Q99FIl1Uolf9aa4Jjrw0W1/klH/O5DHgy4SAr/lT5+lhQ2iyooXqcnj9EftZrqLLVdsYSznZM23h
uGtZV7sm/1wwZYe8jQFv/o1v7KpoFHQ+xZFEZsO3CRXpZfYTawyKSZ9cmnNfqIrRfwvvfjqrMh/E
DPzsSqLDyF36G9GE7YM+KnYq5KLAH9ZwHU0Aj33ZJVQrYt2Vn2gG2gMlvI5SoUBzj0p3L/k/WGdd
pLlWiTSpn36ui2LvEWL8cJogcXh7sJIO/IohQhGFYaaQWmVniCNRzgdOGs74v+m9C8ps+ppfKzue
78o4S16lK7SYPEqiVAStf8x4LJqMCEoUR4YYXKQx8rCSvfr8qWBhi+Sb0T6uxbvfAt/ZvhSKZyA/
T54Jvr/AtQwrwcDe7R+u7ThndHWK2L6JPU7ZP4RBJ3lYuowTGak3lQirFcrP8GXxmDVyuToZGZi7
MBZVVRTQoZ0Sl/Bwe+fXJKAQKIbhardX9+O3jCGX+r2tYOs9GEwT4jxTHTSGfQ0GExEziHOXPL6I
QlnhCXoVENxwKz5tP48ECSHPXkzeIfJ42zjistC5tf5jB2nwZUjNlzn1k1zE1LJfwUkxYxU0OAXV
tTDmIs935CSDgmdGX0mwf0+cfPfGzvI95HyDQXdx2m9tvHB1h2BGMsmb50ZmscHZYe12oozitYwP
G+8Y3obw5713HP+Ab1g/yscdxhA8g/Q0rgAovTszYdWtU8OI4q/F/pITUkpd8XLS7WUyuI8Guhjz
tG7QkqxAt9v6SDSepOHgU9wPHrMUHqSizS82TXoA+dvrXO9LP6LJ2bkr1h0IDgQFWpGAjJ87egA+
JqcXRE3gnRlQA1pyhQrvtG32j0ffTZeD7vBo/30hCtjlSb4qji2ewu4q1dyR+/c4psrmAuiYKql4
iZGg2mTlv4xHz9h/UDAOgHkc/h7POFyp9Sjma3F1op/0Rgzq9yFMZvUeM0KLBo2TEBG4dI/fK5hK
IPRWtoR3m/ldF+gH5gLmDZeJxeQT9V7FEQ3PYsYInk/C7QlFGzntLHwUvyaPXiaQLl4+uETX7Bnt
Z8cMLuUtxN09nW0duOulQII2WmW/tHRQ9Lhdh03iqUwVkbdZ6xN9ZAQTe/9fEn1uvCMPDLeHHRfn
RnVaKSxYFxCs4QF6aJ+cmeC0vR1DIro9iCK1BP5nq/GISgHMT3O3HzSP+nW5VJWpkqRwxGOAOVfi
Qo9GrZcwICL38D7Bp7dLZqVcf1QN9J08nGcAmPuizV6yFyyyjQ78q9m8zDnLhKUhcSM5Riynj3IG
lQbAWoYyQ6U/HoziqxwOK/xQR0TUbE/Tvl6H/guMHw26Cj/knLhSUWieiwYzl276ctbdHdiJMvBa
TY2AyOs6xszgi18jI3lGc5pzgcbuDYzOypoIHqZi8wMujzzhTvxDZb2NFFjHJABK2OlElAAF4XrQ
Vfxf59MSOgbDy6Xk97LeezOwH7/ueaIyersS1VDR5owjTWSdo6uVyzL13Y0TL/NsMbEWH12fDKZb
bKDB2zYZjM+DNeb7+S6lqIMNoUccqoY2xqd2pz9uH2Tv0993J5h0PERdbLKeGnGnW8gPvlX6pzRI
g9j6gaQGhwgP5uH+9SdD5XDFKpYFX3yPXCDuTYwECLRBy5Z4o/NkZEUnQm3ybemON7J83ObwD5Xv
/zgad5eEjQ1+7969HQ6vd4bPmsGtFSZqNSzR0q60EpWLqV1BkN1oiQ/YXufo3YuNicKmudIHVT/8
e0eN0FS24w264qd0NmKGbIVCLSCuM90iqz4vzSaV5CBf4RVo1yH6z6ReBJVACbj4v1acilXdZ0ja
cMSyosZ7YvvCwoOYkGMF1RaeNy5jjmWylbMo863kO7/HbremJvRsnwu7AMDf5xt+w33jaSCtmI53
vwTOnAo8vI2vQK8jYFXb+c+olCoEn2ipzyuFFUQdDjzojIAxrj9Lj2K5S2o4iUuCGiMbo/2iJPhL
HcO173iRKLV8T7fdAymq8l7OULWrSsiyhpMOTK5u5EP7k8oB7gthcf/EuFeryL41+kE3aTmyt5it
ZfXTxvHropAwNeFtAUw2SKYqQ1eTEiuTqjkDqwPngzO55/bvF4eaSCpYTq3zXuJUtBLmt1SGDTEH
ltmfhiwA0e+ZKnxIu3ds/qrLAMy8v/611AfxQKMdtI1OAITey7xk1ErWtudRm/5AYvLc1T7rI7Hc
PhBapgcTbUq2P3LPCmn05vQOqGUVBGoiajvjBoeDaS2hzCANERnawPmYisBhoRC0xX2MT2LxXmnb
+J1kseg/aMf3nJbl4i0zH1OKixByTpe/pioPvuxSm0Gu+VdJuJ6dwtHrV5U0VchUpkZofqzAhBjd
O1ZBq4F+aVBxq+lZEFHuIF6Jsd/pqgBvBUW3+NiXAuLgmojp+qy7b7zUo4FQ8vR7JfFI3kuYJdXq
x3Dncm/z5XLlI7yIqj92xgHEAWe/lE4UlW4+R+7TR4Xu528pI30TPZPMLeGc0zdNnoYagzjPmw+y
cF8BYs1ekhD5qIjnb5ycQMUPnN1d0ZFohD0+uN6x+J4tL0WomtWjgXGMOIRUdTX/xQ0D1ve7aR/p
15/BGijaU/P1VfqntJrPJWPyLX7nc+sT9c+kVEDP8pbcRSrQ7qE0gDiBde9JbAOB/mufi3/AxA/3
DzQz+zexnhjFrz0DUPJGZlnQk7LXnDm4I5mYXbFNYOKMyFNKA6FQnm53HxdebvKs4MHSfU1+trKW
NHx6+hf+FOavkq0RWs3Ds1LFxHgsvH7v9AKDQWPrc412ZbsQpgpP2nRbJ4rPxj1sj7EmjcUNKOeo
htVXXP6Mq1FZgQGgkys+l9R4QrzlPOd+kXWG6K4DVQ2jQETBImGWnRvh2oU6BieaFlwA2/7K84BP
QLizrakMDVT0rPEDs1IPA4+ikUpgpYMvlpiTXcXEzP60WIZwdgJs8PZ0z9b0rga1jUHNuhVYhRJh
KeJPME8auhxwM4c8MzdeiA2h1fCJoIw+xYlKzz6iDZKZrz1ObHTzMpjym+DhWGtPh9lnx2D+CaZR
U1acVfl2nB4SfW5CTyo3X0PsGd21yvc8DTwcRU59+e5kj9Xbri3L0/QWgEMPGRnwyUizu5tjZBwN
tlXZPrHXkLv739E/miBFw/IgBrdhHXCa76Gr3/9l50lfFumG24ljCCULpofqCynUfTySZfJ4JbE1
GYF2YxGpFJVPN26xnK8lp1zrYU+yaap4i5eucYvAJ5weAIcMm7f47SF36Y9SzBkNHchgsTS+t2od
bIYhS/AcfvLQxPDY3is/8EhOyQk8IfwyjspMvZoV2G2UHDaHjC10PVp27nUN/UOE0VmHrCtb1Def
PQIiNPcY2SmQeBtTiUv1tFerLMqwNGOObuQJpf97C22CCPUxnGR+ap5cGblAwT2UNA4lCEFEh+TS
zkWeyaIRBclwy4DX7psr0H7WVvKgVSeFA+OGlRomp0hF3vgtHDRlsXbhqg/ERGhJfR2GaRgxa1zb
zA+hGKX4CyQkZKqUbqmfmfZbcpjrfREdLGoj1kfrsV5N3/6LfmTb2n/V3f+bVfXHsJnBjedhNTgf
uWE7mNgj6rMzWGoTlTTpI+cWQRXjO3TOwTJ66PmMdjaMbSqbEWOdMsame8jorkR/XHvryKMtkElF
nAY/GbS/8sv7P014qkqYmDJYvvNWjYJa3qJw7MwDPVBa1QWvhXnS5FPbKFRbhRFD55Huy8GRr9jQ
YZY/ceUjEOprEF8VJpD3yiD7DAOqPGh96FhTvWzFvqe2wEktRgD6VwyzXCL0pdyuw4D9tecmbgli
tztsZgwLJbP1YMNnlAlMYdswcI0uN4lcF0DiykcPcob/e7MK+SUDYRCPA8QTjZsgJVPmDcQpjuhc
dg/PVRo1oh4v37DL9XLvzz9cpHslhUQ6Rmlu9UfSuhpuKb10ggGjvIGYQiC9gmYOXWMOmTP4dcup
AtTftZYGohgXROs72Ggcp3jfHfSs0iLiagNVR39y+t0q1AmDeFVV9hPlIB8wsj60iITIrK0uBQWJ
ukDFpzWMcPHaQhhKjBRJHnCMUHHw43fxpSE6RtJJj3LNMEbqp/0bI8XJQ/a/i277MbGrBqSxe9Lz
1Ok4S2NLLOxcmcmTn4AHQOGI7AAN8cML4SOdgsi1GLzGDO6+fI2SnReenok0tghyuEpueoshdZ+E
IQx2B5gT/ETpPCB/CKEsqeZ4jtK7+P7bdD9jmhbtu/FNjDd2/ijf3ZP+KhT697Ot1T+omfpazMK7
7a+xj4Q8TSA7VatdJD1tzZfDVqa5xThhB4aQXV+ZV7DtMHo4e2cKg2J3Z92LHDtNv3AVbGr+3fGt
okU4O+8BefNZ2YyqA7Punb7PhOipoYKcilHUeQsda1G2Bn8gnTvT5Ct8ifOncnZi0u3w8FVK0HxO
1GIE99Yzd98brFoLcLRVld/nHA50RgEQwalH2Dn+6XAL71PnIVnCODkDGrNpDj6CYZuR1rtEZ34X
UtvUTNB9JpIPIc93p8UL2kYxQKNf5RD8BcMrQrWamh2JqVNLJX7jcoBsla881RP/Nj2iBCLXtEXN
Eoug4ZL9VfMD3TLOiYxEvdmLBHQbXJSM+Szvdt9DjbGCpwazapne5j0zWPrhVKhjHyA8B05rguE+
12gCfY+WUj4FlXmVPYik1z9WD+OEbYcVfZ97U5E5zIhGI+wCnJy03ekZzIqOPS71tfw0qyheelNA
kpL0LQyNoVcFjWEg8h/Ey1gK4n/8UzrNrICpufoe7+cHQ8J8eR55lVPUna7rbnutSTpY6JB9++BZ
W6URTnPjRUHWRpzSUGIk9OH7v4wqBzsx73hYeV4GZMHR48Jit0CT5RkZXrOMigGSsGvikGZ8Yyqc
xWoykey7UVBrJm33VZoeRB1R2idoJMFXjOWwpHQGpEYhAbN4HK++WWEA3Ze1otdk3ZjKVmje3wuB
RZg8Y7+qmQnyjVFVfvIx+6KsM96ixJ7xON9jdHxtnKaDkwcpB3AZfJ9vbcuC+ifj6Bd7kN8e9C2L
DHUbmX1gIHp3QsTd4+LWqlz60j266AWtNRPhztEmoaSnAyCnyaJVytYTO8FmYgEzRi78lMsBBY13
Rgv2Bi5fcFOzXqJR90VzcTyPMEnVv/22RORTU2DeMiq13Xcqf+W4HEzI01Gbml7Gtq/SaFGnZ/8L
m1AVrTXLxUFwt0gt2Vr+YroO5sFBJl0tJoH3AWYCqxP4Mr/eFE8ngNv8jEcYDcOdxvQuMPDlPTP8
7lx6gDjwKszl3UsfEPXkaXMcoYR5Hjv4bwfrEHdTm/C03hEGOmIu3MQIfxqt3GYNJqp443IxF/Jh
uknrOHOiUmRuwFmgyalQnir8hjQBdGr+kbQCuri9arJgj2uupYH2dZAYMNYcKGmbacw2yZL8pMf6
IsDmm+JFBccWCOyEs0Sv8I9wOQU82/MuqXcdcoMU01Hjhi4wASB8vDkAuQCjpa13GTAhqFD93Swt
Wa5nEaCfCBOrHi6aQ0Rn2rC4Kds7yTcSSXZzf8miz6NXYn9VxyfZS9W+PBjsC/Rx0q3EQyhieg2S
jGlipCrTg3mQ+BtvIFExzIjxa+YEozEOo6LgaG1y4BZhLzd7vACc5LKpIFuBS6r0KmXKDsiDBfI5
Ngcplh+jd+/GqcEjewPUhsc2hM5ZnuZkgmnR8hrYNDXLv2e7eYSX+ZD2IDO5FCCqnfFzUo9o5E4p
P3hicXqMjlf9d9FOrCihdtd+ZKki9/ynnv1McW0KPgSk4ce7HeUt2s6+pecRE47CWi92EriioasV
4qV4Or5crN+qhjukbQvv7d2tVaXIs6U7I74uljvy8A8Kxv+xQJd3RYBzlpUBLViadLnYi/R/yiif
OuKYNoCxXbMZ4+/madd55oGfkIOrBbkC59gvsIhuUNErCNbl3W0NoQt/YqYcTm4DR7bdZEPPfSd8
eLsNOofZaLvihiR8N97nXQtgwPCh3T96XLsFC9aRjigbM/W+afqKpvPXjZqVnm6MiVhfDH1c5NE5
aKY+A9tdpSaufvtvqu4v0cuh5VsQ017NGopsx+GdGrk6YSZ7A2HU47WuFqft+W8SF1jrQiR1ZYIX
WdQixs+HWVp26eAWgX73UyykfUoZkiIDmMPnprC5devIQ9UDsqkLc3/Hq+q+M2bW8dmsqix70VH9
SW9VqeeTYs713Qhk6ttnW/00Om8QcUZ5SO4I+y+/9Ssev/4GxMkaCd+mRhPb+PMlnHTFiN2pTn2P
d8GK20EUmLwQYJVyU5Ej3AT5p9NjdbIqZiBr+oKjFOZ0UfeSx8cQsYT5aw6bAUed0yfmcWscnOFi
DYH6onw7bZwuBc2T0vEojfnUHdcnXDCA8WHBl6IOQRnr8YLr/A7eeYo6LbYuVbBj+DOb1jYg5Xhp
LFwxa5BquJ5nT6tiHORoEIFHSzJD+lY9H0tLlaLFU5rGtPTpdJD05KJhiWe9Sm8Wx5LM7/kig2r6
+88/dJfGdRdWsa8KRz7bYL4B12RopTM82z87MrEM8d/Pc3kCWKKM+G58QWZnjDZOepQvEzT5NJSI
oGPx+CyLUEgIW7oB+84tHuI1+OLaB9QaanukB6pT/GGtKOYKNADnZBYYHvIJlq+xZ0jomcFrbwEf
R2SX845ZYRNd4fppDVqzE6AmAyFrmTE5zBy8x669P9iEtVpoxfl723051LqdMXeNze6PkQeSLYr5
c+jSxMPbVMusxCZc3U4xU3dtpp4UBEF0IlxHKla5BvLt5u7hjrrUtbdlx7VjfflCaeqeIAvYPoEG
UUsS58YeTjp1KLdrgnBX581CxH5/MYsPmw5vwQ9Mbcf3CuqbuD5Es7QFUfoxjpa2XFRfkdoRmqrO
T83B4ZoONm8eZtOS3A99x1VhV68Enhec1cKShYqcTRiNM2VgYIwTlUqZRQ8521v0RFdLvGJBZgbq
sICV+k4bPgSLh3dPrZUH/XJvVxQxmPhi9njj14xBRG0PnQUYCJjFOuZfwijm3MlQUnGhr9TrbLz2
DhPFQG6rFdwP5W3mEbvLSX1tzOeLJmxvdHNH76YeU3iYDNoCQirUh17ByZvjKTPuloBN1DHGV84h
i6AlFErQNTp3P6Z2qr8jXRcQq5D0KatxbPv21EoXPTae+JMWvk7h+Lo0rvDpjaP5wXPvYTC2T25p
AekucNiobGpQxlgbL+xs6cMcBnWMLcqbUprU7FURnrGPjADCU9RK7bcuboinlrXmhtqHBe/rxktM
DG+kotXublVtWev9RjiYYba9e3f1ULy24xAnt/6VEqhataDiin2d+pu5hEoNGEfJFAbzVi996bhB
5a69zEfThRTsyOXhuPU1dLqY3LZjFcshjEierDoSlQcYytk2gsZ9pOeD0tss5RM1UgtihrOyXfNf
C+4gdSPVtD+IAqRhcErC7HEy6dblkK0KxL2+GGGomvqNBEfb1XTGHvD9hWHm6Nu3Y3gY78X4fUSW
8KbPOKdrAIYADXQsnvRWuREtp2kGQeAmHO0LkWKFOdWMhLtaJ0wwnAdOWKWveJ05IWsKvP4I7OlV
HIIGBkZmgze4v6Ax5eXOLreDexj9a7/UYda6ZMiuClNxhv+niHQaYMFTCgsQNCjEvp0SXHS55ehS
ybQ8L5kfwQgGXMNLFiq6v3NBIHZ2daZ10eC5IEEeXsegpIRVbgPrV8QE/LUJ72s7Ez634n9Lu2JD
qyQ+JtelweIn1zzMskdJiKmYAc9gT2p4tNrkUIPW7cmAwfIksYWNqxSrKL5KSwZKIhNpdUIUtlBe
RRK+CoIQCX2NHmt1qmfroExJwN+o/ShfSxi5bTpQ37Aqt8zojw5Y85SdieTTw2MEVSM73Ipa1p36
lrbRhXQxzvOthe+rAstWlXSVxcr1pmIj5AWw+MuRmeTffpfiAVAMSJUHbIULpjv3cDouJK9u+tHh
voH+tTLFOX1rg6VfxC3ZeMcfaz6gcwjP2/Br7NbXNmYbDiU+cVQjZBNfWvlGNHVU7YB+AFBbxqEP
GCcE1pEPoKrm07P0sQpUhI6FvPblobczDQa6VlXEaBuNRGjdObrqTSH0EdOezfs+HzrvMCC42SeQ
2yExYTHe9amo08EFtGFCMDE9hS4Zpf+Fecbczl67VipOEnIptVUgOajgmkCDo4N26TR6XpmmWmGq
bjhOhz8nQIuy0dZeV5Ru/5NsfPvtzHE/6EbKKAbPbNiy9o5OqMqPbUdnLtJwm9AIEyk0OiZmsA2L
Xs0Q4jj1VjbPHD1zjj9dFP7ebSjgKSwDfi7cJA2NQtPN8anwf7krXglXGa6N7LJKnUXBV3uAk+8u
SbxqAsoi48uXqbbQ+sYVkUOsLp5QzNpLpf1XlKuDr3ntgG0gDaoI7m/szVrrmjYWC+wxZszvUrhs
GIB4VVL08+v/e2gNBUG4H8yHOWWguT0iO/fI7fraeUhA5MAUq3k51sE/QbQhItzd54gUpRMLw2Jn
gDchwH5p91P0tyMTGKtMzovsEymOrcH5LHFC0bXn7vDjTOJ5keMoNgNc/M2wglgKuEl7D7q2NuVC
5u8RWgYD/SQkwqSN47/2Oa3yGRnABvqX6pnDXukBQnNc/VzAvmu2a2vGjGNVV9ODiC9iSigqKf7c
CAzZOMmhmOAPcDGDtvoUMTXE03WIYHf+TwVNkQ5br8rI28Y0pvO556zw18pIhTh/Jo02cf9RTAEd
BEeeMP/qJrNrYT1m2pGRl5OoEMd3qCQjBeeNXBRtcUWll3Tbca3gVsIpssxeDOlN9uLLaNrBve/n
Y1wwzRgd+7Z+HddyYcFW/38YZveaS6wJFxTkF8ghJDgXtJ5iuk+4a+sAWooobuCoX88trh1SWpZa
RexNo6yt/KdaQ2WyvQTBEHCoIeoseLh921Ngx7oMYQrn79tEsi70EvXncCHkmJf6BshEAvOG4mgU
hb55YjCXcoCaaO4OiLlm6evnowxNNzvL/SYgCHMGbAY7PPE1IcthqHxHJJGHBYhz+wngaiq1k1f7
pbfSuNEGuxuBaFASDjuca38pbYZrj6qhtAs2d9TNO6SEVhZSzxN/NVRbmy/ohxJmSBt+rb5pcxsv
BsvK6OFp/JgY2PnB4T1pv991K0MKLV+HOwbVW8lQTZq0S9PcIJoe1A8qWleTMYgF7E2dc6wgmlPG
IXziOSxoaR8kzZ0XOCqGaoo5vAohnapM6NUOmqVfy4R0IymhsaxXqFjl4fscKEM9IcExe20NMOvB
yhghgBPu3cUDwSsN/JOe2WS0P+i9o9kTqWMztgiLlt67rpJC+W+Ao8Kpd1GpVvxZUH4M6NF3sDxl
WrOMuEE7Gella/ScXD2pwliuCXHh8UMxptmMxpTUiK4gFydtHaT/P0dyCZXygZ7NwyWKLs3FFisR
9LSARQXyAu4iDpJuHROGFWNoQlkQaD6z81X59kDpJwLzfspTidARtaC0PBb/CTOlE4ON+noiYVc5
gQzTLAqSoREOdTXlVRWey4qHchS/jMO57DMhBv9LOcupLCROcc1SB8N+l10eJi28v3Eq5cvvXggK
gszYXEyYOipNs4pbk6GivmHCDY5oL8H5/h3TdUm2K7oDHueqaEh9H8kZlqEGxiP6lg+kV9FEfuKv
O+mkGvC08cooFBvV8Y0GkvA1eE5UhFyLYCBZSrEryQq4e5XMrT8I+V71oBZCNPfJvL2S5r+FXY8o
6YrDa0pd3QRlUOLPc6ZiZp9wexO23HM322NO62TAtHde9CNtBRF2lfHdVn7pGPVT9h9ME6z1mlPn
mm5ZjSZHnysoTRP+T2GUAxw9Sju1dEtwAkg73w7dOHuLvUbaYzn455s7G9SRkL+/vJOZW1vvMb/3
j+RfxRfwYG09kbBZL/kcqTdTAcNAIrvNtnZxQcTYZVLnqB9RelyF8JiwSnNQV4ucxDsrKFFMGMs3
7On+EukV59AIoxWQfhE4tOVcRT0QMTrr2ZjZmOFU4bo6vXY3Tvz3p8EUwyt89awnQYr9SPylBD0n
DVG7kefYXV+QxgHmgqOxrD6JgifHPFnqtMKsAYfuQ2u+wK44Gzhszm0iTZ0SegobtFNBeG1bjnCK
TDHR6tzwPkzlIzBSZSzrOYyAAEVjQu913GvTUxy28sGMqIqesCuk90TzXiL6dGZRppklmos+vvVB
pz6QMprAQW5A0m6qkcFaz+K9ldIuuj6Nd+sXC/JQSo2V5tjMu/yGk2vzSJG8q6gLBjWjMQrBCkez
UZhO5R4XmSirGhErjlckl1oeyNDuTqndZwcqfJzIwKs59++iheRoKtkRDgnB54KsP5CujS/nOwiP
O3nJ7ktbTbq1SuMTsJIldc5OavVMW6wuWcFvO5KJu33BQAqDERbEqhfgfoDc2QbkmxoaOkxE2EfV
5hwZehuanGWiXqj/PhgrUZ/wvArmGGY+kD8xKWbZEWig1ass0kCnnLJaYB0RAzEj9xOj1Zuta1uX
5pfo7UydX8UyVvBpziOFepKPgB0rlBO+c7Osr1ZTjlo0XicY3zSu6ulTMr/+Aof6sZvGkWrAMjVz
1Psq3rkYcIFXp2dlrA8I4jRXyiN+7jMSFGt5IM2eXdu4+69I1JUfW5QuugBDFguM9KztUfPibAlu
qO2uWbreB3wdVJY/zGgjfKMRVyfLblyG0WEBllyLTyux5o7kFNMmglTPNpusae4QoXThWdK9cR+U
g0KWJeeh+Uk71rBlwWK6jbM5oyHFFwpB77ss8Ps6SDnSH3knpXzs0h++qFWP8PQjVRNL7LeoHs1R
XObRa4fZkG7kIvT2MWBuObuE0WNpUpeUy6auGcKVl0xnh2ZTV/qH8EbaiZTTuUb3iVODSVRE9aEL
B9qdO6lsuRGAPbo/f/K4oN/0nPXTZbwhd480pJ4MuCInuOBDq052Nv10DPI1F6A1KV40irJNkO+2
XjSqFsWxJDp49w9cdFKA6ej73sY0p1GXW32LtsNJnIRX3OepTjz9CXfXxTRzLDjWHHr9NrZpHtMq
RtR8U4K3tPLcRkmhWuR1g3wZBU79B/DOWGk/yjU8cR3qMbTBgXZEWf//faS1TNiNmYQYaKxsPkjK
LvPDFKVAHg/w9KuPvVILayXFYDuexSK95OUxeOxACi+w1Y0ZgHls+twjfxGVWSLiF315KDjS/Msz
GMhG04wqiEbaDYFRGUWjq1XAmCYQrTqtoNcvALwr6R4fXLRZ+82Lat8PNh0P7pHGwep8fNC0O+F8
QY9UU0jzD+0EuxdlOAFpCZ9YqSA8ZjHAaPW2ey/3MUbEocP90aTXGRJ9be9VgNfuiqA/18DtR6fL
9YxsMkTawABXam/N065fdDP8VEPwFq0a81ofrDTPIoKMVPf889UujKhWU6MOmBrNBcxMo9bsjvGk
09/pBIpxp4FxDYBA6xG2UDHfzS0DEhW/LRAZQZiJW97o3zFKXatI+/yhGOg3Yd+izyipUwzwyBhv
CVPE7c4B7msS5DcdkPrLi0dubUweoUxPLUqUHDkFpA91rXWRC1wNlzhwVx/GLRlQ9ggFWBpBuaA2
E1cYjxx6z3JWnJpy3YWo7lmQDZ4XNBE4bZDwjMrBieKqn0cJ2JM9oAHIcbZvmKFz0M4I6eGt23vI
jAEiTm6PvFVz/LIG2vytkgL8cjKpmXPhM67XfxqvMWm5GvKTxTI5vV921tqvuN3pIv5e4zywUu8R
tDpUcg1qgbhCi3qX2wAmNZdPIlt0Rvx7uT1VsQS27w4H3d0zhfKbu5vqQoweeRMXXK3cEA0B8E3D
eBI15Jg/BOj9VLfMA9Ooq2DikjPjxWZuM00xeReYQ78OMoeBu7EZssdnZAQVLTyigp60ukr2KwZ7
KTZjX0g2uv89fqeWflst/xoK9rLrziQBoewGaAQZZYvZ1QItedLAga182ThLoWKtdItfNMoQQmWj
4F4bKbvOETJ6EglJZtvppa3YKbSfwJyrHm3yzwEYZacNwLedyGQCoE4wgfLnOfJ6sz3oqTy/+/vD
VpaBYt+d3UMfTlu899WAf/PaihX6XNbVhS2TlgRhLEouUe9iHYfwcZl+cq3Krwznh2EET38V+owv
qSVywevi5qJ2xO2UD6T4OIMbl7GKjW3OCAXrQR/sYCTC6EH70VZVv3YejzsLWmWtkNDgi8T+Asho
6Tq4o/cfvRbegpBi/TrwmTi3dgLNAIQor9OivMK7vHsqjb64HtA/28KmoHanoEQJgQfyXtHLwtFP
5EjL0O44q694+muWnSc9/51/eAx7KDWbfHZ/mNz28UvNlrnIKpACeefHTxdsRJzGNM6nMs8QWNcK
h/EeoigrvDQA/r6Au+Ha5oac4Q8ZZCr9MilvbPLorWAmKxqX1B1RgEdEedP2nc+q0BeQfrFcFFTw
eGsP1IwVN6lWrptPCwPUZO9doTAnsreATrBOUWM2WxRValIffP8h5fFmygzPrmcj0msJkY6miKbo
/V16NmKm0W7wMKeSwd8Nu0gufwpKx8W6NV6XLp4IbQbpdOWdZ4fItNP4MIN0Nw5MC8FiEe/LxhnM
0kYcYV10eaDVRQ84oWkdkk08stpXdlqVI4tv0/U8uCo4DkjkOF6hAAVQAATfz3aWiyJPq1MAZie7
+KvWTVhzm057d/5m9yhxhM91hOhyVgjwpnYn52i5JQe1IWWZLtWPAGeBlRe0W/4Wt2II7wLvvvbp
Xs3tPGTubctpYIOjHUuVHqoFe0uojHhTbJS89gVSl+lSr2WuAtPlebAxkPlQfSJVJomutI65+qSI
jdMrKJGcE0P8BLDCXYM7aY/fPYS6TYDirrqsZ7La9R11KhyDgqeAoKqJxpV+LkhovqJgeKZjOa+3
7ZmDTqdqMuygItGvmoVMGGplHnS4w5whvzgmH3yzQk7rMrNGN0v/MfPHFRcYUbZw4fFhuB6UOjOW
Fvcv0hsPCGBd+kLK0diwIYofUZtxdws2QLwVKpiBsjHylQkx5K5lrj0UA4fO3OXJtQI71/DcaoCo
02mFEDC3R0dXde2Xqj6/NC45tVFc24P+kyshanP81rMMtNQnMSRnSMiivdjMuw6o+D3/ALqUKmP2
/NHojxs/70ViYW8dXmdYZK+eN8evVlccKppxbSr0wZzuCS34IrJrjluBhoDeHyNT1Kj0I6ZD+WR6
zqIhdzmUddMsTpCF2+eLePFonzk+C0nMnpYk2Jpmv0+BBz/VjqcAzQCmLWL3PCRPyCulbH2dtxxl
4IAPuGeZHMnquaio+MCH6YIpmfKtWeW340VztcFSUEJ8y1sc3R2Ljwxk4zPSmZWWo31XhWE/+thZ
MaJkk0EBuPSNUIiDlBMps/Ok1FnGAJ5rKOcCPZpu3m243aQrC7KY9PB15EsF/Co/CC0p0Zss8TUu
OCvgNVGfkna0+Rjb7ymwyDCWmnzN2hjdhYpw52f7qoG/GcM/FxEb78f1WZiUp4LGrnhhQNJ6bKD3
XpS75ZTpxxR7jBHYdSHZxf1/5/2BGQmRtZmd/zgx+7rVG3Hvu9qJKR1eZNw4+jbyHrbFqw77mWd4
cLOleFilra7tB/bfB2zYLuqU51XKeOl7Dve2BLWUX2KQdXYLaaWnEmWU6BHIL7QOZnAVtcG4+EFJ
InbJOIOiWJBi+gcATGPE/F6kh0SEm/I6rHvr4LfrHxBUfORXOCx+r7c7tcw5Bkl7DkW+RI9S9oJw
MbjL6pY59JM77wf9hgLah606I7uli78LVngRe+XfgMyuHMhy2ZT2/iLfWzLjZpeFhuGQN8CpAYQr
skAfGtOO/Wyyf0S7J0GAPJbEUNECz6Y93z2AfaPuyL35cxgGA+K5Hx1qXcNR2mBNkhVxtbrE5BCf
54NERbfV8NLdw+Y8bkjIJoNkRTUHqzdPhnOQ59hPzd9BFJw2K/9CFQse0xxsjZ/Mpl0WrWQGhnDu
I0gAULGEtBOMVtX4QztQaARJrudnXybndMtNEaI1c3/99ids4RmTrY/6zjQ/MxHg4Y668r31zItd
mixBpzfJNGjnkMXY8qr9Z+MOJbpZyxP3RAh6wFTqBEA/tf0KkInryJ8jB1IAYPI3Of6ZPhZuzTFb
GD+NPQrvdebCUGtc2KIhkadF4l+OsEJ0dEMt4Vll7xl5yGrdURerdjUlXTIrLCDTlGUBsYTgZFH/
wUm0HqUjnnL78dardfBSlaibBTHkU+IU9sBXqMpAeG+Y7AAIqjel9DIwAnbzxDLXjgX5gPLFEgQF
PG5YzTPP9xexqHF8ZlQ8UojWDur/sGJ+Rzc0OAt7a9AZRNyArv6OLNP0VdpxdpdXeBuoO8wsjIU7
gLnBsOIx7JUaZUndFM3OeCRavq/IbaPGeLdl3ch48gaTdXJDEIs2A0b6OcW6M47SbmS+33FUMQpJ
rFyLR7GMaLPlYozQ+GaYkiZGwQbZ4XrGWAcJfhslft8uurtMCXfVrQh45SvMrGA6RSnnsuJpricS
hbo05oMcW2RNbpDyEId8vK4uh6qQzspAu1nWzd9fbRMb9jtqx60V9ifhZSp5Tap4lx5EpSAhd7GN
WoT/mD6QT2UQRL8RaTd6Y+9oLqLJpgizY3QpVs027SnnBvgeD6owAEicv0F0AM1eGuYVCXTYXZHX
7IDaIWVPVcMq1UijdvZhclmdTyoWuebTRJxEzZeElUNnNrVjJKEPj2eWBmUfE9oSm/r1li0h3VAD
LJjm3xthV2inR67ADmY7Y03Qzwy41juh8IPJltsjOdwdIEioW+2FgCG+FFQcPhHDdfniiyu+4mZf
W2ef3oU93QZmB5NBQWITLwMYUAPve+d0BgjV6S/GtxiKiAUQUKq9XEtwT0ZWVMLG5qGhwRwHjGDa
flG/0Fev3x9kLlgLwxnCYljz/xrdteuSH1fFCQX4XIaSRQ4kawJscufsvl6sxJBKrvn55GZfj9u/
tT0QhvIrcYPPQTOyBnP7LmtiR2qpb/7ygtBVoTDU9i9m9vY4ixdq/6am8vTRmG9IgSgy9dyHh6Ta
IcUNkHlDAPP2rgm7awmwV6h77Pa0j8h6boHwpvl7muCRimy/HUsJNykgALrG0GPzV8UUXUSRsEAQ
ezN7w8oGUeeLrE37mzRspYqEoriOeoGChTGrbSNYRIlrjDMbDrS4MGMPESPi4gw0qyxEdMq878qV
xGNUF5A+nw0o8rpcWypQZsbzn5kvBuxLZiYJ4j589jFSZZdLXimMQ2gwbveuXESHme+A/Pq89+gH
23B0AVeVo3XbWipw7DJ+KvH3AJBOmNV+cezlGjIHiG4ilbNTwZwIl3iNVedaHIe6yFp1p1QDeaft
nqTeGFXIbKMmQ43YgpaBLpddKGkoFjN3KcUk+fF/dpHbZw5gwEQoNF0J4ooax/cQrsoKGQBysir5
9xzjTRw5YWZicghEJdICD6EtpouAJvyj1kn64s6kPItc5KljA7IYeB+AbZ5gW8T31xvva+3vi9L0
tqOzwdagZ6WTmlXspHevNy2P9fkW3wkI1w6dIC9hkNCQrUsnW0mNmcwOWxHbIuHwCEwO8c3OW1ha
+a/TjC+8VhjoDLpZYA1IRJUitk9eq/jN9B7YbpX4CvRNOHqof0e75ZtEMP1Z2gQ543IZaccMPIWH
RWud3t2mXauoJOKkZFIxRED73kXqUnJwqbsWLUN6tuLN3QMEfQGTF29cWAA4pHjRbbbxg87T6zOn
slYu9jKx23x7klt2efRXPlb0UNz1IPp51Y9+tgN3rhDENgHiCkNm8is2KFnJpp5UAFDuoMirDN3B
mJIp8JF/rynIfqe3tPLXpT3Ba7+xwqc1wL8O3tzPOhEMm4rUeaUaThkrQrFdPdTbPyYz81B8TtwR
uDBZ3hewGnm4Lj+/+/cCyR9eL8UjjPu+aSa+gXi1eJCrey2zj5lHjQ1DccHcppID+Wmc9AG162a3
G2//UzIBuNHTwO9P6UWWCRZfMeYTrj86mCc3ZWtRL/6JGnU+KfOLCY5PIoF0g+WBpttpUitA2619
sdTIrfp8juDsEPX/EE8il4Kri9PJGqkLFxt4UB4kcc+5yeweuIe1ALIHsJbW4u3y+KdJLxw0a+6y
XRHcdV7FC8chizXwXjsKVUcZRtnflqxBXy3tBAiqP8INFZGZ9/dDlK/2qVqdMT6gpAaTw5MjMIO6
j47VtABV2J0kaeUJxxpBgevD4Ggjsp5jh5kZ8p+GyICvxwzJFjNgcTba4U8Ec8PE5fyeN1aCmMTJ
cNpDIDwOdDqTBwtoxPTll6rJbnFHli2OS//qs9aBqr20J3DZYApYly42bb8ZIf3SHqZ1jLVwHGb6
IjQ/5cNFw7+ywJy+hcH7OcwcjMsgdpJ28D9WQZmJUOaM3EfRWODbj7SkMRJ+e9FdSgTC8ACPN2Kc
dSi78pzu8V4mwbfsgCXbglBZCx7doAI7ZSFCw7o83KRZCwtZiyVcw1buTZyLTijf+iaLwnJLVSbV
+wHBguZpUYMvAaCng/SYM42Gc64XSqrbtZaFmeaLicbT0dZccaTuYCjj4TvdV/cpfPU2aAGIQHDT
gK/SanqM+1X9jfkGnteVCoYeSTp3QM6naTzCxkRFz/h/HtbLkK1aIHWISza2sJP6VSc9vov6pafE
l2T5tThfuuaZQX/PSwUo5JSL2xfWZUC85oWnvk+Wcr3aiRCQLEYH+KhXAsz8YOD7Cz5wZyikh66g
9WzHc5BJpkPLFR/Nqnl9Z9s/G0suuIGruza9wOnSjdz4vgx0ILHG9evWBct0XC+Q+0stMDZ/mdJ7
/6w9sRsPrbS97AyVz3lVNlkF6ggRKbnCJeqaOT1iriDCGgUJVg/qqh3JDqftUTeNM4z3XhCG6kZZ
FwSm5tNAA8mKpxGifiF2XFqe7FLdXzaJqJ8zgXAybVuNUhby+3a3/gM1EcKaKh3gMEWxjCIDJdMs
OjigtS/v95+WpRjC9t3n5ADCCulYBRP2QR7Ji48vAsrmGOPZHnS6y6gwQZ7/Xd6SPIvWQnSWNZnf
EZAZjyudMs1q0/H/V4AJB4j4LhRsdu+DzxDKCNJaAILY5tBTCchUU+mpqyZAP1tjU0RFqomvdypm
SF9Sv+p+BxhJiMRJBrK67c+V3XNDaLPCF7KSmwcJsNkEW9j8tRYzjBe9yi4Bju+yChwsJXrxW9FK
3Ram+LBsW5hwkurr8p6hVBssnLYhw7LCLa8bhSkMn3ZC26Dt8FfJQwopwmGQYWj5QWOKJQEr9VQ8
hnH0P6XJJdZI1Wl5+YhtlYONJlIJbCxwCpijidY0aDYsjGTiN9D6vNhn3coiZCcb5kHpWcxxAmR/
eud6b7t0XxWUdixz0fBqSPjwPMb9iu3FWDYrKyPGEO/Zq4340finDPI53OR/NSvGzjN8H6rJnwin
iERDf7Tv3UNK0RjTHKWuzGPKX5Cryz3NXrhCDYhgbbBCKSdCaDxfi7jDcP0UF07GYMyitc+uJZSI
jPWoDyxWfISVKt43p/Ngn6TjsVCQBFkeaR8hWEhTs9FZ2gLke/Q5eKfHmnM9tw8ncukk9iaUbEG6
5b8TODqrRMlJ3uUfPNpXvVGi7vRKt/k7GDx3dFqwLpE0LDwjSuwq5kenYyleWaNzFS895pxQiIXR
l4wt1obG6dsqzgnA+0whVqVFvZa+9Bt4ZgmZUv+Lqz74F1ZB3boEs7nXgy9+qZkDu7nkjEKs37hu
5E8HcTZc5UGkRrpFXjOlnL9nF3c+s4yuA0Ua1SiXNz9DCdxgtYMsO77VJ2WmZGENsEtGaDSRwJUD
eyMVlLOgpmTgsqt92+hdUMDg6edDfGsIA04ru8AcLfO9EGn+qhdauFS8p8Zc8V7U7yHtgdpJWFy9
/o7pcTSeYTMhIS56eTHL+VRapXFn4hFYcYoJ9DT/UIoXwDvMBFW6fIPs3Og/IYRPxcsj2JLXNnY+
dOCK1IUHEdxivx7/dYa7qZWxsNn3CuPhLKfh6WTwJCszvjEjkloa1/ZezUQn4EnaQz08AXfX67c0
0sfnkeUW19gBV/TI265EWjnqYADOwYM6I+d4FRH9PL3wzxMW8BIqfXy/f/XgMZQQGBSI61/V+uFh
g9/OH5M6hgkYc973jgloU2D6FteVkfMBuX/cYFstZxX7Cfnb31DLAKU+OPsSbHm4DFa5ON8x2nDb
+2+yLl+v+/kw5BZIzdNt0+KbiETWwblbu7bUGDKHV0Sztn/R0qDDCE2IKbPuCh/CdfjJEIX+r6Z4
WBwh8BI8SxfVwAc7OOKiGanI2Se9+xral6Lt1ZALVfgDkaeNLRmoq89jJhX1q8cdp9gShs+xm9fM
nGVRDrSjC+Rmj59i7/xFPFN54ISf2j++4knonNCbyrXdip6+Ulq3oHNl5oqZm4aPBjiky+qsUCCL
wKYFuekTp0+6CetPYu7fBxGoQg5kY6W5L1sY1GIHbJqgi86Avb1DLS9ZGz4WgOIPQw1eTjxs+2qQ
u/OOs8m7wgAibJ6Vb3aec+KUz70vduhGyoNoXijDQXwbVavvytARFlL2Xr4yG8tI0H/xH1XlNcXl
kL5vhAQEtnY/OgWMiUGjzN/tuRmKWojHzzP4Y7Hni/+Dzq84ZsGtxlpfCAWL6z19SDvqrCXrJAWn
/bpgdUyxwGtJ40jQa11lubaWPTu8xbD5tCooDyZxqivu+YSg1ms/s4yEUi2SjqN/Bj0R4zdfvOOe
JQL4QY3vusa1LZR0Lp/9q/Pjf/yh3y1lKjAo+fJhjR5KyhTQCdmjQ1bzVFIpVlqySE6NuCulu+4t
B81vI49Dh7ZLTXLSddM4qxG9o4XeX8pe/wtjvgmyuJCXtAaoHt8ouQDGRX2A4Lp+fq5xRzx1dGYZ
Alkq2sEf/RdJfAhgBZEzerioKE7yZko/ICGFBBYYA0BMpQwKj+z+b4I4yZdn41AYmCGPw+3pn3CJ
EFxzrXPVt3U9HYuRXViy6FHVRyx6pp2mncZ9hIU71Ewm47FXkwmhDYqr5tQGcTp71VzXQH1JG/tj
e4LlvzdCfLMDcVLiP4x6iKi1inq7bJxundzfcJEzZ/wLNm/uI/u2i+R890d7w7D/CqhsOJ39n1Q8
m3UE/XTbNi5lb8FNvVUbzVimAUdRe5/FtZOITUhxihWoJ7OBwD4+yO5PAi+9yVfYa1NgmGs2WnbE
2HRfTnqRnpaMQzMr7Sk2XGkUPEXdORTARAznJepqpdWUFH0T4UguebctJj9gbSMthS+/Xt+XTPna
wqlaVHnM9+nqefJFzM6TKB95amNeVj9osITFhVFXSnmXMVv9T1vrZM9e94foBbXsnclM8o8vX900
Ue0LkornGcTi98INl7NQmdm+vhwaRk5LlLNwhK6mAGtLq2qIk3gNd+2/J90453p7YVV1H2bh/NUg
MbakrQcfk9xyjOQ50eTeQt2GXdPX7LoQgxc4ooXNerUo9ll0tW6wTu6WzOPeQY7wDRRHSK/s5FoJ
b/fEWN5n0JT88dFqLLx7r7OxM5cNN+f56UcLKV49QES/PUNoY/dXsFzIczTxAbcDu0NJ92wsR1NZ
Q3cTG6Z1NZcS+Ri+VpqOy2pAlMfjBADa4eBwey/vIx8CBQNV2ErF5l1kLBVo65idRIROb7ywEKeO
jxvmwA8G5mxQwkYMITtZALGPl5rI3U5Xz3kNOFxweRT14sO10FKxq0/vAkx/6RoJ6xMtU/WfbURz
DirPagsveixFPexxLLBv2vKlMqsiZqt/ApgQFLAPKcrZvDZJpW7KNwOXib36mwXdVKP+rSYQS8yY
Kn+5ceDij0awg//5/xBBEJwD1FHzMIXU9rNt+Abr5pK1iLdeDnpqGoCIJX3PykTfvWz4LqCVcL9n
gGXaFcpIpeohTVCgMGjx/d46lDVoP46rGTRDNhTg/My/l7QRc1+XIAb+JMxIG32AujsyXL30ScPS
BowOdYxcjcfiU4Fl0gpgAJ75XjtMmOEKWXzMJL2cA/avbRzNVWiU+Lc55gHNlu7wzq9elYV6oCcQ
jDhBDrKgzJ6XtPnqju31nxFAUCc/cq45vOK7NC2DFB2gb13orKOU1vXYD7Ath7Pb6a+hZkO4/ANs
LAQ5eXQGwoKo4ZqvlC4TfwTngrOjd2ojCSong+Kyt5oXwYi7xjVWQFMd4gIt2lUQb3G1WMwcPYe3
kU5/h0Q0J7pJqqpGtNaBsubk25/Bp7Fhx1IeCSW2OMC8RAecrc6kPkVcP/1sHhDlwV1tOrJn3MuX
Kx6a688w+cdW5FsSgEFFRbJw/sJEFwJbMj/qSzRE18Yfcr5bbKy0IVSqht6yrOqOOiC5c5gqMLjs
A6hGwy/0zFtU7vqrzjSjYsDhLJOo1IVY7JfzC2V7CXn/tu384od579GSYGxUmyMlPFBODsbLHpRE
eSGx6zFokWeNGEkhaRUk/FgMS/iyigD4b8cwZQ+2wMty0uzvDE+9WqKpKHODXxamkpsh1sEt483K
w7jWxzpfTNKcpbJZdIQvFWq6yFykalsD5yA1cbMy/qqiSgqc1GPx9qTdvgmvK2QCg7nrgsjPmYbz
8HmiAGTMVZsXSdoCCxMzk2uRURSZ1qwSlUTTpslG+76qbTda4id18zvZR0VxKtKomlS3mstOBmRL
P66mnEk2wvGstnRzNRL6WvwlEIVMi4XhADIX2UAhKg8pmMJ60Ir1ISsdjXK5N+I7VgPPymexklaS
vKbly8nEm0Ricl/F3a84gHzhiLLiDEqr02UDsDC8oebuqZ2h1OIZUdATsdl/E4WVW66BQoes4wW6
kGKNjEk+EUDr09xwrDZUwhxQiMPnMrwEXZO/m2DwsttCdlt3JgHhYEX/1LRgqqOMSZgSUvuPlAbJ
laEA/lH2fL0Nn6SfZDqObQhw2OPzS/MFxwHrXKteN+6ueRF3MJ+G7ia+AqJNINKcmCREhEa2o+Lx
TkM0JQdYxYjdY+D4DTf4b5CBCFc+S6WCNyDYop/mDNqsYU244dkSELrO0OwDXOoPqi3g3B1qatFL
mh9Ngl4LX6e5sLQSeiWxE9tX/Rieaw2exGboDx9nQkq95XP6TdzlZynMS2tHfI4A3KRUJHsITXsR
TgRRNtphGmFISFtNCn7hx7iSchop/1LZqGnol5RK4KCp6RZLlKPu1f9jiWXA1gYNbECAQu0yZX9T
9RfuDK0yMfzsgpfPT3bNTqwt+IaW/dFMMegCyhaoUKfWHTAZEx38SLziKLV5IHdVAPMd3uwSyFMN
w9TePGq4i7t5zBLab69GPXuGWz2B2+NbXZnj1pzYI4v58yeRwm/vNwEyZkNskyhRzENkK8fHu548
Y1FSUNTUx3a2yT3g1VJrG7Y5P9O+eybcvKuwYxByuUvD/jcHcAY6KYPeyGMzPTnNMgaWSfXX45pD
oo8Y2ATSt4GjkxLUm2f4VjmNPbCITviokfvFjqlbHOJSKwqsWJMbhLmTrfyZwBSysut+qyC1ZD4G
E2qns+8B2IJ+vjHP2gLdlK1PNdYZSvWlqWUGCsAMtoglG7s9arJb3N+PHzSRhL3+WMkjVGTzHIh5
vsaeo2hp1el8QAHujGc65vSGKSVYrGmzFX6hgWp8BjMk6VWKLpUUQ31h+WaWQNaBJQfePcbmB8ZQ
rb+Wf+zhcYa4OCtrSp0FLgs7m6gslR41cNV3aXjwukVwwRfN5cOMw8x6Kr2fQZpkXuxP4Xjhnx6h
wHj72WJrCDcMzJlOKTf4vUoh5Jc8DBJS5aw3J3/jEvU8i8Q41UdCaxq3ai6ivRp6oV+qz7PNd8g5
aidOp1bzwzRmIpknjTcuRiQrrz4OrBgifodtsTzAE/tDzmhqxq0b/JZGLu6PFWHhMNdeGMvu+SKj
mE/o7kuEzLcaBxxJefJPQzehJ0i/cNf0yjqrH/hkcac6Evd7xr8a/vXpJNlTWtdMlAPnnzg3eItd
5nBoeLt+AoAUigjVxmK6vtdtvPUnq5G8mH74JqY4SNVEuak3mYX/4+EvuX8TEoSEKqcYrZOIyHeq
ReeHp/3wF2l3ulcQimflDkelhpvZ7vburQ7ykacxfMxfLUdVJmczYMuzRyvoEWLyVSlRoe/VvgCR
yv4affC5Hh8bmahEKVW8LPnrw6I1u/zycNnpMztao82A0KD65SFzztwo+m5w2tWrPlzWwOMZ4J0b
PQslGHh4qle7u+/ZGjuvYq5g0LWaBWyaxCK689NrNeCEtdM3Eln2Tooiq8a8K4SVWsMw/PsbD4xN
mKKnan5ymIJrn2Q27lwbHK/xFMtq2ke/ZsbO5d4tudcmqqtI3vRF6Akoy8zs7RCo/4ZxHb97TMEo
VoonP/4o8+Ard5kBoasYerpxLqKMTi6vLbkgdNBqH/PN5hxSjJlPEKw/OXA/CbmoUmFgkrnA1WJm
+Zrx2PkubSEJSOJgh+IDRj4ZPNPE6JI06IEWI0ZCSqo+w2fRLbTM0RpcIwhLMH49gFdPzmbxdJGR
VmOBSRnURYsn/7zUEESxlF8aoaXN24ByHb/BeqNsP/+RzGouFNMaPWsbjzCZ1xYACSh/4iF1JPem
UxxCAOKKG1FTgEKM6TFCUTExm908M7nhGnnGKavf1ZpafJ2FjYRI/GHs7y3/cb5I2GIY34avNcWA
7El1+9CAj3wp2GwIXiSadkkguxdnm4nIgUNkbhbBRc10Rcq5GhcGzK+FNLBefTsVL4cvl5wJ/njc
AuMUpnRxhZzIoRbYq7iLhCjEC1if/hIacd7qVVeGL/vhU6sJxZ1gJadUcJ/vCbcv1RKq6tDyJ7S0
SMoVzlJSdb22UoSTOQp7HMVALiiIhQuaouvCxgOBDeHCAjZMM9DNqUiZH4v+D7aOARwFU0pqDV7f
t0sSE1Ib3Qfybh3hSEdBecqpefeEH+vqhPehALIkbyJom1XdCGraX+4WgXLWO83nPaSdl38ez+lA
W+w6UhvS5828dk/nwZQPB+jOSSF2Ocph24gcpuq0q1vixrHwI87Gb+Lj2S0zMP+KRqw8+PrSoogK
+Vy1Xur9LBAgan4jgMQHit4jk589sRNVQhA4KkuE1iZjVjO3ZtUOzWJ0QnRAeyIWLnQabyh4aoyp
8sS5sTtgbw7NPEkwy9nLGnVp2N8MaJro5agzgsrByZu7j1+WYgYCnfl4dNmtT2yY4FVfsYjkVYYj
QIfp+a2kSu2HmSCODYC04k2oNKaeAmrPqfJiUfEXvTptauEE/qUYRqvAkUtMU9NR++9C1X0UUJVp
NCgz9htF8wHHJ4BgpHH+5olh2GFJvt4zF7JJjqidSUJHIYK+6jtrtI6bGIEpG8kPTVXbc169SEXk
iOCyUjJZB5W1Gm4icNmH4idR3CDarOg4eNKe43KwO6CZtvDRJfPf2JVGaZrfMXhMf9480ysYZ23i
ta1pTC71U3WyvHax3AzXdjrCnbXyxUhIJ6LTW76JWzpI0ACX+znYIopKxopit+cBgavBkNB9gTYd
yqMkfiX7Qb/2axt64wnd7YteLtV25e8JlpNqGSSh1Yig/5KpxsA3Qj+QAxXU894x5JXGDP8kU2PA
w7ovAINHifIBrVqP2J1zoHYaLHbrwP5Jrh0PtgMp63HbUtrFAgwTDHMDLUyH7Zay2vaPhQhA9Q+T
3YCzUeAR5v9Xt+YpywUlNeDpqr4ZuM7O+/sDV9KYof/yvI2v0kubITxfO5+L6ITAns1XseA14zte
l1N2Aq1CCEARJhHIg+JR8bShh+2KdBCXH0IMhF+e8y2/vhj8uqkCp3zYrJcUsoQtdq9/Ssk8Txgc
YUobHed1KNiQqEHnc8KOg/aGi6NgxDdzKLYe/hbWb7uNi8iBmtDAwJwiSIeB++kB33UY4zgQveyr
pDz1Go7EUtNv9wnXGsUb4PUWLFGpcZqpWSZSitO+1cw+G9upzrPRuLyuJ+6xu3l8km1lGmIotD1B
NDNtEzpG+DOIkqMDtHLlNEzCkplKAI7lTm6Prg4HKlAxyN91ZTNzUGOYGwHblMrYMimEECJNIXZA
eoU8CclRYTdwYS/M0l7200cjGM1g6Iwkx8vJO/GhZJ8lwuddCqmuzy9yFwZR/tOe0dkTDFpHYnAu
qkBbgsoORPYnI2ujdEPVfJSmo98B5gXawu33DG4xI2wuCNCXwLskWXxlPZuXj4MnzrfQgJDhuNl7
J4Ic//RlH7y24NAUL8WkZ/CyrSBDCg01aS2r8gL3Dy0cOm3IuBIrxNCQ8HyNk1rYyXcgUS5Dh43T
fqX4/MZwdNopIyqsDOG2Cm3PAKpd7PNy22f7KVWoqz+Qaa/Y9ZpY876Z/KTT9sggoefMzyLl2Ok6
hN2zAHHwDUcRsN8fogc+z18ORup/WcKYEap5Ftt59efhqZCUZ8Yb2QUtyQI+yZrmxWAEzH8IYhM7
MF2nT6tOxK2AQqY0gDfGKD87O0ZmC2oqa6vucbpN2mzze9zLp4nM+qkxrHnCf4mABY8cUvnSCSOv
KdVp7twGHyxnQ7d86W+MqqyEy6MtV4BbHEBB3wgoMzjeqlxT5WCZgXewzUnRaLXMQof6BSBs9mG2
SZ1d5mD8LP/4FWMV3RATPvdI5CrF52YwQsbccEh57tw/GbRgcZbg1NefaKazSnooCG7HB77YMFwm
yp99T8Qr+PhBtdcmjBgNbZrdUXlcouKuc14BRQumzreGSp1kwjfo8+TFk6CumW/tNQRihzl+v1gX
eJ28paqJ9dXJYzFan6nH5n3KZ9R8EbRiv3rPBZs07iZup0O9rNCFnc4FhUNGN/EDeHrtSajHQkgB
xD11fNiFTgax0S/vu3yE20myzuZmR76A3BO25JDT/Kwn3xUBTmv9W5YyZW2Bsh0MZZdp0CmsvFJG
1Jp9UyNT/vx0rVmtsBk8gSC2kjXUIrVb2wRsDZFk/d5falmLRJ4k8anuUL7GgfTF6yipHrI8OEUT
rXU/2kGg+yQ9pVYp1HY7Bg6Ygm6SJ+OksufKzv+Hif6P4ywNd3QjvJ7OWOIZJzYeEZjxfEU4iBEx
zfrkFAtlHkscIk1bWSyA2ypn9h+z6hWntgy2Gq+yhsfsYRwQ2asXzdDTPPLo4F4TuSeb2Su9aQcb
jxgaZMwJZ+qfnJ336bUbqpaAoufXvqlZo+eYRjqKTv5xMHLSH4aOPpasjXjlAIprll88bc7LGREf
wNVCT1UuQXOuCj8wLZp46Pw6R3J9u/GxT9Rlt6S60oYqyO5TZVX37s3CsEc3JiTgyAp/n+txhsc5
f87A1WQl+ZmuWdZFfJZ64qn8edNujH0schk/iFVFiER3l1LT1RrrxyqULBBU3MUiyrbfFxtuiMCM
5ijD/L49Z6iawR7/4aGfnuOEb0BmSxut0YnzMMxB+7dNJowsz+He4Wib0IpfZVQihDOHsuCZb31Q
bWBKBQaM9GDajFP09DgSaaRcg7x63+y43UpKR2z1VAL5J1plcV5ScHYf5zXNhPZDW5PslUxEii4A
DoEjiZ+9/U+ov/bIag0eTC04AKvYqrZokcfFXawnZEl1xSACaoxaLfbDZwMt4haayHICKZKVQ9W/
2stdMfD6xLXmq4+vdnM4BAupxqkP/cEpp/UcfQ0Z0ln0CW4GsCe6d9h1axIHEefW1eNuhwzbn2Fr
2/j35WSIHwdFBolodpCLDZO5y4SeZ+9Tqw3gQgTJpfXg/5UQHumIpUaKVFUVW7Cjmq8huQlL/NIF
cIhBVngv+NqSEf24nLSIx8dQ7SVO/yH77iXCtl8mowIgQAcDCf5uSqdvzALjfYi3tKwbN7HzBgXR
Wxq1KbteBiMT/xnNxEzoHJX4UR73v9kzbejA7yHYrHvEOwbqYfDuKuK3bIrQJyxuDEEkr4DJvtky
pnSKGZo7owNArYOcv2qhgG2gZyP1xvi0/HHJJZJi1fuO6U7QoTxBR//k8qEt06Q221oymnoPMcws
wCOHpBKYo/Fj/efUQyexgWLQGKDs0bMUcvraqpPyT1A3TzaF8RjQLmOCiZ6toZYAfPwZSyUquc/8
/9shSRgcvx53X3hGiQrfcRNAhYU6RgeqrnOlA7GeMNIPdXvHrJD8RqmF18n5cRxN+r1YQfaP6MXq
ipr9uapSK8kgH4j4koO1PNDA75s1iAi2VFLBmbb/NCjKatLo7jZrMwPNpmepUTc629ELu3WEYWU1
LcsLR0YQDqrSYXcv/wHVRuDF7EU77cG2HNzR9yxTVjUHTlQpsy8YOmIhwhwb+kiVATmOz7qC/CS3
ouucteSMs6aWAGf0vy3AsLXA/ykKRcEHKDHypG8/DFyPRBntD4Y5v2F27o7K5z6/cHnF2vvV97++
lzz5jPfINXLcX8Uw+gtrjTlKqwBnQJy+/6Lac0ffvziUwDzLgYtnsuZ2ZdbciJA6W8Hhx4VwPDca
ByqV0xJzCzqFJyi/0riv8WvSS/aNNesmGqDueCXOSo86on7B4efYQp9g8pw08zOV5XbCkyDFXY+w
21PxACUegAyaPvD+o5wJrQG7hXxGeaIqwtLC7EInmqsQdwaN2a/ZWf3BBDKJXqzjFC0ajZBTKmLi
bRiSfE1N7/t2tPOc4uuOWC1SIPP1LMbjl8AzM4GKpr1GVEKjZR7yzSsXM3YQ6K5ywP7loWj8OP07
lQZAqWIo4Y/cEjFK86i6MWj7rzf+MOPduyAnI0dR4Z3HrBxn8gV2CgCbYoBAdd88DW/peCIAi856
eCq3coMLPncl6rFDQOfLKD3C9G/Ks/a2lie+7DfuQjEGt8dbdaExUs7PsdkqrgECbNazkkrLQCu2
AJWD230ikduIpK5QeN27mqt0RWXSsAt2Qwq1yR55zxnxXkYvR3bRVrobbXgVD6Vpuk1foyrRQOYi
rZYI2agFKKsIX4Jc8AWouwFdCnB6AnDn8Qz0tlktw/KjMpedpnU5KF1oMffRMJwupqMNejJCua7F
hWKi50kbw+4lFlHw9oNPh+SgStI+L+OFw3VB+TjravuRbEPwHOqhP1nIXCZedMfxbDzpcTY665LJ
BlhaQj18nLvw8qOxe4wAdMwssevljSxifo+LXAaE4olEGJCIPm77VZjgL2CoTgMdiEex0lpTOpTZ
iV8Lk0K6R/4FfOHT/1BImOIvrnyCAu6TUSJcPgQ8SsYuB1zF90mTSZDikMCRkDLY9fi6LXMMjafQ
jmV38qPWrpVA7Kvu7AeTfyackzEtRjdWy1wVg+A9OLjKw6SGWYjJ8zolJWfd360vslvkSJMv4/4b
sEUTpucovsvFiVdf9IJeZCNxqaNk1Kt/ozs8UaED8EETtT3Exi2y50+oqSE2sNY4F5goNPc6pKOq
dvpmn3Wf8tF65H5yTeBDhej6np9+fTJ0LlJ88rBCxElLoHfwhO7a5fQnwg80kJcRwDrZinU0IYGm
4LwOgs3ZxexH5EhRcXndW4uPEVOT4ep0/y6noBexw4GKmQUORZgaYgUn3+b/6mdtUS3AwAjU9UoT
5mr3rcjRWdUZQhFUbI1VZ96T2Z8UTR1LgQCZiJZ/ahgFaoBkfZlfiNm7TJR27SBB1rTdeTHuWEMC
ZXKjZIeCqbSNrOJNl9QqYuQ5QEvMQBsKC7R/bOh1G2OTj1XA/mCwdHjak6qaZPfqr8vk9HRxul1c
TCSqXR4fOf3/He3SAvY6QAy/xQDgLTdCOXPsRAKQbYciig8NHon1c8snqmggJ3p4MOrNSI+6w412
r/zYn5GMRoB10hiIVcpycJtWyYeTJ5kJ/b4tXYJDPLqNmYGVSfJFaEiFfE2Mu21LdoSeJHTH7mRy
2mjNctOtqq8sJ8zu4P0gNTWY1IxElH3jE5qDKLYyKO4HZkcScTEW8ixtyr3QI6uMmRuZ2sUW4/zj
S3opfdAKaLeRHrP9QJnbh8MYEnmzZ+5hw7SGJdboPmiL0TED+w3lc9CCUIgUyv8pRa6FFgKfnlQ3
/KYPYXgBDEg6RmxGc8FQ6lywcGX8aXGuGu5NL313XKvIkj0aI7Dys0gUWFXQFJZEv/o3JkBOfh1q
Ct7qhoAGxnOkFAV6WYPzgremOtQU0WCpXL0cy1WletzpZMWJT8LLsPFyNxwqOFiBO1yQXjw5ZCJ5
gvhonFGsGoWLACluSTewcAOa/K9HHQAx5edqevrtD3gfdks5qbRxBGIxc3fpppH1U29zf5/OxFlw
o45jT4GCEKgd2UHgz41NxSxc0ee1OHbQIzhbZtSBvZK2H2SAOfY4qVsfa1vmhUd0NlRuHvuQZo0c
053B/oJCNyPijCO9MAb3mbb95LYDGuzD8OUdCCqZ2AovVAsNTDityaiAai882DqWw914L1t3Id0v
rZ+/RuMVRFfaifI3euo1WR+j0Uqfs0rt4uegeukWcRl6832JvXWeoUvbqOpd2zCkW2UAVz8xJ9JM
9o0gHmsfxZAwMnEONZD1yH0Tbs1FxxXtEpXR8qQTr6zDyW/veNBSl3ZLgInc+cL7hY/15kW8Cb51
CioNM87mU6YVltGrgaIN0BrZyCoy0vL9shRu/cRqXFxPwei85+G7Y+yHgZ+qBvUMlRP6iaNn1Ofy
PGv7LB4ZevIvQ50jY8/q+vY1oKfbA6if9ZgSGtRGJEudYyjUfGKKpaLFR4tEb8jDCobMrZNOpSaA
5wQvWldAtBp0vkR1m0ksdexOfn2wDop64H3+KfMMVq/QdnUTGRrTGeG9pRN2ivQI8LvmA0Hz9rI6
62qb1PbbJkVe6nlf0krr3bKBVXIQrXDnJSiCSOW2XVjqeSYehHx5uPm2SWCZV3SAlREe/TqDxTCV
F0AniqC9loYZV3SulNpv4JawrGin9GcxzB4CwqY4WXccIWI5gMzgE8JSuw+XdrTmv+gcCqJjUbbF
tfu4980NkWaqQUD3pR7LjKcm94xpsxhTucMtbHRqI594iOmvVJb7IDtJRVQdIT+8nRwR8CtFIHNy
IFzw7psIwomAC96wMNFQNcSUe474H3DvblivCMV8dRr0RFvBkXymkMV3aRS3+pDW0SYB2dfdQfEq
ZNvBr+ojeNWuFyAhHW/XeoHIejBl7e6BfeYt0UaazgiYI1NjtGbbrj2QOKax05NVEhvirGy4a+EH
0p1h5svXMjlOqH59LGn2Z7P2Yf2JA5L3fQQJ9fSnTmBraxTb1pTnidOi6/kCWF6ZPzrvr+WlPfq9
BlT1i/b+ynOablh3I2sb7tIYWEoXoA6nwrGKPx7VkdBaILj0EJNW9JH6Oi14BBDc6Ggetl10CRMU
YVS9A/G2nKHg7KvqGkqmu8Yewk2Js+8M//EsAkdKvanEkxVfjVyYkkoDTJsFGSfeW9fByUFHND88
mqWtPIL88PBLt+nTcZ94RHqJJPADx+oCrY9DmRQe4qpiNp8OgU2qIp9b4/SfyO4edyOQiu7/IWBM
I7I0lBIqBRpT/Mi4umvHkZEXAWUJfsooFZEpy2nL8WdHeB0wPP+JEwe6RL60FZidJwC7AMqFmQ61
9JXwx9Ya79jJXDemSQldAbVwWPUU5NLQFAbiWBU7akL9z1/pfqgbpfoTJiSNnlLFak8MjxJ+iVWr
4NNaqwSsDeBzXzqE73O05cUhDd84lJuIPO6cmeQpIK3/Ybu0sU8Q7j+Y1pJA/NPbe5mFWousIy80
0VMkK/PCf7G86DYYXqE9MXQXpph+8+bql1y3YYz/E4l7fP4uNbEdHgQBm7g82+Wh5hJJPOFuYtrN
nEuowkl8+foxK6/AnkVxoonK5R/NOEPeLKj6UXcqdJqUDXWhe0R1xkagqKfQJ6ZUr6KTB7yh4MiW
ik8nODCytBu1a9L+cGgBne3vkD6ZwvhXV5sWBsl8HUjt1ADPXwbJsuW86AzafINSksHSSuRrDMCp
47Ik+eDIUwhBUT/3PtaDy5KQPym3aE1bGeWfas6Fa0AB4LBrvy53yHkc2OOzyhk3jvnr2bu7806D
L0m9CPprSNmVqFE71/IXjoXlW2FcYvUGy+MGbLvDYOhe6iuJSeGGUbS3t206l01mFnDDpBFN1Cxi
0xdeph5YkCMIeCD8smpeZUIuXzOBDKOtV6VaRKYH3SEmSRBHs2tOdOkPvTNA7PXbrFApjKUr8Y/7
jc0EoMKZbJ2YMAIyeBd7GsZJWUhdrLLcR1cTStrzdlH/UA14JJ8xopLFwS58mxr/pKfrDiHR3cDl
dq9CFoY11OyPhzjqUnR9sFT4ciKpYH9lFX+cn0f4BIXSn9nVzI7XoVevaAutBXPXJtcUlqPc3++y
7CoIDIgLHVWovY7Ccu7Q1ttKurcxDu3lABeQ6jRAv62a94fRQkj+aau4VQXMGF5GcFU67hfxFuk+
yvRtTW0GOPiUEdwBrTBZDvj9N1rM2wzNu2CUopltkA30LwYHBu7wLWyyBueheupdrEy4O5XN5XDC
jqAKSbNEbnmbp2ZHgiyYnzMV0pnjrEH6gaUP6ZuGwsLYkO/eRFtMh69HtmXzJw7mIqEOVeJgo6Z7
7FMlN/+vj9C42Ti4zGjmSqMDbnrGqofXNGMIFwmMOCEbP08/kgtm3AJoRvk7Q05qJXNu4x4hkPtt
8r/fEFKcnY8CMY9g9UoiD2LoAvI9K2/Az1qgcMws/RlkPcLFmGeWLXivdzwKdkkZ2oawO4eykG7l
wvTf/ANhShFQf63dh1W6JvBn/G3GpK5hBW4OcBtF0jKRoAB0m5CYP4BEPMUj6KeoJkK0uj0JuMRq
kqUo/9Sa/4YaTFWuknG/yTln7G6l6mmXOVu/KFP4W1XyXZ1g6ZMAtN4fHk6+IPNDhGtmat5YS3tt
5Zcx40PQoF9CRx0Qoy2Dezs6xDFdqOq/CMBgwjZqhVAQvZw3Hi+3tOsCBk4gDEOTTBSRocDqLEAk
Cz6Beg2U14uVtja4xTFsOZAyKd7wFYxkSneWh+pyy5YFCLXV/1mZytak2CKPPlRw2uXhBRK0REK9
2pUyODYY4/DPnd77fZ9mtAo1TADx7wiW1fpnSYO+ZWVqUgiAB9XvK02wcB+coo9q3ticEtumxfFr
V0gYIEAPfkN/csfqXL6uPqV5qi6Z014Tev3MZQG/EYkXFTMqxmm9XOMTvTsbGdxoZVGsR8BiWUCj
6abdUfbW2c2S+tHfit42RSbuIAuJO8g3kOFkPzk6Mtxr2vVX9bBsVn+oe3H1kRvmJdoM89Ccyk8i
XL+Ut/E07FcslG+fb/n3tUZmLhXWjYAmw6Z8TgUp7DE2XSf7zy8Mm9qyi4JC7ilqb5aYeQNzASrE
xR4ZepVl89p3SInUHzvAp71UMbzEU6WDzOhha9K+YPyQSfmRLLPJXJ77y9uSv/blXmgq+iEBCBsL
Hy6AcKWxQnewfmj/Xcr2L1ghEtSYLLtmlOlx6Y15wJxwobjhNrKNazp2GC0DV5hVkU8MOCp+hY0j
sH9MjolTIgNYA4+4tl70mL/IGeuZ6PQCtr/qLL26k7jTYuFvMHHHE7uXHE0jdG4M7CsbFgrPgIjq
cO4xHuDIXAcGJLE3AOxtW58KgoTiKgP+U9eC5HAVbyVWghvN8t04qC7IwUBEfWfJrWm4dTb++j3D
qEUbu8Ld+8KTqu19jz5d/JS0tLUvoKqKBnpwZBaNGT009eNzrlEixAmKdmtGPQDVXZuUqNBu6mzK
uV8eS5MZ6lM4AbR6vJPzvEIqeOg0SmujOaZ7Lp3EcouB5a1KWUVhKNXHmUOc4t2tVsOw7X0mrYV/
dWnur6f5XJjhBi2hTpFSr5HOr0pOtRPRPBstnsOb6/Z/litAJW0cdU96tFI10JqfkaVBoDACOQtB
LC/s/NCBiQswXRDrM3AUK4tf75p3YCeQXcKYAX9sA1HMpr78hG/7YN47N+NBEKCmdtaXYPqV89Pi
d8WCKZHTLNDLnIVAsKu3yFDQDsPpmkqPClR13dTknmgg+aJ3Zkt5a8Rz6YHPYCUeIKro7k3nRQ0u
QFMRX/0cxucJHPxtquFnP0XSfTlq2LMCwMOzBA1oUzymEQ/B9Qcgzcx3VdklD+CR/pyxDvMqTE5o
BIUtY4ty/YCC0XX21XuvMPvpod6kOuN05dWGl97bHoxSPBlKOwB0rpCWuGigReqvuoETt/TaQmoo
AQN7Y7Q5O3NqoD2KRQQ8DE8jx0t3LfLJG/hE47bpYu4/AEd1o2UOWZD9g2xEEDLHY1m3qtABU4Rh
NPDYLdpSEd5i1P0wUqw/k7V09l3PZTSIRfT3bQcYCQmaAH8N65YIC36pfkb/DkLd8NxA8VgQM1ud
iUKsaAgctAZLwPr7/WEpzmZM/LDCGjo2/p3Z+KqFm7lICxvqqr4amX6KD487F34z7Z6qYpzmsYEt
Ng4oZmpoY1sOtdIbZWaLs6WVIWaxodni6dVWcANmTCYRdV9iVTOM19UeptRfXV6ohp6qY4YspYCY
zjoNafnqRt5m+BtcRB5fCZzB/zWfy5YuE02+yFSAHdRRov9CaSZMqym5QKtRP0F8xfpp6gtpbT5R
q4f+KtdmIyGdc92Ow6ZS/UCMU53JxccBkbd9yQhhSnT705v3nUnPZ8s16sfVdVYgjWIjcYFlVCaW
4JvONO7ha6FC9PlSG76APqrLxO7moBm1ZVZ8rjNjF1+srKA2EX4PcX7zUWOVXxIsUHkt8S0vitbS
ag9/0+tWjVI0Xpeq5H2pNPA/WNoaQIEBsLUrNBgrXUD7QzotAxihX7+HNDXexd0TBpbg6j9OPUq6
zdyotOGVjaeY9Gl18YAp3y1+ndoPN6D7cFbkdlweSvduYmm5B0lyRsBhMtlUZV9vtz/92TmIce+D
OMkrB2hhdV1e15p+dN5HS+ygxf/Tbj4x2Rw71Mv50z+N+vcAy6/v8pkRVLbguFmCZY5BjunuQTPa
q+uEPZiU6MdbD1aCiR+8KkVLwWATAub1T2CRnHlMinEiEjBLnYljhFpIwUcKGXyeKPUBPS9Km0jE
zyacERfw+X+yrncAFyNrx8WSRIUz5m6U7cGl3O8vSWYwJbsICEefdcqCuSBPYaMAK8UPOwLwhjHC
EUFs4eGfGu/oDnZpEZzN4jmPX7lry3aGQXgCDX+FjAEcv8Jl8v7ss+TaYtmBUEayjDQi8K4Q2sbf
1ggJ1MkGQBlQOJ7EB4xnIKPpi7/1ouaV+6FXOk6zUbYPwsHOKOdMXAb387mYyMbiSs2SY6SD/BcA
UaFcS5kQKZRLdIjex8FwlScjVsO0NkNKaKxhtuhmc734sJFLK+0Pj+MIw3t13RpxRxdMwsptDVP0
PS9K0VgX7plg8HzFVTGxHuJ0SWSznA6NKNrs0KGfSCwVhHHMyfqVMNrRHw/5VyM+LQDrsGUKqlwZ
7IpvnkmK3kd6g0S+WQUzF/wLOY6oqlOcOZjrEUydvKPZg3oqFCXKVJE3Yn2CaxYk6dfMFI8ymcNG
h0lNdFGKdKqCAFAuzo/nM8M3A04/UtFVJ1vvOXEXDJqWPvLFOqbVM/V49NvD0/+m+COqU23sOXJD
JGqS4TgXCh7OiBRGBFtSglnVmyX2zuDvYWZCYBw1XzWkgjD4rSxdNRY+hk/Ka1nlz22J9flOVIv9
MfUcwbtDAcELSaaXeLdN8o3clw68FNXIITyf3vHK4z/7VSYnBZ5JKBWTNSgMMqYcMd87LP4SXkne
Uwu/5DQConcb6eisxQIp64Z4Q7z2zugmhABL8P7HG7iJraqx9bwdDkWSSt6a3dZxWcQjrjvRi5+0
ife+P69QNlXod9s7uIxQNA7T1T0SXYCHprO/SRHg1XI2k2N5MyRxg9dAl0NCQhoCurulAYwhgq8k
AxrIwtG60uPao+p9j4X5hN3VUoutlZ+V60XdyLvFF9jFLBdC+91e2f6bkYMZnKfAvOWq7AuLHr6A
ZrEmB2bSKw/M5DqtkTeH8oxPMJ6KLzC3UNNqcR9Ru10bOe1HdP9+4Fw8TYbyOKbBdQv7yBuZF2oQ
lCmYpKs2j2SD8MZvKLcKfjtmBloahcSy/ORFC4r6VXne0rBsGiu4p2EqVSWYsnY+AzuWiGvQXbUw
uHRKEs2C5WtM/4oQo+cAQs0r8vn9PdOpM8wYkctMdazXhByKV5hmldVXXl56QJFR05QynoBnAtMo
ZnVGXyNK1CoBUyQagTWZUtZH9kMyqR5S7wWR152nVuB0HzVflCmaRIF+GqTO1+7refPJRULiRVUX
VY346N74yuoQbdfmyFTdGMZwNaaWJufdC6cQLa5WXS9uD2vfSwBk8lduXyo5CO/n3ZtrlW02rhNh
gFvT08KZ33zf4oSPnUV4ZxkjUYtcsAu5DEVcidAA7YvrEdIkXrUvXtX6Z5I2Bv2NqzgiNpusjSjg
P1uhiMa4QCS+W+clQOBi8EbmKtfxmB2bhF7fxlEPVaGntkPUhgI2CN8mPzxU2QcQ4Rey73omhNEJ
P0/SR2AyzoHshiiT5DlfT0/lTlwZ6l/+FvWgt2ZOsha7H7eFVrB8pQpxQeeP6mI/RszLnJuz0kvi
GGWgT4mOI0hTWIctu0dKetTUZoHXx4ILLyB99SXHBCDBiFj9exNrRm89NCs4l+wL+FUrmPF60dLz
jnHeYBtLsJfbTtRbzxg8BsrCpNogaYmHEID45IkXUNCYBDd29DyoJDkzXiW7QYmPX+Bmsfqud0Tc
6iJXZDfQWpS3ypktyyAz9gsvA0l6P6Eds+nBn64k4c9aXtfkKAZC6Rq6apTLrWpYIslT1dylyZ5n
KKs7KZHOcEqPk7WA9Aa1I7CONjDqSkKmpAv836wUBb1nodT1Bu7CXC9rsh2YUr7j0/UuoisgiNXH
GjAWtfOGeyQXy81jvlm075SP8OPKsJ3mtzyagex1XMmN7PG3Nf0D9I5jg3LPVASnrt4ZoQxdC6p5
/emNWUGElXoF9aSijYCLSaMmNdn0vvTkQ7KAhnc8+nQfGI7rV/6hKwKR05T4SOBAXVNv3WB0ozLN
SLosjoxQnLXm0sc8kJEWh0HgkZ0BifT6IPzTw6dUDFE6vvWTYLCs1if1othkZxRsC2STSr0bLUdD
G01iYucfUeTl9XMFlqUub+w0y1D4QdLdir+LeBTiLR9PQip8d/BgKWn4yMbUNPoPc0Q4jY6rptvV
WqxNA5fV/cvHQVXIYk83BPMJthPGNm/Xsx4gbMJXFVPRWNoPJZPK3GO2SWgI8rQqGZirTpW4Cg1g
VE52zOJ2T80qrIjw0b6KGAgIDDGO3A0XsoKa8hDXfPC11v6aDjsrc5RgdHmNu/p/cisxM6VfhHDg
WyV7IFqzU1FKqF5HvwYU10WI++FTtgOwYvNsa1OBeUtpSqaMGX65hZf0royIIAwthsEeNTaCZbBB
vBfK9JOmIv3nsjvR7NFnDDP0Ztg5AZomOjZ2EWAzLVX4L0wZGkIAySSJUxKNZkqxH7x7WCq9DEuY
s6WLUeg/2ue+mFobbqDRnAqykXCQU7EExzeNMEWP8XKrBWAv5FJQukmi+clWlXl1URLs+cbOsKeQ
odFoJUuNH34LU9Hw2T7I7G6WEKXbqXt5LlGRS9KSJWauxLFBpg2mhg7ijyUv/+puNLyaiARtzdST
4AKYGsZ0RQvT5EUPU3opSGmqISygY4poBwYIeKIx0YI8ovrDjZjzUVr9D7UKYWGGfVJvBD32ViRb
5TcGSvssg63m41Awjobl/UGGZxuZ2uqpznT6Qdl6Os13mfqzNbaJSNLy4mGsGjWB94H6ei3nFw3A
+0J37X6vp/maOoF9VSWrDqIyNqrQSuuSauacJah5jawi+HqcC646RDDJw2HXWJt7XFeSEYm+ojhS
Mgc0svdwbQrWavR4ww49S7Js5IOfekm7Rwet9+3KVZpqcOPeTJLOrl6C2f+HX0jlqUsAgUSPkXx8
ueKOsAMbQ57/ubElYYWIZPqU9GsXNfguS080WRmI0Z1fAVwwmv5jOLjbe2TGQpNkC0EhNM76rIkQ
6qTR4RX13iQyyRwbAvkQ16X7ToP+lFkyPPpM1jgvmYr3Q0RtYRVtScpAInLu+Xp0lBokZBfzuCP7
6tRxijImGW/yXzjX7NDc9DSf4JjmMj3POgxHyEvIdL7TEjIIDgUpKGeziX/StF1IpTfO1dH5lZJW
USqORrkY+OfXUix05iMvhUkk0WP0m2aebd4qErxn0plx+whD2/4lks06cWhhIpAXHK+l+VohdWtt
FtlFkvOQKDOFmSrkNyxz/URHgLTLC3+c0yZUU41HQp5SHhqtMaBCY6xszYDVldNdYDeiTLcpTxs9
HLM2A9ri8w2lBl6fR55P50G2rwENhAkGYUOc/2lazGNc6gJYaJn8QATWNxS5zGksnv3Bv3TgvpzU
S6gz2EzWJZo0tCRStg89zuH6W+zVoZZNGoXToyJx0THHisz6BBF851GMVHjXsF+lrvjtTF9ildD6
b3VC4HtrKBR+GBHs5KWahF7/zjODlUrP1niTRjmwrFWtOW2s6tK0Ahe6U+koFygHumZFlv5dG58H
1n2dfZrXfE40oVwCSLPWilMoe2RT4y+HLvD1454ep8lLmqE4hoEAB/091BzH8x/eUMVjdpTkbm34
BNeeYSN9of/sV8mCRvVD22qCmmReK/90yqTmhsHwFpYurUC5ak5UT/cmHtlXEQGtA3j1uA3dhGmo
eGp9lbU0kj9JlCzlh1hyGUwTTRBgeSClRegIP6+gyeVWW8/PKHyy2JjMxc4mpSZWcnS+YfTJvwQi
LtfK+4jZ7j7mqLXle22eh3yzlBpWcXnv+g7+Jh8SYV8jTn8tBqBpKCzDficPW+FPsM90ABj5MK2l
Bimp0whPw6xvpfVneeoVDnaV0YyXEFrnWyXshnwqcxVd03OswQLf4BBs3QZEW1MNKwq4+IVjfsh/
A837/ZloiDmYMmzw87ru/JDKFim6hjff16yNSC2nKmn4JY8Cigr85RCX6KYOW525by4X7irTokOo
+vPxHighmZ1y39J5B5R+lLPx14u+H6IilglB6Ube/aDi0hgFHc3HG9MuPhxuQfGSQhBJXpNrhhAD
OxVUn+7djSpDiWCk3eOG6VupU30MC+vDyIaQ/rgy1nbiLjdSIv3MS8Q5PSMt9o7CqP+dSzC3/5BN
VdfhzEKJOgzpFtCJt9XS1HQn5ZXx8v8DvNnoOJg+9HRj+cA7BVNezCj1rcTNdCHz/6viOxU3v9DL
cmUbsxP++VrYNL9numEnf1zlcTaYV6e68B/FntMwg/IXlDxLZKRpsjY/YDUKVY3hhMG5+uCHauMA
D0m4SLxkS1Zn1AcR84Zzxr6JagRU6UpfEtc6y6IgzrgB/FIpqzyv9hqBllN4uchJqqV9d0Hlm/r6
dsevpDzqof0cDDo+xu3gi8vjZ6UC/1cy2YtOpspiPBCC/Iw2EBn8ew8pUfcxbvU4rdQ3munY8tsR
XZjR01NxbNvIa4vUdh45zHzIwMRuJBN6SXGwdnOCvm/Ohq081fZuO5jxDP+YNZqYJW09mvcoHU/z
Ap5/HpRc34OjXB8YGUyS4/orV3c9xw7UpF1J70UM/n4u7Z+5S4f8N/Xd9bA8kw4L7GvOPV/BV3Nh
YNUH4zoJKt17bXsPD1W6Ji2ojxr1AT78Vg984l9tEhN+IjTBZJhQ9r/26ggRf6az1Z8zBP6C+yW/
g8UmN+1f0DJsgovQNJ3WgsHU3+rg6x7/oB7JY8ldGdWHLuM/DJLz4GahjEyNS6xrlcpHRiFBJChf
UR6fbiEvv3Wf1QDS3SDQb1fFt3bMdVbUaa947smt0sh2/5+B5Ih8nfuOy3p72/N+PYkqDvUaeT8m
REz/8nNKvqjNmGQsf8Ii4H0qP6YU2DQ7CIrfJwgvEuEgqD5TFF4rwsMhvrc5+eIS3yz5Orgv2VI+
TWMEA07KTq5/Iz4+xiAK+cOPW2VkKt9d8xcJMwgE5lNwd12YeUggRxlaoaoVVEf2MdLIVrAg65n1
IRwT7dbHMwvmDsdkpvbiPpQxJqEqhN8xH9RjHn2U2JqZ+5om3A3foaeGZtDGy/FruCSgBNvkBNCG
FETpiR3JrrT24wn6mumIJIfL7oHfU4eSO49mWMTv+aOJ6znA4uM6+TgwDi1ETduWNuqcF4Axnl2D
Xixbqm4kVMNu/aLEVd9uJnVnnd0Doom1suGB7yVbwzG3BieWDtrFpdE2dHgROlluOP7Mbl2xquU2
Pj885DaS60zJmA84ph8xs8iVE8RtieWRvVLeHWGv1mxwGKAnMACOMQeKWS4yXrE16vFDCYX7mY3X
JGPyf8RgRUfcPVi88RGQvj4h7Z22XUA46qmQuivqjCrNn2+M+JaRpiTl2ot0qCSEZc0CbTTz9tE8
xKUBM5cGEHSuRRo+Gm+b/V57/mDaWRHPeVhKzvf9LnMxKy+JiaZl6+VkouPSNEteh4WWklbtQOAU
CaypON43hijEqWCRvlAMF5TASERYvVW2RE3IIAmEl6h4cF6z3Ed56MjqOTDmnpeZFVXKEdZjx/dw
2XvVjm40DGwWu3g1pOQRMcVxGugOjkJtySwOjRm48ZZZ+ze6RKnFKcCkW0nVL48HeQN+IPtZNAJ5
34vS4mZ8NajQAlxG4/lkw/JVnvVlHxbex68C4KnBUE5udUHCMrw8iwbhgCDykzqw3Leuhy31kZ6n
/o7/3OlbZt0snAMnvKsGBV5Zz/kM3Mw7Jv+DEFcomUuYGO9s1GO8fbbLLOfNlQUxqvYgHasrUIgZ
wJ8gIODBuCyzUA4PNV2wkHaov2LTlAWyaPuWzTCJEVEUcfyLt/vpNh7CXgfUwoeayA+93pi8yt2C
RJyUOFlzNd0bqjoFlsXRUofKhb1Y8SlPXGrfFLDdTd2zPSgMbGkaS25DxTz68D/046Gs834Qlr4r
NlC7q6jHh8+uw3Xfxl7kw5MU8Fc2ofcCgPd6jp0dzqacoGVX4t0+P6pDZtOEnwnDf2RV2YyGSn2J
uqNVjXjPQQPMzFN9NrdYR4ohRGHXLCMRf7sepF+gZ64J5MQoEp0Dc6/YxohK5AL/OHHOAY7bUAnU
cPprrSjoF0rB01Bkxz6+EWYy3QT2HTlroN5fV1LhKBTGH6j/yVTKC2877xruQGkun64DMuR9unvU
OoC3LtzQgsDtTxpmlOV3D4DDc0iDf+b8F7ZeWpWUrdXLwhEPncCmfgbXzo5B0JoR8Z53LBnGz7kW
hL/3J3sTtip9tGZPx8ZGtr6WUdKLTx1xBozjs3DkGTUMWg+Vxw5p1Fvku64QRU0v33N/xxYEz60A
RD1wXgRH5tb8/qbqFDn61gTLtf7y6Xtwd/cKoSMAGQbBl2fOephobFo73T8QFvpMY1OQEl+u7vUm
VnsOAaLYVL8kT9XQcI/6YYRytgri1i8ZdaB1v2EOhmEydh0liTa6SOrNeokE9KTswmUaGT6chvbh
0foGzKuiX2G72h1+BbpmCbYynIkY3bBX9k5DQLbnU9rzhEa6TZ+5dG1klLZfcjxl1EJGnlc883l+
Jn2o4wDBMf8vOVZc67sdAXFOVQ9w+01RDZFSTulMsSzvNPejRKpDjR5gv9hQJF7pWT/yaPCP7qu7
9NwJ/qMqOCQjKzeaROFp+plUMJXMuRZtUtimnH2+yA7VGFfxWpLbNv1qygsV5Ln7c8QpPeGaAcft
B6iXd4F7ny3X2IwD+EATPVZn4R2FYhHp79TeBwYUmKT/cjdKeJFnl272nhrJhRyYboJ9oeA6Qmpa
RsjZdiB83jZO3r014qeMcdLAzbsjPGQ2J+rm/OEOb57GJkGTlZg3P/Kbrt6U6qS1+AA5MTcqsMo6
JDUclRGOV2cJBfjBxrcUNErzpyyl4eHOaH+7L4v1Ugzdf1d15zG0ghKdFat8+cqu2GPb2kRWxEra
sJcGoLOTWicKRPZFjtBqbviDMIWxaLpng8eQcbWqwIxyS8MciYm5ik/EHwds+6cQT8xTVfc3tzo8
t/CYDWpTCmok8Ci/gGJImVPaz/JhYa6fFbVGqncqyHmAR7BrSlekCDnqmUYFCkiCW+vA7phOfQwP
JseyeN/BFiVTvRkxyCl9/SAEcfiUAcE6duPr3zQvD0S6QM6uoUyJX+8v0c+JClX0g2vf9s1OFpeq
dwUKRW8HCn/xeJOzOykJZifMbtBZ4sNLz94zXJfSEG0Eh+5zVfYILSZEBVXk+wuaiSpDACoYm6ji
R6aMXIyAgD5Uak6MiN6Et1EPQbhEAFly7oPB88lmQg5X9d208sVP9nxWBtwLU1n/kf2We0l+JfDs
BOemhqf3yJAHg1GyuYyRwZ+qkoFxvGEhJ+8sRHuiN1rdVqEv1y8vEkThSaJW3cGg9aNraBHEfEcQ
16/Tc9zxQjC17vPMc1lXHsdZE8BiS227ETUnNnrL3f5csF/oqmlU/ravmZRoFI1cNKpA8UK3IaiN
dEsC8x2nWXjwfQzeaM97Uuubos9Vbo0lflR8cykPwxBJXJU217nRLXZJf5ga+wvBbsG796FXiBe2
Rwt9OpPHgXzmThf/SMPZRXYKWCF3aT9WoNKyDzpMHl0ZWyNPAHfs8UAsQdI9GLGTkJAGuC24OoNe
AN9f6xA7cMnu2bQe18KynfojhNdK5ct+LQLcgXzkdmD20sXcWS/9lmkfkekxX3hCk7y8xW7UJZM2
Z8EqtERyj3Vwmty7NNKB3kNG8xUfYlsbGFJ+n28z8/xWBTqdVjum6Ncd8LsOTV5raK40D3BhPPq9
lkEzfXdemGMg7rwoLeRRmYYU6EFvefsHFD64rkAby9bGJL//IJm82ZsTlnwDuPCMeNjHyagEPC68
jvU/bCeSgn/lvAfFLYdT75NgNZd/MMxCorGOfiVt+cFx1jWO6qseqW6C+LX1XMPOfwKa9jZ752+3
oh2dttEOj1JRXWjChXC6ccmYMVjovq52eA9q1c1efbSIXh1idIboXJW9PcFzs6wvtmNqAi/4/xU2
AF07BSM39H/fY7Fe+FTZ6UlRRvYDRIujWsA0Rr79aq7jyBIdZQ+r1CalHs9hVxA42tEr332V681o
1YOsitPUjUzFfXIWoZBpCKkLI8A1MksGOzNEhGsoPQEEEXQyspRo+DHFbGCGosoW6oM1GdvwG7NC
y/3Luld7noT/gnIbmsYR2T3Ew2k8V8Iju5Rlvb2IL4HtZUaRFC8g3kvhdfSFWwhg74frs4+4C0vm
8M3ti5rBvrwsur6SrV+h1+8qjwaxYevbUB92C/krBR/RYIudOf7frGDshybT6WQNuNYx26uLMYvz
ad/ws82Ks8nDlhpyqSZwZUyrkyzJ6R2gg7rwvBP/UiNUP5Lxrrev31kVeKvU57BNG06tw4ekEjt/
pYLZ1gBGetV/DmBmvwqWgFky+CDUpD9la4wl6CZn4c+URi3ILeO9UJCZNzmxjh3XhW53zHxokT91
1r0P/tnMiDoCbU1YJNMc9zpxXetykCnSYgfVkykXbW6gUzqN0wpqaU7UfiqDl9GhE4aAp6hFoIPv
MMhQYqJaSKy7x0TQ1zEHCdW3oZnBtPK/O1Kud7dNt6Tyi6SaypjC5/NP6M8cPHtkMjtmOEDJnLZw
N0kudZ6XAK5mti/EVEOWvw6tz4/97LTkc/coPaHEWS8HHuNQJ8jJXoUsdewA+IrnH+8MfPU0W0Bb
Xne6Wvzkbx8CRKtCcq2sPl/DgL4UZQKgtFC094KvPvW6eddpBe/IFXyEXyXDm/SBYPgMsdTXrpXq
52p7JNB3dp2UT8vbZVPKwTRevpjpXxHSA1kyyyCo/Kg0PGL9sIb1Bj0Qz9WfIG7g/4jE9jPZ7Twq
zuPsAJWwFnEwdUW5Fym4YMjdeU8rTpeLUWFUyj7NC4xr7k2G9eRNK8DmYB80fjZMeRnQOQKRHDAx
ud+kKKoAzSzzoqkgfC+h511CbUoThroNNuuvpmEfhhNylcZEVwhJKVvnRhA4CapL2aNRa3EJvAO0
pF4gIgqgsAIHv5J1ioL9EDpvCSpiRhoJOsqiH+yAUGdtLygaEBZ1kz9uNJ5Y4rdpRH0nGCFjTezf
5pZlUv1SyTbVzqiV5gAMzqOuQmMVCetJ1ItjNxoY5NkKoXOGOIVqJjZZUmt/Xe3dvM1D6267DVxV
8LYboJF2R8p0om3ANAcHiLw3ukxd3CA9M7Re3kS8kikgLQsDEbz9yf/9pXbsFiil1MsGtf9u19Nj
5lh5cXcAJwcD23gh/kcrblkN7SuQ2cEMQbY2We/uBuC/5+y4ehwTbVfrKB4lGzKkyq6wWavrOohd
sTUXbILK8YDsZI3GbQ6i1ecF/WZdJVO7vP7Uv0RZbPRnrc/gTWfGofO2lwu7miVytRUCSOJmYUfM
nBzpxEPiHulwWdXTl1CJK/7MfidLLQU8lhhNVuvU9V7VkSdujF6qtaGA9mej/IMpBCJuOfr6bWth
HVpdTKSNphwN2BkyG8J+5de5WPWkulX0IKxad0+dStB6nC1542Zk4Q7u/dcQbMPNNM6UskTBPmb3
x1NIKTwsoUB/0SPnorm7fdIe7B37S5zSQqCcFlYkvrHqyuY8gXULQFkMApBu+KgdWlQQ7WvtYfMf
2B/VNQUQNJV/VJwjCxmMMoTyGE6eh8Ixgr8/qyMHy3/veMW9wyX7mYkdl/mBmIw2CPc0EF6YKwPa
BJuWSMB+R1ol9dQ58d+CuPYfmagqyaSgYYXhQAqqKpZj8IDp3a9POGhKfnm8stYAxLglFiC30RVf
dOPPTc6oiKB29uBqKaVAdF0d4uT75SZKUEpUYZywpRqtHO+tP2fSKlRKWvCDU8nbG9h0wAv8oW6O
ix3mqb6Zk4LfS1g2KR27ES6njXw8mXbZIUKuKPojlpopjjCw0LbnA6qvH+ecZYW0ylso25DE+CSu
+Uou6FTQUqVmUCtJt4uTwW9RkUf/cii7x/yAVyCCchueTEaUCRnL7yzmc2sP1x5Aw01btIwS457E
tJHCYMLdfxFhDw7aLbb//acLpJK6wzFvU+WpZeTh5V9ZRZChTeHLgmULACL4ceHk32CPhnWXnlXk
FOQSOK0pgjxnHedDGX4BVHruRx58w/o2atPSALVNlYoQUGj5fwJyUNXYsxTsbrXkFV064U5f6kkI
AozSTGargDjIZ/8Ivk9gism/iiMomOHXwQS2e5Bu72bqV+AleTqZkayJ/DdhAcfARjG11HHspOnm
EHwTXLdvYqoIjOVBcnxfn+E95KaAm8VzNeTLd4jE0AjAF+ospDKuDXlMb+ok3bycOqEMA1TBvmC8
TE8EIK5OJJl2k4SmMl8QRlfqXJx/22Lginn3iujHh35MGcx+4MJ2vguWzNnWEcFv3eiV4ew/LOOw
tEC3+mPW4wrsU8XqLy4n6RCKLByZA0+t7ZVfUzWaB88TB+AsJOhsCZPFyhq9cwunPf/N42J+N8dy
hgWQ+eRs6plrHJHWvvKdRYfXsRiW/vhUFLsVXqLNx9Z+FcrevOopsaI9ktNHD6EFxPLV07Xa4HpS
G25Kj3WVEAO+yJKuOh77XTvOvnlSYCdvREODGotsC+Xf3OUJ2s2A0pn/zMvq4GcftlDPsKxmaApk
mjzMzM2ReQEauJVrqnX0DDIv25kb6laGDEC8ceMt1iVcglb5ZVXua+lC5U0KeJOPyjLJSel97Q59
BaTLQFq3l6e+DXG4bXN4Vt1oaW3RH4q9MjRWDiJwpKuFpQzsqNTXjRA05U/3z7eiNvLWbZUF7r4n
jB0qAfouw1xrG7YW+2lSP8v8022HwHjAS9IBcyrUpkOQat+XSF1Jcrs8spu1qezQpmqOv2jlA3ZK
Q6il9QPTYXvkLqOC6LdHFmrYJf3KaTQmI+9Rb6iB01AiDmzYEwOkWdJARroECjFvKeLAP5KIMExO
jNbJO3odM3BtFxuIi7kRh1MNReJHktJzD4LXKePU0v/VuvRWAD0Gqv0mycCpjvJeNgC+ELGq4/fR
Pn3ssS0kX6r8SMQwFE+HUFpbvqrUQiL7jwlWw55hEjUce1wiPMfQ9ReYetG0WLvzFZoSQCeq08AL
9liWCCSDKYBAttVwJ+MQxIGcY9/PhuBiBFT6WDXsWWNiD0rofcU0IjDneCJJB+rEyZTvU/s8XuG4
nphzB6AL8xYSMhHBMpDHTRe2Y1uAqg8oJ6xi4k9vNkxyXOXEQeadV3heBH4LM9uIZ6sxj+KZWJUU
Qe//XNzNOrcfEcPV8jmf1I1C9uQtGe9E57+4Va+NHGpb1i76GLPvEZvSW9TfCoTxAt83+vrJq6P/
zT4IblzfPeKjB58yyb2fCdgBdPJz5bwCa4sDM/nn14pEMyMGOikCGfVtiM2S42trXhhO5B7QbMkU
BXJ0H+ZC5VP7FaqrAR2Mq6EWKiAm/80yfLWGYgcK3cZvNErq2nUNf6vEFVnfNMTte+JdI6gB9Jv4
OvN5D7yGvclq9+0pr1DcYz/URuSV2gUTor8e86s0nmrsltUQIU8Znnm+n5vqZ/wuu08vszVLQyit
89w97rbisSf44hRNPtgiRFM5lpLRgHYETAwKbbq1iQnzut/FrQS9HLqRbTIQSPCSHKz/99P9ycrk
j4eLPMajAAF9dM7UBQLB6gGkIfk4BmFMjn7yK+tWSmtWiBZY7wcWWHcr9snDTuAv9DgSJWTBaGK0
zIFSUz/68yeMIzVBw4PZhMB/V/3KM/Y7Kpr9wRbo/99VSNK4vswtlFnWatcjX4fqFy1BnyQKli6c
B1jxKUGyM3AmubEtBLSWgXoRy7n2Rkm4zJZoH3yq0B6F+bo1tQcWGCcLEYWystQmEYT7Uykq687a
ojAWFzUtFmQoVIh665f1nsowaUFcXHgfnDIyHZa4OLpUX3dlguy4mDocz3O0p82ERN2bLJ7x90la
S+fpsJPfPzkkpXAFVCnc0J20MRyAqFt/Rnu5Z+K8Wqd4iFEz8kFiFLybGAzJ1llOlnY3pqG7/jDG
QiEafouMycikQgtaNjvNPC87y+2iSF7n+r0dojHxxn/6m4LGQkZPf9O1ysqFwkjCa6X1oGc/xXva
bW5zJpUloxaMNsQARcPZ2+4DYRXRiOrpm9d4WjJaApJLI8Itp+Ttx75K6f10U6mBQQm5q7R6K3Lp
unTCh+tevr2qDdWxy3UHQedSouOCIsSNFn4w77d58lGdxgKNeFpx0epDsnL83mYDcD7SIEzH9kj9
Ig3m1U+aJmYF/IWuBEESW48ODPavKKCcWsZLY4AVdngN8dEbDwTnL4A2M582VpRoESlCrkfVnhJY
dVzmxUeYFEYVsty+SbIufYAU9mQAj4HsC2P4N/NDCoiSctobBXVPve5cijwO5fUyjsR537mPaySw
BJG2lJ8v/rwCaNzhseUHGEwrcMSMy4Y0dYx+0Bx6y7CaqfCnJuTgAwd+CduoAiMe/Btlp1CvP7XV
IPUIWhv0DFuoCwhL8YtqOcDYftg462Gk0mwRy1l7DtflHQe5zhDXCdtZ/D9li3CguZUd1HvQrySy
XJSC+cWM/+lZjov952JvKvOrJyujuN6pZenkB2LPq++vlVFlqXHWLR2TvDrrFzNV+Be/YW1JeeId
Flco0WrF3BAwOzJ2aDog0WVUDI7Y4uDWFqqgCb6inzjH2+mhmRkH2Njmn1yLYUM/+xuKd6ZqNyHF
ak16K6+b+gtKgCG5pFe2ZREAIhuHr6a0J5XR2XtpqtPczC2lcVk5okod72vBx6U2M3KzX1hARxC+
fg7LqCGjSf3uSWrcm/kY7AhnI244L8m35Yb0ld7wtpdhgHsYd3obs5UJs80/ZlQBUocIg4542ce0
ooYlXaCHH/D0CVYWocx3dfZmMC8i0pdDIpCw/AXg8QuNUtiepyUREUQ/9wNsnAexF3JFD8lbsr1R
iTGO8JaiBwY4tWxhes626f2oi63EvokEx7ZrukwTQp8GOTc64XWzT3dimJ4tmjplztDdRLBIpYrp
IYlE2/IAb0QEHUZpcPMUE4Q1juXd0GGpZNvLrrBl5Vn2cCN6L9ahnMb9CUAxr/w6Oq2UuwJQJXge
rLCFqGJ6j5gEbEdUJMO7ERU74abzoOa+AUypnbXQVZ02qzBHIDDtkuUegcwBnuGqUHzXgf/L1Y4e
dj14vW1p67Qg1FyERJqAaDOS3vf6XhoHLHEkyKYFfnQ0dOM8UFImFUbdxuGQBTCBBp42nFiLWtlV
igpGLQ1v1//1MypTGLg3DtER2NcgF5hWoWFC+JcVycTxqr4qFc1+NiRfmUzKNX5GwfQ5TPiPngha
nFIS56QGfTH3xn6h1xluUC0lXUM96lp8te3g14arxMEfAcPMHOpUSwo8w9RAh1Fexuim7oy6HQqx
xg2xJz6HD6b8wzSVE3IAcwff+jR2z2DeOkvvJse7c69w4ZDiGGEb3aegJVcw8dv9dwhZT402kqNw
TpWetVEeY0kG7ajdvPpAOrOmK7SBXowTX+oE1YgJGhCJTu2Bh6etYRv3oiAt9713hSK0FEvUdfUv
njseYDlPjcZocYdtVnwOXoEcV5Iaiy34pS4t0u933wUH64xBd6WNIbHGmBAWqrApXamRRSJkag7a
d/wAGf0eqlDM5pZenOpPeOVlUOYnXRsIZPODuJ72pFV3NzYTFa/fzYvMLXb5vIRXjKWD13wLNech
BZ2foei+eTrxqTXZw8GS016dhINVigrXEpghUIwyKGMUgYulhJuIJWif764WjFXXuFwb4ZsXTG0W
hm+T0BwRwBavRphHkV9nvBWitBuMmkBkJqFEIWJuZT+xZk2CoGlYrchSr0g5p+9plBv9yVdgai+v
f4T0ZFMOs8gpzEd+/UnyDc3GjR+1N49GWfubJouuXwjoAn7RWmbnFdLEuNgz07s8EAzOBqLu84XB
nt4TSehsp8Q0jci58Ib/MUUrPqRyvmdXOmUo2NpPafegXEynN6XcvUo0fhTrFGMEywjIJU6tyrgk
7IaPX0+3G7XLYdtfB3cBzVnL7KlS1eJWTIWc/Z5YQGVAy922brXzJ9iviufbDAojgWlC3Dy3Eg5a
LgxFg1a2e/hb5vFm+/ZCPZz50DwbpqffTU8pbC4wE7NcvEf9zWSCO6/B51T26/36BIQy2tMZ+vyW
1pC0RWRUzgLfiKMtHWSmsH19WWeTtZW+CEzleRiDRIHaojqlfhkhrImXx6gQUOIzDVA3yWUzPW2/
2qkreIiPykSv4YudU768JblrivUplLASIHfC8T0e9dkIr5H1n2EB5rVeU2VLm3UwJawrrTdFeOuD
oOVJJ6WSGgDnvFPN0X01CdZlgbMOth1cPalDIe2fhkw6QAzzZ86bk2P6h1C/QiTKZwSfxk+mh8iL
Ocq0UQ7ynb/93SJVbtlgupxWV1V9VdTomDl3Nw+wUauikAV30y9tSF4Af+SAiHTSnCrT8w9Du/+v
LvI8DKX7PDulaVPFg+AkSflonQ5Sa0HnmUjs8Vb3d6YiZq2wBGeYmJiyZwiF6zc8mL7OapgHYjFe
D3c5m3VrCCaRg/WXCP5SJKt2lU1OrPw9t26Snoe4+kamvi24goba4Up1CtmOPGfwyhsJYPkULci2
84mfzSzDcmNekoJuIUzG3dlVhvxVqo/e3/m6nWnsR6HVq1jSUaFwj5rgOHPFRptzuEfgXaM+w+ar
4Gc3UJa4c6oe76uY0au7mHrkQHKhgNCOuWoknlwXR8XIQm+BDidUPdvYszkR9+yspO1H9xtGhrTD
UZkZpmuxz2U/Q5QaN1PvuTzRmt+63TMWZWkrDo4GRhydekIqfG6o3zZiXqRbvQoRuAeq8L7zie9R
yaz0umhhN/deDsi5uhB2Qkn/yn974rbEhG6gRLAONmbNHxr3SUSa15JEGGnKBMwwCfe7c8O7oj9T
1CSmIml/UT6PjF5VBlGrvIXV2VjRhEYH3S2vL05a9ozlzapFfFfewh5SrV0dlq+fPR/TWKMPZQ2P
+7iWUGCr6DOTR6ecJr2y++1PBbjDpg/8UQVI8dKsOtT3hU37NSe6ndoYJQ8JUB5DCTC5LHmCSlUY
6MVi2vxej3pXSuKSOzwYYPfq9BIFy+9ZWmpekBi37izDrA9PA/tVpW6XebJu0y/NrOVizPgNcHRQ
DrvygPw3VT2DzkCPqu9WniveWzQeWld3r+nOX0Mh6V6IYWjzlh/9IsQtXOtCJr6locuj9sVCglAu
OFSusuUt5iNP0DGS7x2qqqbnMlOvwOCMEyvGY8LzuxOBacanVMG2NSm8UDJbFexCKg54AmkH9vLn
JByW0p0VlXaboPotDFYE3Ic9WD5bHJed9QuWOWM/vpIuB3+31jhlPBOlVzjbFyDtGqMhC4CoF308
wDZQP90Sn1ekzHxKxeweqwSJ+7jB6V+eOFba/+vN0VCc09hqR4KNh4UeZYZYrwWEcyVdUWkEy76L
zdO+pWRlsueidO8i6whJ4Q+yMR6prV90UjxlWQHL8KoynJquXxYMiJFlK0uRmmmgeFFOOjF1DkRh
KVN+46qRTkwWW3j3ruGpN/f1gSdg0MX3lIEry7Epo3Jow1GFWHKnXbMgCeI4o+HAOh2SZL6KAxM9
XwD+BpQuo+8OdVWtge/VXUo+brOayx9cP6KY8Ox36B2rhmeRTSHEp5Zf2rUcooNeohbqnC1PE+v3
qGnjHlSAW+HpBurTpjAG3+h+rWZ6+dermN5HdUOaNouC/Cqf4BccpTuZdEKDi1Ey7KlpRmIp5etr
FvX200eX00D+MTgVuNDs/s+vtWw0LaooLlVxAcbk8XmQB6OL7+oeGDAWCnlRbky/D8dqPeux7BYk
Rb+h79tnG1lTI3sBDlFEvWf2Y2dUexL0rDAZDNyNdHmwTqW3j9HxqI37B2gFov4CilYYNn1R5lha
Ft5axgKPTx8OLKKZ0bc1p8Eu+nuW8vk8WPGREb1GQHfKnvmf5h5bApzU6OMy3vXEk66sZ3wyk/r9
8aH2RrKKHIA3G2X3GdgbpC/WddDasbhGcZKO3cF0SQJ0SFmYt8AWaXIGWzknR1Qhp92InvFzpac+
YYRQU4xTMdCLXAnQ8wGqGFQ2E2dwllXYY/Sb7WWxEVzqnk0F1EC9COcb9uvkvEI0b+i9KbLWenMi
vA1TCdyGQ153YErWCNNQlbEHqViuGgmpP7JF/aba9s4/am5yRuI0Wnv1hp6KzRzhY8h5WnnZEAE2
2M7K7QmSY4eZOhqFM4sWBQvB8vrTL5NWGA4z3ku3KZzK1N193KpoipmjSRjewz7aW2K1/FryJYV9
Ga7j7ApuQZQIF2RmxxQtHxqrTWuluRPjtesOHLPkusRWKl9D0GRuPxqGScYKEde5zG3zsMH1W1U/
U6bBdqBSZ0PzGDR6UkEVkz5onrNeB8OXYSKAu2yd2UExHuhlcRk58F150Euu4x1fejfUixut9WGB
/XIjEqQo5BfgR/J0PnQfpR/MN+SFgn6jNH9hMIOyxvi/gz3ldxqcgaeI+911f7DvaYTakNoCH9Yj
1B7tEx2HSWcJfiYhgoqPbxvepJHmPTJsTp3dmQWoHhp19f5nb/WgDs0fzWMtBShT76anCM+YyAIL
5ULlt0fu9YX9N5m/Vx3VYGp+8yipiHlG/bWUQUt4jRbCqYkf2Ea6b0uXfutcQKyqfK8khjaNNbO9
SYCrBC1czUc+ax3m0Mw9wYBWEnVKCvTQmZpDKomL7R4KM/HDykUHHG6ZYzpdCfMvHxA//dT8/D2I
R32rI8JZoMMlZtsBm8pm6Kkbl9q1HLcs0buRMjjtuKl75nXFspqqaawMdyL4sT/YKD1A2h35EOan
mwR7lmZKxS0UwueRt14krGVavzY9zz7efTCh07+tFIaEoj8PVvrTy5jMyL+C1BH14FNdOlZT5QFO
OiYZGUwG6hL2pDSiRvZ7YIc+CVYFKGFV+SkwGh0uUI2F/3Rre+5DCjcK2AzI7L34gQ346lohpQ8V
GZWGIrvIes1kuYI+KryoVRL9xJ0uUhEtbS6DdNVULAD6ipW7uJ+vwwAGpjsx5uuM2zwMVPWzqSn7
bsCv8vYa1bCLWB7sOLKk/btDBRzBoLtvKhN9b40S47O5V7JsSMZ7kVD0NONvBIhbmTVlHQ5QfA2Y
QgQJLxAL2wSsZjeEYWulrtTpTYu796ItyiZOBtBmW6wHYSwuyVFlz45bWD/qIsJUyVlxyjxl82Ay
WDtT6iFfmclkWQJ6Bfdok+afhX+ltf6Aamf3OT+Y+gc1bJlj/INz+KlJLP6hpbnuZrka6y/w85Ze
QFQq1q5swUx/dkUgPZIu3rJuSN8TahrZzDUM8d33k/Yob8tY5RYSlDqiSevvwMkfVKx88qiVZLtR
eyPVV4V/PHRFrO2eyR6hOtQPh2pjaQcNnare+ssjbJpe8tK/MuBfpgrBwEqm+ZLQMLdSSezUOKWZ
iV4c4bbrM9o0CvI8uijE01YlmPX8bNMIPfEAVEG+8W60N/N12T2DWiieJh+iLdnOyNCjdmO8i27J
wTKXHRyOO/TXVAXv5MMpRc8ppjolPalfZub4EKwfVe5kwUA+7ujSAF9BeeNDVBOk5OSS88Rmp0Fd
wzazUcq7/S4PqKBFZzGbJBRBu2lTQdymDGfqelpfawRUgLKae+AhA+ffHxARa2LcLLplffKjivoi
w91huoUhIyLqk8VSOD5mTLf5xsQeHNdT+GFSTsKO92rG2k07A0B+gkptvMqOySTtg0hKU9iu9Dga
2tli1VZM+MFwt+rB3V4B5a46Py7EWGxRSsylwqMXzA+sljOP5iM+7ObrRq7KzKkMu7GxyI6bkx37
6WDzwni7GA71JSLZSuVHQmpioBAZZVMfaR/1PqvOxMeLG7oNhUaGZm6EHG6kkwR8Qn0PDSNN5fnv
ZX35N2b/mdzO8buXojRAdkTxFMOwCggYj6cDwZ7zaPbI2IRACVNx4eftsPfsns6Uf3VTQT4U141n
57khySkZAunnvAw9XM8pVQSlmzajT0xZcfycTOJdkgO2swnqK6rBnO2gNdVO/ejmN5VlXjLx7atl
34DL6EeUdtOIFcBohhS/2s59YNa8luHC1yMpEdtp8r9YBsgI2Etk2eQyYDEAZzxERNAxyZxfKb/8
RKjhNR9HbHyypaImhzaMMmY1YbGvIRm2rnzHli98qxcrwmdGUOFoYUMT2RJHeGSRipUCskMTh3lc
dW9pIGavYNr2Ot3e5Kjnp7oJN4hBjtMvgDO5sH46UIsmkMWa8SmZiX0qAzktUcB649YYiHF1Lz9n
cZwfICRESyhO/RaPr14yFIsQd3wylVCed6vLYEnvctpeNoRyWp2BNxDTvefq7Wtc0cW0w14ulfgY
4z+CzU0NqVLMSVsBAiH9n6mx96G4ZVpPz7AAWpFkA8ZdZmw9+R6AhW0sgl/AlNHASWc3tP8rbh7S
b3hycv21qJmJ9+qF+wkW9u3rHmblS/RWB0dY0HlBjR2GKzExxs293XEvfMqYzTWwDuFtmb0W83Lu
Kh6hGg9B4Y0dR6/ju07e/ovMtRlnRcH1xHfX9sS0vgdqNmEJSdwrsk6yIDWqowv8CDCeBLgi1xO4
Mw1bdqwhnhQj0xB7qr8mCOazmr1BVpvOaY8RKJUQoOIsNUbNI4Eo1tprhmQFD2CFh8vNZXTTo2ic
a1Mq249ISEB7zIBzPDsIG/yONJAbpznMTMOS6isA9TLru/ob046ERyrkwK3ERm9qOsxg7QTU9fyI
fJ6K9bqUOYEJe98kmuoX0CU9CN+iGuYkXPk2er0qHri8tVDQEjb4z0yvt1CyqFQASBK00Nj9nXHD
Noma0uJtPnvmwwmnQCAntHaGVuN8MzHWGarjz+wWnYa1Qg8vPY2E6PLH/1YkbskIQk8DLI7PWwje
6mWHKZ2eKyKBq+b+KIH5LawR074Ap0XsgYN+/HXZSwriVHIaMwd2H5vg/mfsZVSU6BUTbxyj0uE7
zN43Wa/tOEmw36IZvS/ycGhkSuTYkfIvQcIS5AJMTrixTo6UH/6LpBt//ENh5vfgA/c85vHiouiN
WGwYeSjuKwjoXGkgevJB3c+2L+nGczURiBd41LUJ8nKHSSnA7Hut8xeVC6Jht+fJmHMiq2tnbN3b
HI+Ks37j61QlSzcCiN9UQxvpouXHgYrJ5+8k8bLcQS2YtINcAWw33h9DDeiLvVSKXaZFZBH9YDjd
FEW9KZAQGe2LmxbD3zYPBdDKknXB5utnlLWwon5zb385CklaFTaOM/9kTGEBe0hIIRDnlD9XlujQ
3UEGKwU3N2XbQFer4QPkVNOQ4Hp9xZacrH5G52/fOvkZz44CIjwamtLHMHOPy2fcUHrtc7tUHmH/
VeXatMOqM7acZ2HO5FYt0RNQrquBEsXnNN7ZLs6R0VLiaJJzXz1zjIZ0n1UZS3Dq7J1SuKtL+oq5
XiYcVkLKXbO96YXokqYnQWkV5IbsDjs6oNgvJ8knp4pvbIp2GMDhUWOaP+H388jdrEFiX1IMBnK0
o5VjGIs624S0bffRcIVCAw35Jgni2FUcJNJHsuMT/KxrnjWfR2T9eARgEndRhw/NPqb+sRWahGNV
Kl7pSwwLU5NMuYLjIwRAvzP8d/rsu47m2RC0DE6fuAwWl/UbBrDNI50G2R9Y0zPgpgIPIvX1Nqwd
0AkQSIo7ArbJKJkOdixMqWJHKY/4ubzdzCHKmPnJuCegt6mzI++rNAz/qx5EL+COpYviM+YFtqjD
ibgT1uUbrIemb4CyX1tJJ4qDlb21I41aof5+GO4xElKZFaEYAcQic6KMy3hwcSQypS2KbWO9PQyb
FCkrefyDXzjRaz8MYWX6CYFyKID/lllG/2gaUtsZQpzG/qS4Ws4QThp2zsABIvcuVsY9YcxWsNIn
IMY7epA/vAz2hmg8GfePKmUY6i9Drd0C1GNCriAAVc/oHXYLBtfbHNSzfG1JdQsQulhXWsLE5A0E
ZbG4d2mjawDkmbAmlu3ISGzmR+5WaMyPjzMUJoYx0UBgIXfPc782YEb1gTRM3dmrXyhEGMAWT5/U
8CB5kQzrERrTnq3cLrTaq4l2HFD49PcN7lqo5RKREik2igZ5IAZsY1WZPqFnzepn514Bae8nugsE
zxJldMGGmZ3pxbQoFNenNcQcSgA4JdOX2FbWpDU0861pb1gXZSbYOPA0zGxNP1vy6HwTsugaoZv1
N9aLBl3sy0u/UJT19g0CUxPBZUl81FX/jDMLlq9AYm5lOud0xoY//hxyz1ksYxqhebBuu7Cf7qxE
diho+D2LeNOT13EDBJ8Txe3Qa6lYnvQcamaeRc7gWEfYPQDYJKeLvuiDggAPXgInEWbdKq+uBUU1
iNlxes3Ag/eMKyRQOIo2B779Cp26T0xaGl/SSlEh+T9uThN2M4uO307CQ4paxAF6B+Ue8v6RLRZI
C6615+vZNEExlnH10vSALipJ1seAKYFuvY+QMyEbxGRAh/1PLg8aXSUmvrmxjNUtIUymVl2u+pJr
LAxHpnE6ERx5nF+CnrrrAVsEer0qfDVvstF/CEjC93uFQ44cAkvPJw24LqI4kSFaHmh4kOCMLfmk
5CHF2QEgEzHm7CjgwZ2+EWaXd5Mvq2utWITyaCK+e8fQx7haaXznAQzHM0rUf7UOxZj4VKfsxNIv
rKz6S+kEfz8FeYMdFXiNH/QwjBFkK3P72l15073U3NytYaBgapjS/DsF41PzLSHtil11AhF2of5A
62TB7HuP0AO3LEzmFlj46b93W/arzUeJb5L1X12mHDL1eQT6GQ1BmIxA0nYbnKo1dcKnlGwx2U1I
55cvDeWkVgC0XRn7Oywhi6j/iIR+aFdaiBg2pmcJ5X/8MbzF/jhnqyKX45vsCc4FXNsXa05bBm/I
nbZ4NEwVDzZhuiB2Y7wSNTbQnmlAfsAheC9+I7M6WUqmDAgroJG0yW0/uoqiUj11dDeHy30L1NHV
A6TRATYAgfOWOc4GHAK7tZouNi8DrXLK6krT8z0AfEG/iUgwxna53UGYrKdhuU9QQV9YDJWjCKva
lghEB02FFfIK9/3i6ByA+onp5o3J2coGCi4+j8XkUmFeDwwdZE6yHSLbpkzAL+zKyTxzUWQPEjPR
Cf0Fza9x8ndeCJ8Fg2gIkWG1kIHBoAnfX5cX1BxvUpZpnwpdDQBODLhdDgsGn/KbHMZhYRFBPGtY
GiPqrdtm5mFv7Oju3qNi+ovN4SaaELhfTjY2ZT+gXfg5iROpFhGqxVEQnMImZTWaUFgsMmBEAC+i
kGgPmyNIjRXAJgSy7J4fSTYeYQFfM4xoYBi1ygJt3dsfDLh5C12N1QrZMCyUBRqE8j45Yh+tQX8Z
bwjwgoWmwkGAOsqNiwBy6cAeDcrmHfIoUoKhlmcPfJ7EJZkPNNj9cS41Asr8VkTNLCDZYQ7nW2N6
JzJADARUYueTPosBEg/0KFdyyke8oMUD5pmIoMktHkbwmCHCRD+bPguVBM66U1fklB7SgZYyuh7s
v1RzUJxtbd/5eBSAvIgZMgGWJsbuwBz4L+AZ1FJ5+O16bj8HV7zw6FNTRyYqizb3W4JgxvDuI8EL
vjOpqEKFRRERSSVcd8URPHEDd7u4iHDl1aT6KoHvBvhvCLFWO2cG82iIYPFXRZuf8jzYuVvSX+/Z
Gp60j3aQDqwTwNTIVuELtaWrbmhiuyuN3NlgGAEWdXpN1fbTZq3NsgORyWZpC/UcPUy3h15UklT6
87Cfs8PIp8PIIqwzhFnRB486knxjHFEkZALIdN5N2eazS+I5wK7sHAXu7s7HCZPu5Uoy3dq9FNol
M/fs28R42Fsh22r8vo1nfhKvF0oOR8M6/6pzAeNUCQTKjapzRW6/4L1fGBFle2Iba8DEcJT/PbDm
wrSzoUwC7qDqKI2OiKtR5DtsH7/EKNwDIicdgv4fFU+sh59WbiqIhHrnzRuGzkn9N01lsp032/jH
Y8Gr4nWJa8ioQrarEoyyO0oJy41GdZVYLRqCKAlDUyc3zdqVEsNDZ4oSfyUUe7V6ixQKhxD8YsKo
RWekgC9NoeRMOye9kKNcHWpzYBUbkGZDwRfTBG4o2hVNdnrRLmJjMUYybBgku6Ld7OHPFHkfW+jn
Yyyi0+7/ne7sI59wADHHPI8/M1wy7dOI0sT7gbC6DonM+z23BGGUHxX5XBVoOVspRan/o87NeeHf
4FJzVDnhfhCUqhswfEUjM8v9S9BAElwy+wd9pnR/T3oONhENEIHBHgD5h5Mv2Q0pQHqO5EzI5CkL
Oay8F4vPXc8wpVZKCIjhW0kWMmzD6M8trLja6On7amKylkn4y3muTqZ0s5oavCxsuZ8A9MC3uehn
6V2RyaDsaGTHzocr20ARUJDC8zrvXGuasCRH2K5qVWLBtf8y9h4k++5073WbH3vjCGZrd+am3QK6
75A0HykoFYPNZM9RkDHQcAoO45xgd8CnMYPlkbho15ab/tksrDjKsU/jCyuCEeem95509y0x7Uw0
bjSONNSuSOI2Ezl43nkI1YwRJl5tFhs3WeFxpBNgSGPKuVsOwe6dlL2T7TeAI+1OJWRe5Zz8bkOp
fos+ygTf5s90rz3Bw8sYcgaDroTai980pVQFxPLbFLgcahVI3efZppO/WgCK9GjvsecvUb/vY/aL
T4EODeD7x4h76Fph7a3EaXahCcR/4D2KtYvXFEZPAFndM42X2UUwOKkUFPo0XIHnDRR6EjnM71pB
/h7bXKEG+5/xmin3L+E3m43WhxlTWpmjP7Hou4KQZXa0x/hg0RmYqssjjvlmhV79nfrnfruKFwRX
e/wDPhg8TUN64AmQjylZLdUuUWDP98OOpM7HfOBX8H+aHg+9wf8K8tSGxxTksXytZz4zbRIAImDZ
3MPAJEwqtN/1ggIw+xAiysKbUo85bLu+oHT03oPeOiPH54tBeR0ad478aOUeborH5NweXIzAK3a6
kxQcJOyV/b5/JcZXqMc3r9vyld/Td1BFv/Nt+V3ZoFZFhrMmFpUQehtMN46661tWIlZyD/kPtSPa
nC1ka/eVwbhaa3n5aJtRid+1GhPGuvZcz6TWEZ723m8Z0np5xwxA4RHITctpBDJPuZtKAzy0D57K
xqj3bp5S2GHYEg5GmuUiNoF1ZDOPBQj8HJbojYO6xFPw0Q3bcYM0p3Cujy3lQSwL9DrwkgcJhFgs
VlgczTW5kStRlIJABSidRvoC2pAGJHCkAo1jzaS5gSzowGSSlWmPVNNzt1BCog7xgrVQMzsOzgsb
F5ws17mth1n5W76ZdV+oZB0OmhjwwxsQu/3uCC3yJFroKm9lCCKp34TUciw5YmOP7eIxRn+rLec5
RKs50NthTI5v7tbiUT2qDhI4HvJucwVWayxs0PbghwwnNwP6DM+92XYhL7wtiAs3xdJGXwmLC8jx
h2qwfQh4qGfLdHbBxIfZD4shEC1ZSNrEHSX3Eds0pFX7baxOdbO3HFAuS/wjkGQUbJTmDwI4g15Y
+6WNLM6R4oVxP2JHCOEzRfmjTw6JNK8hxkkPVgjyL9FTRVG0Pn+Bolq3U4Sei0uOMlxYHN0NWi0q
ZgXOgVnM4Ver7GCW0/iYsWxuaYDmRbOf0d/P3wNEJfr3ndDcUiXIXM1zPvQmvw/noa/LOoJdvaNF
ntTd2xD+qgGDbMA5iaq5E1gyBMXpCycHGZLjdLg2GY7rw87gYYicALuKJJDvSUeeHA29SYDkhXVb
VMoiirXC2TUEq2aLqVy3I/zxPXxMAWovGhyptLy36Rc6yiOZOkuUUFoQ1FkjGHxKtH309kF51Kk3
VxX8Sn1ch3p5DLYEN4dy6mBjeEQmonLt2BXgQG/kT2KY0IXkWjv6Ns/eBS9bR4AsuqYDV0g76yIU
0jbNYhn20h2s2CBb8EHR9I5Yo1Tn0SOPRb5TYmpp2+8XT5sIJJPU1umCBC2fpOG7Jxs6rJZGGShb
vSnBRm1I8ZU3VmPJV7vU9gHRMJGVr+qsuTSxnNjIQs+wrhRSDIATtm4K0dW72z61+mc/2hU/PP4J
l0owYTMjcG4mmcusIOM/M3gnUGa0QZTZ2jiisSp3YNKj3Onkq31C6zQM5zVJnfqobijrW5Ys2ysr
rVTdlRtDy3ILd9KIhQ2V0vs7KmS5uFSto5xnYD6k5IoDcZ/dSJ79ijAXIwjgNaFYZ1tHlCRXUwba
4fIJ/ax7Hg5c34vtEanHzLaRIEtyRZSJpn29iPQ/VNYGa39fQPYJhK7ycTrjrvrHHZZ0ok8qnG0i
PyP73rut75KFdl8r+qAkyFo+KCzQaVhm7PKPpEg7fO4yUHgeocWDM9nIpb3w2jfqA3VBoDMnJnZc
3TVjbknFbgiQQeR96RsRMIWznWtpfjdJp7SwRvwHBOK9Mcm482nkg0eWRdh8ZBXVsORTzIJzmrss
xi/JPMEOeCQibcSsGQ0+OAKh6EmXf8GUQRrwURx/upWnpnutd67qhG3c891wT+Bo0iNMKmQUIMFC
0ump8AdcFRPLz2AcZb1LukYMpoILpIxA3u8CxJnnu+6caOR9aKNc91gsgsOiL84tFBHqqLiFMe2T
fAJbL+bxXPP495Vw8X94Ue04Dagy5ZVdTQuVdDOgbQ8YiqYbpDZCoHqGjtHxcD5xzMfeOs4gggUg
xg+EgmMJhk4AbKj7SSdTolbMlOmidiQjjRJoKV0f/rvtbhvjM1UJiz4j1eYXLNR9C6vgU6hEZRlq
2Im2GSFUJRJneWLvw7TCH6cP5P32ncEoFdCgyhIrsZxqfnQKeRHFh2WNHfcX1W6TKDsEH6SMMN68
ggXHzyI5f9Mfb0qUq2cPHU7NVWxTOqQnmFtkSAH0Gp5I9uD9/ay6U0v/Sv04mHM6noTDUJD9K1cZ
VGZ6JIe59aoyeqhje0JpZrnUDsVNwuUm0ec2TXSFPeeeAVuv5rhw/cFg/xajxyc2GQnqHgmEYnv3
ogw6Nt/1FYwqAXMqsLs0FSbG3Zj/2gbtReyEYEx3bjuDeejXqOTYyTVEnCpIHZnbylWgSO9TzvXL
Jv7jDiKdFIigno8W/XFG0qavXkZl3Km6vYqKWvH8fanYgC+lGplaP7X2jXVy3HKAwGyEWMYJsTyJ
gbGt9alwDCqUWFAeYi9PMkSNMmRRkKkACLguZ2D5WsVpOgq4TS6gMEFq8S9WFhOQfy9OhaEfoZg6
C6jxFUddwj0oGzS7yVZJybpF5zA+KeEMlYLz52Tx0k5C533nwiR/HoTcola+mhY6iE7NmhHmUMkx
6o61dUkrkh7uC5CaJ6z4onFpJrwhmNRKugUEXBXJ75dcJ33gGx0SSlNSD4cCqTF4t1Pt9hZccc0t
4xeE3AlrwCEvm0cefaA1h2sO2n57D42U6HGZq+fYZG8jMrHmpLhvJR6ErPhg8+gd5LBxGGjjqGQS
AVmXY0ClkuwgXEtrjkHPL1BWEf6anJ9P8PIaiWpVh8NtjclmC/2G5PtY01nd+1Je6V7AkBxPAM7K
yDqxgf5P7mbLekSR2+P+wbpVKKND2lspY1Jia6ftnCaJz4LHKaa0SjkT5Np+ib4g9WlaCBl7FEm6
qqqzSx+wxkOMdc/Cq16weMeabx0iofDzaCjtoz9FXv9XBWeyaxmQI8jlkYjxYYHGB/+s37/TcMPa
uCxSWc/woz6+bM7C4wDZ80Q3d43hyG02fWC1Q1Bef4rAYycAwqs+seKBbrwln6RNtzdRUVA7jSu5
WUy/q7jDY6VFOQaJ5AnLit8MvyANXD1XhhOxTFsKxj3pCt60asQmtL1vyZzr+jfSdwX7IB8iLAPv
k0XLlL5FnfbsNBlk7w0oZpHFLEtth7CnXQRyoDtSAfvjJ1puUWyZNpnS1ND6y4TcWJK4UzyNyYLl
UAi5JySlx165mXDtEerHNa8BxXxU14aab5eoMBpxfvmEw+0ZV00fKahgJxTP9DmA6LoGGRxUf0sl
FKhLVKWaE5eUu/IvzvhpLH6VIqq/gB0vJPvndUtwt3MjrVw7pgzlOy4QFK4KDj2zruC6oFkk/Udv
m2AtwrCsxk+1ZlgnAEtM1LWUog868SpWoZ8CCCcFQHLHEq6mEMUB1VDYsj/3DTeF+4qpEjs5sxj9
Czcvn2vRF4o7VJET3eLNMlS7dqLgr8P7gk9zIXRdji2RYqx7PdKTyJmnpcYp5GBkqDnS0WDJarbg
hF1qoYEo3eq7aDLAiGg7o4VxSo2HYTHWSXi8/ILpD4ZSLi3Q4aqnRkAe9UxUE5biM5ZaLmZu5TBk
3ogvOBVA/ZzO79I+7g569OM/D442fxtjlJkcI5AH+gj+wINCx8uNy3y6M47zr5FaH3NYUo3ULUgr
FZymIKXlY9bLdElCpF0D1UWfXlC5Hp5EMjid43oE6e/nKNc5RrMGPFVwDiUom96HNB2SSsomFFTW
w9Mt/zbytNE3rvUcat1AnqXRlPECegtfe4UMWIdlO0X0pjtKQMsqqZgQ4AwShYNflczX852vqdqS
zq4utfwQDnXinXVZJAShSzcCNLufJIlJKKj/VpiY3egFi4A/M0p782u3CRJJeYmozYMc1xaPVjSg
TIodySEFDZKVzPRFkhsZdTZp1h1Kc3xcUqrr6tY84cMNCu+fXsUiScQwM/5+w+iuwSCfcD7V3VrW
+OrSq1Q4p0EtSnMf/An2TKl8ZQHLZytPBQgKCok5t4M/NoWhq2jgFVp9VyO9cgTNG7AvFAKB3z1L
4PoB483mvxt2MiNkFHHz1Ih+VBqzhgSF+pRy7madj7VcDX7c6ByLx3tDNV2XeFievAQMmKtxomj+
t99u6j5tAt9t0gUnCCdO1j8Vpst/+RRGQay7rvMw768jrosA0Kp6kw7dTD/h4HwqJvEVfLvepz4q
Fv/p9Y0yeXw/qlGUoaR8Vh65KFQ1fVRtCZE49YosSkjTJZFPcVBGYd52VWPgJ7WbdNT1uiu64wPn
vzlHETm05I28MGGTbFjhv049AbfU07jyl89zKBBlF0BF3m3ABkFzq1o4eUe4dyTs1CD+k2/mehp3
AgYUKU7HpcNBn1D3V0/CnUrRJB5j0sjaTqrz3qs3OSl070AYkRU4LwR8mAX5VZrbIiGUCNt5uoGj
n8XoKN59du3pv8kqg1dRamgl6oGnQf55LUr8b/whTXCNjM1LwBTY8u1v3p6bhv77D89IbaPjzlJs
3Qvi7i3NYHwcqxxukyDIpsKqN6qPso/ZCWB6rehHUT0CWPEdePejTy8RTdssM3cTdPRTCc5oLpwo
G6SRP9jRu0N1c68pt6GRiiB4xgbyn3Gg5fpw49ltEfYwo76l4vXc4DBFyB0CeGhNV6LCSTBP5A/I
ZYuu+YJ7mDukdWJ0msx9Hs6vltLUuYvsBcGFRLR+vxsr4aqK5pDXHhJ+AUCQsr4xhF2enb3W1xDJ
ZZdyOiA+26io8R58DSaXC1CxKPi57/5eBKiX8UWZ1vS6o8RF+4ieNovRh1jM6qPkco7ppOjB/rVu
Ona4AFRBkplmHVSLhiudLk0Dc7dTWRdN3+BncoJe0EwL2Dayq8hqeD6XTz3516Wzob/T6xpexJNY
DYdV0VibHqQI8MViKSM6YIb2SNZtQfHcf2Lrta9cEgj69rMoEZ0zFObz97m4EkITHPzdTN/bBCr3
TWxcqbhJBFg3bDx6IodtBSEsVt4dD7bpr/q1wZuRM8cmqUVhLDu//VqSMUZnpT2fJpH2yKr/nhAA
XW3+HMveKi/iIJ533nEUWheHkkvOywNYCLAHJcj/V3vTeryGPWq0O0XDSXFgl1rYglH2wGrZfc3t
ru5m+EWa4Jjeuwk/BcLcXR52yQgFw3zAJGswvUoLuQzx1rIvytyjXjRPWEKwRqLR7M2yzNiG78RD
XMr0P+faDId/6ANiWpuMl7riHBROnphlmww7cpi8Fy0cxcGIvsVdjT96Zp0JUr76s0p1+H/orYcz
8B7uByR+e88vxI6eaj4QfOZUHT2C3Gy+OGQeENCPm6lU4HzUBu5m+wf8yPoopYVfbkMtHOVZOyP8
Qc7+0hlhdX8ZU4AhslBD8E4Ts5cHp8RRpODKn8BP7gxHyhycsWtV0Y8go8qyyDqjklI6D6DDHVib
t6dcmi0x76FN3XyVTBFI+MBKSSiwfd+znXCPqlua0GI3d/30sbojsTADEgLJof974rYj6shtWYXP
8QPwNjZ/M9KTVl35NwVzJoD5D4FQv+Z6/wwcSXRKT/xI3v9U2YPN4yc8SQiIeGLSVurNKjQ6zKXh
uAbvwWddnvefmEeOuvShsXnSwhZz0aLJioS3OAoWh2Nso7TLqntEr0oRKgH1munMcxu+ESC1aCV3
2Rq4HXKSO6HI2bo7p0rk3qBUwxD/iBcFUSOX6pE+Tr58E+LSoezPRv49sZWKV4TLtO0dDz0teDm8
zooWo+N838XCZaV0N9F12sL2nCOjNnwBGxzISIYflrGyiDEcazQBkcNkwJQkwGx5ketr6rCGU33r
DHJiKh4mcxMB2tdA/oFvbzHqLiiiqJyTTvh6Tj82bn7Da5sbbyJVoCNHZyVOXoU9iqUlRsaSQYPL
nydbqEH43zgKPUpGFt1EJGg9O+AJiB6Y8re+mKJ5mZ1vNW2UaMKu1vdWiXUJrIQcOGEBX6Dc+gaL
plMfNOXIqK4h8Zn5G9dU99V99I5Y1Q/+hXAKOfUp+zVsq11jTQQ+SIkqIM44HGlIK6c/zhIqnYgi
Qa9eL3o3qIU9rEdn59C2MfRM6qFJ1mionDk7nUWUY78fA2iftAfmu9XjbSEtzbDCT6PTxn9A8rIl
m1ulbXrTvL9pWMDh+hAkR+HKEU9LOB4Gh/cFpD8pbF6j3mJzBXh8ZuOiMY2Q/LSVFvflstChLqcK
zJp6CGn9oHrahfy33h3VL4UiSxCaNr2rS3jw8U3jyh5IolKULpvNcjdZvtxkkIHDW5t44ge9U9+z
hmRnxpJsKya+ewogE/W1mvk9B7k/mLAxaELJIeXww2Oc8eCI7m8iZ42Jh8hHsIX14j7YKgUqVpuy
QawyQfi5OHZn79fo4I+boSkTKtoiafzATZFcKkWIBN1Bc02noJh6Kd0JL8OmjsHHrcUU613yQbT5
ZwOEOmlhQzwZQiaZnLWWYOiY8mWccfUGEZsSGg2XeCYAyVNoWh0ZyjmQuugY/ppUvC5GBsPKTu4h
bZhLQMz3ILNXnbbWZOYH/674Z2+6XZhzmrhQZDoFPSQ+hRqWPB0ctTvMHG95T0zA48pRZbyoERgW
1UrE6K9yn6H07PU0SfQUis3bHMIXI6fKW9wIP/NpzCQm1k1pLVv2XEUkAZSfpN/vK75MFo+PLHib
uh2rHeslxsZA1lq+u7tp4enHotqIw457STHpFZFY86hvNKNIRksDqiHfyWb2IZL9TZvoOPjwTEKK
lE4G3xH7ImTC5di1nm9GjO9yR4U1+klyFb9Lf0CsX6jlGnbBbSJbjUi3DhzoLwxBCQ1a07+Fkop7
L5w/xia7S5p+vrIntEegtauptErDFIb1CtovT5MMa3TcZh/YCgQr68S3DDv2BlJ5PCHgsKQCwPi7
6NK+EmzvyHfYKQEQxoyvWWe/VvKkI7B7xk6DAd1hONz6uExSLYrEsruud3MUkUveJmFnr6VlnPom
idPh9kNhmgmqjANMt6xLS+pPSxibxA+NIT68LKk6iwCNbNLFOsQwh4CoU65WBPzCLPhWnLAkVqXL
HLrscndd+O5PnzvfPm8fpaNbgd++zmqD8PuBcIOSuekwq18qlcYf3jwXU8GDAJ7YwczP7Vk0Ce32
kDGtqsWsG5FWrYcgHTTtCFeJJyd9ra7vMJjhP+brX891YbgxOhnzTZskQRxisvHqxBC/rDV0Brok
mJUCB+id93ph+criyyYQFw0PPY7VS3C5n5EJwTVYcFzPbsUEib0zf8YjCFSD6dUTQC8ZosBXF396
jHrWpAhgJiol6NMATmxSG0X88Lkw0PZZOne7JeF9aaV4GUt/botP4O9zjfohmqlAr28MVeDTvQy+
bbCQg42tI6/BRjlZwyzYrFZS78VKw/HXL8wU92mKjzwDr/A3TSlUSSZq3DJF2Ny9dYvCASyWCF/a
PF6+iqAbf6UTWcvwTM1TEgdgpGz6wZHCJYnNbLh/CJ3XHbrz4+Xxury0NPAMmXgiASLPo1cf51Sm
80GWftQ/hwnP/dTkrXxImbMMZct0Tg3aUM8EMCKIyUAiALx9J+mqEcFPF6Z7+tb5nSbaqrEJxnMM
WnPPMKKtNogk7Q1D3Vw60N4/X/+mldUKQYGNuJiKp4RMdo2YaWUhQzPYAw973ltam16/OD0f4+5t
nLc/f+80WEKWixfOyyXQooILnakiMjJ+mH3F7fIrs8+gy6khNAMAzY1+9SsWGtfuW31Ur3bDOgLn
e+cFuyeA/bb1ISgmIa8f7c3ruKfoz4EMmax91pru/pOsAIx45QV9RLjqnUzRNPvk4JD0iitW8BVu
lmW8vG8R5np3spsRX81PNYyo8sK+Sqb0yIpxL1SvtGAYR1fG0DX8ipYaDcI+JWCWft6F8Gojsx15
VtMKVT13TwwV/IfoHh8dyq2sPM5BxKEaB1KSuL8/wW8lQKzS0Bt6kKhgKJXS/o5xvqIQKEscRtvO
9yCMPbsCnRUV2xCGc2M8AZN7w3hq0Bbc7xwq931dtNaumxBgl9SqxkQVU+5p1Gc32hDLdgACca0g
puVv1OZqdYSh3TMWTUc8SSVGO00aCVlGrEFgPO73hZ9gkBFRysJ0iD0ejKdZxsRnUitIbooEO2b+
6hTaqdllSoOAbC3DENQN3QTdtCGpUd1yqh0WI9p3fdfcoyOxKI07cwxT3ZxVSgcpqxnnET3SL5B4
qS0R5K1nTuscbrrDK1rSZAo4ReB4qibiCGl6769KLpeSOnoKUovhpWSqLqlUrkc4fFzozdii+SYp
JpYPKdMitkUNqbCpn2SOzT6sq6AVxRZFvzLEAbrBq2JKJwgjEjDUJBE6wWP0Kk/QPMwnO91d31zB
zP8Ts13NzNqfzfzAIZiDtlWLKAtW/wKTOt6ibj7qW/WJ6aAIT/bETc/xgR8xaVpxrIlT1W40tL18
CyqLcl+4QNs/4T5GjLKn+HlYm2+Jvs0PHWvoWSa9xwsvEO3HUBjcYTSCEiEaLZDUqLLqdj72rlHq
OcRbVQex148rw9DjKYL6h5bkR8sBAc7n0pLfhPENoKcvH5trxX8jz9arnfgdqtbEy8yd2Cd2R7q2
z92AcMHN3rie+5pQ972JQE4gEAfIxNh2FNy211CPTrWoIYznFmu2vDZ7cfb84rMuXOBjbuZCnkbR
97JJMFuoUtnhHqvK7hTo505sEB6UsppjUz7rEBfCSd1xW71I1haBS6ygxVmcQrbVQ55GhVq6wB+Y
VF/S78p84q1Pa7f0HcKxrZZyrkQkZGliDdisqyz8DB6PoMhmm3kbSJITH3FWrRsSJN0WtpbaEDAG
tIvpGdxyQPFpDNiZbBDVDO5/3xt9eI7SD/FVMvihHGgMbMBmcS35ZdWylgk0qRanM2epSjgQ1jC7
O889dIlsogpjin0CIygv/AfYNn4tUx0pYv62lsT9p7QR4Utl2XHDko8dfXZLmn661RKTY7vWn0WM
k8T+J2TxNDMnReyrkKcmTKugdC+bqdq8MfY+SWVkBmA+m/zKj7VRc4Kk5qWK4a9ww9Kaq8KKGKNS
DI6K+D6g/68NAUfUihvX8FXtJ1goj1bjC2tvxx/5/hHwXhAf/7YMjpOT+Eq7kra+xO6YznGmMOFB
VqAj/dzOn7ffV8J991I/fXCkzmw5SyULwOBJeD7qJsBHtyq1ZObDAi53uRXL3pNAyLOwApS2CFag
V+OLwdIeWuflWQWF3GI1wlVC1ZT8ssU36rvf/8Da5C94+hM0UYmmAusAf6DGSr8+a0MXfpE+0UtH
BPcRlRcbxUWZRWe1Dj4bxOvzNbnqo8NOZhe9g7pRaoveKsTd+GUIsJKZMMfl4m9usk0teoPxmfn2
qSc2LZHZSzL9FJZPCHT24mW4xU1VBjBAWZWqpvYL3UXD96aOiq2H+BXhPpO8mc2WkLJNQ0RMuXJS
ekmNLBLJwftgsuMHV2GzIJG+AFO2OQc2CknQjXh+HAeXMZgOEt4rfZO5hcLPcCNHOVbnlDE2rsPB
+gMJztExexAww2ZPafi3FLQZHPzgUX7Ay0jyVxbu6z3bW2q5ZTtZdZwhO32UNqx6rhF7JddSvGyD
3mKy171tSQp736V4X/SjmIlM44c7ovDJvMots/icLZzNVvFtCf3a9rznguQW2YmP/ph6nMOBY4oI
e520vpyra8LJarpjPgM7gnqHwSbo0HSPRBVtO+X1kD3XuBJ1f7ahV9wwik8lPK7UwJcXPP/VYEGA
YO4P1o0m0eU6tLt+q2GKGMNb+Ax2JyXy9nXpluITxX5ZCcYs+U2XzZWrGROns3Uali75MUt5K7O2
y2JsxH9Pf5EYdUj3LeG1ucnraPpxFauwkY/KcXGMBQJ/cXL+JvS062/za664KQkTiyRJaMTmTiGg
wC7XXO/qu9TWcuMs/gzqwU8B9OD6741epYWPyjW2GG93uVip7V5jSvD7lrwLXS1Xfep1U42g1EAE
/qj0kQ2YggsZDAd1/gH0yG7NLf27eql/5Ejk4s2lrB+ko8KMHuVSoGw98QZlgb0WW9nxtyCuDZH5
ptS9wGDZY51JKn2ryY6pCxOlBhVdrHoHPFKN2DCBKsnzi/L69AiZsmal+toDOe8x4cBUvZQkTKrk
80jxEw5tDV/ubTY+Ljsl7FjVjSgXoUvk4jOwchQ3Q/Othj6n7vCj0ePXNsVupVLqRhu5x+xPXGPa
5beQnHqWbxsdoV2KFHovzUrjzfRHUAFMilIzyoJ3FYCEcDDJN7dpTs3ZFFYSsx7KnH6JVcQRn7UT
aTTFoRotEIQLDpG18+c4tpudtrWcaGh+7/S7jE5NXOQFhhxmL7eZrtUau6nyZYiMAuW2miJWC+G0
a8yinvWF+EMXhCnRySweyGnojCqv9czZNnU4vPcaggzc4qn8PGybEqIRwzW+R1dC3M0XoCPv+Hqs
T6H9ECoa0+UwhZqq6V+GzXkwZt7DM/PbV5Sv2fnWYsdCSVmqY5MttSyewP/uM+ml4KzCdyAS7BXU
wnX4fWvX/3BPJ6T4BJAsa02ZgUJVq7qz2DxiXbaM5BIDikehFzmiI3bw6AylC2/BuuF2YnD2JzD8
3/xw7bkqPb3tMtV66qrwhHvw4fRvtwUizfHDapBSNs39cfAUOBQcNRDZIpM9P5V1h3LfH/OSOB84
Wjo44GHGNUDKbCNL8OLWQO6jeRva2VIGtvVEA6uK2rQFLDNKWsJJ99RuiWC9qEun2PKJ+BmkZ1Te
98KeX1mK5vXpOmonF5arNja+UBZ3t7NIjWZs8py6fqt/dnA/Fo07Olu86olPlZOch3Qv8KXf8/6m
Rj3HB82mxHyU+OJv3ap1Cy1sMQrUESmK0kieTOYrLYr2Zo2IXfxemSwLYKvj9APFyuYYRXlPKI81
hPbxY8Zdzd92fU2EjJAMqfXyN+AoCHRyy25+nmahPMjZY29EeoIz2qDtZzGcszMdgZ1L1qbjbiLk
Sg/W0eFJ4XnaTYqs6Z9rLj2+HfKdgGgqDmkyv/wViqA4qBOHmudgnDmmsWUjjRXhGeFSgd1zzv/J
4gBu5aUGt/oxSqnUSPR04gjBUrNDUFBhvInP8BV3/mPdAMJaXOBLNlB6ik+J6/CUKSruMMsi2UgJ
Z2cFbnHqCCZsF+twd0KAAkfI5Frcb+/eIeiZ91qzSbgYrAFVLgVdI9d3EIAkww00GAT3QjqpGxWm
hND5IvPXWtwd+xErZMt8Cmp8ocmisFPJBpXJQ3TFPDmM7MI4UvR3Z55Gprfhcew5ijWGZva7ZGhO
Ya1SlCyrekkxqESufkDpfo89Uk2EJNvLOgSTH+O5MbUahW3ch5QL3a884E5leCRFl89cnHVQNAB2
/Cvyy/iCXgdNYaoYFQ/my+eWYj8zU2PnoM3D8RhHB5eXzsgEF2rsz1k8hUkPqOsz+ug116OqGZCh
bGgLfpq7lj0lCBl6yHmG3DKv4M7NAzNCqXRPa8JVjko3qZrN1YNqs63Aj8BhHZEz5itdQrswVUBd
5Igz8Vqg+SEvEgquP1sr8kyBQ+xHMZF7gVA016CZhi52ehjGTTAeD+OrLQhUgjTYKqO/ToY2cc5m
k9BF5vfZp/QM+luTuZejQmCLykwzSRft/2KjRu5J+zIV0CZGpCZmT0aL4at2P2J/RKOtVL2LkkSZ
4npZqus2UaPmJICGjkWDk0bi8wTuUhsmvnEWt0gF5zJjkpbcZDySbjaVzcBBZLhtvu8DllgH9jYz
W3aMAr21Z2Qzgt/QRBXeNXPO/24T+fXSTEaH4wKzroEJTWZtMb4WlTr7Nsw4mPrEDLgpixcT2Wzr
9OoWZDmiOZPJpZh2q25dyQuMPMhYANqMkueqneTJvgmfOLN+scsZ3ukUCrtyyuVvnbMpJ64oZhe3
iqfafvgRtFmYG/HxAl5POoGsAxeB1e9t11XfjSkgjb1DBi6K3Fmc1r2exlimE1OcwY92ICd4PnDM
QhcVqNT8SinsxNF3L1kA18J99ste4y3PqDQ+h2eQngFrH4PG4GSVFm6PiB3fUeIxqIC8CYrEGb4N
EX/JhVQjmJBO4KGkicZHEMiHpSkl3STISsk0u8lWSZqdc/pHL9y53Tf9JNoxkXLmP1p2Hxkc0Ra7
RccDSd+5O9o2jOE9Ye0dGrQSc9TW3HM/aZy7dS0Fu7Cfcp1HFq8H9TV3ZazyT1aEBRGUgUeN23wS
IHaV+4BdB8rwN8upxa9/ezKXiU0bDwrcTqU+Ay5O9kNfWOmTxoKsuRTu75z3bfxY7hKeC7wONf+c
aO+wuZWU6Mbt8dZmqJRzLzRkxhB658EP12RKraHEzDLJKepic3uY65dwwsRWz5yiGeHkKZ3F4t/A
+AwwEu9pMLqKt/D0VBEONf9WAvSj//MP7sk7P8/k2Ki6RocC60fiL4Gavy1EC3dHT33mK+bDI9UD
ATpweo24YJHpkb+wSIOZsBM+PR1f7u0NPSKER9qsPpynEsQhrBSmCWCoBUQUXhSgE12D0JD4kVRF
nU4ivaC6jrOYgq6x1oYmYFwcgQgwWpDfO4R2yIRtWbh7LxDTdSv/C+sm+csruYxV5VxeVZzYhjcu
4CmF194b4ortM4g7fB1Fk0bzuW7JGNB1La93DuVRoPKW83Z56ue+odTVHaqcdA6YnsCats8EzYc2
6zMKqhT35TxgAZ7tNWrgagQYz5JEBnKpT1OINu3MXwFwKuMu0sivL4xlPRap6fZLIkMaqlABLoi4
HuASQ/4I1shUBaC+D96iwfqo9+ORrOzPpgLSxj0e8ibQ5de8WJ537vkP480Dz2uunwM6lgaa+qrj
Bc2RYzEc64Q5Fz7vuD94+6wnvGosaKKpnwFctlPccNrj5wOZTV7nMvIAqw5LoplF7JoKOFX/IZy7
DqgaJOkwj4hcSHgG29GFhYRulz6eW4A3QqBf84dHtO3ksQ2Ml0oH/93mW4ki5eDndMR5Pip6hN77
gCqX4DANVeS7YF0qccc2RVdDU6grQJhVR9+nIdtS+phpiwrcSrgFskYLf/iHj71gcT42KdScX0Ht
JbeYBylYe/4d0n9WKJ4mQvLgPMXw0xQ5fEYEeuorIX/teTPiFGF9li+n58x4c7Hr7T1seEBeCLpV
t2nlyPXa2sN7b3rhXV1ysSwI66Qh+LOH/8LGdh2Uq/AvjDnLhWOawALVQDrYGiBw8p14PkRAuyND
OHVtyT1rhct92vm9WviAi7tE/tBrzic2XshzVY3rGUBZsSCSVqRq2CMz9aZ0va0JZdTV/rnuRHOm
QjRs766yxDGUWTmDfyjP1yo+6WD2AxTjw+FnSEQ1KpS3C6NPWBlSIw7b1s9SmxCLyeOhvWZkl9lH
0kqAfvDvDdHQgtjiBm1C6DQXssmw+sqqyjISNLpGLPFM2vQb2jTX+rU75QFq0zACsXfm4EkddJR6
SR6y4/fakBp0YsE9cLL4DJHl7rMg5HejxNTjgpqu1EndwymmVwc8uvpEICulTJMRgT1lOCsfDEAP
iNZAA/AWiDoheyoHP5SuVHGgYRkLH4ZEhzhhU5YgCeeyxabSfKaoBUqn61CalTfkOzBs+bXjaNXb
BNExvgChVUd/lhztvfbWodjVU5crtua0EYPU7tYTWApJlsBDNVxfUA3eYMEEf15tfl99XFnIQZV6
C1CnNqEuq61eJUisKEeQXbeODUw7tvLw31y2iy6DfhY1WWU3rBwJYQtzbKRyS/3pfR+EZXFXH9np
3lBLKCYKdSbnZs/zjO0qCxgSxeTo6UCHowmHgoJ3NYKq3ss08hpqN1zWr4Ij/zLA3ZjEbJylbNB0
T9UQuRWZY5QnakmvBh5RO59YUGWyEeB7pZD45n7Fnt1jyP2b30Si1X3jGuhC40PkRgdgd8tnnb3Q
vFscqxCwUfLEk1CXFMrts2DdLqiwt6hOuuNm0ZvihO5kQIvJjmcmc7eT30gtpr4+kgx2qC2YJorH
FoFCM86BjobRSn+1eZoMOPvhjhUrep5uT5w5+uzJpFEkwyxwb9sMhHQAWHUVW3mvqUzKPiLbZx/u
g+oyhuSfZAGTYqr2lKD/aOXJ8gTfHgayY7KQfCA4zevPxWRYk3hc8mgBfihH+AyaRgeB56UDyxhJ
Fak9zUnMvzU2+09vsjjibnPwnI+/dM6rpWikzGhWBvdQlf4g6mAqSm2pTHbBXdBT6b7IQP2wiq7i
Ki7hFY8V/DL0VNwA0oXjJBOkqImjQdJBFINAgdP1wfpxY2Rp1zgL9t4uph8AzFB90+qzqLsolkma
d8JXIgJ31lCOewlTGydoLlzD/1rd8r5cZvQ8Eqm8UtFk6ltcGKBo8qiJnVY63+tGS60gnmn+pWx7
97k6S3qTrn6SVoRG1EM7uXRQLpM5y2DT9Lyuuz5xgfXxilVhuWaH5g2TPMVpg3rkHgCIvmxsN7xc
rX2s304H+IMacBmlrHaXlo+K9T3eDhNqosjb4CasXbpkPvBhSnQmJD0C+7UYisDmIEFckDc2tCWf
TZUnfvR728I2mWTAWZwAQ7UGXgGXBpsSdUIxC2M6nlsMR/by+LlNvlR8wajONV+WIQ848o41eZg/
SCqz5N5Yj3yjBfMExAkFU0wNn9hiEzt876PwI4cIE8hwbOmvZgqVxcwzu507TCmNbW2e7JqsCDE9
nRHTsOlo7a/JA9u4PpkBgLaLLY0LFd2/ZUKays9dGifXUZnUXiadwKq+HQxnfj6Q3u3jMqvYF8mb
mtBkT9iwklG4cti0eZbEDx9spgDiPi1Yw5RO9yFOSqLEh9XN+vsVd/V0gzfc7CLvgiKCaQOl4ZCw
u5titTEuVo07jNImMwXfZxR5PWAtEwbVzuUYUjtEnNI3eDkldR+Xog0sgfuyi5KrrIaZ33vALR2M
3L+Q2NYK+7jE3VZbfeX6PGQ5SO8HAUfZ/6rbENWMIpdOo3OeDe8vad3/dM22HXKRthMLi1qQfVsQ
j/bgJreoqfLpXdiYq+6DyO7gROimbX6fyLJEHPv5mQwpM759Wg4hhI42WQSO6eQjt8TvmGEkHTw2
YLoI/K6gLvkFIxr7KOgA4f2HwGtIv2KJ52yIsKQEyK2R1F8B2trVkqAIEG056vNvPIIPXWJ6koxM
qwOoD7Dkuk5G7PQ+5tjzAOyysYv41XRhejJpx19oe2TOJuneWYANDT7l6qt6Pli5ivlPM094ZK1s
W3SCWEXdclwEdcXI+X2HSjLoC5dExG4fXXJzEodN3TaUSYCO++Vx2qOCG0KOOmevBdSe90r6ftXA
5fqK2zJ13fdE5f/l9oTFJkTJ/JQbD27F3cBxERYzbLlFebK9q1zjc8CrPZvGUWaf0k3H9OSjg/xC
+CHLIjb3cUK3UrzYHjQjOUVxzCTbHKn+4T3XpFZAh5ZssG+jydZEh25gn/OqpDCtTk6OnC7tnICe
LoGFfP00BFceb+bpilvHn91epwgneTPibGPi4CK1hiineGhbW58REWoFrxqMM5NygfYdP9MBnJ1U
eRVIzMRp7rsfsJ7ggZjVU0xCf79QVca/O7sJ8ehuMYXnSnJ1wkyppZ+7hNMi76+RP9vPZwZOMBQg
E0YkV9ebzlO15iyu7K6sEambHjYwm/I+C2HqcdjaxIL7EMRxh00CwQZVa2C9bW4dOe5CJWLgWKKI
ARoq58F1y9yN6D+hAc0zrLf0lkprnpi/my1kVpaJPhIFiVjLovTbfFav2Lg8PhJP04PLAzuUgczj
nMXfvM7m5gO1tdUcC512JT3lpZEPEChqmxWh8/QRZzgpnnztaIlLXbj3jRfa62HphaicxnYVGJfO
F2CT7oqY2Va4Ymw+LrXRAnrDK2Uh7ThN/sPzY6A43nJDL50sxvna9mz9z/iIghXCnb5kAqgN6hOB
UIGpsAz4M7QCq8gRReNldQuC4RfsnTSKG2HdNiHKSmsN0ty8HPxyzv5SHOgFCcdMFoqWECNrRyCR
odSw6J0bcI9fUw2fa7oNI/5EyccUpY/R9pPlvOIksmtyC9mKW2y0ddIcgMPFvBM2ro6aR/lZYmPd
QPUK0yDcfbTdj2MRTcNU/iHh+PQ84HsZIGVIBr8mlBlS+DggIYPXNGLl5hLnSez6XMsBFITn3oH3
CVGegdGUpbJDxgI9Yx5TuU13lpjJW8S2CqYMKyQJKowz4WxDHBKBACY6h8UsV1y/I/QE3niWEVfR
jnLFNIpJx3ZeFwcuBGYyo06FdvhE0+w+3PoBMacBjOJ5WEo3gY8scRvRXT/T31LwAF4Dzo34HnKL
06UaEsCxMsDZXo/ic4mYVTJaQFMkxt2rMu6JxFjuLe+PgzV1y8yTXcC9m/Y4qqizixDzkYetTqy6
MXAjb1rPdamoykt5GDhpaTfgIbmQQKFME7KxIbhCk3dWD6mEwi12BJ+sL4bfG1nr/BgUusckmL2E
+v2N1mQHVddBkI+D8C3kUiRS0buu/uyb5oG5E4Rrf0H551QAR2YOZwsdBGzd8yAUshkQWva98nDc
WX7oyWEAnt3tnHhO/zVpyMeHA0YzKMBLm9207DQ59ShKiW14GZiqwn5xQix2cdBSFJddWKAZLVRT
unRrPgpyfpORTzsZHkJ3z5ORq/q2AZEe3dhAzcCNT4UzTCvatdsGCwTMy90twDRM2FNq9av+sPJ7
XEBvvmp42DAYmK4+N9NUno7LmclFmPC+txEuBjRI3ufXOcBkSaLTsVl4jm+y1Y+PL6ByKsAaT9FR
XjL7chIGDlDslT2kCFxIqNrC+wXHZQzxOqLJchr6orfkBdfhFh6FizPEoo/V3pMYDB4FKaRUMIUi
REHvzMIfJnzoFv5wquY/8AFqQOJ5lRnyC0oSxz569FYyQPnCcpMnbL0wpuP6k7x8m63Fsy3ozV7h
/9fJu4+duYsIkwYSDKJ8tcPrfocyVCfBj3V+k++DZbtDf7RWAqA8AUidIWzabtie5XGCDyB7k4y1
eH6p+OFzNOD1dy3wT5QPOnHHM+HZmln+1J9O3JQaHv6ekjmWdD4OdyCM05ePeXN0XLF1msDzRw3U
DT5Y+72zUBphYiq4uBorRryfibj8kZEedJeNU1zmL2xWZBcuSlO2C3pWK+C5obyl0HuZ9AxFfyVw
4rgPcf2EkGQ4UVPQQr26h0QBM8R1Gg7XCHXboERyYessAoBMAeq8COTk7VoCZNiKJcrkewSJak/l
akJCkvL+2CVHL6hzTHrmnVNaQvlziZqJ7YtZ2nwGXw8eqo9fYB0gvfQS+OiPBy5yrQhINvBLkjzc
oPUUXNmoUjMlxZXKD7xY210JYuaBZmWpE369RGWJYfDXR/gXfWcxmakZ3ol6ZK2t3CE/GQ21NfWa
0ASMk+j1pooO2acMBECgxA1wJbOacuchwXg/3vd5haDX89xoPhat99U39zTt2WRu0OXu7ZIyYOq5
RUjbgAx49hxhrwFVkFBYE5w6vLEdxPyhLmVdKeE7XIoOhmoDPiQkVu/1EgQzOHawcwD+I83vHHEZ
2pnCtUVfTa5elJfPIS/m2/YRHortSdeG96L/t5Nd6JiTRm2VGjRruNZyuVFXZ0f0yu2pvkdOXZH0
nvejY3YAqzYNR1uf/2Br8+cYZ4IY3VxEYVClbWRiyBpspKScGOm2fJONaxr4FMglHGezPGiVibJt
YB125DnnW2VVibtfVc6itvHEAaHvpWjaAfilQJz4rEw8JDSBrQjxvzyGGjMZz7nWFQVCZQg3YF1v
aMk1DglGyrypIWi9C2GrntyC9d27nQEvZK2cCZI/7C8t1wZ05HSBMgFBEy+cIsPH+gXZ60zEFlkK
CS3QjV52InSa7UjwgVYWp4C2z6V+3+Vi6jpuyoZ4/r1T8OPfA27RuWdCyxHHowyaCWUiBr6C+HPl
m9nbylyLd6nwGRDfEmldAgOKi6ymum+wgmaM+p19RClMIG7YUIn6EWX5NzSmU90GcSLBF52fhno0
JmK2lUzDbtqfb08g+tHljPeKRh3e06oM1QpqY7zhxcSwBN3qCQMxPg8yFACbjJM2wcTzZ4JUE8fD
BCUNjXOQLTfB/ryCy1OH9oS6zdcuKfoP3IOIrXbdAvpCXArZIc+HYncsgG7VGTTT8UMDqh+yRn+O
1MW1CC7d3DJF2hWPRCI2Wf90HHGq7hV7gG5NXhvum/rIbSVK4qyGtXNVvDoAlEWmN3LOTRafAPf1
XPcbZaKcx9oQpH0vvAFvY7mcVZClD152XJY0gd8AC3kO4vNXzdtx3mQZ3C+9ZudM/eha/NQcg8SO
eOIkcWk0v8Xg2qO3rNFHZVGV+XcaSv1p0GfMkj/o7epjzzGSscY//1D7pDP2hmFil1dT1x8d8gBf
khHVMCxfjSgMzy+5/ohSzRvGzEFMkeUmDoQCJSzQ+SXhLutjukm2+gkJH5mulJuRwPDLGoXWqFNi
vdt3uDkgGIMlNeVWf/HiYnlHq5rpArW0lFlrtpJtDDjkXrnAzUxpainDqg1TcnHtOQvzmX+Wrx/F
DzpIeZRxrpeGNniNjfsnwSoAFPS8+a7mcv0bfZUm2B/rw2O+o1+Rvdrzo05I2BQeiHHnOfh9lihS
npmt89cL5OWovt7tk/7OD4/lQr0ajJTrzVMx6Ckjk3OcoLIM/kJwXLCDAgpRP5yCMx/7C/Ja2aYJ
N0ErzZgAnD06oEPgr/h+3mk+XoDnBhbsHZembhwBpxE/TI8eUm26SbCDr4UVC0Z9Cq/fKQOHYta7
CD1x3a0AlEdHGbSz/Uinf607EorZ6uooAYBVwU4P7oD6WcdgBPln5EIBS3+TMH/lb/THo3raD801
ODSrptqmNriUlO4CtxNXhHfcnxcmKr+KeSI4Nwp5d9Ta53PlV8JbZwfy6jd0RjhwL5kbleBeIg6q
2eDW83Zg/Gu+D/8dh1CMlCH5G9twjFF4t5/2n1WQc3Gcaa2j2tj+WQQLTjPd3s7SCnhPS14yvcIr
SC2hbd3DS9SRH2tdi5C9/RaZ/ae4tiY89FbKOpIRqEgXggBJ64G15AYuAVQpiHmK+9o7EMtZOzDJ
0F8jDNJya0kghcHp0tuhIBHBgoObGfl7xrj6PVRy0CS19V3l8mZLL/F+i0kZD+9X0KXPgwi5zxUU
bDeu5AcsuC0y5IoyoqPbrxpAYz4jxLTuygodsw3TR6BKe3emMhu2cspbKhV9BfQTR5LABwHro5yt
8fygbnPPOZoZQJDfR8oklUVfUAcWQc/M6LUB6bN+gmqJ1VUDVfQQ6Nxl1jyVrAUmpbohtYYcxJJk
Fj+XpaRgJr1Amzu0pe/l4hYIU2UOde8GmtuvHIxU8hANzM6Xos0lydVwtThGts2MOQu9rh9rtCaI
PvvcYA8VGqjD+MtJBTXerJrdlUOFMyLDF+C6KIRKfbyZeTe/JJ9MJf1C5dNGQQR7DLHhdougcltp
qjYVK3SfOAOoOj9dIMgVXztqxvEdl8MNuJQwKiQFWAuuQDWOhci6Z5Do+ll1fuKsaS29QprD11yC
KsXC5wt+PAqsusFj3OiSoPEZWltWQjd0JEpMbpLzZb3zPkCRYWJ28wgxolxnb6U9RPhDR5MonLuv
gfGaWgSrk9T/RmL/N421kiM2C1tjDXk9QTlUv2CByltBYPvmBgUUDHp5AZJShxiNHhJq7NwrYBhq
l0tAG52czxEKsz1CRz086l2nq+0Dwm6CT61n8o8NJx8Gopr8MKByLx7+NCu0ExHuT6JWu0Fol8OG
BfVM9agT17TBnMNBiU91zPCrceyFsbX/YZ684nbEKFdDwwLREnyEVCAYWVch/+xvMsHkCjW9KHcI
x72bTjtyyrFEtCGitqlnboQHFSTRbcxxhhvc8yUmRbiivxJoGDR7MsjGEGM/LXgthlCcXdqZzuAJ
teU6OjrIcVbE4dJwR95X9lE4Mnd9Z08yodBIDmCNhe4OQGWdL8BWB0Iuqp10onQfnLZXcF3+cKg3
jC6ifuZC1mEQVmoAaYNWbZGFovAW/IYLmGWz7M4n+ULNS6HIw6mqflzCHtqOBSDkg9Zy7A9hjtaX
bOMWvLPW+580EHTY+xTWgh/TZlJS3Ma7Z0/FP3p19buxxcE0UNUVZ7845uRNFkKk31eB7UzPk/dQ
vJ9fTAGuQae/2dkQ/CmBlQI+rcHPC597CyKSwOPjDhUnh2GAoNrIGO/o2qDBtNWA1b+wBPmsqHQb
02DIjGe1CcuFG9E2qzbW/uKT1UEUZDWSgyN7G6wCBDEYMhMC3HY1RgD7/lU4IhJlol91wA3TYu83
sxOB+yT2kDICtmtbFmgKeIRam0+CHRJYJ19FDByavGKDc5Oq8kgI3u/sb/gAjGdh1gSecguh2uJO
b9DhULhmQy8zhnTrKpxKJXcEbhejcbCqZWNuhyBOidix4IShE6DuA68G+YFNmmEXsINE+S+fw2GY
PMQmmilwTlsiJkbT3x9v8U0MNp7V5F20A66rkw7lMDzuYuyVLowT3UUH/dAlQ5NYJK663cvrqnfe
b6QS4nc08rJCrEZyc4tWfcij/3jhltjZws9dLziBgfdRj20vHRH20ncc58y79fbjHP+Am2CvzR/i
CBKwktIPJeKt9KBFI8TREkXpMTLiPEO4R5m6HMgws2/UHRn6CiLRisORn1+iZk2eATYYdTufZBkf
XXdMyuFlfHujrZnBAK09tIUL5SnlBwdQEsViNhR78jqw19Y5l/gxPHAdMgz7V75X5QuiiIDNOUXy
UmHNQYMBWTfTIyqvECZYIzdWvmBriC6LPooW64fWY2JA90Qyp+UU5CAeAm0j5wmT8pmv0uVP8ydY
gTEihgJmQ8DTck+tKFeEHgFzLNEyMDUXMZz7pwIKaml2q+BJRrMAJPI/+1JvSjVEUhMV8Vw9zuLc
qapqot13PbTEBVWrqJPCTP/pIegXaZlGbjcAEAmCI1NcO0gZrmVshfdcajHB4qbWiNCYmUnNZXrU
WsZo5ynMkKTJONyCXI7B5O0yiOvKpbtVxtE+J/Nmhy8iiLorXObf+FV0YJqMIIyAuYqQtcmOFAte
WpBZur4Q9YOhkhlvpo9yzjSu4jXLg4WZsrbMzEViM8HTlmBB3QSH2hL/LF3dknbgf2Rt7cT+K+Bv
jIgriSAb9CeE0HNF4zbsey2HNb7N3DBrBm2HTlJM0X9CRtJWBQGOMUBqJ55mKW7CkZqVv+E/0LbN
FHlRRGtnKWGHsa2sDpAb0ZF4wixNwV29itUCBDISYdZOiSy17tRBJ162Gg5OJ+jPwM2F72KfeLVl
IQlt9DpXeiJcw53IQ14y8Qs/5kCK1egta+OllcnGR9jlte05o7VMFGLccTMhpn4nE05Cy+LyJT1c
udL4rE97urGoXNECXUbhs9Fvlbarg+RgnHiuXMVnfR4EvIB1CQ7z10EicwQi/VIT0EIx21Q/lUyO
TTKvPqjd8LBJQMEf76C10ic738lyKNWClKvqAABfalRVlekULkA3P41pSsZXM3CvNzUyboQE0iEX
6qliPJEE7Hmre9Ym/xXT4E3kdC0x+IW/K9nyACWWRIiIFK63vVykqlnW+oRxryR2lHZoq63aK9Hh
5a0fNn8XZL95QUeMQ1r5YudEbjabdXL4hxHK/DcqwfOFZbgES5ZYQu8NH8DzeJozesdNaP9SeWbe
50xsH+LAiRn1q3aSuxC3Br/Kam54Q3uSNlMZOZcs09y+yNEnK/1rvkwtk6pJfAfsAB9sAsUa8pBF
qIB3/4zzrHUGyCGenaHrLfyC1vG/0cj4YFQly7tEo1LNRxGKlVZKHkwzfTToPESNkhGEbGNZ5xfj
g1wjSjhjlbo/nHVj9Ir01ydvtzWuUvsiZgnFKmoTdB0bhRlJrCAPUoPzFBont2Wn1DTk6ARtVPKa
ItuCIqXZB0aFeY5Hu/mtZm+ZTV9U+OphlLIotorkrFkaonqxVnGNBaMePEmJLqc6Jg9s7ZvcPDlt
TiJws6B+zVg/fmZsONxKz65SBF/IE5dIYBIVAtAeSrFjK7Cc98MHLwtIQ9/Px7eZH3j8Gc6TL0mp
TWuGPgDRgNRT/s70IhGdJ0bfRfF04mqyKbX8rcuC8jqs2EkJ3ynTq3zFgi9+STXHDq4/CxBWvjHA
22PDHdQpd5aHVzHrjio8ip8KPP6grFeclXFV4BhFInNDzhES4qwcwME2PhxQFurseGBo7p9c7KBr
5U/sGB3bG0vqyETUJJPrjjeLNfGjEm87ECkGhgFsm0dZkOKDpa7mM8buSHEnA2bBDsNpCjBUnUGi
VC5c415SAG72//WGcOThnuTc6utskHIHo0wi512cya6oA4HsOUAB4O1bJwwvergcRiu/zBPHhvAS
/vmj0djKS8w6FEzUATpB+fXfvtvp14SaUtzwkAQ6REMetQlYlRcNi3um6FuEcI2EXwwjvxK8qLz3
LS+HHK30QwdEs/NNzkkYPYuElHrNQ2WPPdKImR7YhkLi90G2jOvlDj0WPhoA+Y9nv+g24fq8/XEq
6Yn4FKgmTjKj0D9if7IC3E+bR/IxSdFL6Udut51umq1qVrJnzmdw5HOFrCp3h7GTS/w9AOBicbMB
YCE8qsPRycaMXm+p95H26K0gnxeucvmjQZiSo0UDKuTZ1ujcMM6Eap8msweYutP2D65gejlxnY0i
WVOINVmzPorgTqHyMVN7v/rf94TkP8omxhS6Wu4Cl6CE4tqvoZclJQcKpFmnqtPl7NRe+l+tLP0j
vSH3Si5CTsKosjY7Y/e9pHeoa7g4yZlyh3wgSW3FCbWJNr1RqKB1yLOdmUCgjAL3LQROnNq6hBwh
s1e4NSXqJ0E86aWQicgm5/eSc+v33VU49bBu0Gjvpq8jKdJI9ss9B61I8PacUpiXdCXWuj+U/AMc
t/HVHUh8LolKRZhusCbUBwnarDmcV4SM6mLYVoiwXMI+35luVTq6v27q6/G61u2EBflJL2xAjN/0
+MYtceLdZyndyrPxWu+THGMuQzQx7G0E4Y2oxDgfFF5sQNUBmwdCgCTvLLJobsbW4+O1VsuyE4+L
Qk1EzZBBtOHwfebN2F1GAfnQNkGA0Uuuz9zoadlZs3/+cbDxvKjQqyfndMehzSDan7yiMoNQByGO
as3FXtNNmhM/ORJxw2nnrsvdcpeqTV1uWXbWdHMJ2YfYOuiQY4Jpuvl+04+Avs4DuQKDrCysur9a
ozRh7t7RvuoYeKcpHNo/skjVNxULrIDHYlbGjU/CIp08j6zXfbTg9JuqawarAiSIVNTsqDNZUvM5
jUF8kFWnm5CfF9N3cDP1ogtJWps+MSCc8D6SuF2zDIseFjGW2ybneZ6hApJYvfkdE9uBtKlQOxex
vRXIAweHN7rFwQWI0wonxssDQjkGIPzu5z5xarDjgjbLkRFvaA8+0PyhAJPd9gQpbZQoshnb7fHc
oQkdlCFF294XPgyI0uBdx8aLAuytFWTYSwm4MGfQXQE8rj869xK0Doeyou0oZZUU6Am9/apQPdDd
S5Yr+8BdvMESa1OdtRTJkewUJ/lGwdebqdooSz5ubfPZbF4r+FoXbW3BINs3z824iXfyn8f7xOQJ
lQbQbjFsMhD+NegmRK+6XhGywYLalAS6hdN7GFlzNRkKORj9B+ZG6dkDw5nKaAkwu565WoyFjEku
QLuaQ5IvvjHvm0T+1VVygVZ1oErmmZ03z5n5SBN+pW7ouL4tBOaEs9f/w1p+j4tn+epFNGNcRCwc
CTIj1Xsyy8RUwqUkuuPnRu+F8mWeKx5b2wBvB8lL11MTldlSPsHqOsdZJt2XoPk6ClAcTIYM0/9d
owNDt2k1S5haNZv21v5yLyZGay48m85d/8vIziXnSjkl4XVPqoz66SdRxJThP+moW6Rl0q3LnLIT
qz2GXp//D1eR/PF26H0ANklzyRTT+uEbXComE+3hw94F1OCTdfZ+XrAPdykucQIUPLl5hDXvnFm9
DUIdmpkq9oDuAncWAFMOx2hpaO8Hp4TXOxs+xRP+ohbX5n1jmpm0rnuSXu9A7g06ng2wy4NCYxbZ
N5vFnSuTqJBGVtEYOHk8z6NNVI2xlwNcJWROia/SYQvbDIERr7hO1D3OeQ294ao5L2ry1Nu7T5pJ
YNbaik10q/6JZmCCW2+/SMQpKOpaptobz/tvQV/Zob30IBgmKv6th1Anb95ElyWkV01fe5WwiOP6
7/B3Ry/fx1alidFiV/o1KTNBAcHHkauoGnGHn5AfoBZWqs15Lg/3VKaxqqR9lX9iZRU4ysAEj5cX
/vUM6yFHydDK50Kb9cLnoqHxq7ntjeDFQt/jj515ZZjcykW1PdrPdCTlVZXjNzy71AqsilMIYUUL
uQQg/jL+5VXk0Iy0TG6EKpvhsFpOFXxvmnaiWU16GkEmnEav2B44tWBRnXIXXOa+CaHCGDpKakS0
ZEuu54U25dSyQJFkCTdr6i+Eh/tKD07einaKNpBeF8VgTdPq3I8i1kqDX5uPGRFB9RZ0Ysn/uYon
h4c4Zfn9h5JPuKPDSaLNS62LEs7FWTMXZFWA8rbTKAbCzOItz8ELp5MliTPo/n7maplinXf+ig+R
BqSjDCC9U8kgHwzdRIVXfWsF1iKtqXOzKJmw6N2plj1//qK9TWElqhE6hTWgYjXU23I0fwnS7j60
RHT7qtlH0NO/FikJ83tHfGEEvTMSb/OuHCDKlg/w7Ee7dm54JLLyOkQfDx9Jsa0GNX/0a0RbjDns
pcHXGU0Ym74LMHBQkYecoOtPILgSau3FvSVyx6kohhY3B9tqIKU3EuSGUabYF7zqvv6i9pPMRkh9
8zG2NQJubURkE9H1c0+NdP3YHJri6SeMWXsQ7j3oH3xRLIXdYD8ClzGhcZ1fzyFKMTU0J44q+uU0
NjoQr6JBG0kr+vPmEvT/mqFTP4RCiwchtib8gBWTjjSDjqIh9WFxAqAcb6BAlMJioPXDPkPQtb/g
08/k3ewb/RmYczrG5mlFic3SGVSqcA8QLwsLy1cTp3sEBWKKiuWrhh6ebCazweA2Oo/2i9rniwRM
ytp0oDSgM5kGXmomgzMYuHO/MetSHqeDu+ALQx0JTtR/LPL9x9Zl2RTsT3fovFSMoTnjI7jVb2wy
XsQOCIp8lQULhNbaaupAEbxPEmCTzilZVpxannflceJBheMXkwvH5HyR75uy0KHjYfIyVpDMNDF/
MWxR3+iTRSby6Bo6Vwmv1UqD/JB1orQdqnuMiR0ySKqMOJTmpAUEZZL4Uk4YxUrXs/LJ7thon8vb
Or+rk3IGrajTwNjaHkAW+iMlIXQPGcKRf0hQZ8hFvHBZuSnM8HBR/qDRgHRmlRqbSAUD6ZeJxI5f
IB8+JS/jLswwmO8C9Rrd+1jAp9hHJmc8AbSEecSdbIKY++n9reUDK1mZkh3zXLTiTk3L7TuTpRjU
ukIek2FWri6kktP7qRUjs3gf42A7pJv+eTV06Xdp41CY1Njp8OZv034BVsSJ3ev7vxDM+FC86Vhv
g8xNYoB8BHkqj+jmtomox6OIrv94ufFTNsDZ43kV06nsi7PFLymTbqJIyADjLnAsbbB5ydo1xBcm
/5nE2IJwOqTN6/0S7qD20ALSsKRY2zhOX0x89SjQ0v/uTQDIRUgRfECRjcmEVo4xVETUKizAMgSH
Gnh2qtlG/aabkgiKGUeJ/DVEPA9P0zApdu11bRAxCY+a1BxNPq2tYOBSWukQ7zLtgFeyEu+qNEl1
gojsICamwXmZc1zfmD7fgF4BeP5J4Gqn0K60gm7xghYr8rZ/dNMbsx6WNEGnRTj1Yu95MtVN9Zm1
oHOD2QMt40ThNJ+vSMD4Ryz0UAp5wLVoi1Po9VkMDN3hST2tnv0PxYUAfG6XL59pFdwJz1WUqs2o
2pnEL813k1cZQ09ryxGdHejmNBxseKzUQw2ZgepVrZ55fq6El/DJnO/zU+On1Pug3GTB2XKroF5y
62OG1nEHJRMHT4ZLF4bA2feJ4yVaN8mD1BkN5kZNAjVjyVzk1bFWideGl+3Vu5MhbmZxInJoRgM3
ZOLZf770HfAwxP0C2y8104CkPf2Wioaz23pJzii/qpu3zz7DKajFsEdaEO+TQ0VnDyyz2IUWzp/s
MKpGtAXj0pzrWZCDiuym8N2yBNY0/o65pp1/HnA7bIVnu9Tg8yRQkdwdEuK4Sd5MKkHZAV1zCf5o
2r4ixavcPLk6rvT1BabKmFwsXbCYEWfCYluetSH6zIMnEU/QM/In0YXmJtPEBO2L8cTsq1MFWNLQ
0+42GpBbhoig6Ef/lFZJLKdyDUvAvXr7Xum8OdlibD9eFgXpm8FliEOUm95U6WwtcvvmqiubZL/R
mAQdg0lNtRBMpxN5FFtIoc+2sAq2YKA6YW1RUmon9GtI5xur+YhKhY1j/nRLfEhqb5IbWh8pu3se
npt0jdQOBFQC+JvJjkLgvMDPbKqOQTLN68OPYiDGkPYExWmWRq/xCE1fRidMXZKDNbL+up4cFM+L
tiiZIVwohOg98WywyJ2iXHtstHlGVvTG7L3rekdeg5KRBkD4fTMyV1nLpy+3Hdy+xN0J8ziwymNv
qLJVmlVh8w6cSOCiY68xrwKuq/FqxnT7R0wiDxG3UnlnVckUOhZE2WwSmakdkEABUZXgdosNqaSk
U+fcFefwBJL0/1NMBCaibQ5RsnAZuEPPqdUOEPqp8x3BeCAPD9jFRhEgBowwEmoWY86hDJO4xk9T
3Zo57yiJi5HeXozsMc8UfKjs9lXY48csqTBUWQGR47kBjWP5A2ThXcQFWypuepYUy+5vt4ZomiqF
ksMMtENgvxPFke26nqPQX34ZuX79YfKXwgdzfwJgVVJkd+EHGEQtB/qHOfJ/U9A1r3Uu5NsTm8Jw
g5DvLd2Km0cTRTBCuHnGXqggJ7Sc9cfSmklrT/gV9Y3BNVCOCQFUkLYW0EkiPGHB2gjrpmkQ2d5L
OZxhEPpOLARlnjh8KdrdR7SsghLp26xKl5Qozmokg/5+D3UTOkCivg+T+lrL2hBg2UAesKNeopHn
MaT48z8VhOrnBi0E5kL3E9iPqzBi6kLV7zk3CKFNLBApd/ZzEduHZSOvgp2GDecAucwUzQ4t7/Mw
ZG1tK+eMfmu66quNPnCjNooDxU2+6d34Kr5OuCRFuwUWAbYTA2ebCqNNyT3o2CpSURgmKvBx+DHu
Cbf4SCVGiQymTFoP5C4hyP8XwRphl1Ij/IPJfT/XjThJbjLRHbstHmRALtgup6O0wpVX/zjGXvjw
LF36lBNMS16RyRIGDBTAiRpdmlhb96fq5P7ZPNsCozTxwwY4hUNQ550Lb+s8I4DEC3uwTacPEXtu
+BqJbm/F3388a2A/IGDmtg3lBHGT/850+MHtIfuDScJhPJDKthQDSVzDcUlFy+iS7FYrkidFxd+W
1cVgfK5qbALKw/skyc/h/ysNM9q/B0UyJnMu9X9jP4Xvy1pyOkOasBOXaDK1cFj57Asr5xj+MbYU
qSOdA4ko6wEzVbouNvNGJfm8834Yi7n4Amcz7OpZ4lADoI+AzMXZgtnminIOKl5CEwbbV7YsLEs0
KfauA0odKrYPA12F3DE+XweLg4pS4YiAeJWJs1Lyu16nzfb2v57OITbnDLAO1DussQhnThStX7Xh
p1ytpQo4kXE7ZgWeM/u+6VDS6DR4xSYeCMMR8TRptVUXxhEmWKpe/Iqs9jsDdXaE7mg+8+z4F2lN
hEHxag6YPt5UNC4h7bhLsJ6OPnT+lJ9Jn2ZH39wSgvVbbmmJopv0WSZ5l2dGDk8FCP/gEeV7LyWI
EvdCJdPI0b7keP0nnld8Q3Cy9vM3YCvsrIF9w8icbnsWHzURD76lC/6r2KQ8OlyVnt8ieBE/JtEz
Qmwd1c/B7nXKZynfhM+SpmU5UyJM+Y2PbTDYabvU0Lz41PYPja1QS7rf2pfJInwf/r6ZcaqsDxYP
UU/No/z7QwELt+68KMOOfqtpfNz8vmV6yw2GdkCfxlo9+jdCAZwmITDFLRCdSjYz+iT0LDiyEUYy
L1PUQKWfJTjmqyRhTffOSqlHKLcpPYYvmO3nnvkfJ6WjfaZQ+MURtKvfXlK2V8+3L4+3EMFOvB25
sY5+PPKD6i7Eusoe5gg0VAUo/wcnnlt3NVH9P/9CLoSnXBUB2RMP9FEuY+yYmtE0rp7aB5qTJy4j
ZieAVik0FJKZGLCqbQGb1LNs/N4dbhqA78AOfGXT5yrv7JuLooyN/XBiqUyeuEYH99AI9gbti8LE
l2IIhGBMuB4q/wDyRWvUZVjM88IdmzP5sI6rQKWh7i9Hlu3kVc+zSbBNvUl1JkCM6EahgfyACJsy
wCmtn2BNejAV4oEqPcFPy9zUxWpu/jHwRf0lOIOBNwB8LbEy3cz3IFczoo5LC1gHtkdm4jk3376O
XGQLxt5ByRsQlK850lRwaInbwLQHUzopaQ77Ji21qMpSOHN6El80kFjF+ZMjq/wWgEEPbCuUN3Ut
iLErH+VztfEI6xOo62fRrk2kbqOF/2+O1hY0sFDp0K5pn3ItGSeTIfw0Hg7o4xGSCuQWfsP86u/Z
t8hIZkJ+dOKw95xirlHAvnpmunRxpF/3CeyjsBaTFfeP+xb7HCkkK/0zJPuBrRk1bD3TT9JfXT0s
bb7Ao2QvIEV7vgIJ1y6eqXurRdPEW7lZTEl6X5jwDIDe0ET5djdAZEsS7JoxNOTw7y+L3e3r7PJM
bv0b+XC+X+y4GcgLRATSbuVCmGjTMQtZNtQL7hRkXvsUSxebQQEGGeFIAMOw6LND8TU0VeLBxnPn
zrDh7SlOXouLOG0YJkFAVwGniK2hxSAEDB4d9Xpv+83kkO+PBWchOrrubYNzevmONAMr8alq/udx
bRhciGVXf4TxAgRFjLcYwYVf0G36zEQ8SXyWZcjD51gorx2MI2T6G2eU3dqjMM1w+PMPmBv1rv6Z
678Bpewk3RICeUN6dns6LbB9a1otrqkS0c5S3K2g87b+gvtUUdLL32HSqpZ02ZnimQ1OJk19zg5c
B0QhQZP9jlTjU+qg42zUDIJyqnhLWay7Gcul0ouENwBFNzXzCOTdsi0igIRBLc60gs//67SIoOkA
qQdUKV5FH/k5COxR6w+91VAfhW6brjdNUz/xKSIoXnF+gAhnGVctfDLLi5ByXr7j1sTntvPGITgC
DDcmb7/gkv9CYIyzcnEEn4EPzt2H4LZPiM+IDTS0VUqbXEoOid6QPKp4NNBXOZQkIZwRdTXirQdi
6KMJKsKYTEpzs4lKGmixRQXye/2eLqhPWE8GMPUHW1wcpj5clnZNtdvJgpWJD51GL4/G99PH0MLi
qHfyjAI9+zCN6mqPoJATXfzAgzw6APXGQp50QBBKhgfFyK7lGHTVqgLOU+qTRsOUkWNLtrj2dLN/
F4phzvMwLy1AtbKDckpRg/7d+YJJP5ryHg3wPrnnhMTbKK99JdMyQdJO1g0iugho+ecSl/2whDqc
zyyoXrwCGAgTxaLndCKRGhH8WgV5atYRtpL/5kfvIbTcm+viVSuqc1ynAJH/1OBlrmJIzzyInzzi
lmp+vpVHfM0xZJ28Cv4XhDDcGceHDWl1BIFFmncGM8ndRYxzyEksmqZfW22mzBp3Tzbpgso/A3in
bvwOGl6iynPOqtohYK/PKZhGtBWG0UgFFlUvhKUFefMogXZyl9iZciCNyqh7mwLUE00fv7oYPsay
wHV9QwsvLZxXXwLrJME2441C/PnQwEcMg4Mklsscj9ta+3Xiz2hmpA1tuh1uvYa+6pzeb4A0sHsM
VDXt8N13cJjyhIULGiddndo66SeEYUnIT5rI05nHfR8f0zJ2hWGZnFC/Nf0QmbwERw8CXybpoJBx
uKSW14tj/8ffp1qN+B4E0cUExZg2PiE3eFI7lYbk4y75xK83oL2DdZe3JM8OoaR/dqkDd4sjOCKo
GCH+Q2zWLFzQkBSavHGd8DO6GqdqJvDWUk6vZIQQSmUBq5vf0anyWU+ivPQhBQFr0N+Kc8qg7Z5V
EeX7CCfjss9BrKVBB3SRVv9vg+pVAfag9Wzz4pCvGZ3tgXBLJ2kzMnYQKKGHIcQyz//79Z3N6OSA
fOun+maTfLb/VRvpLV1UyBJAxdQQZ5pnoTNksy3zk/MA7mhyhLoSvy5+Xzkqbf7yms9M5GTLH9nl
18vn/09ZAzIy+59HXsu5scI4qmjmMvE1StbNiXf35vyh+bTUkkgOHhcnraFGstvIXx7uxHVarJ8e
Ie2DG8YP9E4KBLcSzsd0yUqy3+Q0QVxnEMFRvuNJg/0yzqCMHDP6AkSWr8dEwEeKG9Nqt7ZM+D/F
Zdft3K2H0yqMPeufqQ3u3WcGTvcdCDA91TKBxgCJ0ht5zuzrY5lR5xPRAgA6RduevRBnXr+ws9QJ
fDrDrLnK0pm2mA7DubB6qHlqzmG6PWCAHSDXPOXqlbe7KkVh5UTk8dLBiXCC9GsdB3euPVKLFG2e
HIzKGw7ziU1P6lFKGKmIm8ZlMTlbW/LGceRpjLX8A8TE6t6VJMO13w/phySUnwH7x5FjYt94IS0D
ykdXQWbt0UuHziNYnQGs496AByMhYMqmy6/HVCUBwmDSFCrGnNUNcrDK/XU3MwjiLGXGj8y16xpm
sqWWI66bBaZF9+8yoh3ygZdWlq45zWlmpRn92u3UHA9iAEG20ib7JQRRKxIKKuJJ8Tu8THHKBXxu
/cJSlHwq3a+6u7JO1uwaPxn3SDw/kDv0HBBDdYoUVeJal0siuHjyAKYOFbvEvoZ/Igug9ar0TPv/
52AB2K1+aPHQhleDqJ3RP18XwZowh0dWHkudPnDL4fTKUq09H8yysHE/0L32gEusU26sf2I8Q5fP
dyPcHorX3QTh4hU6BzKFZgwPbG2bCwdEnXf2tJAsod/k1RwliDhNk/bvDLZ62BuOp9LspLCLVjI0
VTkV+S0fZ3TIsEbRUljt6geJUOp4tiJr+T4Q7A3hPLVbWCjW9ahKmVEVHi1WmkSlzJdTvZKwTVan
7JZ2KczwcIW/Wl33pE6Y95q3iiKnEOBywfTgjlc+3kEPzaq3CLoUs+Mi2RlekuslT5f6ud1Wywe1
9CJE1Kor286hjADE8GRjd3Ofpk/tU96rYID7OPXj/hLBNpHxF71uDwlg/R0UJ14keko3zoyfJB0W
jATPUHQTjx8NX+swshLcNlMrfIM4iSdsPAnC2LUgqKTxJ8DGAuNXe4IBlRyr+Bj5BdBmdO4LJZtK
SFk6Ki/nZmHhcoeVsCedu1Q+U7FwluoT3gBzcSlb+kjUBuw+G2oJvd5LPUnP7euVxaFz8U2JZo2l
Ivt5xTv39G13OOl/U14f4qx4nv0Hv+1aCCNk27+vsP9+7yuqEeQ45ppnjGXTpYFTQrdAE9pNMCle
kjUoU9gqRfr5Rr6PttFfvl4gTTUMgc1nW/tfTaIX/jBglDEyekfjEq7CuH9i+Wqf4Huas/lFnDRO
05HiSC4MdB3e/vimT43v+cgGoBjnCrTwiERxh+ZJ6ZeIEzNgWVFbe8BK5oFwGtjwvxkm39NjE9pK
KUDCTiSdVm39pO2wQevMU0xG/Tw7tHR4RuO4IX7pFdrQtfBXl2+Ffj+AF8aCI0KBkP95swIpwsbw
ohWdyTKh3QSPEcip6faPRHsI7yV7JQnRCyhosNIJqvHfPcYcFkFDREo4YgvvAwK3uBnPfMSsjJ3c
oZivnwxQbYq1ajaLYW9Wu8p8wZT/p3y7tJNiIAd/UcGrXVgeMSTrnBnwyeOrmq5M/dHXnxu4osea
642y7nIUcB6WLo7smP2ko7wx1QCvcENrWVRtHz6ZQ2SHXWLuOmtHYELmErWnClLkP0iccJIr+jL5
o06OZH2llBuH2zQho1butWc0zso9ZgIR56N2jYUFXB3PACdQ0I9d6wt4zQbWqZXqL3iktlbktV/I
QP6vLYugjpHuOv3g/eqoAaek5q5t/uzyuwN3COiBR1PWm3FrPh6pScSq6+bPOJAg3LLkkSdI2cke
ZaFgls/BwcAG6S2xy6R1ztQtZDGxt4+fTMy4p9wbaO03no/nSsYISV4o350lRC0kqnYfx6TNt1WB
JdF3pODMBg41tziV7BbUOqnwORkRNs2EUwuONsZlm8W33AkOJ9qsPRR1PPtoTDZ9r2TyeTHM2YHH
shvdp4ZplN+ma8xrANmGuFAL1nxF1LdeY99aeCdiI5cH3+1bi+MBXGPwdyt/GC7jvEntD6SlG+iV
LFEIQOGWR94xFWkj4PmU8YlWUm9KuYbLUJMmY+WmE9vkMS6QKlgKq3Lu83XPMVGhplUVAVWXJxP5
VHtvubdfcDTdj4e0N9GwufsiCjFMnJeYyxcoCx6yRzXDRGJ2wj9fAIt19w5VzcqivmfaSYZAYhds
byqkNNkFRNyeiNPp0wnqmfo3nel0GsWh3fYOV3Q6gA61yWTsvxcoky7mGDEI22ufgULAZrjUIUnZ
Z07GuG6CW+iPlNcheoUjfVkYLOhgIwMgtRE9TQUV5/Jrm1j3OST+/ZGpViDLzLtcas4qihdY4K58
aRsvxWD+2CHVbSoiGoyUiXiGcQf1Cv+H+m8huobbAMiNT9yLH+v/JCAGEk16D1n/e2mD/Aytb0X0
wSCf8Jh/F5N/9W3fVPoUGb6vdg3N3BkLijwJ5BxsfuWAPFqsb7jnbn8rW8JA9AbnpHKqP5/6AjHm
zBtRNCzSA8S8dizdIGR+tun5vyZGW5PF/HBspO5sCzmFhkVo8wZoi4rO0CzxTtOFt6T59sCpLrry
W/lhnt2XDkTFNvGNveypdLXbFbwkm+RxbKcvjMrszi9qBtetQzOocFcOBWJ1FF2LYpoAVlwLlout
Qk8u/rmqK+nLYS/StS49dhmbuZE+2AFacE5AmV2vgB5T6IRfoUF7kyeI2CGbUHvJzqH3OMLwNa/H
GMGXiBYql5zeDWdPNIm+6u03MkOCG32XeAnm+fp0dPVCFG8qlVphQsqE7C4AolXFVLoz0PEmRVtM
pp20Izv01iowKhTItKxUQdXrgVC7osnZLbi9RBOt0sg7bLYaWr1NrSEE80pwsscjv1tUe4Qay/Dt
Zdk6ndSqolxWL4eYxq7BSO+pKpvXF5Sy2CCH436h8kPGEIygj9r/MA7FINLuBPHJNyd8fdCYrQ6s
JLP4Ds8H7uFwtrtNjKlXkFxPHyQvZb6tFUm8foz+UvSUQjfzVFVFez73nuNGGJaV3g2XcTpzddxk
tc04KdHXh0nWQJUnW+EvE1fuAMrtnmkCQWuxqgUilRtgekQ7kgXRtn7nKaemVDYdmr+KCOFFF+uI
MMC0VA8ji2d4jljsyoe5JBPR1weOw2NOluqYavWTqkYbh4Wmw6VXN4lwVR3ennZMLXaG+dqDQl/g
b6W4QT05G2DnuZ1bQCSeZOBep5zjgCabEJMnwn6jg0OZ+/jX7VbDH6QBcHP2M1K7nNrTMkUUEVJY
nmoEIPV4aFm8iKfcMmkaFro2QVnbNEoh9qmGQTXhLeeo21gQdfADsZyus+WgPrONKpouc4hJCSRO
1AyvOrMjbebGfJJBgOYiD3fPfI9h8CvaKrGZdpJCHKh3pv6zIyQWbO4JiSzjrpUdsupuO6Fo0Ig/
a1ycvLAnNtDXbXcMR/gkw0FYXpKNtSKNNOiU2Br+uOMiEaxDqUx8VtQrpbniXu+80Bd1+CB4g/Go
D9dUPe3VdRc2tWH8no/b92mf8sbmzwjLAaVNBCEgchCWXExfKG2BP1g60YQfvif/uUBVaCSyXMoC
+dIHAOzLCIfCGP9CrOsoAe6K3nMiPxpnOeoAtw7D+/aSC2fhvupFPitCwxwqk742WifuafrycdyD
spX0TPjm8pEt9PmspMBqGB5J46dYHufME9pCdYbxmvg63fOMxJWrD4P9OKy7qb+yCg8PewYykx74
Q/r+FiIjcRVhypkNbV5EvZ/hPcj5/zYso9dDUB63PmYn20zXJbC9ij/laLtGrQnckwcgrgaMXFvv
tjDX//rfb5cezLGj6KsVG9Iz2fWcbRBa1gb6ZlKPbimxjRy5mROrvmXOI1mFeuK0A7Z+3+vwVNn8
7M6iugnrBubgGEMSpQ3xT2PUrwA0K5OSYKsLEQL5oIWw0Ppv6QSdUfR4DRmK3D0dyxS3dgo5luBo
ozZA25jpq+luvU3aKndT236R/ReBAk35tVS/WSl10rhxdOuSF+qEydLjMGEjFaEZNF83KjnFuq0H
WoHbMNQSab3pvx4N6tDb0B+r9fF3XWB0FX3ITjOBRaALv48yFR+VTaTmtwYM05iRCC55lMPGHKtw
igGrqL/RxgGTRYjcolINywcHDUKR57aM4/5AvBjdtAjzKjidsf5mV2LyDD1I8FeGaEJMWStKh6CT
Robq640ljshvIox4neqyO/i3N0k1opDl71eIFo0dGn4UM9e4GhzXnrALth+wAQV5gtfVCNO1Mi14
7ASvwRm1zQ/Av6FsBSjbDisk3oRNY3NkQZXKwZmQksAWpSl2/0yFcs188M5ms0veG192qyGGYM+a
0xWv9b+ojgv6s+8E9hpi3fewAN615GY9s8WwTvEU4Dh8XaKeqhnLUrK3p94VV5ojxiX/KRJGvhSI
cf0gvOSYFKUZGJNrc5hxM+muLzQwnfHVJXkM0c4Ah/PtvdnJNXdaNr2hqEEAoUCNUntKZjiKYom9
FefOZqBEzgOz+sIw/UzmjQmSyTe0MYYFO0cuyjTSx03ZUe2lTgoJo0PWw46lK2oyjXeWdJ9Rc8dl
MI4AorAy0xaAIj3twfF7imEzmAVfmfl4YwO+NN4V+3/37KBzVxcyceLWUpGSbkG3nJUf5U+aJLLE
LU7D0sotY/m/4mCZ4+tHYHR+mdmIzJETUE1ONjXxgJkUoLOJJ+qUU6EAKm0mW0pNF+TohSGWg0zC
+Ltlxo0XbJyEul2d0Vyd3ECohMmT3QGEVQ2Q0MKVymxeY5uGDDiiSls947VrjGDTOIWtIJSdZ0P9
ftM0zuBpcHFhKLpzi4FVDFl63vCBlQbX6caUBzVIA8qz40NrJEvKjwEPGVnrhFyrke8d5YpLpIiY
3VulVzhfWBNydGGLXUfZr4JAxRMCTiRtsCHvWqu/XOCosdBA8zMNzSOPPrXeU2fy+7SefqXoz2gU
2nYvSWJrFiBA+4H/mCLSwFR96JqQSFYtgstoXjt6vV58Y9vGR+MKvEOR693cjHtmi0FYfpGq528O
9HU1DM3o5UR1lnIhXjylSm6LTRSLo6QW8EIQkj2S+5kIw3sM9urneN4pNshoeZHgxr5mLPXI5C+e
2LpXEbqPSRrJySHazUUm7OxdExtbblPOfiCtm53aR+Qf/D0h9rSq8+iOVobdaJFaksMBaBylKbHV
AEyav3j+GtUZECAGsk78wjcyX6o40h4yCHy/gZFkwwnakhec/c9IGYXZDjDkueAhYPFVooF1RYaZ
pDi+bszSJ3xldFBhhiHlvVN73eyZtY/6vCmzJIat2nZYddceLyyZep2RED1htFCZL3FnucULCqri
3knfY+ONM3JLEVzXssD6YX/K/hYP9partYNNRzMgFECwLQlZJq0sh9WMxkY4j4OPoqSI1eVRD7yk
fsuR7Yk9zlAPsDbR+rgr/C96lJqjiMrGoUJ1UV3VOaQvCfdNhFk6dF4sEuaPK720t+qLo6E+dFKr
SvDxIbjgpm8SitAL628hvCbRDBtceLV/bjpCwLrDQHXuiZdqD9ZF2pvVZ+KnXzPmTgFlSXXHSr6v
GBV6yfT03Q23BXoYYmOIFzFR6RCiFAjCkGOaIYspOOV1qi/9E/EpHtaFbAUEx4U3XmGDOj3cU7Eo
MQTWCclkqf97QoW7UWTgPDe/AMfySCOy+NZon19kn/L3nWEVoiZ0yD5Qc+7uk5eN8yST444ZkzT7
ClXhOg8aaYVrEW9UFtbUxkkcOYsfR5Jf3We/V7Dnj9ZMjnjV42wRCthOpvRnMDreyeofL2PnpRdH
cgGVw6OgYNEIwEMEzTIuWIvfLQNhczQrm8BtwHCHSLUD6tcR8yvztNkPjdsVi03B3FhZxNjpHria
ptY1wThF13Vb0a5Hin/aer7zq7WgKnFxQ7SEe+PkmQ/rmINIEOgSNqOsM+xPcHgc5Dz3O/ZRx9CD
QpTiW/nx9FSo6Ut0iopg2QlK63cRQMKLRzZFFSZL7itFbTIBi3SbHMpcYa5E1SCmv6xBI5/1Aqkg
+RoREiTOk/y0Hex0QcIfeyQ/0jSwgkzlrTQySXHWOggNveNOUrlAkeaTqoJ7/eKDdZDwM8To/T7p
eTJ1V7VVgKk40k+GeiRBIBPrxHw/AbguJHWcn+GigKn4WsUIpiJy0CCx0HVBWoPokQMW0RQoVSLZ
0C6VoA9ZyOk92XkYIMFmaBJw6CHYJGsw0SvGWX1Um4o9vpMeX3zJdF9QhcmWUko7+XdClnNULil5
xtHRkKJeYNH3mkXnkcXDOi7vHcEsyAFz9InlcFrykBd9OjwcSaHuHXfZ3ZqdPiN3Nsl0fhA6S4xu
tylPA30cUgi73rTk73IAyjB5VYNJq+sNwQ9/ZaOZo2qM5tMyuAVpcAl5ToivgjVm2p7/P9FzT6Pi
JgIxW2ycbOgywmXGBmMIYPosESjggGaSrT3L8OpcLup+IbCjo9QPFisFbfUYgR/Y0jdeJw1SSAc3
0m5ZnddBLiPrQDvrfIZBOo/wX2Ub+m80WgTACDdvHjRWWSOz+YnCTIrouXDe4y84kNgNsASfrLMH
+JXGn8dtIV7DK0g099jtQSnV2a+KkodSocWqewJS2b7rAwPKB/GLaIC+IVhPXTw99mydN3AiAsvc
3yeqH9Gf/Kj2EPndTb/8J2XLKtG5b5OX4n29uvg0zhStxd+gfSjXezlz0DPL9bwTvTvPNgHIXtY2
dHPw1deYVF8hFOfKSx4iSYMnFKYmheQsmrYVdXL9s+ag9BjvsCxqdR2vnlypIxTLyvirsH9ERYC4
lYOlCqFEghZDWi3iiaTUG8ziAqYSiN6TAAFUWEWzH92P/uqTeoF6QzBJHRbqD/as/9MDUai+NExE
jm5C5txj5mry0wpmlUhVLM+a8EK7ar46SCwUCOe22C4YOBKGjTREveGMOQ0bcYS4T5y0ixTEHfXE
RWYykKs6c/dDl7ws+XsEtOlddtFxfvruivsaodJScLEuWSTHx2f2Tph8zHuaD4TAedlm3vDUk8Yf
II6RsrLB5PQFcBRGPRABvAa/TLPVw0lQzGROU86mnCsWU9ThnQBuWM4GqdUe0Oq5oCTodhSdS3kS
sovg/AKyiwY0HQgeQbnGDk1lVD8AEbutbEbeBrZGvJnaAtkZK2/3fYB9AoGjyaI3IRT8LiUsuNPy
K3U6WpYvdvF2b6wD6+65XAFr/jgUoBnk64J36vqbQNZKgb69weP32N5hA1PIysrccE7gQbUj0lxU
fFSQqxxSqP03n05re7kboXQJcMz1RsSASWHmpWbGbIRnqQpMESISaHMiYldeDqddN9WPQiNR0aGH
d1UUbdH2ammZpgApyCrRvGeixabAJvMvN+ORCAcUDqAIn0SqJC/4cLXE2PiMLrQALwJ0zYNV+YmX
QgPPFRE/FahJX+Ut+L5kYGYB7oFZoyCi5FWGmlCDtVZr9swigPT3zuDhH00xIF2ZNQEh7MozzTDv
vzhfNdCw+D++iDL7TebAWXt4kjo8FUobUjGpW+o/q8FkvEi7/G72w6V1WhJoT5kYnF5lECQQhaNB
wxzP2S89kSkvO9HKDMB8+qfyq7hSE96eXlplcbtefYB64svgAGv9I4aPvR6q4VJNcRzMbOsRUe9M
kSbaed2c+mPAMDK05zMnT+7+7WlP5VmD8klqYuTDnw3dVFZnWyUuzNOeWqOfOqqgexZ5Mmn/aY8w
wRh9Tks9h4kzLKg5UcjQpXhkpvOELYoA8xVKmA2Yjnb5EGbYNpoGi72bhyZlUOCQ2Fgcr0sNLvDe
32GcVfjVVycB5UtjwlYBIiOOJfK+yK5DGDnFSZBysXinhCo+yY9l1Ay1UCovpXH+nEit0B9zbyLp
h45moN+xaCQWuv2Nvw+y1HhSbgKI1xNhjIQwHB1Dw3CEMcTV62zvQufnbQPQAYPk1zpF34ofYDXE
w3EHy3BvjKakSIjXbydlUpMPVhlcfZoZrHzuRFSFNkomw2FI/tKj9vhjhmQiR7JKWiUuWV49iD1X
ecUquVgkSsSUHqiw85cJ8QbZL8OS6B5gWgNZFBH3zQ/kUYL+JgIceILeqqSZryPX8za+vz6+XOAh
o9eJhXy4IYVhROAGHvZJ09f9QEr92jyoULzgXdWdVM7PRP/0vg3hwHzrZvVmxhLc35qF7Sw9OLs4
2uQZvpnST/QMFBMjB2lVsZW+gEpkdUrmKqE9tbgIPQOy443FoVjmpsb5Agmh3S+mqcdxbRDYhr+2
EtuLdYK7AZ5gWyPNXeXELYEfWlwC+bKh2jRV7/eAAySLVjF032c8t61QT0np2eX1t41D61GIcn6Z
5jmXQ35L1vImflgdXTGzGkxGgrux9PLymptInhUkMfrPMVpmLGaFjNhTWiYh2YEYbzEVWo1gO4VX
YJXRAKd/npivrIJxG/SLiAq1RzbBN+QYaytycB55zS6GDrBRIO5owxeM3CsloT9nfpYaj+aVcf/j
XNYYypu4orfpfUsqNVKfOi0a3GLog3g568uC2gmw7kUcFUpChqmmtX6Ajpr/ks/R2jX2fH3a8SnO
6oW8DG1pb/mBkfoCXIUMlleYdYK3IkAMpRu9dqKX+EsgrMOtgxG4ujzixYFdsiylbCF9l8rpsWr/
ZxU0WTa8LaZWsqe0T9Tnjg1FYrQUurXsGB8xaxObNUOLfhW6CE6RBbbWoitz7P2+M5KdPES0mckO
JzWj/YXwnDcWS384knct4+UiQ7eqLYux8wh1fgmzLjGJwxZP9lrZ4Tv715r2OBS6vfrGLFLnixLe
u+kJ9Ao/JX0l6rWLo9zvKiU5XA8lHIosujcP4WFYDiuJ3SEp+zOtX4IQ3XE+Y37Sfbv05mAWqTFd
ERsc6pbL8g/SoXE0BXhKJgSajtfwV8o4ftLtpD3FAEbUCwixEmZTnUJYtL4zlw9SswsLQR+wl0ay
rT6sgYn5jenVedkFxKtwRyykRNhok0AzQTdwotNodF3qLZcObLaEpDwSB/Nn3VXrbXmrAEjvA9bp
ID6R0jmxWm0CwN458VkQ6+JQSXfdnSfvj9jZ3/lb9q1EmIUrgKbWfE9KXWKKBCbNUCuYuzXLfEwH
UqZj99Tg6aZROBy/UiHbJJ4SYU0aso0YoYEavmxSuFdvdOu8fsEKg8pZqoslCm3NX30NXS8e163b
XIdU193A+IPa+WLDv/pWO4Kx7YKqWpzpWVXq4KdWzJOAmiWgrWSkR1IS4Wp+V83K94s9Fon3mppp
riwFmnK3EeSLariR4XXgCzHq+grlvusVq+kmukHPXLiFqUKE7Bx61vY+4s/2BVuOwU5LcaevHdDs
AXdJTyy+cku0ynncSt4jybrmVTicBFz4DciMohoEO5vAdsIh69YIjKqkDDqi6kR044cU9ov/eoHr
ovf0kKB4Dy+AkVnXCDxY7JXP1qTOEiPd4bL4cnEE/YsDM/qBwlIkAfcK81XUFUY6E5BT2B/EKTnP
UBzO+b2oJink23NWTTQoTEIP8jeEhjAhx2BTKBYE0Fqb54X+RnTJag8FrzsN7KWf64TzeMjkDd3n
powbvO/V/TKZ/2YOh6jlNO34YhOMGrfkUee9XUA9X8OdPai1h2mM0FNCRr848yHICtuQGkKLR/U5
m0MbTlENoG7pAas4+Co4XcSgFOue90l0WMQciLk6ISrygp4iAyOLB5SDIfEN5nCKF8SGwNzbgfZg
gKDQeF6uJXgsqnRTe8lMzMo0HHfl4tN0rBpam/wAeNgZAqGyu/Te9LkL8q1ruxAVmUuN6x16B/ok
fM/eyO63QxZveU9YAm+A/Ku2jJ72L+7erx0QGcfS/8GveY2QfNT/HhoOyoaKkdMJ8eEY+52Vnt5N
TqSdbbdHgi4On6efnQJBmlshqiphP3Sph37mjPupao4lv7l39vbNjWzLmgTfboKyBItIljg/Tev6
jPJgxGGN4vJJeLvEW8mefwUCoNU5PGFZ1PcUSyqfx/E/fV61t9myzMdD67esFJETYBU+TidhI2y9
v7MI+ow55GW3FoOj3lPDuSWYmzBTJTbNWXfLdt/88txi55BUVCNH93gffO70D2WDkqaF8ILSMwlM
ed+upw47wBBLGO8UwEoZSo5wuX3vqEo7FIUH3xz189dnJqXV0UYKgqG7h3E2j7DjyeFIpBS1lzls
2osHxW4Li1m8tGc0OdcWatE621pg4SNECBUubfiERQMtH+lWsh2tP6tRtbsY80ZEPUDlWs/YgF/4
QiT9ngiLTcmadeJ8MdFcVOE6GIYCBcIBsr/3aMecj8wOoPCgIUG9f+myPucqzH7dmWNPNYCE+VSA
tJvohru46EgCSqqs/HY7L2Y/PylAvOH+H84WtxRsB1ZbSMqoiXP4CF+TJP3zyGX8KjMNFvBOhgCH
d/T88qgCKBizC3sNcOXqTWf2nOuSOL7WXeBsg8fS7Q0k2SLVPkG3I7yJKxGtQogiNPhDX0ae88YY
/JcVplnphEPuHG4o8696qJM8tZ1JeeMU0cEUPzbAnsQbAE520nn3C+YQ1LlHFlX2aWS8EssSGW9H
gKIS0c0g6ZxJV/0d++mVAUTHQPYBT+VYHuUhlKNAMxmuIzBc7qNonz0fC8jahVfjGmi2P7SrJxC3
LXVd8TyAZVe6qGpoIia6JbzrJgw31jWYA4AnMm3lJzjXtbl2Sb/K0BwXo3S1aaB2VwJ6i/BQZ6vr
C7+TRoat/1oksJ+MaPzvzbhpT4j41sQgiyf/7P1kC3iupTsnZ/mrqcgN59u9nTNjBI60R/BrFtms
crDOYts5AWFj52hdvxCDQZfQoidiPHMZnMvqXQSHgG0BDCPcttWSztFtxOy1FLT+yD/FyAizM3pO
RVNPS3kpW08Ksu43xa5Jl72E7rWf+c2u0+EhiV5AqruVmbOeP9ot00DG8idrO6C8LMyIZdAve//9
gjw50uKThHzYEITDcBu70UTxithYlJwsaFAYgFwxgiEBHST+vEWeenWuoZMPrTNz74/WkmeVF/Tn
GXgK7zqDztxFvU8jHY773pnBDpJjkxyPfYO5RsOEPIrGt23iMQ5/J457SzTICiw6ISnuzWDmloG9
UGuxYSijDLWMmmCYK7P2gGcX5/2otKJ0YHS2vHrIKgDBxSHVZQQFJX+YmT9vwyyXEWm5WridR646
agUDpQt9l4ddA3jj4SjCBX8CGXpnF6AK23oSs9Yj/29w55jlA4exzRwOOpRYKOZjFW26b0y1ynAj
epJymQToo0tq0HqvM/wH/H11JhduqyZkRTe8dMjpC7bNlCPFSuYq8uiqkz6abHLlAIW4rXx0d86q
vE+KGOZLJjA3xoXy1uq/pCeFIGve/m0ehZmjxDeejHIiZOZ9Cr3cd+6gxOz8aSKYq47dYsd/qU8Y
P0c7WE/It4Xy9dOP1efqmFoUAm8fdIwf9wLmflD+UhG1TDwOTzwo9ovZqOb68rkYFDOq6E/HRq1L
3o1ZQAzcu95K3kYcEtsFmQ+gopslQ7b1fsxPL42XJHU91AUgukHPuHZ9yFlYIAqvpppofmEL/Ga+
3uDHnXAIqeGDsvxYsjgcEcwdDd7xpVlNvaKoWep9y/yAoiysxafqOZRn1Q7JGkwGZg5oCsIFTMqo
eUFvsXXSY3PNZGpgw0+cBqgnmOaGqmmd/2D1OMxSUbNMD8Xx4/GzO1NscwtWqsiCKDPslJoOaYe8
ChmmqP/HB14BwieUPGEiScdEGIZxkGaq72st/5nKbcu5VihFABp/xQlAM+FD/T4fUjqwTAQsVnPx
aZzkHPxg5q72UAf2R7EmNt8ARSsjh6av60DWNr9J8qxe/cK+1SGNsKlKY5Hx/ukq0FgQWgjMdl1T
xvXUy3zVf0M1mvnpLhP1FhsU1827hHhUovfs6JHIII5F20r5QR6Ylb3PiJPlpBOQnMJodkVmcLr6
Gx57/a/meFj9JiwB6huKqfYIH+Atb6GscjkmQCAOhlpxxzh+LPttK1KZW3TOs4B4dT4ViANos0dM
FccyB3LyGr6nYqWsfcb29el6iOrnUFCKb0IserB1s/U8KzPVm3Onhw3CGwfUniWW4OORui/tSAny
5garULwWOyF2+LbhXZQBlgZXRu6IskZiWHur8KHGme1iixh6PZuS4e3WPmSFczcZhvfWQWjSH4GQ
5vRQrpAPSPNgoGhNIl7QCKEutaVcDl2vk3X0opxV3FCWd1gI963ox6bJ1MDAUc2CHYn2k3viGgdt
yF+lbkXGa9mvFXvHY4IrqDHXvPoTfT5pGvxPP4WXUst7WrYapex5Gu2jtzOPC8kiHDYcv0xL41TH
gHgqWkyON2Z7P2V+j9dK6BmLa+H3Jf0dBoCMF8ESbYThV7kFm5+ufyyUR4Cw8HWAPdvZ+Eu/jlol
V6b48f7WzqHPiCIcmPdjoNYHWRCM6CjBQSmb3UiiPM8rqwNehIZGQc/RBqYe0KaNlw8F0lZO03Se
FJGMlAB6DHhOFZlxb4FnFQceHQz3XTA+RB8WNgjxGcGnIgFXvuxB65f3TfsqWiZWgYBIjzGVdEYd
N/wAwfIe15BTLlXrwJIUXY/tpnqSqvfOzOg74gf31Jw71vFD3BQ0dmJZPUJdnM+IFTPqSkzRpoo2
fE49LbP7BZacgzjYd0qRSW5FpiacUex2ct5B+ljgt9UkmZCsQ7dPFLXsvp5+0OriMo1WzvKaL9zp
36RMQ2rqAtCO6tT/Uhlxs2FzF7cIBUXdvNG7d6WEEKp24/xSSQV+BoxyHIMhs02tzN0BdLkzoZ93
98gfbXGIVquaXtVU1PLionaKxpfdIl/8wgSmxbFLpZEoUJdOTWV+yZONVPeqWgQCcy9p8M5xZG9N
mAA9dC0TP9/MjigWnnivtyCzLhoyp8TfsdNh/3q9F6qq5k6O1ToRmSxO6z2oSkZlkZgSxkZ+m00I
R5JQN+11pF8td4khRlAA3Gn5Jl/ogUz85ePoenh/cWBzgsPNjFT2I3Gq004xDaKdnpkdal+LKUY2
/64EtwgzB040TkqdHkaWckdwuauijwVEef07qP5/GOI9CakLtEsKmnmPRTATC8qGYYJrtUJSpQdr
KGcwQE7vYrHf4rpXOYhJqPwe7EBswzcBz6R+hkLxbNLPcHKh1Jjn5Snm3UuaEmsBhLgCuA+c/AIC
r9YLra4NpUNVCVJUg4sHWkDt/qKhTScz6RH3eeasKKyNGhp2Y0xGabkci3A88vUV64trdplFbxdn
N3n9Z99rdPyJAwwSawoM1IAYaiCdSX7OBwsHmuhX5WsqeEiCvDDPs5ZfKj3yhrNzSmU0i8Ni0vu+
QsyZz2f3HUF/wShAbkTtNaU1SaX0FkZZIlnNrVvphFFfz0PsVgV7CsR2lLxAhf6F12S6uXgbaIQq
YMz6/PfWCaBRTaOfIwBVK5MSDKxMs9PgcT2IeE2WLtze8tofWDfxqiZpgvZ8evNk3LW/YpDqU0nv
rhhoDkbnZsV7/zu2U90sm5OcA++T5b9jtP66xCesSD8L1exa8C1IjX6qIlEJdimKMTe6YX3/3h87
/MZza6hztWAG6VuRZCMbpwV3RRkGK+saVmGTciBVL2clA0exqfoIsUgVxbCVeVhnOlur7jChE9NG
P0WjvO3a937BH5iF8UkhP6JtrkGeu1+gQFcTSrcyk4obCYEzSdVbaSanSCCMLkbU8tWtXriUvTBc
qv1T/MyPhG2wi7T1gvHw3ZdKETQ9JoDVMX0zp4KskReGQ6Vl4SzBltXRLwUf9qOLfXmQtJu76Qyy
4dycKuL5HER+4/dnqrSKTY+zr2dblU2GXHdmZ+gDRrWCKefgSlXLjjvANTbN09c+DD2axXA3PNbG
Jers1kvkUVj815dU8fmhSZC7CqZOwes+NPa31BSAQKt1j1vIM2jYYN+EhJThycvowGnrg6ezn2xx
u6xY1lPrpNsVp+goFwkdyi9Unpkzgd5wYLdli7mKK1gu+Sw3xvsLY67SP7ssUYHwprqCLTAStGRf
es8+bKMFgO+8UpRrLdCSmqxraQxgsFiyna4u5yx2W7UXVTsdpfIZ6NFUImTBqaL30mtsZHkG2wGf
lN/Il7gDbRQJr8wo8r2fIS586RAn5ols4y/kxpH2uJERoenY1i+vpgcTnTI70YDeIXulzwJncI54
qPrjfwfC4Cwm9imzg2POgLqK2xCSIa1VibJETAPnTKIXKj2Dbs41EhUeJ/L8nEpH5Pr8tgNOpZL2
L2GT8gLKTY+UWSWEZKr6qYVdz+qrQs7qtUTcIfabke4nsckQ0GO9TaA33ImMAz+wgb7qV/ww1IWj
G8bhTDyeSeJ8oKh2VOeH6LvAXjLliBBzGW4Kvg7XTELXZlIVSh5mE4anVzdmAbSC5KapG+yKR8Bg
rN/U9i4NajwBC0GOdDa40wwndOxe64GNUXL0gfDP5Zu8INJ2AcJvCU4EldDUL5sG2VWxIn1/Y7Jg
/vLX5JKKG2Bat340ZSptmWmYI9wrQ3isOEyxyZBGzCRGC81qp4aZ1hRb2UWcEAw7dSSkL7cINwMj
BxDhFBKwgrIA9B4xhS7mVLpLj5PFWO7SVrb4Av4FtQlUZF3Ht8yZjb+vYLhJI/K0+A9NLV8dpgRA
P9DModlenxtOuvSZFne3L4KWL1aRGGLGa5L4Q+Ypxc/4BobsaI39oPeo3ftG+HOu7jLNRuB2FzLr
xCkvbf3lNZYrQKXr0ND8pUHp44woSTNTUuIM06742zm6kZfLLkaUBNq5xJwsGGPPQVsxyUN8b3my
/nxr82A3vBZXVLhsKgG1JAKvzH7SpXCmp1qX1aNKqu3ORRWLJK4/9n5ySjHfoeO2+w6vX5q3YMph
aHTjic3j6WCE8yrxn7/DyoR5sZMfNM5c1UEDUM3VVZR9YUlj0pb66si92Ss/LYh+FLoBwiWqTdA4
otn0Pqp35miiPZ96keHGh/ovrUVpGggmjfvP4V/tq9o/rXgWyTIsp3DyzCymTV4Ryz5LwcIVj6mS
GgCXAFqtF1NSTTyyBFlW+LKPRky2oaZQ4lScSZ2XdL4fFqRRfce6vufkL4UyXVh/c/BSzekUdZPf
HEv226c5aLLPa8Nkzcwiv4FuEFxBAmwaV9CBxZW4W9yEPI49GEaebWEfdfo9G1xCXarwUMotDQ0H
XXHtuwmlPjUuZnZlYYUekGSZw0AACmXOdrVI74eHtJTL7hjasGjCqKh1sAkGlOF6Z2E9lzirvTBq
+f5PX/lm6ELs8nmBsIcai7Y+sZkZ7f2UbQ27ojMYPvtsFrRNuvbQ/MHUEir9DzqUFCWHa1ymvWHX
vsvO0Honsi8IFbKeo874ipUa7HtTJcYMpuJaAnY41yGxnC2VPfKA4inYRn8kak6HlPneu+Qdprw2
9NS5oIcC3HX8x5TIjXz6lZKeg6Zgz3jIxDq2n6d6rShY/0mwJ+bIr1siCx3XGNsGibC2OqHAOy9A
+JwAHtWBhrWigTm67jMsMLss1TssDOCjYsjPR3KKo1JRnn/Quju33ENHxTcK2fP0lDlrsE0ZV4V0
0jQZs+x7BAPJFYNXU9Fk0iElxW1q+GeaINiSpGWHa0rUMPgih3uoBPxT3TNaXNNfh4FYWG8+GOUA
nECPmFGZ3NICpvfGGV0kQ/7L1JtPxV1dzSz6GVAeFErVWUXWKrrlol+eJCt3fsb2pf5fz4UBD6rb
p1xQB+IgtgNhnQQPTmXRkVRs+XZs/sCKtqlhAOvIpvj8IM9iejXRor6pAsPCaviA1IjZGSLdDWLf
LmEnijyUH72xSa/BPh88tvJznS2ljFLlTesXMEck1wNDMtIT4x4Lrh8XyTZzHk6eaJX52axRbxJJ
i8lgiAnlg3ARy5HRMPrRjcHAFSSLNqlgtsdyaD+R4w4X26fxnDGVVGX9LOAz8N4rEBbiD+XTOfBp
0Px/iwTY5M/3LCjg3tTmaxxNT3GB8Rwm1BHHqNXf87mvI7hS5Li+C5Ptt+ZnZlOQ6PLbfGD7VKFX
TGow103wPVmqwbNiFYStKyt5nCzf6IWmMaEhOTmreldTGUWMSVm5jWIziyIg7BH31uXhxQObrNvQ
obU6WtDio8E9KvED5alWWTlYx51ME5wG653XpkAar1RIzYM8vtm5ukCs0CEDIx7kIPyXVinyKzoI
KC2aU6Ul+2gsr1eEHTasy6IkR8jiNFX/9Mso30P30SIyEotUdbnGzcLvlIspn1LUvFRih9H/nWI2
XfyRSIE54Yz6PdKOs8EdhHXlx93v2D4GrqTnohbmU6DuFP2dZS2bU+jpUNf1DTlPIc20HH2akDTq
e/Ap+jIAYMc8U57GwOTL3Qj7kNkeEM0KFJm2cN+SPouG+DAriLurh8ifyUiDwqMxK71Lp9Uf0kpS
D6JC29bTj/nkj8dPsDDAXnF+79Oif5rpKpZLtt1sGxb+tveTNF/Rkb+apO8BAlE+tq6MPsUMUvlw
i4ClNC7d6RlWPKrMBHnzfQDob8IuliR27LR039njUN00g0onnW6fo4SrwwBrj+15nQ4jqJtdDOJH
FqkZ9RdhMjEkMU1YRT2eCGk/tl7qwGo0nDKyqh5OByfNx4lwjmBl7IAg6wEf1CTOjrq9SQdu6/a1
sodULoG0YLa5HuAcSjUnnDFim1917MBrwaN5GhsKP4nc3YPFCqj381IsM5/U0VyJQr9p/N2zPf1u
fgaB5GlnwmrfonWE5LqyUIHLMbCCKHB9mOICYtrbExvSbFAy/5nVdZNlcku/UoRt0WHgHS9fvmZC
1F7kMKNy0cIKIIw1TXetDuaPvdGbyTXpBNbAC4cUKHtC1mMOeOj0ObEEUmA9V5cvunZarYIcvvFI
e5mYKfXFZs/IbAWECCmxbITnvoJaUlNVHsi/FVcrfECV6nXeJ8WLz8Jw4IAN1+pYVAymbhxaAl9a
jz2zkDt+afWgXP5ZqNEwlCWrhZL6q5cdKSV5vSQn5aaV26ZIeV2Lh38mlte2PsWStUYXbM1n3e3g
S+eFa1gCxo7M/y7yMPjMoENKm3SPLojkzYmpe+0CCDbokjPdXl5ZClTFuHiqDE9KHbptyuFw4Fz5
q/E01KG+zgvokxi4BUavyfr/OJ04jN0tKu6iaLvlAkeC7LAUr1pzD0QZMcddAkwe6B6Tdk6xxjMI
ujNyhcp/nIf0IRWAELxnXKbDFpgFCtl+VNLB78mJGdFJo2NYSCQDT3jnbNr1W6uKwoxt38OiSM6f
Ns3J6PfyHBmoZgEzdaD3gsGwjgls/Wsr+oUpoBXwbUq5kaahTt2DnXeUsBTcFxJXVSr35SpCUfr7
9+5Htjpy22rqvZbhfAkowpH2FptGok1Rg+heyuB929j5Q+MNEDtenZXpMf5AKbnxUBB1XOEz6L3d
fOjVfMJCCoqGVKHz6UtO4vKw0HpfOTKsLlB9Y5THHpRimd3MaNUWQgCTrhsRbpv0ZCJLDAVS4BSR
D7gyGPzjTJxYmGUtaUWC4tNoNgedcaUJZgisWNoCobfreV1xabsD5/0ZA6TMeOSFbD6H8/ujVoxH
ivlb6jkn0g95iNgFo35/GmuYdyBOWVA0HmW0q17edOS01PAYgVBSKlf7le9vDK8H+MIb8ccu9fBM
8n4pR0RTZh0i1RBs0WYkn9UJarPDSpbgMgAOKk9ZqLZnTiOmvcQzBdP1sYYDbkUrIjnQ5zqUy1dv
o/k7fsLBlvgh7XAJ3mJSZMW0wBWBvE3ua8S1vmssH8oiEtfwSiqj3vVMNbrRMZVxHSoVGHroia6F
L+MTIrQdiNxveYaGcmYd3rdhVl+iK+1DgOs7G0x5VTqUM1ST3GiGAlKIQduOI5S3q5B4MwcNLccG
YskkYNBExJg8t73nfQa1sm9h++NfISpvH3xRfDf7TNkxX4wtuydUAnZRs/khlZexg6jqzNtQ8zLG
Cuynlqh+GhCXil6lag0ZzfpPF6W8zSuIS0R9+2QlLEUoDx0PraMvaOVXSPMIRSTd/YP89Wu1dTtn
EIjDTlw/RYHjxzmD3imKOt6jDKGZ1DIq2cJU3R0ZGbuwTwlgeKgxESfniCvXXsjc+uFe4RkKlzPp
nk7+41LBA9bTAFyPw+ybpK3ql6E6lOCp29K7XI3l42QB2pjSa/zlGvCN1ZTP05Qpf8I7kaUQDmoj
73Gg/PNpFp8R4rnCeNreGanKsnnD0+i2zxC+uHSCWpiqSWpsn8gYes7p1FlTIupy19MbRAhQV48h
g9CnV4HZYwDc9Cty93f6V4w9IVy0/1N2Ycnymjw6yOgqpiTvn6TmobGSoE6EH+l2aj/APjBXa9/M
EDid6+zLPqGsKgt3a1Do/oKvPjq9Ty3tYlXlQO+/HUIQNaFizlc+GTedUQ23uR/kEExbHlKTqYWy
f4IChQsNxhxXna2dN88qTXMeBAShppaq0rZeYRvzRN5wv2EPP9+AjOr1hDZYutjWXtnTrrDC5DRW
xROrVsA3Yh5uTGTDnb2k3WVeiU7tjVxfAVg/MZjlP2TBuQKByI653snXWBJv/DlAgK19q6kF+ApF
6Xku1APEWK4cJAgFTfAqLtdSsGL7IIjtBjCZr07aeABfThkLd3bCYwLE1OmPhXdOKYeThbvi79ir
SScTKccTKrlSjXY9Ic8bFbaxrzlhXU5c6Nb4eHgr5o6xuTNMfnmWVxEQ+pfTNCCfYzDymoRRrbUQ
mbsBhNbXYfFLxg6ObjfckEcKNZHQOk1e4+AOwX2vFURNjs+SPPD+C74e0WFvNydwludWpC8VK4yG
qpa9frivc+2X3UH2yy7DzVhiTi9yyoOz1bK9OCevlc3KKSs1MbrzHZfnxb6oFuJlnd1mefz/tMxh
ENUkdAX8wn0D2f5ukg1vwVDbUPVRimAmXJxoDr1XTEcnICnCZjmre3SvmDsoaKBi6BZrg8xPorof
vcbhFngKSZyohZWmhk4lZPGvUkn6IVk/9PnPtB52B7tm31S0d+l4ZeTROA2F9FEan0czWWstU/Tf
09GVm8S7c0hnsSnZqvwrNgrK34roDEwrBCx3/mqkYDEvGVBEO637opsDn7mldJHV9zgS6a6qo6CE
7MqoCNc080yIdK5xFx1tz1oi8zfWdosoFgd2khmlD1zKWMyOormG/9DI22O5iraadEv2XItcTivB
oTq5dGuau+QXpS46NZEL9mY65a8P84Lwem/+XbOux3dAmXaAMqRIIn1gYH4U8WaRGU9bLViwjGvN
fihslQr0446Z6DCbx/2PHkZp0Nltdx0jmHyeVoNU/M5JOGBhmQ5Mr5sjmHuzXmTR4cWBw3EjJ/VO
OrOXGL49esAStKlVvRjU9d50M/o8tG4NYDDKzo+SmC490FSZ0ZA8O/2DybVbHDG9qp20787eW3qT
6Tnn7XEltQ9aFqGRNsY2c2lCLJiwVJ88UIKBpqO6Ha2Tq6LYvCwfV6pnqYDC4PJM2wj3G+dwfxAk
k31KOFx7Vsl4rZof5+XBLw6kc96iF5GbWYXMY+s7sxgHOj1StSMfAJOtzl9voNcbDwEhcGqA88F0
KrKFQ0FUhzEWUbfY5msVfBspLx1afzFfAotYZu84D/0CzSMFesMaT+ZY8CADC1GWQQhAFbO8WXuQ
UjXq5EJXTy0GYjziI/BZoCzyyzWi7v5NS57t39RXdULZ0S/tN5oClCltSHG4MMpiuJzQ/iCCgmVs
GbOJDWem9SOEZUw7HOgXMACNsoV960hAsUXcpPLMocZET8e+MpOQYSX3aZrIzO9Z07YTdVeQJoSB
Q8H5CeGpEaPVb+4rZO+QbhL5pttGa0vQHCwNNWGKp86WfyUuEju+1rlfwKC57//p1jUtwj3TGKGO
9tOl11Jw6mK/uB0W4kVp9efW6axLDOCFd7Ru4KOv7DSbs1zwXFT5Lv1zYokw6GriVrQWneeCOZkl
P5F4HKrZmxykwsqaWEqyRJ5I0vgG1n1VOEZJM3CzC0jgsaduQVqYrV0JdQ2PvMNDGZWYmCHWfeDT
ATZscasmL0/6LwOJ2ST9FBzDXlihBVplv1U67SlEPd7zqXq68OXGFoI3sovl9smsmqFh2nzGKM0F
ov5wpVSnKpouNK5UdhtSQPWE/IXEZRzVNaxvK8RkfOxfDrmmy+mXke0ytLwrfsbiIlu5FYfBQfjI
QGP6CDIaFVrVogW5sV5l8/KRw7OjD+R38IQ27fYyvbNtNeWL6wP89hqUt8Ub6ouL263/Jc/f4Zz1
LNtIRMmutuk6tuPfYXDgYYhNn192ELm6YPQuzUSuuVkFn/YUAEhLjpI24IV97312netZ4iBiRyx7
A9Nm2sXJLN03PTf343Kqyk0qvstSzDH/355KnNBEyYSNyhxxALL4a6XYFhWAYMPCgH/FjGhFSrTC
f/sngw6AJelXgnBXeuQQBy9rEm2feXKwOF+euwCFY3QEJsX25RPMwXYQJPQpRnTyxhm+DA4kt+Jn
8MZXWeBipbSlw1363FJaojyhsTrOTu7L5j8cJJNc5ZkHWZuBzlYmvN/fsj9AkjekoE1IZSMI2/Jf
Rk4jFbDDqyZpZCmlkkOl6LQzuzutgGBFSrEgHNksU5SMJsxML+VP0QrxUdicp7YVptZojOuVwZf7
nkDR5f1IC3yHaD0h9rSATh1Qni2+u1zPwWJkMSz9eXEfB+J9Z7JZmQ8rtb58Utqo2HNzuaWyavbH
KBXcb+oSX+VHt7bZXZW0mo+2p5erZXKvhaR0C35AqNZg5b6kKrU/uaL8+VI8Xd55gP7rTVgEMZI7
8aDDKyI2cx/Lv9aO2+CPms0l6zeAE3ahMLpXMxDUa2lk5sE2/kQzSH+CofrsgjoUUm+q7rXYQpb8
MBTVpONRyXHuR4dKBBNXRfoztcavJvdQhmVzWMRmyMng1tUKObhO5+wOhDqd8PRcWumpeEYaDpKG
jryQ9fhUQDFILP6lYDPVukNnQQr79iSXKPwqBEiPBpEfm0JPmhkoOBDOFlI/Za2cBRMKi5rIWUil
XFmw1EzESN1OHmRW/AfxoJ5lbpqWQBIYayndzQZJn6GXaW2THane2hJEZ3aEPe0YGPPIzWN3VGiF
m4JKVZl8Azyotz7ZBm0h0MhjEwndGN/khB8cDABQuiNfUkAsDzMXBcjHVnMaVRHJOubgi5XemOSm
U/JiGkUdcBwVghiEvWZLb1BtsvAOwXGit71r+ZV1JM/AlqvFiodKwd8dUc8TV0DUhP5Oib1XHkme
dQ5TvyvC3eprAqZd/s1jV0xoCo5CweRozKKz1T+KJjTZ6ZdK1e/6yHBRbavhIWWNf6hIUlV/KWIT
hlbLR5WpwpnL4vrtm74r3NzEBbpg2OxgFZ3qwwHtwb/SqQml1BSGp6J3HOOgOgarqYUWITjQCrRn
XqPAO5/nya5+z+9zjnnQpF/UbCe3WZEi13dytFdSDpbc8pbRYFqSoGNt8g/gUnooTP1/IihoZ7gf
EsLdIlSo6cOvVtcJpYf8EXrSfqLCyyFjNucdsU4kRpUWcf7h0v7hBOSm2eSJwFxXxQ4jp4V0bLSr
Hj2DuVkwkXkz2bvilBu8aBRgWGao2P93+p6fdOJsakOTgaupWkUpz6h9A51jiBYQs64OItb5w1gB
GRhav7DZ0mXF4soKIJC7TcrWRuv1Cl8nijd6r6j+wAFKFZVYzsdLTrTu2VTpX5FAq78BswO2MnWT
lsFkL4P2zzBaHK81OodcEwkdjdD1+ix3GgcOe7B4IS1fwLhqHWjHNWKp1/PiMRBNopICToysNw3x
2AmHqTa3MvIHr4eNX3mSsklyDqpV6RW6MlBhkGn/oKT3/ef+NfYQqYsyr6nmOhZ97PLRAxhh8eF2
45VGmI58ynQIVXQBAxkxuGWbV93pXGhc86V+jNvy6cPJoyprqljyizd797wa/Gqp8RHFZMtNB73w
aWG7NRvTSmLcXIbc+ocUilTQcZy6i780OHo1KvPaQnOAriAsgLdTYtvHyycr2hNcj4i+7MbqPr4S
HKy5N7GfQm6kAW/V5FRMF6Mre1ZmNpArvmoEUtA2ioRRzHVh/U5FTR4D3eDIBbdXb7X7RG7AuhTF
GZz/fSz5gDuDpr8tBpvSY5odg2Ywt5mj6s4smG2pAgNzwzZIcWqQDbZ/lGkHICqBJjL1Po/CLLIs
gNhxA5h0Bi6s11nuk17NSnk6ASy1SxId3ZdqWuF6rvVcY2DYGXeEAtzdKoGtRjoxVSsIz7lB4kf8
0SMbgwRYc34OznLQmjV9FRiR6iUEU2C9P4Wt5z/jeSenRKotOoHe/Q4tggWnyI7YW+c2R3Xfk8Ra
FhrnDzaSOSx827xXHCeWeunWHf9HTG8jD+XiyDtm0sCkX2x42LXz/VZcV8OtkGXDDLsgaR3FJjs+
0CIMTrOCrq81CFLBWBLXGAw9kOFE0Q+nRoHpzjZBdukmv7P9B6wzuJPnO+FpISyhhN4maLznYlvl
nH/e+h5+zrSFRQnjoGOAxKCLbM2YcsqZiNEWXWJ9Na9h8eIkWrbC+bfbvKGDZxND9OukezD//oFd
HBCN0yaioxV0R7CeaxoGtSghnsYmZGLACtZWDPKHdwyQ+UMiB8mC2exI83zQKPTij3Zh+0M6KIOG
oU3BWORkNsFA3odKGEC6jCNaMYXPK3Bo82G0M8rdkwmuCgmvGGY1/xt3QQmFfZhcVOnnt5SQm5pX
ZtbE5A6Iz5Y5srtIFar3cyd/kYD/3FimgcrVI+rLOr4fFUiCmqPqYo/1tLNpkZigmOVFCgKlfAs+
Ms6vjSzFp5rXyR1jd9wQLLh/gh3X8VfIxOuOExARwqtoIQ6ggr3KyFkF+gpf6FWiYoabtosivNED
Hy4MXTqeJSX3mF/4NQ4Krcjq98VImuL6atZkqdLdwFqMS0b2WfQYM5SPb9HuIpORqzwRnRbGN67G
EigHf81YdKKDtKMlCP52mw/yqTZ7mg0kjgC5/2i1NSiRKrXoRU6dYbaxuJW4n2jBcOlWn42Amigq
ugYqm3lzbmNC6okBTCHmbADl56No76Sq5JC5j/u3QSqCCe71sPgl9R24AkpEixXQ1h3I1nwhqog3
HYNXBrY9jfXZA0sK8YhpSOGaQKL1m08+2XI7NBuyRkJzfdht/L2/HS1MOb5flfoOsaQp2lHUgP5m
BHeKldU5sOekcz1DclKtz9a9oqldC9eqcnDvRJK+5GXK03yQb0NFjVoWRsGBOZ5xobimGDWKiWNa
FHs0vkyXbKVO/MaCbj5rc5iaUBQq9d+g7aHAdx7Sjignvy83GBff9ZyQTDJxF+GgxrOkubDsiWgO
6SVTtFJRMi4OpdwzDQST8Ak5bic4be5cmnMKIEsp7PwdhYLP3UuAS2KDifrKi//++GmrWX9/9A8V
GeSeNQYWCgNA4Ix4p/rl4h2yR/h3K2hCCA2j1/SYSkJAf1oMpz7CCItPQqdRKIv1tk8sb+xMkiV3
HsIFPC7tRJz6VeyD6Jn+knwXrIfgCvNNkuAHakpsDOGO+PZ17m6L4AXCipoShcabtzwckr6pgvMq
JsGXYbdV1vHR+usux+2grzOX/eYMP8cFYoxbvN7OdrVocxmK7/hoKt4uZ/tQfYwK4K7eCPgQWRax
aShJy8vfS4s6H8uk00MzykPsZccH6ghU8ceZLwP3GWY6HysaxO9KkE/Tx0jZnOT+QYbdeW4UcEED
7/DWPNpoeS0qrcBc0/2B0JKTvGBDQqzg62MrFk7M11+FlSZzX4aXGUL2CV5stwMF8MwpTfRkIgh5
bAH10igRy2MtewlqG9aR/fQ3Cj/rhIRTVQyAeE/pJjO11TKm/chxwNFqsz5phb0RNj7RIUlyvdlq
x0arNsaYF/llhveGz5P6+nE3V4IqVtXX1eTT9EjTRtQxUl70q2Ts/zowZhVYdFQls+gt3Vu7/5a1
TBwPZqFfEqH2OIgLZ36ae4cWIOB27rZL3lzSMV6EEDjx6AjMkpBDmuO7Cjq15vQORAbKnqCcaxZw
CLGON21m2PbZ5Fn+NBBhPssRiSglK7aqSCZh/J6Devt53kgSIl7S1eNsOL7ax38k4L63dp7u8Bol
fBDOV4pgrJ2qpKk4wQuQXgkdOZhG0bqmRG4qeEhjNptsVQV+S4BRWmnWmVx5vOwUDWU8qETOmdEs
MiRRKC1HPZlJC3he+NV4RDhPVXxAlWBU9RPvLJ6ct+BSO3kGQxLFU/ONRAYPF8G6ruHJ+abi89CS
Hs7Frp7fUSJzNGiKLWKXW+UKWNU5YSyf4QB3F3zi0hrmdpVCzZZhMfqaSNAtYca1ist692CVc9Zu
PY1gGfYIESnt9tIgJTmblUPp0rmk0W+v6t++iHH3W0dMiix5amiDTY7V9X22JmK8DO5nqul3Hqv3
ChLsFdRmMqpikBl4wap63I8yQYFBttlzMZyEwysp3XePXsZjYBgYJjj66rRL0WgGOAGlWcX85nVf
L9r/o5oRg7L6336BqA7o4JUkp56QOk/xy9wPan1qW9ZYMZzftZtDgEXJNHiWaf5UnDsNGq7Py0iv
m7Kx4P0R5QTij0oUs1jNoMbqwV62fouAaOuaXpkHEOpYOTnrtKFHBlm9yS+wCM/LSmpzudcL+lN6
VJ+D7IeC2UeLWu5ItBAAmvb8kpHr5mDWFlumu55khgLgac1PelZCDTl8N5GosKSeg0B7/VD5mFGC
D3xTyAvuXQjg0FdZ49i5i+sgmC6tIbmpbLFN2JuWELdWWyNCvtyXGs7jfhXpy4QQ71J6vLVl26VT
jzqCQS1MA7zmepTIyFgIj3hcNk3SIgD+zGjXSXhfJrM5kIo0uqki9ElDLTnKthaF+uaCvXE3jiba
2Hde2eOCgtZMbQ3R/A8f7fKJytbauPqClbp1k4Ullo1tdpCIutMFpGjFd+ZARu1rKuV14FeKYHZh
EE2+OGpeJWJswrceOmQ7ssid5fH2wUaNgm7uGHPhfQS4+ZKIT/TwtgFI2/qBsCEaa3Q+l7l4Rz3D
M2psemQu1OAbAVJi9Y7zp/GZHCp12cD0IUTitAMAWJJQCJ/bGS4MCa6yxsmzoLnFKzQmKcrtddsB
0vtGDc+wuhaOT3xT4pOOnq15g3MvvbsYEHALyhfxSnNiLBnZCmXbr669BWJlDNZbggVChIhQBfTg
fBcImcMKcEwfLHXSDFSL7ZaYYAtKa4r7Tzu/5+ZdrPqkPU1z/z/hk39ky05f6C+jFfhc3Pgqn8yX
xW3dA45H6trHLOsrA7cWu0zRtRMN3GJMu6e3TBjdRb75Vtw+6Wnaxl2PpI9RqrBZkaeJl6U3Ot7d
0j016CCSTC14+6V19ujIdbmPY/8OUBySGH9GOPQ75gVSHiBs8urDQQBgm+s+dBwRDvxpWjuwqlwj
kBOfdsF9GyBzzMd4N8CqyHhLfVV67zgeOLbUuWE44FZyvIl0gZb2oT055xhou05HDGLPBvFjHA92
6LvnqzLgMT2PKjRjIaENiIom6bslkdMwh40E1EXBu14rvt1ULtXcVkEsZwhGXkQrl09dWWFeKdwa
5b9r9Ow0THc04Qm7oTbCFpf9IUmbIfJ0F/YkKm4M876zFkxaMBgR+XYtK7OlpQ5TxjfzpPpPAtSe
Nft5XYZSNoD780+ksoWUR1Enwq5jdYS1Eq2jmXswK1gswaZtXEa0nFFEmnYv/UqS5U16IVAKYfl2
3BKmYMCC8wgabwHCYKlF9j5WhkSa1vRtORG/yq0IaZFW0hA6pJBFYCjTy0vHU38PVXBwtgtXJMVm
nYJrLCtSc3bI0t0Bt2qsxg0rxDUamyfgkSebIHCA6pkZZlM/M63Mqn1w/xVOtr3vcizgQceeCtn/
MRSGxYdoUi4iBOW8c92+Yf9jIuKTuw3tIO6QqDmjEtUAT9s3/xSv4FrHUE7aRxXghtFm/rIDriPz
662zW/uY3dIw9jdjr06x08VHANHwUqqh3bF8hsxdtkkkfRI23yuqdOk6biiGVJjfnaG1vCQRI+KL
aH4OBPLqW8XORWJHjO1krJucyfQSY4GfwEMHAuK2IU5dqBrf/Qr0suD4lpOSxgAlnyhHu7JXbn3P
7Pny3V5AZe6pLoIaX2FVEMUAyXqAR7+aWF90ekLNJsSoqLpUF7RBab41hNasV6Vpp6KAfLjY71H7
ScYDIy3Jff4Az1QbiJZOY+x4J7NOakO9oyFtXlDd7Ha6utr+8u4J/Ezxh1lcEWB4ouN1bXLr7E9Q
jx/sIlPCDz7/0H73Yg13ImtjFcSd4CQy2j9GNzwcK9tRmcqjv2RSln9d8rM0bIluK0EPlZJK+TIv
4vKA2N/jIeuk9plQk90S93cnVBWMe8Sv3T9oZYln+2jfmO+aHTQWz7nIWmi256vIsA3hTgnWb/wI
i5neVETBXgycb9OpHw06ewbFENHIozSMMUyZn4e9JIGvVcjqrYXjMI3atx7ukF2cHFCKfk+kb+OZ
cDx/eO2tJd8IKacRaj5GRoU2B4dv0ymR6qOOpD1FH/lvxuB2XbT9qDPUogoCuuU7K0E5SdtGEYWe
o+5UbIQBwDt6QfL32Z63aLIBZ6LlB79MbGpsaFhWeCF6m8LUGa2lirIZQdwZpXvuriKt40TIqzmL
l+1yzcHNmAIqvpEFBedHn4X2hqzqSYCshamypln2ABk9GBhANHkMZd1VSYig9pgWZ/wzZYu/3032
tk0GLt3BVZT680XFrC1a/QQ6woHytLjxCjsZQUlFVNzpsXh18wIMJctQEeJ56yLnBKHp1Qd2/HQe
b/rJxFPbftgMZD3U5tvZv/UjpsWXdaVFM4V5aiK5U8+fidOMSajAhTyfaJ2iVlgGbpdXSiXVzdL7
qyTz7pXYB8NGrANNdnJ4/luV5gXu13jTt82ABCn1yqhOjJFI3fU9PJeHS2qL0k1L04QlOtd3bFo0
MYncTT7GrwswhlBL57lv3Cnru5gImoXlroPVyCQUWgBOc7nnH5Xzu2G9ylI5zHuMvOmjojSmO1Pj
MRiWwdQD65xeZwF3roWu6QPLg5fW6NA8F4WUzJKM/1XX25JC0wEN/J0iBJ0cUZvyH2p/w3v/IA4V
1+o7Ydgs5cd9rqCSuMnlgxo/d3ZugiiyqLNHj5E92WH7//2gca7Ymjty8wekBtOR4dFhOf0leZ8y
m//Sm+ZrzRcG14OgB4/i/K598MM0SEsDgohn08WgYtXacRsDKGyiZN+ywcSI/PoPgAugvDe+7pO5
QI+6qE2HmC7brKR3+40tGCbuv13ru6zRKQCT8rmmgJQq1n1xmzLIevIo8jTcpiCAdX4OYqRmzBds
qamvhYMyKRW7McKLjnm6Rvl+5MlG/HNMkdtVaxKqNo8eVt+UBgL6YTz2/aW2CPk3X7LqDjfFGxlS
ulll8zokYeBP00s4jK5xh5/awE0bhNvs8rza0tRkWQ0AzhdsaWxLJbGzcsUPjz6CGGSGIKd9BmoI
/9PqGIo7Xnltkm8abH7n3FPNaBvtgGYECRBiw40fx4GPRZfOLt7kwVDdVMC9oupAfksFKRE9Fqzb
AfYZ3pnzpMx1gSUNtUKJ01gARUpJt0YMtShWvH4lnr2dGlJfSydSEZsvOAtQse6wRFaWfhaH2gG7
wPQR4g8uRWgCSh4qZ1L4NSMry5cS6Te4csjejW2zgAUIG2emhI8MWS8eRcHrvPq0Rm2iGgcEUe//
vJc9nrdTz5WrjX7nnl1uM/NOdVek5b+YJGw3b5H6XDc0qgirpwlmyBsVOofvL23cRZDdtcUSEMDh
tEskReHZZ0+CW4MS5n8f02xG4+UhVSqgMSaoEGqD+M6wufLijOdgUHiLcD0BC+aEKEgRbMKPn6zq
hNJcPfYFJWmpIZ3Gry1nisIqP0DsHxCo/stTZS1HOmoI9nOm6mB9vmNw1egul4boMGhIBrVtb1Ff
hfNdFZvSX41dmvj1IRazO4MEYYZaH4jdubEhBQxNNiNEvAI+o6AAAtZpV0rYZOfWzopTxqhZXCU/
0hVaRERbOJxR5Fd3iRyXPtecEIEOV7PYplixEPahJ76H4i15j1X9I8NZaJV0D0+nSf1i29aX33Qn
oidO31U5ViPZEzR3nNBHzyD0mEjU3o8n9b84VhjBtqa7Nu6hzrTKu0hONZTuD1QYb1N/dbK8Ajjd
JsOSctXrnm6MY4FUvgSY41FXBMojI/Fh7Vutc/WLrnKPwm8KYuPWp5K7m5CwfGVwhfB6XrAlAuHM
MKaiP/S4IEYn1fTyVcBIxmalEhburSsT7NAIbOAPTHM/JDG0WDmZsU2vsN3+KCwE8EtrsZKAuVA8
oSSK4eMJW3JLNRocz5A9mVs7FrVcxkMQsiMxKg2n3p1P4yox4mKG8H0OWWGVyB6qq35O0bUdhn82
s17SYYUem9GsUAKTFLD9AC5Ldi8Fm+vzM9hxNNANwQdLSfUae/bTlzHzSs83+a/t6rdiAf8pRfRc
SFy2O/e++F7rBpkE+NU9+E0bo/LUDjUjKXs1YZtQIMx74j0ooXfp1ds3/qP1DOtIAoXZmM5PTS83
pEHbT0nJfPaecZgmRs2l4tc5ygOkLYdtgYW9oihdv4OHg37shinFP35Q7J2dOegP1lHE9XL+ieKF
5CZu55tAfjKh4DPIYmyUG8UY7IYJJfjxsMAjknUzni71+yvhEQ0ZdY1yCp8q/UTNxPeR6wYx1sYT
x6AKRz6jlxkmYB4dZG1aLgk4VLCL4IvbkeHTsI3E6xoxw7WVaAN25Ob2J+3n4G37j2OCi5//Z6wZ
WoQdiDGgk6+szGyJXp2K7e9e86Z9p617/vizDrHG/Suw1EZRfcpgpliRgWSvU/WOC/q30/yTQTvV
A7VtKtE8T/829MzAR2Jm0Nu9FS8VPIy/lLwn9/T96p0jI6dlBrzNXGPmcvUilqs0F3bwCRWSHW36
2C4w6Nj3UE9djXCmqHlh/L/+9VIfQwBGKCkmwVGdLAkDOgQBRgk9VsX9q4SdfVJApewWSyKMRg1F
20W6P8OwvaKmOdyZX33MHr/U59Gh4n/hGXnCbPGFyAdT4Ju77oPNhVxecvEH6gSUwzrQNPxiBi5D
LoL++I6jFCzLYqsmosPRbi3XHFYI0VC5oQFU/JesbVruOwnoHl1DS9azHYjEo1mdmXygaCdb0Xfc
vZuN6kc4VDX1EoPcLt7x/FBH09a7hK0QZU61qaRhS4Q+Tzp51kidbuWtJ7nGkJHh3GhEimu3A9Ye
WNnvrl/twieuzes0hzImbeJgyZ/tVs7iM/T+aGi7oM2/9IuTHCtsv+I13kBJPMhNd/F8mllGmuc9
2MdMgrND5X5iZ3a0Au/4X/1A1VCqUxO5OsbWMObzsiA4ToAd5HHPU64Q44yM3NKdtkbt+8FU7bPs
CeJ5DGrhlZ4EEzJD9qZepaHRtF2Dez5HIqxd3chRqiKpJn6UFEowwbzsQMn+KrSguv4jLfgTPxQp
RXFHjkJdnBV53rQEuRwdD/r7SOmE+YM6cF178XrI0l5Vbbbn3aMKWQ4PJsAT7obkNJyhhAtOkjtV
VfWxHQjYp0pF9XNs1okFvINTK8MVeZqUIjQx05Rk4wnU99RwOjKwQNPd3L21yDN8x+k6CUyWSmaK
I87fncMjk++MjTEU2X00AzLdQ1Y/63MrozBt7GxSnBbHjxBSUqHdTZ32VW8sEaKsL+3EG0wfwMEa
yobFCSrcPQu+H3DIEB8esA3U1YhWVNr5XAcoPJAY8jN3s5RxqHbCEvPDbQli78d9+1icOWgnwbZl
lNOciFfUApArestPYxq4gL5FBzJoD8vQBgb4KXv5+7274KigOyO05ns9HRw8G1NmMck6FFQPlPdu
CBfImF7VwiRGhOXwbTFCzeSjil0kIm5KPijFi5qi4fjIqHrX5nGLlq+yl004Rgty76OH3WSisODq
3Thcre0bj/PybVDZlR651I1KPqZHFVEhk8X0QQ0vHklEp7TO93ZMKFF5brqLoa4gA3X/OwdbFFDo
eMeQSeHbx2eKog1oX5pUIvvlWBaRSxV4O+3jHGF1fq529ySwO361ZVTyR0tTY61wVN+8JIs3hsW0
3XB/WiEPloZYewAd2qhVaR6N56tZDr+LOJLsulQPRAvlDeJ5w033GOheiti8Ax/mzF2ktxOc7lWc
UrpGPe9z7WrR28/zN2J+OOYD0hmiHjKR8u3AdG5vazvF9iVupNvv95OM17KLf7+XKQjrf4eYfnL0
QHN0s+lD+X3mrNoQuKHDmLZRP01AsMZxVKlk2VUu+SEukK42q75P9tF2RofXSYu7cbbbi11c4fKj
cpztkXpohpcpnqStxMElMcrWZClv+VLrMtecZ/1h6jPbIw7SD6PrYI5nCzu7McDYaQmWYwK8KmWK
w6q5Q1bhcmUKPW52fFxBKtwdAUinxR7DQAcwFOK69vUVOiZh2A+dhEAL0MxpBGiTYHxoUrigUlp7
wz9SM1JToExGeKMRrPCxyrjkxzDJogYBXxHb/XWJdT6tHB0MPVLqqUV2bne2OvKOrlhRAd58oJBv
6BTWk7B0yiqxEYOzwHJoPw8BwI5oZ8/oR8gY5zfWFuTX7l3H5hfaD3jqrkoLfkViTxnm8DRJQRYQ
Tw8SzhlUHO773IsXLCPRTvoWUQqBslAq2+wuMiDgQtnYuMRWqb0a9n+V9H/OS/JIpqIMqUuWXlYr
ylLs1tkUsU4BHJXXTfXBSkU1N4Z3qFZrj9nBI1PGjnnsIi/eAAU1OMTrA97COWCKreRdWPNFemn1
30McXNWdE7ekUgrV6YuaUraLcDYqfcdceUUfN3TI8cl4FjzeZnItYs9Yow6lc513DAm4/g6bpUBc
fwda/UVTsCS30GrXuEscVfJcPulJ4X/jREUL//yd/69fxZBJdp0TmWHJTSKpiMw1nNoBFcTcR5VX
2Wb6IDa+z12llhDJyzl1rS+4IW03HGrZdRxtB4IfW8iw8hzhEiGSSR0aULxv4wT490xx4NWLPxYf
t5dIkLB2A7vTfVWKdbRRlRpQQ0OVAtUJN+h36mXLQU9KAev+ZjMJ0SVVepi/Yyd6qZVd/zv2Tn0K
A9VAw4CURCLeLBFloM51yjzf5cuCwSYWpSkIKdCg1hozSL/8uUHenKcEuLcqXHu3ns3dPt7UAKHw
CRqfEu/6Z8KDHZ9XW1SdpJ0nn92Nzr2YYTInfuz8r7utm+l2REtieuXh745YMBqOlWSNyMye9J5W
k6emZb+82wtHuap5yK/JdljdCJeOfb3qyM95DCSgReC3zTdRTVdCYHMMBlPi0+Fr5Y4ZEyGo6EAP
Q4LLcpMFKn/lDm46O2ps9tEDqIELCP9Uya5HAVEuSgv5vwxCQYsBwbx107iRgfBYL9Ck47SSsfqq
wMr9N9pFlOd72sWlpLIqx2AEnfHbqKnv/kjEWbROX76E3nDEZS+uysBIqbGDFMwSiZoBC+Qv+IbL
KoWFU0Ej6oorz3Kpsg5XJCh04zU7dbk41xLHZzbwACnMk2KeNFTkEEu8Rh3bn85tRs/uWMCL0G0f
XZjdjv3TOj3wviIPqlFpxoh8eJNL8dxFV2BSUci4WLKfl7akOwKxt+WR39xnDBTxPmwfk2ZGudvL
RaH+Q0jk9k/iiDnZ6DC9u92PjfgfzWxYNKEU1bKlE0lFKlTRrfeVOF56vkqtFj0ezEEAaTHv/Zap
//T01TutFx26VhZx9roLpixEwicXzeF83Xe6sMXW11np58kA7LyhTohBO2XwctyX4FEOaobJrbZC
tPMLO4ECUocyBfg4INvPRPlQpe9OOJS5M6n4nUPMkcu737CfpVg7IULhPNj9n5ho0WYFBQ/RlrN0
pOUnlVCIKDUM6uyfMyZrNGMPAUFEFJMmBzWoXuKFS3jHI8UZUrB5X6yVl5fOFE/2wxZk7KqHuYb/
uR7vf/LOIwqtNc6aSWTdHl5c9WTdSHPf+dmAFohx4Fvv//spNrG3kx/lUWS8+81H7qXfGOeyBHsK
IbpESQpJQ8VAnqvg/uw4ln8T5Q/9IPSiruOTb/hqhZotJmMojV73AKQyWvt1xOwHVCFlwuWOZS3k
TFj7ymtfVS+HwKypw/nmOXWqjjhW11afJ2NV68yi2DJqOg3kagr2+THN96J4ULmydv+oGC+1Rp1e
USnPrF2iFz2oVLgMnjqEQOR9bM1gmlkMJyWCDPQKTkQ60hk4K2UTVIisp3xXirYFvKOOU6mbnYen
GoaVrlDaUNDf8rFcToy3ug+PlrP4hUYnvQ03tIUcB+wHjQaqPEPtnqKEwwpf/up3BNDaUC/kCt8j
yHbelYz58sinmDhd6J/PjyZiPcPoea3vLYv6TBZn5IId7bFYfD6FZeELNSCcZM1kZxUxW3EPKvPw
OaVKudNA9vfiA3LTVDpreZVeRl1HUWVITEuU6VrgpETN1p0efO43k4a6f3pXreaR3iL4/k+L9KOi
Sh0snl5VhKPBE1iCQvoVEWEBbENdT4sQZ555lN1xCGWVsTaXqACptaj+FK0Jw2BZeIMy9kBxvPU9
meS+FvzJo4iC2x57AKI6FnsxlDeJw4K9K9HcKFDaDw8APKpXciRorkR6cocPWkpr0OwORDScTbhE
cZN4yqMRS1tbJwYWVLZaJLqs1rsLLkddPPESe9RQOzS8Rj0CpgjEo7sgqT9oViK7a/tIL5Lk+ngB
xme00j88/nwz0XIOOsh2EFMPXNocK2fFPCmlk6ugZmAG3REZlGNUQmGscg8+Gk3K5/EHJ86TUT3M
Zy2XvmsJHi5aWo/1L36cRDohTic524YOzyYf6IgYyXEQZX5qc351HAQYRCtoRYbIMxxwRbf0xLjq
jv+rNAeOMvIGQeJDkDD97AmiJr0dQowNTKhNjuzyD6ootqkeaRxuEgqSSFTbzxuRCViLRio+/eto
Hunkhy2sOqP/qo0yACrgKOrt9idDfjQOCyU1iqBQgGmVT9VBOzTwegOKdmYbCYtTxe7gzNeD78zX
Z5WPhIYFvvo6aSOHEs1hCZE50eRPQ8psvKZi1qyubdqz067PQpdHusY4unoZnaSh4MsVRz5/Sz77
peAUPGyzfETFLzwWFye8s2sE52DjLbkPynf110P0jxsVSqJpSIeUv9rKi53DMQbl0Civ6dY1PFgV
7sASTEJp/Mf8/kZLoy/IJTcUmuTmsOZCln21VvzZU/bUCGKNsIkyGtyDEAETlbfQ/EKE/zLC3C8Z
jY0mkGY1y9CndbR0zYAt77A8WlsWDKobLv+i/+p7+97BEHqyTuoLtlq74Qcd5AC+qCx+M9lDjsaY
K4/yjE0QEehJzzeUpbm0bX8QGeRbjTHUcziOwHoeKOYGVFvnIWRlZLJykQHVUvnIIuJQcIglb8LT
o+r0DjQFN3ms5rvIZZLRrttOV2XKbK661wk4d3XwznTQq7xxLCmvAYC76awQMUKmQsGCS4Q/WqJQ
BFS+YwT03siSoaqrDsc3DQiQ/wJ6PEhzEPYPXp/lqCMmNbyFTp1LGKCVMImk7clQtVQbb9ufwtkJ
XYupjmw+8ftLYkAY4pUgvP+VMdz8oN6LI5X4Ub1BQcSD66kYXBEuzJyYWtJDCxFc6iBg15byPYZ0
AtmOEv5u8irCVMQsY9CedVNNDTbV/5lzyLQ6CnaOeM7Hd5J5mS4qYebOumhN/kwnno+d8jrtsqw5
gi2Q52lCvAlEMGKGIDMJnbJ9RtlTjLoOO/mcFoY2iZC/eCf0aJcz9SPbHQKlVu16WjEacvLXb16/
qyBDbvtq03SgTTAGf2YKQbhqxBoLcroamaNTa6OI9IIbWb2iYdIttkAgDJFEmpGF874nFwC0Mqqh
UrgnAiecH9nP88UxFpCIx/E/7ULxouO9NMGZgx4f6Ed0ahbz3VluVPhmByWqUMnesUJIbkto9QX/
tLR3hWtp8M/7Z1PscEkf18/wKoJdR6GDjZEQh9jXRNRYF9WAjMOkXfDoD7fDeCShr2tHmMG9ZjAi
36/lNLuxjBGYEDAmjoN9/h/Zm36MtG4v6kSK+ESNE7viY2eHEnrZoEnTUp8D1Z5Xw9MTXGpBM2To
b0W9mMNu67zmH3RfYQOuMUTYxGrJPLixEwbrSa1ywdeKC18oGrgK6ERx8AqSJvGWQngYUmDQsOqM
W3i+8Rp7qRyOrynD7rIVS1J0L+nKOC28tZFJAsW4gz4bbZdGAV82w73vPAPjTnIFdmP5omqsgm5+
RjAFTBWu778DwYfwb8jJ4z5VtGvdAvf9k1zlF2ggnYc2jO+utgy6bdgFqapAfp4FBHjxWUOcrnaA
oHjnNVbSrsjgOtU0uazywXVNyuyxk+GAAZf6eeJgnKOc0hyiugOTV65rqTLqwBQwiFxBo9yIRn6T
P2aBEIAlJDaSgDoJb5NsrrdfHHaYkKrvN+ntFVUUYJO34Vq/SuhatvYN/LregU+esU+eANS/xfQa
kWqD7i/WnIU5crvEz/gPfER0FFWLtEVli67Ufiw8s+IQ8HCVw3enYTxXJZVH7t/uI8U3/jJOZINR
j+nXPu0gYZo8aE2VIz9G3G9g+1uAGJFP7OUyLCcbmx1A0BOa/9KQ1NHDC/TeXqINVrFbPYaMjiWk
6+GVUKcxQYk/CpaEwnWJMHZIsBEJesH/QbQCNAMtmCAzAIpIcnYNNbq41JmEMDyhKGyWCyd/vLIL
tBxgR8jPGnifRnueJqTMjLgIjkrFplDpMpnxB0EshDRb99wyMVcQr60gSqoLv6dpJ8fTVbrzq7z+
Vay4kJrlSejTwDIWiSDBzU/TDxe3d9vF06xKGPkiqJ+6E8DUrQsU2HoKikzyL5n3SDu7JloAvAoZ
9byZU+ubruMPH1s3TAjuyCu48UguYM+3TS5G9/14EIbRFP9TuG9F4Iv/rQoyExg9mtENiyR17+iJ
d7otCdC2cLZZMOkB5DBOSWHlnkKHHqtcLrm/GYgSBjWw8bmnODYnozSe9glQXvCHR9CvzGOs0k5S
Z4iZQ3tuVXuLc2BFpvRic1iIaIo7ZBLfXtIpInp+GUKbt0zxLWCS+mh9G9sBrBh5kACoxBY++fYY
SQ8K1vsVNm+RIsM4LvnvFO5ywCg35vOQgWqRKqw3Js/wr2t8Pd4lpZ4Dnh3uFS52kdsntoLp7hL4
l18YQ5AFxMSIhj7sJTn4dxWN5nSC8Y4VHEQHwMGWCj4VXBpOc1AJ7gkoV0NAeN8TUXZYq1k2xA5D
NlZ7n1FA0cJm9Ls40VFz2tH7C3zD9NugNfmBLFEzT2qyv6DfCbV4jMS8D9nesHwelTll0u6z4JNJ
XxJfEHb7ohCXKaZxrV93U8mBPDDzuDcnkZvvuWjwNLeGeBK6Wp6w0xlVAo4/ws5XI07xsg2tVNJi
Y2iY8WLc8WZnqLHL8LH/7XN6W47WrtshtDD/kXD0YvAb1MfiK88jB0P1uiMvKM4ILdTdibCyoSSN
GNcYbH92KQ24aZV+/q5bPK8bNj2//KQJLgacrzVN8dfq+bKMDQi2rJa7dU2ISvP31vQJEXloQx7y
qxeOc3HD3A0hvWlQjmjivOaYq95GZmxW4q15Woc1KtPYZ+QTvx9qmbT1SWZCb7jFKCngAi2cHPov
to8bBPBx3DhwwsyQKXWKxeceM0sIH/q7HSlXK6JbA9gCzo5LeVwPTiINrBs8Ay6+LDlaMu44Jjki
ZiVBterRcJ66ferrf8oIggPACf/5Z4risv5LwrhaatkYE+Hp13wd5oAqG86oFSJcveQmzWa+vvdo
u87aYC0CNK/yptsawML+62rtOquV48dUqTQhjGnZy8j58LYzersjT+XIYNPwQ+yvC+aYSdDb5Qbw
wml4jLrR8XJ33Jywv3DMzZsZkpjZ2Gj8PbppGzhqJ2QqhSoLNn8zsmgWQThpANPWcLt/Clz7qrCn
y3abUAwO+aUyMGixP9rdt5lC4G0RkQzSKleX8bNWE6GmSQwxbrXrWBlhAt+TRfoEJ/5x8BBGkJ8h
4py8soWZWSLB1DaDmVi1kjj7L+kE0HS1jc4bsEwnMd7TY7m5uK/KjPE/MZNK/0ZaC8HVVomWuF8c
demWHuvkU80bPm4mZptBqyZkKGzOh/ITysv7GzAkLxFDrUvkU+GvatV+01H7jCPAZbcvZUD2S462
d4is8U7SBf2sE1cXQcVEklY+EZf675SpL2yS0I4nRE6bdpYIbjrh3zIcdJHmPdt8Hb+kMj40oaq7
TMU4fAlX1F5KE9rkeZNPAObLszK0agNFPD21lHLrlbxxJlIj+ANfGpeoj91B2dkIpdHFexRBW1u/
HwHybCSVEbukmd6UyP/cMPk91NmiANHYKFI7BBpoLbpQ9dD74ZEGay37y1hXU2yC1vWSpJtU4s4F
E2rjnkpnG/rDV2z0+04UQSNmUaXG0qS3EiGrc2DvamGekS/A8i8aT55AjP2WbNXW2psimGwGj6PW
2bVFj+RDaaQlwWVkHeYIxq3hNlvoGZ1nw34cF+oZCfATxeARsMnz7MtvR8LDsrfl7MfXIWxxtNaq
tHVKWt555xKIw+YoV5QJX4cAODTH5mMkAew9zl8fIGqI0cVdr8jetzB2GI4oEW8/HJCzkSFb/Yus
i6EsqmYBR7U0BAq/13E9RZXt08wtbjwtuocCf3Qt9kzLwQ7Up5XwkJO57qS8XMPXAjdLp8Fr8D9i
6x0tH1dJhxEHWQtDMKNZPm545Yp6/tdeaRsBR3b9LzZMCmR6rR+63bnrG7dAv+VfHUs1i3mJLIqh
IN/a1x60vMuJMO+YPLxJRjZq/Rm/idqQWrPrHaeh7Q84dkQqRZE51+b3ehDjyot5MA/XD3IsFVWA
yXP2LcNnaNxw1lUfFH5wV2GcL+/7/gkv98UgCAKRZwatEYiAns1P9lB6XwFcqvBXGmR9gc4KRvan
OYtpnKLz1Vi+jg5s00U719xOQwKPF5ROvtkZnT2CYHL0KoI66HkIZi3xQt9rIWIIBsoYuSRJbBre
XKg+2pDHwL380TzBgNoBxx04xnLXVwuUkOZuxtr2jjAOOGi9D+5vr0W1p8EiybMzJnXoWh9g5yS/
CHuzcCJZ3Hf8XzTYLye6t/4H5pFMsACpv4GcfErlrqJ10J6D4Lt9oiwoy42fR1fcmQJZw50Y5oFI
DAJFRyuDRevGoc0XBOP7rb6R1+l186KWgm7x494AcgbQx2lY9I2xjGv92SN6hj1RKXYVgaM8HFFu
wfI/giUvq6iBIEVGFYM+QnZi8gMfwSEetcxU92XBD5rJaErF44iSbOkMP0VImdb7qRjS2TAV3uYl
Y7n/z+LMTG/7PS2mVFwF1g4QBwvgt68gBrHdT0vGOsred46lfN50SLlsJ70r078YLPSFTWrwxh9N
vGgobGw2FcUU003DDvyXOKnNpypo4ZAetPisPfnQ22lmw9oYnXSbS/Jn6i97/aW3ZVxD9PprTK6P
K5nAQ6ZUVQlmhmUY6vF4TcMW4yirXSVuUna6oNa7hbIVmXvM3JIgwNLYxJv4nsnQbYa+8eBq8CI0
YZLnVW/zVgLSloIy9AhhtV9mxHT743+3xSH+BIBZpgCMsS/ijzUDquyymqlIa8jOyeeTbHT48AU7
8CfJ1wXPP9yqkgy5peQMDJuBUwS+afLCKoAqriPDn3QR9bMDFRy6qgYhoqDYvE9SK5LW1CqB7xQd
Vx+I9P3lQqRAprFZo2Ae4mVkWp8TSdp1mWV0Rs+fAEwgG36i2oJsE0YWhoUUmeJQFM6JPfGSSytc
hfb6iZAu7won25ufLvZqeZhj2y4hiD9csBxrnN/yf5C2Vb7RwVhEOv7JMB8vn6ERL5aUl9D/4JaK
cbQLQzeJQW/FUnOVGpiKKyhWSJ9j4ndARSDLGXgyuJvp3WRKhDwvoq9hpMVxn9gHYhRUO0ZkSpC/
VRJu2WpaqNKW30uCDgOV6+YeWyeE0Pky4ZNQth7f6J96x14F8X/Pv9M/4/W8F6YgiKTr2edSU7fd
/N+xK1WMdve3NZVbMhG6D3/9EaeYCoGOe4+0mSUdJRINkcmgHgECvj2bb2x1zIFOzHjQx6226JEh
5wZPFT5pM9No/gKxZEcthj/6pcvflqp4uFVvhZTj7Y1AP7K82WLhA6TckCZhvGi71zUeWTHQWH9Q
QdVGDsKni5RuIsWZarWW894xnbIqjD/tEF2Z2kO/gKPsvqoTv4ftl93ZMYGJAGVIotgWhp8Ov4cH
IQgwYDkyq7Yit+jj9fmK7QnFTxrP10DLbd3ew5Z9iX8523FjfY/v1ZaRUEOmP0ad6ymo8JI86gRM
+xiTX0gltdslJ/qHjsrm0RGW7jiabuWO/71BWp/sWKoMYWRI1IiojyhV4eHCi8jTlR6LJ4CQHakp
9LBVJUVvj9RlkB11DYv8ezS4bTUTo4BoaSGQS382x41hMDmtq+qB1/lG15J7rTu9M/eSWslOh9h+
bT3XFw0eUF5g/+CWAScD+3B/MXLEmNJ1zAri1F85zpOOTs+SdLYorkOmO9SXWVOWFFoW3DEDaS3c
5L0x66SjmtFUkygXjdJ/041cnm64itUl67i6IDBKo5SOXpn1EWYrgImaBnCW6UlNWrvl0BxoMbSs
V/fk4NNimBoOzlPRhSW3QUEEH1Wm323bAM86FDCoQrkkz4gSVieAyB9VbAt6z7pNSyW2Y4rCaJ6P
2NOz6BunXeA4IfIL+V0wjInSIZJh5acrZ81hC6+l0iZFYC5SYc3UEYSwHZOlSN8dpNEVAmZgTQex
u8IC4ehhdUNhj1HxevJq/fviiwCqmtYIEmDguTTsIBXJGtSKdFJFLKD97Nvpim1pb9BG1xHKzPNH
6PmecTwQ16S64FWLV7fGdR3FcrO4EE/PedN27tIJfO2nwuIaqwJ5uaExx7oMsZTIQ3Cu2KMgLnds
N2qQg4YYcyF2T6x6Bs1Qkoan74dbPiyte305AWuZQE1YcHxV8sRxPw25sNEERVTs279lT7SivFLi
GIccKLOm+2yQ5IRYd073xyYGrUrfFNN2HUrVGUaSQU+7KUA6z069UV8/i5ozkgHIa8am9D8BQZqD
olTH5979e60/24us8ZBLB6KLq+n6Y2F6MRiyqVwJqR+xRx7nMs8D89zCdOUjLhsxxM3JkARcAn2K
PQHi9CWc36izHrkm9YfqSmbTlQEEJBG34Cz9HOaU+TyR08GRZZ+uDXAJUkV8JhoZZKakgsKnasmZ
OMTWoYQ5SjCt8xy6Dso1OEJlqJy7xodTgRjmsW4ed8ltqB2O6+cDx0v3QlL7HNm55MMybn7o5OU9
63A42gpyh+d0rDIR6NojSnefiZ2vaTsQAWN3l8NAnaUzxCM4Re0VqCug2Nk7M2TLqo4lpygJY5OH
qFEaGWKOVzY/ZOIjWTFlpcoKuslOUaaoOKWY3YCsav8lXhJY3QtkujdPMk4vSx+dLnmdhf/xJUl5
pdnk7dveDOeOLd4rX567qn5FWxoBuZxbCwORElq9m/3P6ZtM1SPHycUVNgU81auxr3C+hhG+fQ5x
zIjaOFFkvCcnq1qwLaECcbN35mZcSRdrNP7vpouBcyE0zazKq0SSKNAwWLQPmwNgzq8hM2E9gGjD
dlVESpX/69mR/k94Q9psesxfuuaxa+Ci11tanp5YyfVWwXPFh2/+IeGtYa6Yn/iRR0r8qL1FIOqv
58/sJ01HGmcae+BjIH5eoBLN4m+4Q3REaT/Xyys6FMwsX33QlzWupIKgVyMgH7LzTclzNbqSyDBU
mwsLHCTvqX2PkIuciMsRcw30FVBjv0zWTGETqhuBh/pfz0AnLMCMPUQzdPFep0LDZRlzmY2cilLF
cuTmv0OILVwFgA//SpBL7RjQM2uOPT7su0k8aEVsm1oMJKqv9HuEBfPgdY5Pa60HlOCmwS75BYfJ
eV2tNK9W0hpA/fRl4+DMaLY0q4+vC/b3srrCHjYbPklldav3pg51fUUCSXNOf4QM6PI1EY9MPJsx
pLfhJB1bVwEPSn7sI9+pzMm2Ulfq+N2oPVpD5927FJ2sYxJwDtvmhj+caW7eeNuRo3bIsN/rwqbD
UYSNiOIykqj8oQrzvF1+nwI/3iZvA3SH5htziuAGHPoADr+EWeSQTw/befz4WUaus23iIY+0RVtq
7s2wNboz0xLht7t6q4+S9ydNBi/KuWXekXNEInPyfZX1K9z6Rjl1zRJURHb2+A7eiDz6ZYP+41Yt
LTNa/z3UrgW9VcEGXMsj3KH/NMh3IexpL74nYiLRF64jLWVq6h/5IC4lHociQtaA3jhXWTEV5a1Z
AWdJGvBizIPx0Qo4V71NbYQDbzLWsCzUwJDyVwa2W5lGin0EsYjuhv7qmjW/mZ7EgI4Iaz/WYLoo
pHt694BA5b1Cwb/egG4ucCE8jboDcCxqbb/ymEYX2+J359uVAsbQHyrHvE1zVX8LGLH4udVtH6Xy
FMjmxCi1rgzNSE409D1hVdmu3IxHM1O9jTxzCqtZFLsm38ppPkDVXefl4SnnpCUydPzOV/4zd/B3
q+pQkp7bw7BRUgsSkDDGSi5heRn7q7fd+TgGrHJnuvM0A2wrUMwUdDmOc3VPVWgsPQ1KqMw6ML9T
pnFDsh7NLej0mnnpI0WsyrKyFxPv9/5dpYrlJU491GzeaUk1vap9xpgYD97xjo++Slrv/jSAW2/q
KvCddp7C/Voe3AlX6w8Pgglv0D6ZdfCcmSCM6LirXHE6afUhOAp0a2Hwnl1rg6goisuGUlsjCYDz
+4dKeUmeVs5YMS2SpCTdzG0D8it2m1bmw32IefEJW9EjCctCY23V1Z49lfvDC7iWVbOfuPp25/Tp
5Ic/qTzjcf3/GyBiDi1E/QQt+c39IHesan6sd32GAyosnNh+T3oXnrOvC378rJ9muxxl/atLJtRZ
/REk0GwU7x/cvko9vqViPsNFJbnJiXBcAVgQbIarude1+u/OPCbYMGNjoSc3fRe/0p5bti8+67sa
1NzYZid0lyPisNPWM603MzB6ggN+EcgsUC4ha0E5GkQVkG8V4bDXaEtMW1JEGn7WchysgeGoHn+L
tKnHUg2AcPxIBDpTQnp8Po0BIfFbxLo/PKSpva4Ribf0KCHhhvJGwEb4HWvykxEb33q0xzIyZMSc
vMDWGPj1OVTrV7QtvJawIS0AtJ6XACZup04q0jB3IjFvvjQldX/pY1chkdVD0W/qV+UEkDrMHRyh
JWmX5m3iH+oaU2Lbbms3srYpy2F9LNfCI5+Knrg6U/EUylmIcFK9o05IeCXt6iDfiWcnZ7PW5ihr
8KPHTocl9jhhIp0t22FMkYr5MkQFpVFPLzijlMmKMWQcNBFVSAYLrFXk+QGjhb3qlTfXudbk5wjG
sGK5D1uTQQXEJKdZwqq5nxkdwJmtAowic0uziqql5INYxF/DwmGRW8aGttwndeXkHaHAJwfscp+F
vkfQDfdow3FXaDw5Nt05q/DkPGYEkcZmoP5w6Gxo6PajbzV7T2olS3PgF++tNLSwwvsr03DcUkzV
yr0Gt+e+duHc4D+FMU196ZRfHN4W9BAuzrYyKlAX8T/w7E+63KxEshn+rdkbO5jHQCcBe2bPj/XL
gL2oLd7gVcH6qoPe8mj5SfgdqxeKzzdhkjI2G6b5FkgiC63yzm6StLItSSbRDJ0zf/zK6gk3/mpw
O825ZVSANeSQou11G0srJoTaOMrZoofzkUQJUxZknB+p2N+0wVoPkHUvAGUdplPPYc7S1CJF1gcn
vVe0Wc1676y4EMrHguj4HFtG916cndCe+d20HP07fw9OkNSakRMJ7LrvkChSOmnJUfG5o+ouN91k
W7F3cj927/shkiJ8KSd4IQh1T6qSxsRskeXPB+Cd21T8LDsOTp3dYaeUdKY/iigwh9VfAofQ9nyQ
dE+nzI9jxhngqlWDx/+gb0/1GR/m0R5yjmTKn/C+Mo3WhAH09u+aMaUySMfoCQp1cj2gMJ1LzLDb
a5Jir7pLwzFvnPai4bEh0xVzfHv2UwlnRJFzhqneE9oVkQHpWs7oouprC9YabXhAkij7c9aV1C5q
5mhaNrZvn0DAciINXv1rAeyslucEl5aTtCyYiOaudiYn3/lqNwiADc7mIN8p+qDJ1tN3Hz40BQ1r
hRfOQf/mso6XZf/xMPDP11Vtzfc4wxIPe/WZ8XNr++grQO+zy2b4C4Lh7jRO3HRItuE0yVsiQGMB
y0nfCvsLcvAwjfxk7PzNXW/K+tQKbvY1OQiHnonrswUWWZ72WZNJlC4ligpXn0GHqxxecw17SoDJ
Oi52fRHi0IEQx3kGYXxfEioOSK7DbC1LZ6efKk1JShSTJM+OpzCfC5P0bImiE7d79VKJLt6NJbeF
mZLQyKi76RKOsdJttJnecCWcsMQALJfJk/2CJA1CsIcWqEWV+tyKoicGgvkZNgIBLrmwwem2xrMv
YqzpIGI19m0oPt75/UPne1RDBPghiaNY4diAON0wbFQQ1NzzucVwsuJ7jgUUMty6aeeUUbfy8Rug
HvDPWK79S/QgeTe3ae1GcOXbpdzFvpnr0dK7ci3CVo0PzxoxE1DnzvNTZxaE4yy58Pal9Nq8II8A
Yb2qLHrt+divmkUpwHyyT6B/DfGFKLYk0nDrRLJcxiu9SC3dF3yHiQufyvkekrFLfQUEsH65eodX
/V9leMyFpCASGrMP3VovmIpi9gHd1mqJfzbi2bCw/eQ0zHi8IdiouQjPTzB6oqk/YsLIqMHwc00f
WIoWGP1hb563GOraHJKSu3+E/Y55ko1mhiJMrATGn92cMIbWmrKitG5n8Xn+9bII+SzOrwzWmN5p
xxo3m3uWqBWD3tbRJYMXFCqzMV0sCM5lueM23UINyNqJ5k6TZ7wfIbg0Kpm3SSuw0ruyyNxGF2fU
95CaDozjmSyAoMvbak5sgPBhRyGUqtruKF5nxkIqoF8bQ3tSF/iQ/Y6GOlcjmXjnvrv3B09nf8/E
KQIAS5EkCM41+ZL49iQcWV1pGLRwvDTvyMdxdGMkJtwmCkig4ka9vfWgHTpDWbWU0UUvfFjJbEi3
8vk+reK2yNUabM3uezsizCckE2QYlgsM7AIX43UDBbjMPey0h/AQ9RY6gZ4CPhlFWBsQY8k6i5Pe
WcRCpAWqKB/VMowcqFnc6D5mc/YnCSmpdmTiwpVSa6xbSv2CEwZzHvzMd/hf+quVcL3r5lJNtt7F
B8YanFN5n3qzr5SaGoX4QUP1xc/Ao5myy7UtF5fzmWXB5+oLN0zUS7s72hsJ+8mioq2yieX3X2kd
d8LLBFlh55gcf8ckxGOk+jNn5kJwYEo4xA/PmZHxwQJ1nN3Pk6Ohorqjv/9YVSRZMXrUgWTDeph1
AnxZYrTfuUQZ9B2oofYju6536tnL8ftyTPb3uQMllqF4ZRfbMsKVA0Kz+zQhG0s2NkVj4Ed6DYsI
SX9qs3mESt3/ison3Sz7Xha821Q0t7w+ImuaPMj39k3LZJD7RginnfuuFs8RGl0gbp3TMb/fc0nc
sMAXmHqcFOJKrTknMZOL4I7fnldewzVeC/h7HL88uAKe/9i8eoiwLP1TNYKzg/oNuYnvCa/mZNYH
aV9+TounwFzI90YjsQiyj+FUVOY/hKxssaLlr06QlJrD3xEy2mZBitedpQL8rENn8+E4xmodneKg
3gM4RBfS/VMnhOaTp0RshsUB1ofREv3/iv7YEmIDqBR7d6yckaVDFjzSrKm0lnMBeM3IvHxRQa9m
qPA3tnytf/P5V0Dy0KWpjVQGcpfOU5dEfIcYotNTtLFJ0eRcWk6uZkXWjhxx5VW00Phvrn23lZCu
JlELEwVB6pla/cO1yFjlaJmv1hewqiWsAzNi5VKPo3xpnd0jPkzZCAm44XQM85E4n4XUB2BTOfwP
u3krBub3zfohmuviMsrmwZ2RhvIYcNe3MuCxpTaSGqnERfNTq3iX+/TFlvHKPCZB/y+qxPaRnJzI
McSVbqEB5K2nwvNNl8Hu+XWi7vl9S/HSyHqagQ8xC5A0MdgtjKCzqfzKr8pWOhP/+uJwK/+DiqMO
O3VDxeu4JvDRQl8zP9uPCjJx7ZcGBpWkU8BgwzHVgCE7J9sTP9klK5/6W62vZb5fqSVFEpFRhdW+
sbtOOynk41XqOUaXACBycCShTHxa9ZDndtZuovykzJQDgrDgzFrKHslDm3MzIkTx5P1gn/jmh9Qj
vHQ9vUoAv07eKdPaiPB8ynuco4fraAgaLVOyueCp6p+bcNL/caVELn5sDxp096oLABuGbXdsQZ4R
euighmFcouBFbE8pqXzVQh7jMkobiTxvmw++q/63PWxcwZLeT3OCtlCRsbPxW9KgLsVy2L7hAT6x
PVJUc8m82kkLItMpGNkcz39gRImGrYbxJRfOA5CLSyjZvjUejwSVAxTpAGz+Zw6bAHRuC7eNsOFO
7C4OoBW9eFxfsYbfwv2/tlxNqWjhZb94t1lIrVEffgFoI0M7MZmUnuFl/erfWbzvVywe2+lq9lm5
78zivdj6VN9ovZtHh7y4pCq2sJUEUvTuhEOc5JbsAZOsN42Y91L/DDY9H+lZCB8WK9ySZi2eO4Vx
ykJwkr1v83g9MgnuRvnZixdihiPoxx/ucCeVH8zl6uzpNeImJMUZnbiRHpcbsd77iNTh6d5CbAS2
Ke49ZAQrfKQzGxiwQM0VLoHqO054MUTXd3KyNUVimnenGjMto15SqgX+dpiu+TDYMqn9x7ib1zko
vZBs4eZnUgKCnMCVze58IYhVv9an1J7kg9qOT7QzKdZRSfBGKj3nOZzZPOplo5sOcLtpVfTbNmfJ
pfIhz1SOyknHNmnVTSj8rNpchC/foh30q454YfqJdLVUXtT7azgqUpiz8slliZ61ksJehW6ACA8k
arczyfm9il386opo58ijRwE7gKKrLHk87vGbNznQIwqxr9Z5GddqTbFFcfFosRAhrcOTs14otA8Z
ldrfn8AEJsF58g95XoVtBf+NcNehp9z36ya8sX9hmsFq90fsahXFmk3vrMYDwGhJe5rHUoUL2TSf
MpzdE1inWXC9ZNF3ZnRgwUVbtPkLPyAziJM9aGVK0lrJCHeYCwixvj1AHZGsIMIUIye4kuMNgN6D
PaAwpkKKy2TZnG0z2HZmlv8aeT1N3bUadjB87BtkWas26pQIqb0FyAxhLuWwxGeggsdyC9bdG6tO
ZPZo7SEWzNw80x549G5axQy103EEX6r8Oz21lvDaumPBgT1qXt6dKhv7MBnNixy+6HBbGV0egas5
6jOWw0DNovxd1kLQKbn2c2YzpHoPcgEJQcj4moLb1CUAoMq2gFoKi4KinKtcEc10IEyJlUk3OJ0t
w28PkSfih9t9LvCNfJ0CfX5fmXi7vYZFrGosDDPvaDfoikV1YFBBIWJeJzgUB55EftJtz54qtAPB
USJIgbH2ckkOeYr+FlsULRmwG9BXJbQtCA/sezvdD1QtZ0AQAOu5zxhw4g7Sv56bOxK/TUIPcFb+
YhgODNBtp4TJ6wyis47xGDYsY45hrr0X9ROL3xz083HAJzdQkIiJydmSnl5omeP0RqLCE49e1E3Q
TO1g0JGEWjEx5eRKlZaA9DW5XNhtfoptuJaASuQlpq9sLmqRO2PIzHzO5FfscMniAO20OQvS/Xz/
4BR3zMZmYwGLPQZ7g2PYt6o2Jk9xRoYvupGwGJ4ILMZHYMgQNV+QNgiWQXevQgIqmWSCjM9QLwD6
9AJhWbq7ZrFz+Xi3eTZ/BGZpXhiJztehvouU52dcP71drA0Bm7fgKw33jFR9JpqwgxZpHLkkY54o
H7ncO6litD3nI2ClyEdnNdYl/G1SI7R61OyWjrey7md/F6fjEJKDUsIbOUIaglJQQGZfPDyIqYtk
acR2Wf8kBUTFUhauxtvJ8I8SxU+Olgi54Jl8s6xjnjORcoU1P9D5Jwg9fXhXljLMIXzmqyZtiMfh
K34MA5cACWIzL0h+vzr9GNmJLJYjNuIStg8d/yj0gMlvTZA/m5RNs4ObPIlpqSYwumQpsmB7Z6Jb
nVcdUdu5tdTb0V4zqXWvSFOKVheo9aZvbM7jiDVjXCXjJSHD8X0Lgp1QejrY8abm0AUG9b6rFwc8
JhNntQyYK7uQy2L00dAfkEBci06pZItjqSa2fnsus7mKMoEUbzn624efSRmihJfoMpjbDmkAWJ0F
SdZbnAn3Q0i9CJ2U190WX4EkFuGahk6h0iT/zyVML8Q/5h9+6EywvkJOIN8lQ/vybSO3Lf/CVYi6
OtKS42ja7LJoH17OZULsp1ULG7EGa/V/WSL2ltkTpYjGd+IMjI73vMMT24sT+SBI5S1suNpudJuS
jLLNI+zA4UdSp9Klnk/m7Nh6koRxSp/IpQMQhpO5oXH2G8Dvx8tjuMNl8oNDKoyNvCD/AyMDeM5N
3Jl65gqBJRVjhyQo4UXQNQe9Ic+OWfZD40YGEmVSEo2AJoKqLqGwnqEQsDI0+kyeADPBJPOwYMcR
S3T1gfUUzay1UN7WaJnf8KFJZEApqMy9uYmmN2Cgjx9i39p+JpzTl1Uwo2S98PChcxvlcTnXRO5O
dnndbunkWv/jrGzKjURvdbtLLz45pkQSAeHyTgRtXG3AxK98Ih1dBqP1OZZgiM/deJyWiH2scHaz
AAUxtS0W5/ox2HbgFA07U++em6GgU+/VrZLuBEsOLtlK4ow3GTYrFWmXSMeWyrlH5i0hiRfiyLmR
Dm3Y5BFyTRBf9BBR/PzgQDpUTKH1J7tUV+02Htp1aKAThnkCjZn4rKlOIRh7tBoQUTtp51WPOsEj
ad3hsgri9SI8AWSaYnAA6w15AJnaHrWtyKQ/VxcWc5EldbpwLXbqS+wBF6RlKseRwTx/RK8CCbG4
Jp11jzAXhbZ39+uUy2jMsDmUPgvSGtY4KBS/7bmCsmt7YcvGElDXocCruN5lE73XNxySQTpdb69G
wLuIGuuRjOHpC8l+RxBWRUyb4g0SozbaaWi294g+Kc08SQqIGwHmmgXmjYPbsC5JsAvljF7LjVxb
M0mqAzAstcUQCd5H5Q+FU4hfhDlVPA9WTs7r3eiZa7aSfuCerkzhioHzezNKUV7d7TaIvl6bqo7o
rKPY8R77rrAeOf49LQHw0QSfm9einlAbZaIuPgIyv1DI3lgEzkU3yQg8OEbUukCCl4rifVzDpzcT
OTO0m2XWDTxrwpozhxGb2oUV4lTH4DYtB1JtbtGIWL6i3qgWOiaKjWewplFhzFucqj9hgLL1hqet
cP2JO2kBvDSCD7OsDQxMamLka5EwKsnqIsAK2H0nc6BviNomDAeLHR40WIxcZ1u20vv0LtkGWib4
30ywR6liCKBipt862oqOsQlwZ5P5I5afVFGrmhdNv4vUquaYDlPDj375ZC9Oji46wt1cpmja0aCI
WJ0cSjVQW/Ko+6dxOOmo/a0u6Ajjqn0r1IKPZNfo3XVVPL0vHKUPl124tSbj+X00809gtj4VSgmc
CYWj9sl0B4nra4/VlMppG9fnq4ykz+EfZE8TWG6tnjaae/hne60uHmOXTjwIBjgoLKV7P+jb9MmF
0GPw2DxXHx6IGyx7JOWl5XpxoDS6f1KAbIJfDvXen8741bW1p9zPmHyakBWFOKqvKmlkJXyKAk8L
li/SFw79IUSXxHCbRgPcYBZlJdyZj2Uu3Sfu5J5NYQmAkLgU2JAnM8WAN+wYzmdtnjqK8potrTmF
/Lv0GF6OWDH979eS/KmoV4QtRSm2P+4NlaqEhYyUQFrB9/bxVGw8/zjFTYeIieZ8wUrNJlzDbh+6
4JPw/lA/YCDC5cu75F10sFSrNSmEEi3C35A4iKnjIWdIWRUbFrTSGAEsUOHJvkJBNhpcF1PGCoyz
2lRvsu4CLknioPfjpGqHjE5e9Ukasj6Q7IBrG7M3LRenLYYMwX7gzlfYPvwEFTGdy5jDJnCV9HnR
t4CilujolQYAqwfHxfkvLT6GEjB4pO3uNV/fnhJ5zF9Ae+6i3CyFPzK1Pkdxknw045nLcFxM82vb
Vi4Cudrh4K/FGCH6oZM4LGo25LWvAwwHCFsLRWtYrHc2cP1s46wGFXlUvkN/quEoolTR94099E6q
vdkeNrz+M+8NusHmOjIpvQ7Q4JxEPumv4xT6Yq0h+6qZWhJnw7Zi9HGCrBTP2S4JTEZRL2at7h0k
xOcpnU1HRff1+Ydza+VXE3/YTttTac3Ix1TVc0wpcKRWw0WOAYGIdBxs2cbGDzFJrGo1gK87xsEO
J2odcBNU5FJy6/b4Z5mtd+Sk8IfDrJjm8kn7ZKcpS1wsupBlvChPRkCdFY8rETx9dpKZ4PO4Xgw5
DKb0WJEkBNIycdI94G+V8xM+/620aR/RGTqiEWeIkwDyxCMo7wIxo0oKRoW1OvbKjCOfvBAH3J7P
/DwG3HZI6l9JEbQSI8mCS4LPd5w4YcBpl2cyYSEQxGHd5dp+43Y0zIBovyJGB3xtkmfW4/QTtuVD
9cYv0mCzLn4bo3W4rXy7mO2ak3VzeBg8uD3JaeVPuY9vE14US0HQza82uPYQ4NTaA33XDdnoxvDO
S5t4qr223l4F1UhPQsVlk+UGqsUCVcSShrXUqR7jRKbNip0OTtSALSDssRbuf1ELqzThFbXl6KoF
w4k0BEEt2PcqxBWc/2IH4UFQo52OcBCDZAz8BkExO1VR6zrvkVVTNXWULhGjFZU+50hoh77B/ekf
9ZOPtr3kaTiLh9jnKcXgV1V6jr3unJEGzAMKbgpr/HB4Fx/+KzDJbFIx2AluG2zy5fTPHw/cVfQF
EwfZJcdo1WEgCbzOTBqkFCrIeufgvAAhKla8fzgm+DVB3k4JDXu2cZ4W8zHdDVT50XWTbXSPv9TC
PuMf5b53PJx6ojMVyHTXRNjv2W6LP57R/1rxpvnwEwvUYUXnnEZQ2skTxiCGfErEPVshRmV8sc4q
OBNFAxI+bKKlmq+ZoyTCc3c0ci/AIVlShgh7osiytm5BSXJ6Q5eQjd2nRYM7aKQtsYEtFjzihewy
DbHS43L1EcXe7ZPRbGAPZjkxFStF5sQCqsIzEK3yFkP3MjJWHo06UfKSjl59oPaAH7G+WakAvzMW
iBnL1GWaiP1yeboOpBAgF19qWQwdEhtxVTb3Yf1dYYPFl/PBhx7nLE8p6knYYT2jjsNOdlP34BDd
iRkl+H7WOmGrz5w2FPdYc7Ex9D8jiJUKa6eXxdsOCfOiFvSe8mDo7LkNFpufRsTPke8578rgaJ+o
SqPjkb+G6mM/YFEx++QhIfQc8ehn4m3RfVOhReXUac05nnDhPtoMS6C38c2FMBkHeiPNu5NNZwzD
iSS+q3ADY3n8tJcloTs0rKCUcDucNFnIBMBpKVdg8WeIWqnMt8gVhC9JaDBdmfRHGT/2q29U17x1
9aElJCyHnroM3sTo152QvTTT/ptNX0X6Td4i6Oh7Ky1Pt+BqPFQXvyW/cAdtjWP9qRVxdVFQWzqR
UqOrTNvvX8PKO75r2CEqLznrqtcsB2AMIVsaCqNw+IeAMM8lRUy0xbC8FTFFVP8Ki0hC1EYQ/I5d
4c/uptNr/V4+DmwIoDk0CpDVXQA892k5nXFQDRhvZcOnZ1y1ySxu0YDmOvR8RagY6ALGQVS1PWtg
Yygrw+DhNwrmgcTGPDw+su3ystQiKefR8cjYKqzTf6+WXpOMiDifv/L6qu/JHicUx8Y3rP8sYdgA
HZBwZ3HOnxZTyr7pMM24ivyzBZaH6q+QQ+kFWQHdg7FNOblrU8qQYfjp2DmyD9Q4HCkaWtxy2Ctu
nccj9PJGbt6Uv0iYh06LPq90XNuX1nAD2Alt+5m9jcubHgafjOQ+o6hniAOWcMIpciFXrvnbLvXO
1WCQwm7ENIc+sZYKQergR26tx603m/gUhC2+sXlAu/6NUnZmgRlSooUEckiRasjdD+e9r6TWLrUk
drJs24hQGQUpNPb9PFrRXuFV5sJZjLYpMJWra0fg7fIOsbPWkOLemwcrJCDl7eKLgrEIg2+Fpuzk
xcC/uK4tXAlcmjulKhzN7ogCAJvv9McTJGidvNCuleLHIoJ4fjlOWe97cfXSSpy8J7yl9TCYofkk
552ALzehT+Wv5njSWsVMkUOoiD1Om92sYll+1Nh0a1nE/u3MzOZhTxyPvrZVN1QGFyjdZQRUCx5P
rb6N45Gn8EMTdSOibk6ARgG9d3+gl77GmVI02KygVe91fiTuU5cG8CQL1e1p6fSFvMHHcOID64QB
ZP2bUSh5+5CEfxirEOdc74Ekof3qa5s7Z2xKdKKXAH/1+SojfijaRG9jm0rrN1BADRYX8RKx8ZFW
ijsaV3pZbySCWFzisCgUJDJHvf8f9aUS8djFop8szA/NIkaq6NIFwOdXPZljgKFRleZoR9eXCH2i
BPp6xZJoZy5/zLYtx1o6SRwWO5sBTXW839AV4isu1uLZj9iWEdfi9nhqoVD1WfQVG5N+y3Dl5COj
jUB3/geuf1lmimxYOMlaLIM8KQCoVBFUz9+Q/nq4d/fBHjLiRsHkVTgN0jrxAFIaLvts81yh6aHy
l2zU0BNHmxIMejLIpHZg3E9xi3v50t1qriQa0+Rdopv5db04iup7uSy0/ysAtAV/XWhNt+nJSoRJ
6IQlABdcCg66V9VYm2cyiIgWh1H8weBXOoabwDavI+rJLvw/StyMrwcsqzLZce5601jGrUXbtWy3
FlpdMfhw858bwnAtug6NmD7UORwF2mW98K7m1+kC7IxMO2RF3sGqobiQJyz9tYqA8V9N3fbyabUQ
vXLNwzs22iyxlyEhXoVYiGCEJrwoB+cpnnG7xudR+HRS+6H7LYhlD5ekxOJD591u1svFXHqOe7IK
iKRU3h4BO7wgFjyxI7+6kdEk3HjXpCz/uHmuZNLTw4ff3CB5ngrqmideOWjj7C+WSLD+U604dXx1
DKTASs0eA/0wwu5YRPok9uFy1RhPFNmUrAptFCB+sL4T/30YEo4sNK2FL1Xm0tz6SMF7OTMrwhl4
aSMvxWX0L2KW8+vcJcg+vQ9IeoR/I1Q/5fA1huitR6XIp/OfTc3K2dgTh009xuIBymf+Bcshzbv9
U++sNNKIwAT5c8EosV8UOnlCjMo4K3HYKeuhaBo1oF1V+OiLWc5L6x26PB8jvpF5I9/zyN9RIEDC
L5L73PqgHEH1BmaKSnHfO+J//Ubsd/f+cPexDiaDqHLc1PN0buj7dhhcpakEkVls4M+WJ9/pCy/E
oO/q6y/7xbFtksuZmc5eeojjj22D/YszCW7NCGYIN5riHP4reRklbtBF1NFR0t2OdIpOrYBCab13
0HJkhAhtM0kXeNmPeoooHvJK03PyBcIQw38vOUDi0P4nyOcAM/PRnKCHnKPb8imDHFK/DSb7HeZg
lilSW3jbz/2Z1uR8HGOb7QzTwRr0G1DDg5INI+jl2/00khhoMeSmZr0pkRHIM2295EerLBxmGwgs
Jn7znCILekwUXg+yjIR26TA41V1y8EepKO+SDyORrW2DtSrl3+hmM9TBmyRWQfyglK5BT9o0nc7b
2KPTY9SCM8ArM3BfFURXTHCfebHBZku1QTqJzG2cuOCTK3ZgyiVq7vNAXGjTJP2hyrnkF77s3UcJ
ZuYizMUpE9932DM3dNGpGMrl7gzd5dZj75FKDqB7VfpMkxAqScXW73eShZGyZ5BLNGYLxmnAbfAk
3wc91YFKd/o3fx76nfdHmXNOqe/ccoXrY09EM47EitEjJNPyQ99RBch+LpcosSvmjxbfW8WbxQdA
M+LiAy7xfjYeRdM5EBYhoI66q1YKMyI+OgNih4hJJtG+JCZSGW8AAijhN0vNvasTT1dzDM4dKcMv
JF6oG0coUHpHu+4JiOARbJ38OsnX8ImaUqabdhSEE7F74ufPjQGpHpYWl4DI/4+ofAh9xM4DOCCv
gnWI+q6SK0QuH4YlMUf7DUvBsq+9oU5vauYw6oLoiZc2AFlHn3az/DrLEo9r1tJUPYyOz7gHM044
ccpXpW8zA21ensNGl7NW/iXVQnpm28dw9w7sClHWLG3lsOTJpctq88mfk96k+pO6/DqXlETuSvJt
+yNb+n3uVEn09wQie6dOeBh51BJCIU2L7c8ykaOSSA2sg+zK5ySSITnmMZMeVWcy0Nw6PEOIkSTQ
/JQdtGeFq7spFRJIdERA6As8rb23OAkW7b2FFQYbwXpeG8zbVCNSrBoalTM2Ne/+Q6qhfezLbjVr
fk8II0LUykpKryq0oN63LfATSX4odQVXV1ZzKNowGBY+TjRUcxGt0EBMeG7GljfzMRz+VO9ivxsN
WWXRdAE2yez4ouyBW7ZZiBWLsmmeWH9/iUhX0sraK3oTRgmyQLzOFsbTxlTSti/jh+EzYHAkzkzq
yKIcwXWLtHqmi2kVV1/AuPhw/8/J1s2rRdHUsjGZzDfpkpsdkwsHC0D5z8dRBBgA8R/BAhUsP64I
n4hYRI0HxizOdOG78K1HFE/DfTdVFDB6uDlEIIdfEFlOha5VLPpGN7Vjg0zTYRwYHjzhjZuT9v6m
rUCi6Ydk3Mmumv8UN6Fo9JL4Doet70ZjK907W+lqliZ7g6LVmKxw+INdvmjQ33IindcdnoG3QAbf
vpZHu1Av3RBkSN6+nNr9iadZkDn1oEcW8acbiLlg2CcNHsPVLT9HLfL6dDItI8BxHvQXay4c3vwj
TgCcs4J5COF91JHDnfe4B0Fy0qrGryve5xftvuT1ajr3TG2EcVev3mc0VU0TZTbBlKQtCCJtq9Kd
VFnssPe5nxd21gqpROWuBq+keSQydMvdQqM4rpHtAvEi9e/f66QVN7ZfPBwNU8KkNkVytGZfNBkm
m0ggaEPiVfmXWXUvOHJw0tf63f45cdj/YA8gxmURT68XOxBD891JuxXLCCJdK+f1QeFMBO+G/E7D
U9LTs47H1lqs0NdN8nM5Cy8uYeigFW7Ot0oTcvV0IBGcWBkQTkZlTBrq485WM9A03fCyWddFeCmc
aI0Yqj1kJZy1ZWW4d63Ned3+wRY7j25j/+0xjATRyGMZFSsXMv3hlevdYyJ8TEBev+ktpX/fccRq
keRFgcu7puX3H5INmm7ecA/78Aapz+jpeLxRyQGjk27UxGffLkJyF8qdbQfI6UJKefrvP7uyoyR0
eK27xSLz6ZAGhoOkHIIV5aa1E2EORlvN5AwfVvNjtEVfBUGTaLrXyeoFHyZfo6KgIr8w6jcUz9WO
szYRAP6MChX38EsF8KnhQF6HnJHYnvgzarqlRBN4kGjTqfWD2uCcs6/cI9nxsYkYbxq02GXCUCSO
oq8EGDKTkqksi6Cax+XMFfcyegPBwDjBnrOXfsJZLKr3hOChqGjSUwSuG/sIqeKz3OSL841CxMZF
tyWmA8sYLL1YmaB6PjkN9Yr/+KJM3uDYcEbbP/BUUNXpO4jL1zSO6bLGn6qT9haW9c/xHuDd4d6z
Dozvv4Ba/fyiJ9Qz5GRucTRa3f+xk4rEg97pNICqxefr3mDHqF+XeQw+nVkjOoHxhbgh6Ery3ydP
CTvvkrS2qv77ATXXNr5TyyE1rYneSTMVlSwk+o/bZHuGtUyGo0ABhoXUYwAzYgu7JrHeaaHDOBUH
o1uTp66IzKB1ER+t/mF7VbAc7LHWoaCjiRkxKp3hV0zYQEHwkExK2YfsJTLHurxxDxcqIBrsqjqT
qV1y1SiDgiYavHl1JevW5bh7XzTxfj9h1xgejG92t/AVfkLmqnPe0m8p+87jWhdqN4zI9JFIdgKo
rlF0KdMgNanmBkPulI1rbGCEy0Ennk/GTGyArxS6Qv3rwOEd3hDsPw3Zz1mKiReNARRgb0jEgCYu
t1l20OTD7iFej21xJLkdGqGcIlY/7ZzEOAXeZgIDN+AZ7YTtnB++uu7WrU0KTqQnHF3S108aGw+m
BhVmuxjN7n5As7z3N0qcPBgCkLI1KrGykIG+t93jIg0q+n+hNMYpOtBM3W+4cyUVNtb0ZX+ltY1Z
FrBv6x3nhXa0YjQskVf0dIvw763+zpBmVGIzc1MxMfBD0z+ubQyJp80DAHnXga1iZxAkriXRTVOM
ejyIy/rxMTWZwM8BLWkEuo3BEqe+LqH9L0Ou1Is6j69obBsi0ngQksSPwIkek138TrP1OTEm2SNQ
NadEkrM0Z3+P5LBuNIQzxsDzqzstAXASKSNpZZ32ffZCbeEgprf6vQFvVYHc+LRTLSUffDCptrAo
DdncNC3c261CxuJS4faaY5X+OFTPh5qkBNcT7SfcFSvlZExvnz46xiDPHAWACbPAutxArqUgf8mj
f2YaXVIT8yfoU6UkMuB8OUukbBGCgYnOoVMC9XN+xO7Zy2/Upu3XYiK5yCXtLIPI+0xlx+gRzrLs
7ufDbA1TCKelyuZEb+wLKvGjfmYtGE2TthfNB338lQz5Smnr023wprv6xXY64WHLhRLFvulbDMWa
YEcR/qrfi57nt8Ifyr2mV895JeDq2y1CBNrfOVAJrRxGqUvdsUECjH8EwbP4kBRjDQgkLRK7onlD
gFPXKuVOOWBaILX1uLWnDwA/IR1/cx/tgrRE6wTwPFotJVJaeDdxBfDZPhoDolYZfZN559a4FFrn
lUZN9PzteGJRf9LNMc88pEbfTOSk/XJ+vBoBdE+YK/Dg8vSd2LtCnfL7nxZLAzh+lajI1WsLUuOR
UOMjnp//5zrxPsNaGAQ85TB6pacAj9uSLTnVDK/xVl6wWJrROJmnziJ1mwWnDdrHn6Q1yDLeVpNM
VsJtFLrIo2mYLx1wvZI9HXAQ31EHC84VKhgqlPfYa+Z46TTNXUqsgcfwVHfFLpJJa4mfCK0kuZmr
Pt9/NYQ1KgOUuNsEuWyxZtRcWU1pv03yrrDJoYt1WNF9+X+qlUPx4MiCoAUKoXj0QpIiDJ5keMtA
1EOweOF+3qJvtm9ZrLq36mOUOEocLEfm/nmTbQ43l3hJWt9nXdeFPd9S0VnnkzgG+gOH89l+q9cg
ryq6qetWVLR4XxU0S1t/DbAoROh71/pWilHUzUSgRHMdyX3ZHBMmG/Wz07bqN9h7s7WxoKMhMFW8
GHKEL3oVPH2dk9TW0tyRaGM7UX92ICkdyQmiqKUfi5zBIZaiORTce6jy839/5yY2TGncBIXRNFgg
ph/JK0h1PfXa5QROb6YVAxHhwT/I4b1Y/irih80oGTcQUfJEmus7TcrULw1DVit9fDOKx2pwfSfC
BI1+jaoplV21a4G+qQHIIhI+ffaxSmD15Hg4yyTmwTu1Hng6aO/X8+bk110aLZHbI1mtBzCMuY4+
ivnj+UYXY/n/q9lDOh/h795cjuWAOCKQ0ilpAsXE2lX92c3te/uj5TQz9Trs5jlW0io2OmCIooOE
ElUk+fXyXPaOJZ2iVyb72OXrrB8D6cy1IJBavC5z5dNILCiL/Z4QgsnjOZShOW93XVY+WOG6aMeA
Dbec9iit66S98lF4/avCS9tAkmIo4OUApKJro3cOnr5GkTDZeUmdkvjiwyqxmb9zdjw/16N3Hd1P
RMsL6txOUcc1WCqpNKyobusVPzQZV5PaQifOe43PXuTd3EnF3jyXbR9pdN6Fzo0Y3ZXBXRVzngTv
VBn7HXQWYX0Nb3YPJPQ67W4SvI7aWmBcmUt2s+x5G8XBX8eCUfDrnpOjuVlWTnxUN6rKHS+Z56sN
IYBSguDQ+F2RlM5nXwDyoF0ud0RzoYBp9ZyWbecmaRmZR96JIK0bzGndVExd8aMpl8wanb+nen0j
YdET6iFdm+zVsOKdMhFx5MeDkQySxfHXZTqBeBhPQRAaD1lFaDFXSww0StYfGgWjyNh2SlXCztjk
nsS9I33srIiTlTXAhvvayRYRqmDBsU2Tr6+PyxudQqrGsvqhBw9CNZDYhJOP5cf+3EoJEQEh7Zle
xq2LApuMfrNn0ZjJer3v03MNODSL1+3eplxU4ONW6ovyRaNagnalBw/HXHPmW/naRaYva+DnMUZi
OMhSXHAJEdE4UJjvF2OHdvydUCaEG2FhVPr+OwCMNL+ibUNJlbQkVOnLuNN8NISRty/Ms5QZBGNw
jKRa8JUkfpCBNSGILamu7BtimtnwPw/PWERjTDHp403H+4YPZ34i/KorM69wkB7gjt9nl5afZG7M
UG7/IVEByCXVyKhZd9BMi7CHyyDp+DteNzFKpseAjfHS26eq4VwkYkjQWFqBC/TkJo0qnhknPsS5
p51UZ6e5caDIxAenO7DK6zK7nOl/XZk2vsyzjthLYr4xdE+0I79irjciLybFXc503Y3v6itWp+Pj
s0JiYxVLjKeEnM5DhkRBglYRx6hg5vuKeIFPusNWh9siWm/9eWRUwdp4yw+H8cl4ScmnYkYPrJbg
Wf26+jd3K1g8OyRzGwBNKq40b/MVqyvuEi54ZIDxg6HN5Btw4kIzsCbW6v53syDFDBXYjAHfqZ3n
hfFgLFaPwupurWLt2b35xW/0Q23oXWoTA2zUg1tjzYzezT383n1/GsB27AEKNVaEs+d0vDgvZIna
3DvO8nsNRkoOTVMlml8JK4xuf+PvK3bgzu5hqyz+dAsa2jIrihpZiGZ79/WX2ih3Rtj4vi7OT2GQ
5uAieBQ46zDNR7jFvncAyi2gQZotX1eXmxbXAZx1bC5Gg3BqN525qO4rUI+rLzVEX81DzGUQNGaB
qK1WYfL+4Ud6kScnldc/UB3dQY8jqY5mDm72WPU1KAW9uuafooWWGDc4Bd3a4DajOW9UulhqcFu8
Nm+gqeSH6c+7VB64JrUWRteXjHTam0AsunIDUrab6ZldLi0L/E88U2Ml455NYMB52sdeINCSaPrH
weT0vdYG3mD3cuGbe3mGxnja+/VWchzHDjLzEWrViWVvLkx2+3uCpO5RMwt/pwtJMnIZsRNwc8Uc
Np5nXF0fe72NqkCt1syJAyIaaOgJLQHaFrvj75h2Ydc4qh4cJHQ2eWtBw5dToaMxPyjOGIiJjk67
fX77vK0E6pqgyEkdTfK2QcYaItlFQGRCp8ZJUQSJS2ui7tGVXenveD2CkdS9v/SGkeVpsqFLk032
lspP8JzlgDNBsKho72rqSrv4ryWypN7C2ppA8D25cLcqCxUXJudxpgMLArnTuXWIC0GDstCCnU26
zb3uObtQsbBzvU/E/XuQBeX2l6LFEdt+ZXHrJLPgHxKgWwsqW07LG96cVB5YlZe72a5++3pNxfeb
2ZqWBNUHuLUakgoLVFyU31eJ7NOsq9LqQGv+EKajLIaTnykVoWP1k8LbY+uRWxsQowybnbfkc6Lv
7wr4q2/izDa8NETX0Cbc9YVY2vSru7z3mCIz2mQALP3lu/YGueKFTS1Tx5eXrg2uiczM/YAx+/Ez
4pYZ7Edr/I3EYp9Md/sVeE8g/48IKLVBZmou1lGIpWgnKTaqiwnbAQ2bnzeElQnd2lpc7ICjotdd
g3DCXNMnpiDue4B+4WSRlkqufq9dKb6662VZA1cU/hts3NKjC7tXPFlKi8hHf5T3i2vknc7Gr142
ffmsFvWdBmJB+hxaVK+qovxeI1jEvnOudWh9pYQkjLQOhOkaviM4NcxDDYnNMzClQO9w181zMd/o
68mcP7GbDvHA4fPfDNgjQvopJtLZk1BwcRhiVW0DlfQOABHeLVr+goPxiuzoYE5hRJxs34J+YDGX
g0NwpRM9wKDJI3l0CTvubT8j/9kmbKRJ9PgQ8Lx+cjHCjtg2dk6WqNMFSurOK01cwzG9zTKtbP/8
SELCz92QqjLbCujGxI/ZKPKu7jba93665QbL4tRjjxp0KSnmlNXAEzh4F0e/yp79w5vTVJjLB1y6
oeP0V5jlWoGaysjWJApWuzzmd6cFWxFsu1SsaXNV3h/wcVnSpVIePX6flwUirxHk0IaEd7Usc/eQ
SRiZITwaB5n7xIPoqIlMSCVn1pkBfvxPhq/AziS6L+HHhiG7Mn8HwQ9yvghgPa+HSz6a3JwY/A4Q
XRI0FDAmmDeVYgbDFIKYX+qKYAC08gAjFngJ8q+vgr47/oazesLUUl93ejkmr0hkD44+QHPORx5x
HsqfJ30Doh3Xt7kkgO/tAiPuVNn9yi5FWf+lzsVt7sj4yRuMRQ/XqTsrHfB3QQUPvG/U0n9T7vtb
ExUQcuQWQf+fzTrk0q2cuRNjhdYlKwqk3lOarjx9835eI7K5lUvFBG+1yz5z/XbfC/kjWj5QGM2t
qdX5jJgJDELn1WcaKHd/s8lvDxhau/xcXdhilXFQWukrPi8xblyF3kacr6WbiyMzMpkdhvhhJPoM
CKa3Cncr41Istd3EoUCA+4qDpeoZCSiIKNce+4Qi8xz2SIYYP90U4Se7FXLUt0TnO/oh6jkHi3hc
ufTGY0sBhiyPRmSxPixLCSE6KARLZ7YoKmJPzVUKHNetS2jkXJ2GIkkpzUeIEIh3o/Jmv88IoKsq
RoHi+kfgDnxpahON39jxM18rrt4Mht7UIT/TGMWCdiRCBhAJuNHZ9AAyTZvEUUO75MHblISj8LQL
0Vvao2G6IO8QqHK8Iam0VMSovTQHx6n3z/bWx/jz10gthmEvZIdOVwgsn9Mx4bx7bOlaxznusiMk
zI/idPB8JTnDSfmfYrb/4kMt3ixh9O+vGnej3ER+sZot5+uDIgVtYxSds/bts2p/Q93Xsxt7cMVS
2XDdSHbHrA1Z+JG/VfE+AonSLsPqSMnxTSr5xR2GFxOST0Xr4f7Xu+/+tJ8QL1Nh+SaUszWXCXeW
z6nRUZgXMhJVZozisCCQozPUVbiVemSaG1yRZheKNdntifqbgZZTbXfk0TztpXqgNNVMSGJ+WmrY
QDgHEmmz7tpOpVJX4jbXnAk4N9Lu6rCmVcD4BRAr040host9be5yX+HZ+OOuCkMzydEEl38pqO8w
ARZ17NkTYDGHk1Y674qVPqwLpvHiGV3yFqdWumXW7nmf6AgwDaTmPhiy6uCP153EzhtXuk+8G6AW
GtI8cflFqclCscHAkt7NGqn02+k7TDZwTn18wohbwx0zOl8pZnO+qkkHFEZ3pKXrnQWv0rmMoE7J
XOABZ57tgD472dKn3FU98SGPq2A07Hr7XDDvwODP06C1gsre0S294bjaFKesTwKmGEbnwabXF2VP
eKjdtND5Hf0dZvaq/+6ruoUrLPMh0o90TXYRd36b+r0eH0Spps5KIJE/q/KH15oyJC6YNDqVUKoS
CQE/asN6+7sEd9qmEh2hE4iJhuv8V5wa9aapsCySsp2xj6lOwQYE/VtWO87z2zXbDb2/hwhyYvLO
6FWeloSPCILoAeTdPXTGwI0MCtf0/fUtmwzmSGDnyH+5lTVWltYbd567GXMz9ZYsFrhStabO77lR
SKjqacnGsf8PTdgCRgHZlrGa4bN8KZw6xSpQeHIAeiYiZMRZdNXZmZ8AVhoINXtGh3hbU8nErR+L
VxMZAhDsG0FEgBEf2bRuLNGR/CfqB8EiquTTabKDBh6gWkrMQikbrwFSd7qvOiGoLomsYqquDz3f
4TqlaPfmPvfS+RYvxxgckah+rQiQiVk0vIZY8n3zNDVmYt0lfQ/x6zeJutSeHQSlH8pC2huRXJ6y
FWsp7RlKDDwCjwMr73oXFI009O0Poh7ZHifs+YtWxU/T4OCnl03UJlPRX4GVX72RmG/kyAU9lQCr
5Lg5tDRlqX+LsWJIl5ttRHm7Tb22DIYunmyyI5VonxlJnV8pujyjbgNCi3r6G7rOekitqDeHbxiR
GjR8lYjHaQA3DI+38RqnQnoJd64VheSLdkTb+Y2kMtViJXwQJ19SNUmOtfF+SG847/szMQ2vW9uO
KCxEF/JdcsRwl0rr2/Xn/6QCTY6LY9iUk4x2el1pd6ISzouJWdSiNcP1DGo9DX41Bw9kVCxtH1QV
/A0GHbk50zqIM7k+Rnck2aBQN5JFfi4M3FYLPhDzZZZr6iabIA6N/E354vld2LMDIe3+1cZEgax9
cDCxxZQYIzw20QU7HVyJqRnDKmGEwTwPA88z5zAoSSR3QrfcRBbVIS8PVnOuR/oq6IF8PScpGv4D
xIbOgK1fKtCCXhhEC+1HECSh6mNzq2uXu6ja71OFrJBrLDuSIj1AfA7cEj0+IH4aWKNDOW+MloqF
cCtKArpa1IXW54hkJV5K0GN+Vz+iVcjFvfhFeuoxUS5WD7xOjLNfHY6P5a/7Afdkof97cBI/+5/g
xJX+IvZ3DvryRrciqDG0a0Xh7TOHLwId1uA7UPv/w4SMGjpxmjZihvYb5m5OZLplQxdJZ71cx426
9IEB9DWUESM1YB0bB03nkxbBD+P6pu0iLm4xP8s5kLXOtrPx49gKBjD1D4nO6gLiNkwNIJTEP1x0
8/NSELS9fvnp4t7gs/wnSE0AEOgEOBld5Z5j1yANRXh6SyTsKob8reU1Ymg3J9BV+O+JJtFkJk9Y
0QZzjFz00cNut1V3IwIIaPnzvmYe8Jd6mzB430bWcVYwJ6a4/cnsFEoRyTw7Er41c4wogJ6Fo16G
IRB/jXujZk7feABvicohaKklvtnWz8Yb5acHsc7DUZa2VhW98ckpoAgWk41/7QcXW4sTDXPYV93M
mPEMrG5SiBQm8WJ1nS02VVh8UfQgic8oJVKtUrWBCJcyOHy16qSxYtxfAOSFJ7KrROaV0soJkWPd
t2zg5pd8lW1jOmcfpGXSI6pvqLYXgq6Fd2q7gLwlZ+qoJaw8kINPFah1SanYqkOHELFa+GYXX0Hp
55YK40WgkI2mWaFPRJWawf+Ju7nk5IbacS+YqwnlSApEm+nUfRVg/R53QYrKECyzN1fpLK2KkGJ5
0Se1eHYrxQiFjPxqgjc1w2YFpiUTUj3NG0oeBOFNlGN25Ub1EKDytvi8N5O1MJmra0yRYk8px4ho
S+dyWPXM5PkU4wTOq1otjsJLnWKH+LuvgBR7fqph6xCLbyf2YR7O+iapxyF/lViewmHOv3B+jpeb
STs8N6VyaP4j9wftGBK1MVtYoXs6Xm+pYPBU5N0LpuiUQckO1I7jTuimyGjj9cHXMBbEeD+OSdkZ
s9ju3Kp9iZ8C/yNCuRsS0Kn/oqdhFX0AB6KvLqswid+Y51+fUvkwpYc++McjE6/iXG3IdimbJBT2
n6IXHMx6wW4TgNmr3AKCqNmDDHLg4ZbF/MO3BzSWf19tAb6m9PxaVdDBKS0fdi1s9ptiFTBIYVeM
wLyVv1PiExA9cGpsBLOzNL6UJMG5ibha1iAYLpODsZet2bGByMZ8w1ydnDE9Kp/tb10MgehdtsYk
TngGMyYJfkUST/DAR2E4gXx05nHBJIYCYxxbkb+eAc7IOw2zr5IKv0Xda7NVQah7yccd8b7JyT6T
NJeAzsDryVAykcC8eUVMvT/UGGLehAhU+SmNcvcQ4Yeaky5IM38eGHAKX+1/mcue1gmQLUJJdJv8
RJBpdBKjY6w6HH5tsSmkKJD8D2DgROD79ziWCm1WIdgIBZy9xKhJM8h8kwEdyFsBiKHA3jCllJEh
ygDF1L2ezhDg3H18eVIzfS/vJ/rHhVEGmhueyljcL6SURnQ3lvPUUlE/weGd+AJbgHWqNa6wBmEw
uUgu3+KN4TfqI/IXGyYlnG8LqI6siKegiY+5KtYtiR+GJlLWJPS58Iv1cbfHUZ66UK1PlTXR08L8
MiQgT/rfb/EUItsN/7ljuG774l3TYfQEPi1LWEyhsHCXr2hzkrepQhPIkdrQBqTq4Gd1M7eOVe8a
n8MrQt1y48802wKXns0si3042fWGrv+AA+b//KM4Q6Clu/75x6DyFT4svyS3R6Ca0c4Sx6Q1rfG2
P+OONZSbpJlS33xMzFKOIYUHz8Q7mlUc1viorzXc5KvyZahXqTUCfIvMGnC7YajZWOwUSmzXxTVc
OtjfPdKvrmO3s3aS5R+DXdUEJKEqzQJigDYktI3LWvYy3bBuxbtz/9K77CvC3y3bCuCiY1XMF1ES
rJ/Qk823LWiHSPaqvd1TyyrJfMC3t9GZ9SXh/8IZ7KdMgR86x5UfcCm1e5tfQWn6Oj7dP4FUqXCw
9gLrAG8aYyqf/gqwbAKZhroXhR0L7ZT5f53aPDAozaboDPEWnDdmPsncn7u3DrEcnbxaTvTzKojU
Cpp5j+6mFt9cUrriEAzJZm73lk1bpUvgHkqZQ/bieRy+nUw51/VAEQ5d4/HMq6/3txbHXabKvl5K
9cX+gNlpZOxSn+uqoz1RFe+/W3ApugV3uzCI8Nv+ncs3iZVVvnBYeuCv2O31Pd1+bPcUYzes5SSz
0LHCoh00reOerdAnVjQ6T3p/s9Urif4TdXStj5MAVkSDiRGS3it9amRoiRFxx+V4SI1xG2UckULJ
JAsxVscEo9n5XeAbapaF3f7cNqVOgYO6HtG+4oxkHPVdwkcrPcFbdW+OY3gU+LJqBtkHIybt6W+A
x2z1hFLZZMH/u6XG92wK9dF3V49FJbK0bRMxsJTqFASyzCT4Bhnz/UDOLmNT3Rn9+2nT3IZCr5ny
QJaKKWhA3Yq1H3lFyKKzNXl5OuCg6K23d4LHlE2q4GM0z76IbSWdIgug9gQQOnjbRMxXSVBdrmTW
hPxcCuYKXKyRNv/dx3m4vIQGi2SKX2hPmcuxu8kqPcnVIIViYrl564J3IW4cfuEamNHAEEXAUpWh
n6OuJPKwO5CEuGXw8X8rV57cvazVNiWNt0qVnudRFilZmZ0YKsamnD2Vp10X48TvOwzurCllJWZ3
9FsOggdX5aTX2AqNOkEvvq0DDuKhjkPmdBYqq3vFmf47pSRswodWFtfvrTBsKqjmCuKiiHvTdfPX
Qdt9qRv8FocxYq1GZpu4YNV+Mk4+3O3hXxFPBxbWxa65X7l6QUeAGXjB1SfZWOEPBmhN0wi0nU+u
EbE8/BB/o+d98DHyKkoHRfWrqO+MBSH+/HrlS8ctobYC7/HxbtpQEPVCFIefVohJCU/bsCIycNqh
zSN4+g0swFOClwnrHAV1+OS9XSkq9/btTwKyl/Sy065W1dTnw2zGoC6pKP2fAL3wW9pxGoBb8QbD
aJ2A0pYXfoO1lZeV0+mLCzhieopJ2g3EEW5+eZIuDfz8HGzS9IMAdfiGSvpotcxhP9xMJpB0vG9r
9I90rcwOJCDgHUdITjNrPCnu9ZIfucRHDfw7oOS3d0n5FCOckpXEyxQ4ib7rSqzWZsi27/3nheEb
E3KF3sHm8cZtGsZFzDKsjg9hmGo6/FKV3Xf3BfimnyCkOMDNOEw08aqA3+h2gHcXeaSH26qAIrK2
ow8zg6/GEoznVeocM/S38OAIUDoDxduwuTJJ2oU8im7PSJt1594h5pL+ArMLDPLZIpp7XppOgqZH
gvzKcVCUHf571NBYFxjKqePasvds3OYLz8Fc2G2evnz1CiM5shuYpTQxYl+hZRAWmkZJqi1slAWv
Ox3DRI3zOqidDYnNR/RtpaJTwSxrzns5eeoOFO9sBUcnpBd8fzQPCsNfzgKklBQEQRhMsHIIMjRr
/Jg+7SadMl4sM1OuIcvi6unYxz6GIW1IMFM/MN/tQg+i9+t0vYWPgEWf3IOrxQCD9h31sN3T2XtG
BhehSpH3jcvFSNIK4E58aNn0zj4pNDOpcnHlcA2YQDXZyd3VGIMxPJQthZcXAfF/kbTzWND2uqmB
/VUfFy3fPjzIG2SnPd34f0m/ZTwk3bfZTuZdT4vwjjCoxljAFZ9bVIVskEPC7l+teBM6AbaGWCSU
5zsRh50oiU5br5oQ/FZINhfbxlfgOn8lNKX0A60t09u+PiAbmcoQBizCvYJoLOtjh+t1M489qX6I
ryUoDmEmq8g0awR1MyVF/Rzq4sL3/KlUhfLI691PUpEbpXTEqM5VzoktoA3UqhxAxacNbq1A7XNd
Eumjn+E8ks0dRjcum3QTdM1wJ+6QpPBCbLISUX1ilenmHzOJaenPKoXaVjQkdPqmz8QkHKfrH60l
ZePMEdHfbDqX5SC4T0l1wi2TLZbwTCZDAe/7pYOlF4W0g3KWbyqHx8WvwWA4Wdtew6OZCvi3q2A2
7TVMQZa8INQbtbedtSE5UtSP/yIwSjHEjVVUmaqgg2xe3qcR0Dr3bOWCBIf3MNIZ0tYTTypptcLf
wpmDKXIxsqzJ9ZaZutTVtz0ptTPOCF0QfT7lGn8QPmWXYUseYkvFnUzSVd6nUl2yDAgdhpXR7+dU
8DRfPfGQBAXjnf4tMH+6wgmUZlpPST0OcEncVuD2Iu+rmhCV1lhGqSuDesE+JeSIW80pcr324Tal
bEo+GTGmbad6KW3QffU6t6rKdv7GE9C6rzfiEZemipjQ05cdpqCKLI2eXeat9dpqDmZqirKjExFO
PJVKhhj0BWpp+XuxjDWu3/0YNuPinwuYZ3Uf3gDPoFXYPbZHe/DqOZjgLcDd8zia8+Zx+o3GEx2L
ctHjmouXP/JbbTi2+osKsq4aTaZiP4VepsQh2M6MdTecTHWECVlLBe7Vxhm/0AUBDwyvXhtQfhb7
kkCKdUygc1vrw71G5JSieZejxh/p29NOzFr3MKIbBG81VdFYUd4Evl/6Qq0mLFTA78+sA3Ha2Pe4
m3fgIRodrZ/OCK35mS++3DU1x2vJsJCfqTCqDzxGkyGESD9iV5MH0tqCXPhgP4fulG/ewr+VWaad
/1wyjlOPBZpPKhVeVZ0L3koYF8XyNtawUOoxfQL8fphFJtuuZKJQ+anydr1SxTVJRcK96lvmSrMO
FdRcMw8EcC+WKbLxHs85sHBO9DnjXcEUmruYtSmnUYgigMfm/oqNAsXFKX73CHSjQxMmlgFH1vnI
CPe+ruvJBPbFXUlYH2Z7AQAJyXpy1/OCpINobzWe2YvrX0KWEdgco3Tm+4qEzkmjq6t1zqxxWdz5
FZ+2S9XQV8E14qktfcHykWMJfXSxqKrFoDTyZE1EZR6/ZtIUITQSJOvG0Zgw+InfvyAJWx0ODZcI
NmNeR8gE/B/9Pkmoor8pAntAkP5fuJMWNkOmI7uM2B6sgadNdYS3LAUVxkUUcw1m1Wjj6MMEJWLO
ymL98wl0rPJCiHhqrl1pdA3P8YFHXJPbdXy79/9gtwNdaI9qN19UKmAM5IaLOaf/ciykMQvPk77q
lNPppq7e3Kffgp/3M7HY5aUy7Aqkf7iMSs8JFlEeiPbleTCPH8/UMPDaXx4xv8FILJPurP4MyJuc
VT/WW+YBX7z7hvKO5BznRg6NNP1I1kDPJwMn3iYJjDRDQlQkGSwqeojmff7umI1k3c4zCOk5h7wg
fv7pyYfO8xMC/OaRj/+cIgdX6ZY0C3Qxj8ODUXugNHjZn6BC3W1z0VA0IMmrt8zpI9IuabLiBjMT
YDoU2EEDq/JZLbF1QqZt6I09KiH6tdwVBmxkQinqYeavcIZcWs2sdt2cgFju6s/cRtEJGX0+dfvX
tGdKfbm1PPIVRVzb/CRfqNbnCuUJn6eo0/XSSar2L2TnarlG4WAbjCOBkqmsKolij9FFiFJQad95
3rwACdImg4Lk7G8zK9LjIXft3uqaIW1gx36nhhe1pHEYRgHI6Ym35eLqkBaAwK/kpC6yLBQZs688
fJ0q/aEigDkz3qTpO7oJfO7HfWejM7Lfx6mYFnrfdrrZY+z/aOyeNe/Qmb3jPguzuCwC2WNIjy3F
vsYpTFqRahP6TVCoX9v3RxRsQQm5eyGchFJhLPmavq6R5UYsE5yFhIGfbkRDE4UbtjnFNMUNdNiZ
knmtQspiOkP4F8YeLrxfehYAaFQJigCrhpp0Z9X7EUaT5jzRFsuJD1NCCT4XJYCPjlXO33EDobtO
MJYe72CMSJUoCvN6GsLuTMfbfej4MPx1kx/2J+g2v7Idmm+u0/6kY5wGXPY5+hMIJnMdOwQCNJXl
B5Esvud1WYhzG6tFy1pH3RPLA0nL1mHcN4Ye3ZOBjvyBXLMsmaECNBu70NqaAttFfV1iTVnIvhsV
8tPVBygAohGmBi4O5hE7DUsNMRwxniry6x+c1YoTlPPjrTE8XX9pUKPiED3NL3msNH8WI9DLBbey
Gwm1TZULIcA9Y07qQKGqwZoP+MxeXiTJ3A3EHnjmtEAC6ssG62fJguY0Rc1Q5SBmJws6ucmy/Jxg
ytutnVbgVVGBEoybVN0p2MXT0J4VbVvjj/Z2xrJ15XodRQy68cxj4BemItT9qkPF7/IZa9ahwLCZ
0uPV2XXJSF0uHqxKd3JkrVXAGnm1M6qwW3Yh1tJT5DPos04coK7t+/bUtzTl1xGNf2CSpbON77Za
PGILKd782n4rew6iTxUdxz/oULvqC9savWoN169eOWkO9QY5r+4of0MXPMBVnCcj5peFHBKKyWTZ
GbJmJ9ROh8GNnc+sMWz+YBY5dNV3594/y/M7ncDbx/N2ICiQeMDU65oJ7jd/JXOasOiSl3pQk+ZX
EH2Pz1aYylG9FQwJYkpW8lHysbCpXkOWJi7Ry0mBXwrpY4bXYiPLWgvn+pqAW/527xrBTVmLkiWr
KU5VnjLUjyTw2vG78dmb274Q75vEFZ8Lq0YGm/G3PDhq+xEsCRQ2Awm5IbCBYMboCzOqFvTgId2c
MaVxtE8diW4YKTJTf1bsKd9Rv6/tBu8bC3CgWVk4noIEFt7fgzkDm7udII5d/P5RsCKBMyCIyhw0
EJETnqD6BKyck0l8Osx+jMZHxjv22irKY0lOHmsFh1vb8RtDRbJ7aTuZ0kSGYRrQfUXuaC5MNvG/
xuNVGRigERjqKZVY7Z1LPqv6drFVXxjRJY9vYq83+cMsQ49RGq8eUCTL3rHFPf6wxy9E+LwovMRS
t9tU4GTeGQ+vCALJTcIY8iABoschjzl720FpHI4cxbDGdFkrY4FFx4wOrJUJ/NbhlXJKJAIQS2iF
lWShyqwEMMUwicdLcyq1C5NkPg/rHWSU9iAdP/zAlQ0iKk8gYFr34XJ/REl0gbt6W2oiLvyTB96w
36g7yFycJJK2e/5RWhkmpBCca/Ih4W159nxV9oqN1JXWkpN2yyH+srnwCuN3W0D4Fu4lCGtyltLj
yg35A+4xDna66JAHZCPuDqHcs2LnoiGMCltm28pCosuQTbT15W7cAY62iBP5VZsy5wwpToUwrflb
vdJdGjR95oB3yreV2u4b9MFQff9IOmIuBPi7BRb4I5Qiu0pdjTOBeVoLFaPellG+f/PwjgMRImdZ
qtz133p3OE8XIqRT/jgvopm2TQevxdNbe2LAOmpKGdO6juzgk9yXu6k9pL5FiRGJNxN82UZ5Dyx6
xCoEXFOUNyc/Iz5B3y7NPy+UmRJml5jpOGRnYkWMIGgCF5D9j7EFpxN2ge5XM4u3c1r+0Ts6AXb7
oz7MRFZiSJLHchieEs0thrqR1DUrFzbiAKcEvktlAS+Fx5uVGq/vPBvTKL+E6nNJ5/IeYv63C2bf
NWVV9+QTSUe/L2wenF+OqpjNuv/mu+9EA8geHlv1mtKSNCJF5E2A8HTkxu/DfofDhwuSWphw3F5g
QjaDmYaPOdhJ7vS7y4Bwk1cxplX7mQDPW0XWg3h2klimd/t/sHIuSbSEaEms1ucW4+uBGOpW2MPP
A2gnLX0Ius8bCZL1LGcfK4UMw5AOxi+uS9kyXaG81/+M0RQsYyvPGMWv+uXx+gRN71FuBlsDZkcn
N1MHiOLPzvvJ9iy+5aF+RDkeszduPQ7Cdu6z/wRaax/ODAkxAlUvOgZVI0MxtFAdUJJ2D83yQZer
13FnUCy5V6wfUqCJLNvhC1cTpoy+5l7RjPsI/IS3b0RiX3CUrhm9VdCt9aIIQPK22sGhkXErI5So
Q0DkMuqV3BwkcO9XHnIJq8yhWUTkfi+C+3AXyTnH+lfWQYPLRd9nMxuLgVTd02Qb3I/Y6mDy7E2J
xr88FdSVKdsFNOor0jDSiMvFtbCtn0zvT+Ae4fkMjQf+0cI5qSMItpIQIqMl4ATfCjLV93reZzei
e9aduXxy/uj2uMEr6NaYF66CYaTRzTzhufOXoz5PXwB8lQieFnIStt5zTd8mb5BF9oFIUP3ZEpha
Pm0CfDIe7Ynd7QCXOONtb1wVCk96HtAYmke4mcXq3x6TJFaYxHayEM/hKb00BjSKLFKTwtBG8QBU
DimVx81pVehv012cUUUiySzKhbsuTy7uA9u7y7I++p5WMqp2IVNY3HMTEZFWh5Xceze/iGmhvRr/
OMaDIOI/1Sa1nCGlkQvmOEVTJ9XJkTuwIH3I8arr2/E+cN2eIuq2Z2oHpVB5weeM2PIHWU/8wZ2K
Q/9kGta4OxPlHxibq4uZD+TbJHKslDL9q141pjptAt2x8w6/0carfquAQSUWAnCaD2r81etnHx3F
wPh3OeKeOZXncM8F7QumnVKH61TK/iXEG/B/wXX/rnu35fQvLyln/mSeng4VhyYjj6wSrXFOWNxY
WhBncWYUU6O+b17G1voFq8sMznNjy0KBq2Vh5w4Ddi+hUCnqyOedDXJpbhqhBEoJgjTotqsE1fVM
Dn4s530sZ0WALNYqBPVvgUWtB8SGco9jxLSfILMXhLOTW1HcDsIUOzbFilYasPNJ3hrSdv8E1fCY
iBLXNpa5qtUnfPoWlq39yUdx6QXrr7pAwWSjl1bw5wVOt5TnRvp70KjbkPDg3iPuNvUhw89NQSfT
UogcalkT8zSAi+mWmUG5civ/buE6sgV9g+n2Pft+pwhh6aWD4aVmuBVZROyLE4dIBroItfSEc1Rb
9vrj+/UzqDLFgQ7ai4P+TTuOVO5G4C4LIHR/gOH6UYejZR25pNZWRtjb+7vdZe644+Nub55oDAyp
gwYqOO9KoNo+zkECknIC9+o5+IxW2iH0hwebD84T/0rzn5AzlMsYyizBLHjGwiMWDVaS4CMJ6coz
HrOd8rPnyGUq7xkV93PQaAMI/8d0X6ZaDsZ1Qn3PT1Y6XipFFhNtU82xGvK56omJSusnhjQeZi2D
c3eck7npYa6RkxM9Cn/DEcQt1s1gx8mFXRqrZmQWaqT9iC8LRtYEiRonWz5/h57HWBVeQjT6165F
1qrzRho2cOWiP5vOWWt3EESb2BeF23LoLmWOG593PssM4Y43uwjX47sLPnPquHdtABBEgR8f/9SM
zVJMOe8lUeIoyaDSubPWAeQXLWTgOWJai6fAiwEqJNL2isPv3dzFBxRzDmZiKX9Wxb1P5tknlrst
tXsiL6Qh5T76YlIO0AXD0jRHIWe38vF9tYKkEiTA3E2RhgBvHN4hJ7Ky1wKID8HzNJQssuS4GlCx
uWZhRteOCflz0jdjQSWCvtA4GoS2cPPjrEvq54YPhxFhzR67/57v7qjvwp13WCdBE0vzWHJEeE/C
CEqkgDN9PI8JD01Jip8cUAq6ZWS/8QKBmLQVEFsdvvQW89xjEo8+3M0A/MRax6POq3i3R7QdjEj0
YIHsl4LkyoU0GZSKCwG2hy2DMaj3W3MniGa0Jy2v+xrQtPjfgpKPpYZOGDm9V6B/7+qN0Hr1XDfB
VF/qpsbBx0Sgj7SZxSgvu3C2El9FKrJelhW9ElcJCgKtoImfkRwucYxF4tq/eoiHaJUMGWK09aY6
L+/Hzg1syoHP40YWZetQimM8W64AmbXFSyJJz4IY/E4scCqgmuas78xKUmXfMqP0gjOYs+cPZFYh
7ycyiDIHMDFnVlQg9pSQ9ItcsZviCRvMKnUq/otLXicaXf9G8kUesPnEJ2P4mroqLfzm448fboI8
zg+uaW9tQ2qj2TM6AVqoynwZyobdjQx/x575rhGsE7WBkiBKwd6k+15VnfS2wQJIgwWWx7JS9OOP
fKgQGeX8fO5Eg1P41bT6SSvrYR88OUhGt9RzD0SitEfUHGNU3C8+Rg+Q5sn5Yx9Utg0wczB8y59L
fxLR1Tnip9EfjS8XzDrKYI6sENXzuQPxyXEF8WOU5II95oH6lnbslYNAznhdTzeFc/m1ib/js5C/
nABGa6RHKO5qSGNYd63HzpWFTIVuCD8d3jqQy0w8T/rnbJLb5PdLBeD19rVr8PE811OhoEFI3MgA
kYa6SG6uZvGQ3a0X2Byu96a9K3GxcfCNdV2MjadSwZ8pqT6m+1C16++93NRFBRLKWdJxBjzgG6B7
yaZoUCb50dRUKsLOWT9GoQsFfmwEv+Lu5n8VPNyAac2ZXLE4dFwyc47PWcHb3IIFlVxpTmceE1ao
v2rgkQRBTVtTGxklDE6pwGZumu89ZrQHu9EOvAguWjgyANIUTkr6Av84NMmv1+shUUQFMSJgm77f
dcHpKWI1LsHndV0+mhIDUuAlUQ/CsmSTanmrJYynXkbzlDDsXayyBlCnLsvniG8NzpGK3Gien1it
N31fStcfWd5ZcYlnyYDte5MmuDK9kpulIly7BuC1t51do4sx5Umm4F2QYgkYvyRD2x9Yn90M5N+r
anX4d9yuSbcqAiLH1X8BJ3rHyOowbEq+enIaiUuTGdEXY6PJ/5fysfI850sN31UqNFPboho4DJkJ
xCbviwRAx8pN1xLSOq7KHSxEiMKoZ27ozZIgu1UQ+7WEd1RMYct1usZ4mZmxyykZqankqu34xR1f
ondwDpRFYIOTxM5JCKUpC4kDe+N7SFRP5PHWeQI4DX71DoqcOYQrnnx6PGI1gxTX9MT1LUDozZG5
SbloeECznVc3sxfOyI++tB/E8fQkMsccPRHvdrSjo1qn7HZnVpugMKt3sY5Gf76jGhLI2kPIpTt4
KZYuk5ZhbniNk1crNSllicENWQVPqkfKZ7srwvBVO1ND04ydoKyRUGOQISCSGk+5/zsVJe3qQMkw
Sh00GDkw41sT0p9g4j48fam/4rTLCR7gOJ0CJisKS9MdLgbD3Z6cRN3zJaY2Un15BtefqajydxPc
72pHcA8Zkii8jh70hfbB91eCfrDDgO35W6ABafbeR1lA+4BBu1PJm84ur6okArUlOJ5fUUIVa1L+
KqtVMLxLsdgcXviOekVBq84VdAQfmur97g/W5cj617ykKAHaBwUCfVM5rzhrd2cGA3s7G2ZH99sP
FHMz6ZtTI5WO9aY0fFYYMHGLuYVgpQa8AUzrAfp1nmFYiOJbopGX97S6xCMJUl4lSz/nTW0VAvwK
mX8vpV2yHX0MfT9K9dHdEI1RDoTngWcdN39NGPnG/2WBKVVz19QIN0NXY/ZHH06PSEYnnk5Go7ch
16rKrc1dwEZHUu8Q9PwjaAPf8FZTgVVVh7xYI/NQJCKA5zGTj8IntEmc5YSlmTkMXezex4lCA+NF
h9dkuHCtTT0Y06VNXGJ5mzzd4aDsk+lgI7Edx7kzygVOFNALOhwg1/HX7fI1bshD7xU14CtK4FyT
U2tLMxRh+Z03AIRbDBQYeUpcwZVTmCuFUrYOk1WZphVSkgXVR3ycmaJ+tYYmRHR7fmn04PwijTYx
ipwPWS72RBsFdc+iJ25A8NZgDs+Dm457gciEMpciV7smuev5PrMK5YmgHjeODNdt6YxoK3YwCCFm
ZxW8+lgbxRhqOVmXf10XQSfeo/67xuQYQaA3U7T/xGz8xNdrzrE61xbVeVKM93QRrXtoXsOyoSYk
vM2jX0VdiiOnIJqfJSsKrbVpP1iAzmVPuvPZ8SZfFAqk++rWHaDHVyf9LyqJchZKIRvizKLJTij7
CI3YfLD1ON4aQv5Qw0fCRM/y+ou6IyS4Lvka4ZIqYcuZ4TrqiucdzzrGRD2eio7JArc0rtT4gLdH
HamOQdYcUgyMVEWm60T7ERtY1bjBZd6fS7x8me1kZq2VCRGAoHKZa8ev3R1/yQByv7tez44SqTY7
68Kb4mAPdRMFT2zdGSUVAytfJsjMDecMp6HgzkCmX3lytLLyD9CC2+s8WaeUadUF2ukgRIIGQdn9
OiGST+PQ4WMwgEWZT/of4yTcAARyj4lUlmpY+nOTiQE80+LekrNLpbQiu6yNCgIDj4dTOGuaGrZ7
qCgQiPU5Rg+N2rIEeXIYjaw/wKbHs8vZJ6iVhOrs3GnSzskb+kMS4zPhTHJVTdV+lVHS5BKYtn9+
bMojxHbqiqAjXhxbFTJVwN7DSq5dQTOQrkeVOUkIVUGykxY1fnE5QOKSnS+RTi1379hwyEs9Mj75
cdpBm50Svdj3zZQtyMIqR7ESIozuGQ8JVA1r3ZEDugeOYYIHRVfqMhn62FyFhjeRS/bz/SisdA1c
eC0g5B4ZqCoU2uS2DiZ8M9Zui37gVmFXycBSb7NXNxIcqLmCZy1ftjL9UJxe95ezCZO6wOhcjL7S
5mZZsh/CXcC6MEx+a/qbA9hAcV4ilsPxD74BfhNrVGB8fEN4LnKn36FY6DVpjKG2Kq1gMxJYQdXw
zGhEvBBhq1bvZL5O78+E+hrU/DIsg8KBlqWRvcGnralBAtVh/4mgQyyVBcsNc3prsPpl+KJQ3Tu3
8giXxVt5BdcdhRIsNeAxd4OKy7f/ky07jTDD2vbPCd3WmJFC0T959NTKhqinkw8DSM/YYKi1y0kf
uih2e8SMrrHrS2awsApR9NoEcH935blgLG/HN1vww6AlJeCeL3+1y6YrpmZdM8UuZu2pEy45SnMA
t0fNZdR6bDjJF/nBnMp4xv1vtduALZeGU6wa3bAS0SVmFmXMrSdMhSkugIfHfbB2KnzTKHp2Wcf0
E7MDo8UGjpS58v5rhQELnxzG6XR+Glbh9HLmNG9WCsePWudwK2Bw03abkSgFH+Ngx9FcCLI3LarI
f+GG6yfYXv4GuVWkLxmVDg/Otcu48AEGzI+Guvdtg6Icx52D/GaNXTydK/YLeI2T0s+/NKz2YE1+
eY72058lsYKdhpntJXsmACa5xKF6FUZMeerhpMBlKL01bmzE6CXuOFyTNCJMOLV6kwUfs7QXY66F
hBGFBjosgFOqbwUHjPE5q+UVUPRhdKNBi/jMKBkCGShARjXjDnBTb0WGTsc8SjHztpRvAoJvvINX
p82ewTpx+Fo6DIav5mtbIjZpV8n5zaDEyZcvnY1ZLJgu8/iP5VuKjiv1ZEkRThoD9ucmwqKCiyG4
WV2Rw0GNt3y/QLLSjiR9d5iW+2FQbODak7WhGgMmXGVFnbeCRFFO0czPy+1IGxHu0B7GmhpfI5wj
huxtoUzOK4+rkK0+AoGdIpScvYWUBv4ofZvpSF+iNG5M/30clIWNDsbptZysqyUNMKwU+2m+Lb+3
uGEM7tCCie2EhvAarmGnqK+rvw7AnqbERFXExsDQE9mJM3yNQ0oyH3eJNa9BSKKGo3iHD2ADckXb
w5eRxpf9RwPmTRTz51LX/iNWUcgyu1u3y4zJDONHI6ZLXbOut3UE1Wyqt/tm3ik7hj6HbSFfLtc4
GluMeak6MrUEpLAEPFNAlCqmYFccTokICGyJiIGzDZcFdARuTiRgqixL/oKUvp/sR4vzWNpUZzqb
Ep6oIvo+NgFCaa6Oe7tqppYANGxaDWgt6I2UBnKz1m+aR33xcPWiWbDZSfMc+NXf6T5vgfkdc2/G
ehv4Ub1+kJEypTbZdv32Swm0IbIy1LimlbkWOJf/qBTdDPgmDd42jvCD+taCaiBSE/IT9SJKQSs9
xsnbyM2AeUUSU5mkgg1pIWwoA2+9KD6r2JDX9EZrfzI5vGxelu5QCGen+V5OhpyZPSWg63XBtaf1
JtDbYW2ZaRTqiaMVK0RsnvsHDM5gt779rcP/3AB4t4mDA1oZrc70hEYZgi4bXV0wcB0BZc+blZIe
r295sZOLXJRW5I1QAIT5vkKbLBGwlvkNqsHPj27NtTDVbP6rCCmdjbqdn33F+UYuLLgt4f+Og83S
x/XeuAp0SlgQbG6tf6E3wBx9Vj3dsumu9IVOgDTIwU4FRgvUGmirHaA1Dg5sjKYBotTwtq6la1/F
GAqfrcDpR2ElDuK5WC/tUJ/ChR97w7rynNscXbCi1SkvXtfAGqB3u4Rbl5zKJIdxgi3QeSYPbqnn
VUUz7aVvCbskrjnnENKxr3MbDdx7RdjdKZ7ozMcZ1CUiLE5ngd/GkQk1Tol5rytZRIdlGqP7/uD3
ZNpy2vgiE5SBCBlWZwQDUmKlxfIaziQ0YNydBbKxsPef5GyYEI0HP3eXTit32s7mubd0y297vWux
dcZeA+7VF15j84xBf2EB5OwKIku09gLlY2g2GEautipPlYj+kj2DPgrzA5NsWbOfB3LZrjyI860I
wfrIX3kRvQ+Srmr2acKUSPHT/tmqYJdFwXbQZsBMPksq9H6d57V/SQtdtUtc6GBpF4biKdqOXByy
Oorjr0ugcDFEiLG3Z0E3vr1zT382aJLuT7N0x/nn4ewmSNPdC5W/FM70woNZbOn9yO2WuBFbJFgK
hr1HmIFvjQnXA1QoBL0oF+L+ptiw1tuIzELE7dZPQRWF3xu0jbsc30Il73JEmQHautiNib9Ro89F
JBoiM8Nxb3xIlek2tTQmpW5mldZnMw6wyUZJGgl6H8kXv5weCzeBYHAPzWWPMBqkZC7+1Jx6U789
H7PYw9c5Va8a2paDE9ljougfNE41QvF6lm+5XCOUdUtNdI/BzXFNHCIwjdjUhpf3uSAmle2GRjBW
glnzlze0ddh8PHCSc+cZGycmH7xqZ7A27uS8vIjp9nvVn9UOyOcD6KbHDLJ92DnR7cCTHzbAza+h
0J5Yu6QlLC9WIPjPSxN9wqGxHA56opRSep4mcC0Hg0ZZcrVcbSBWuXTfhIAMxKLU5VPpMzOswhfa
/mahRIqqgPDABm9rS3NdkrvoLpoijNrf5WIUIkAIpc/5uPYjikbe13FKlWIRQdB5HqNWDDwFMhgq
w6vG7uoBmbJtcqkJ6DOGQHTd48Qu53zAOEg/OyFd1KCEvamAEWIpSA+DBBZqX5PYXedgu5ipgWN2
gZHcs3kIA2N4FLiz/Eg9fO1vnA1pGs3YVPPYr5vOxj4YZbCt3qqS3qm6FFEn4K5VZOEGEphE2R24
fqtirrfdL8sURtRGRqB4YkI5dc8aOMa7g0eoK9dO4Dc3McNd85mA5TmBiYpqsnRA0c727sQYj0Xb
86Q70I2+iHamQBFQ4+DFTfsx07iZGnZ1b8xDqi5D97jon8A54biRJiQQXJzDgejqWCh1yNQRcWj5
G1bjlS1n3hQjy126/8/Nue21wuutixXc4Tl0xfaXvSpKVkfQb8ChDrKs2dUh0Rx0ePS49H9//Gcn
TUaoudqb9nFdexvgLrIZJOEwslDo7ygQXKU0np7sdPLWhnEuhVNBilRd4bvzeoqv9pPRjORdCGCu
WbZ84LzEFBcawCo2vH/oGn+RQekfsMEwdT9QAc+J9jSVhSOlRjtwO/+8qrrMyF9DvrSedteaSrQy
VGChjV7nyvCSdr9LiMYj3y5hLbBRdFJ4FhO/G1006GX+khotjR2gluLGz2WTYLgkE5owx6wR2ejx
DhDGvW1LFaJBe7D0oz/Y244DrGulMWCeLm03a4ZfCsViXuf9h84JGrovzk74RhLKtIeeKbNxVbk5
r0QZlVVkP+xWcojjb1RE1+JDQXSrTSQ9vUs3HtF2sI24NaSD8DF/An1XVOAOk3Y0qQGYP4z+Hh13
ZP1p6msC2L5ekr4ITqQGD4qQwgD1xxAjkTTxQ2ykFh65vptj7LYw2z7b/HOHGn0UiNj3ftIzueNa
TuLXjxX/JrMUZUpu+8S+wEv0LQZsfnOg7YEq1Z4UNKrcUHVcbF5yEIcLpicz/aC9mi7E+90391D3
c76g5i8yLWUkIXLeH+U48lcUb4/6zZ7Ci1a7LCQec9A318MXM3J8r84OEfMl6UK2ncOpvdu85o8H
MrmNxi2KAp3Ko2r5ZvuSL9O76g3XImW2/fiiNZbOHkzX5adD+Zh7n/nokIx+9nwMbZMRaLRThg4r
p1Z//rkInwBjVNd2hPXX1/yQDX1Dg7+GQNgzOr1AZlrcKw5LLB40CQ4qvxERUplAtLRjB2jMeQCW
Q1yz8Z3RYfr1SyvbiR2PcsCBfqYVeFkMbkLniCVPiBuEuIehMrEqmb7a8LKwEjVVUNcifMGag2CH
qF/cGCfYU09NAhi101fgSkI2Rk8eDTrXgXEIDWJc6CNyJvlQXLWRGlzq2XqLwOiiqdRZmpmbymr3
IctLAAL4uJw+4AYwrDfZFnpesEUz8HS+SLHpqwsP2MKdity6psyE+ZjJPhiCdvhUeqkf4NFuU+fF
a1VjaL0DFs/tp1/JOpqUdQ9n/8AFQrWXGo9ZF64W4zfMkwnKCD1XjwJz0C8sknG5BNMQTcXISdWv
tvsJs8ns9yS5F9KqjcGx4C4/gvMs4xSC9dWQMHZAS749d0aIBLTyVuKOHPMP2yHLPPlczriNubHP
bnMCmoJNgKASqH54zXJwbb+S5mW3iKCxhqRaVo6HFErt56eJES/920wAsGUFJ0XJ0wP4pmFWCO42
Pi0cu1OKxIUQm+WCmthpgQZK6XWwcaUYwiglhLhTr8NEBtQJIaPF+k3VAFI8KWW/Q6nuv+HD2PYy
WhE092tZ22PPvei+NXHVOjps629/zHbyQu62cLlpseX0I8MEUc/FOnWpmHuK5N/0wZDKCR3m6vHh
2zv6U+SLxtxwb2rAR/MNFCi4AnsRE9y9rHnag11hkfwuOFHDNfYksGEynRQ467ZTUKrZ8NppKrhg
/9nVsCjQl4e6i7QDewUcnZM3prUc72n9U1nGYxb6LlkhXoMHfUWxhAa8EttfkxTewfqCZlBbu01B
7T+fmjgZZehU/RjhT9CTFjv7bWCYN6L4Md5wsxcx8APAKBQqbhb6YIjodDPWKaOnI81ewAfUk6n8
HJuzmhMP47Xgc1brNyydM2JIH6bWr4qfYMiJx+6yHNLQvlwqFzd5TD6xbgelKeUt2llLjsa4KHNi
fdCFd+I6FRThakFhJkLCjqMmMMqsbBAZHrorlqw2ENqYfq0e01XzympiUrizg3tkdWHuIi+EU+uK
i2cTq2MWzJ0+0jqpcGrmOSId6UO6zPJRXlJDO31t20Y9+GZxw8IQ1uMnKeiha5I1MTltjQvmInWC
d6ONvwCk+OhcvF3B39dO0im/QSKceki/172NdF/syrCJjjfOTvK3qRldPjzmqBqPDb70+kLp4ISj
RtLUxwqEDWm2zy+DJ23FAhwHj+8f953qycBovevpJmostT70kfK1MfR/+RMICUN65XzndNZFlyQT
v6f11earpe2snoVLK+QzPNNMXsUd6z8a+m934ZdgU+njdvzi6Ob17BxM8D75KpXFQEsAHhn2b2Us
U2XINMa6MFyI8NYlFtklzooYxYoqd8yHTHphY9Gvbezr34dX2f8W7AFV68qERjod40tILs0WO5fH
+Yky8Q4bUMZHDu2+IzipoR0HYmOUpHtbMoDagcdISN4i+uYpaDKXSwl2lWCMc2pdqerqmIWzPuQJ
qw3SLAl3AyivmYlMPcjVcPpZ6dOPWOycHtcJPjYILu9ckJzt39JcO49+cuOKubEcvuPo+P3P2SVf
SperLZn8AskvWaKPknB07wn3M3kfMiVZ/RiujGNEmetDnhttuChf/NXxdXe4nP5IW8f7Fcy4agy+
FqQ9Sw1EyV/i+qI7HznAbLJdm6dfYLwfJ28P8SqPooNIlmLZdrX+yV7jh4t41OdolWn+q8jKUM9x
cMf+NtQifdZ3cN9l+a3PSEbtrABueeOpt4RIWLzxBjd0vpqTwSkOxWH6mUi7Ygld6LjZ6ID5KbX2
bMCZ2YON06tELTIkKd0ukH3lax6SNsd/YlQNhZtYJlUL+TBCxeHD4SpUC6eAGou74pLhD4Sbvokc
wt7C0ikrXuylstdn1/1KWbYHCb4dCj+KLU54CiNx8nJQx8QUiXsPIJlegeASVS8UB2Gzz1y2ko4f
jS0me0sxVbFRh6fJI/DOCl/VwiPEjT5c03TtGH5qZ1iglFE91z9+R5pnBadQkjUN86Bjx8CqXpCJ
qJHlaKq1ndXtldMMYZ7CRel3R6RMOaGUpM0ws6hGhot+DRfcsFOyhL6MPX6CaiSLOjot+Kwp2viY
mPe9ot3TH8ruBXKITHDHIrkonHi96wMCmrmfLWYjQ2FZP5/J+SV5NDs82aBnKATh1QWYcaL7BQeU
W4qho5MvimY4R3FNCuCB3XlBxa/GwCnYnEJFwrD458C1anGs+cjkbvOET1UmPvoSAX5B+FKXZ+61
aUilAy8ZeUeOHNSw/U2P/adPZr0aEicoQL8UqHKVwQwZJjcFLivN+7uhhOUVIdJmZn+HzYp2JzZ5
yPkT7QDpZGWKJw6iagXyaGVM+BsHN6VkUeaWNJ1U5UG7u+1PDc9ZCUFDeOpov4LtPLcKC09BsHb3
0AGn18VhdATCvDTcaR2CbDrcAfVo/oXmvBRqSvKSWhYxU5YkkDXGg/LSsIXbOmVpuD2CMSxfGxwt
6VFpPmtnhN3K3MMRLzna0KsCYHiuGRkXuTNh/QduttZ60CmUpRPt4/O6m0JUPnC+tVatmymFt19p
5bdR0OknUTEjvJfZe9JKv6pTm6b5gzjIZq00GovitfSR8hYCXtx5rCIzI0FrsNTyrIjUwTpKGsMS
LrBwPjfFYCQ66SEnQjHhw3QbQU7Bj+Qx5L/BOzZFMOniPj6GVh1om/xQZycjsEUznVUDPg6eyfSU
1DCxKdSwFJ7CcJ/8O9bOqfrWMfZqAWcq9ofj8AtlfA05mFfrdwVga+fuDRRKZnaY9HD6zYracO5m
d6RXI4PlHadh1SxQahN0Pcsu0VPzXPsEzOatcrlq8Vyj/8ERNuvK7wAVz/p8e7b2aN29luS6tfqE
BRz58+tPejec4A9SzJXdD7jtU1U+l5Mublz5cLMZlHLXqzY5L2RYrc9PHCrjaTMOaM+S1tXvng4M
PEDxjk7mmEpr27wfPK9z6aq11hOTzYh5tHYOT+pVGb3mxz53ZUCpkSAs5Gs7kE+jjkhgKqZE09ra
QgrtLmBu0g2HervVEzhNWu0ncKXCdd5lHV8cBxH9ZpzPE5ckCZtgzuSED/rpitHYl7fuzkR1vX7u
qH6kuS4gnO1VWb4giJujpdw1uMALb3sFDG+o77/otrTB5Dm/Z/iNgc8WQX2HZXO83zezgvGvjWPv
kkCCNxb/VYTWsbpgSqJONTm4E1sYCYDPHEYE+MvnGFiYvpw5h8jBoVA5wqwqfrxjitBRWUqB5/f4
v+syq+mG+rHe5elv2fHAygivGVkyOCLlvXDGEtACokTdxvFH7whIQ6kkh1p9KsDzbtJJ0579S3/P
yFYWw3zll5SfY2h6pvAmPLIVJWAZ/Nk2rJHRkqOZTQFpQzp19APhOzvw7RCzDfstVwbb+ChqCCLq
dB1lTF8qKyV/LlX806ie+vEjgLm8LWuwTu+dEFgAgt+vS3Ffw/CeEjBGqbkjHhNxoX1gRGGeS7KX
FPs95/W9M3vc2r7TpaoRlxgJKLeFnUieqaGx6q6iWhKQOH6npvbEQKpiNGKJMmP5LllinW98njLO
Frtnr45yQcimaCsgnd9b5tQ6dTYqkpsP3VSlfL05WTV/adAU7SmhSy2Cu8uP8rPFgLZCzRqkBTja
xO6LzlZa3B/TGVC7pmxz0HZCuieEQgLC1H67z1qDoxvllsGX2ZovWrmsOSsNCMlx/XG33ueqd3Ty
NQE5OL2O1vRMu31HZkcFGVAWNe+cSoAHidmQ6adw09Vb15BrDSX6LKzAA3xWAg9GBdZcZn05AH8W
O7KBcV7j3wGZRiwnDaxg55Koh34DP7r3wGkyxj1Bqqw5ppV6x6FCMIKl0m0QWNw48nB8J1JTGkSM
FJel8cHiygHi9o46UObyw96TbIKwVgrjcA+uZ1ksu50LPURHww49Nw3crYIhS8fxOnpNI3mS/+ad
qXasVJuMEvDmWJPVfnwYTXKYqHDP+W+b7I3NS7bFb9ld3JXVOwJy+Hs9dvXn72t7nJtZbpFEnqTx
tDTkAIO4JeJSfqM5Bx6FA1vg+Rv7kwVfK1iJff9gfi3Zf3wdFY7yMrcTYhLzVa6Nt+vi0XHDTgpb
7mdCHut6GR9/AW5EJP7igYjXyUbxsyVeTRGPLRtBZYKFL6F7aF2XQ4lItxEn3BilCw9ws9vqC1AZ
svSLT5Z3acWa9hrpMIFbCZMDzaJLu1jIxRFJtWcYPUKNiB6YBnHv8+dVmKlJNVvN30fMgvnnlBu7
QX3iuDf/E+R94wbLsSwiQNpGnHXMedn3vNciubUNgMKSBaNw3Vr8T/sIxB5nPbd95sRuFw4FBF6K
0FS4r5FSUxBnhapMA+Ey1D8MvlU6Jtx9yYqiX+VgEH9Z5waYYGWXqR4lggbaNA6vBlswYYJPj1tp
u/yTXIeP675iJHxdIsFhiTU/96JHUQTmT+EF8Y65RF6nS5rqKMLw+ezplIzjh8PS//gMQvoxYwEV
LbVGgBYQDNzP6LnLohCM+BHPbqLd4IXdlNa5mREfEA4bNT9YJH+OeTzvhZCaKQX0BqOSTz9ai99p
ENsheSfFe9xvXq68V5ke89Te9bsVp7jgSvRqx5pgneEukI258xPHmVo9Esx9OhVgr0C1QInyGsbU
HO/pzMihqRmfSaqqn4LqCwRxB/Tzpx3qpbujJ21bD2342ni9n9TxD4JEF+9Ir9TMSBER9fznoDTQ
WXwuTjyEc8wcfAzMTR/Q3C58dNsuKFLwWKxfTB63b8H6cUWLJzuHZVoEPm3PMVeu1Iah2elhu/vQ
c8cMp+JrwGqvvDbWFcDBlPri7VkQQ/t3Gwgb83oqjYK0roeP7udCgxClo+dYrO+lS0Lxt3lOn4BD
suFyoFkFXs/5pPtZHF1E60Ua6zh0OYidw8egUTU9rP/rTRqSEJKyFv+cIdR36QBXwqFyI5vR7WAY
qvN2h1IVUxoqVETajr3WaveSvXuipGXMN4J+qI5smoJTBaotaGJlSL7kKnTnA41cPcu/4gDwvh6G
W4yJGgo3Yl1ZHzPl0MPxail6LMmm0T9/6edgyRBiQi2yaKulX53VZYxL5Oeu/e6919UXTbQ4A9Fn
lcXK9VPHHf4pDvKNROoSgihjH1RR2+azQ6p7CFsNSqBzKWOxMQkHmqO1X7gwLMT1V0DoXZaBGIm9
mKGKhjqIKpYH7joXczU8QlKggRagTK7Oy0RZgT5Q5AH+bzqSv3XC15ApXJgb+guXI/VYlE80CCzI
+L14FQup1um9cno2m5o75xFRxVLlpPhj0CDTGSsxxOLnBupjut8GFbfVX/NZ6vE8NAhungKi8vVi
ZkdiwdCVKPCg55jKX/Iaw4AmNiNxiHoVYEr7JqDSNpBqJfuzs7U19RWilhggYJVlZ+OfVQBkJTzB
1CWVQLnBHxchbufssfCkWCh7x3vQwVZ6eoXuhf+7APeJtzUI3qbUCtvFBijb/Ig2za7GimYXB6ZK
ATOmZB/oqluRZ2cBMNgHVYngdzpgc7N0VGp/RQpJsYMSm8RSYwz7Uf+l72kZ5ByjMHPNkQ6hUi+H
dHGraHXFsLSGAfyIeuQY7lq9YilmHm89MuJ9hIn4D4L+m4Rhr+fPCePywgxdMkvDxYktk91g9YiJ
uadQFEANtLeKhzSTLiMFixooW+dFFBshLPINhy0V+tYq9Rja48XuRcSdSuwV297yqWIIkFNmJW48
0wsMkkpZpyeJcXODv9hs2LTkgEAUqA+UnCfXcs9XB0Vy5h6YJWvLtptUScWSbjs1NJRL4NbgQO6X
YNhKYcmst7DnFUq2zSI97K82gP6smhD2BHM1e0CACCr63REjLgyr+i3YyJyFV7MdxXEf6A1ytvs7
GY7f4M++CtibxdLbOh5hkZWBSwAAfwQemBS8C6jvYWRt30dVvgxWqW0tSPSh/W936ycbHUCpcgAr
AFFet5nDXFkxi3R4+SgPMHSKV0cNEK/lucyU6lxT3iupWkuysg26rE90X2XzGhrRBo3f7ZLW8sSP
SWB6RR93nyEN15MQjKQkIXzhURoi+VRF0bn0JGJv4bBfv6sz+BhUxwVP39cEJURHmbCpL+cp5oAl
z+lb/jAivemg7KPmy+eB2pkN0r09pVPXPu9PR7E4nHPtBplM0hbfZa3VifzWkgA9rj8PJVFHcwlO
ZLU/HSXSp7ef3A3oVU4ZsU9agpLzJ9JXuZsrr60MSQVH/Ut/0tzjd3T7WHMeIbDx5U/tWLZOwVOB
Y105hw43Vv6oeDkwFm3q8hrFb0pf8ytFxEm+LOqF9qXtkD3Y/J/CYFX/LJUiFy2sSjDbG8dJD9gD
LdVC4OZmNcC8ohDqifNs8AO6ngURgwcPxWasGBVqqILYhS13GH4HoljTfgCCP7lYd60ry2MhR2p7
vhLsRS/5t4T1UP1VXnBkG187HMIkzCwdwmMLFRp9AU1V2Fi7cBGl03xxTfAG7MjFC67tl+ViJmYx
66LPbNgp0AiWgyLwddDeMlicrDGw+tqeq8i2KN0KHTuaf32uE9AUPrXCuPr42PMGPVPToGg0XL5i
qx3mnPaM+F67eRCD0XzrNirZdwOO8K1n4VOJeuY2QhwHo36cXGr9Yc45Eg1rRXZAtEOZphRlzv5G
PdqJTSC+T1uJkK/6nTbXtfHZg6fyeGjYTCNsEK1L69hlfEh6/vebschdcp2u67sfIEplmCzurgCv
wlQIm/jnc+3RENwflXJKhKSx1WMDAANuUY8ofcI9zFhB/AAfXlZnFlTG60bVn9tPsfUnbiUJTqHP
kcFhnOENvVh79hemHwZMQgfzSDfofk1hrky5HpCNFbN977EsDNQfanBEU5qYYmwSI3sBoHGw5J+n
J/+3EtS0fUVU1RJoNIt5a9h6ynqZNWK3hn26TFVKLrUYOSEEJ38w/xkxSTOfnxeGhRzksTOJNglA
DlZWBuPajVkoC2QnJBgJ2YVJ0YKinIhO5wf+zhzqQmMLIBWP0ZdshEBTSXkV/+rAFajuRkYiTa1H
1suJTTpn6qte3rpZfX06xLtLloYF7ut9uUNhZnpZj/1U7FuXmShyk63eaKSg6FNCK3rN3L2f3qgQ
3KgWmEx0Apg88WUm9/QoZZh7CpicytFSX9sShbg/vhGoZcur/I8gVDDf/ccg4vh/Pd4ggdlzBoFJ
GFRYXeDkqaCWWibCW5ujTb4bjUO5WqMXJRk4rpU818bZ/i096ndHK8OFJGrfEI1C1XRj6hrfk05D
T4wGdraIGQZ1erwfWjh7+KHDUBT27ZglKhV9tqYbwwn1WcEvNdhbPyJesJlzwzHUZ9ke6ER+z+Ap
KXXFikuA1ANqYHHJmlDHPvKrscJU21rlzen/r527n09pqrmGeP96WTOdKUWZTZ7D0jgcoU/oUUOQ
yluPTlfg8Q6qpUFldZn9pdWg7OFS0fSu5iRFZ/nBZeL4EwkNK+xdPRJQPSm9cq5CzFK9J6Cd5+Dk
903MGQWL2LcdXZgTtVvoU9KPnt/daGkH4YXaVom6HdhNvjh/nN86sMz7kL2BofMflgL/4DjxIc8F
7N8EZY1jkLeCrAC5t66iaELGN/QAIY4kShD4E8r3p6vQaA4P+wrqfoXjJXXGNysnINiW3mlwYs3m
5uJnOCA1artjcXICyeEvCkyaz8ZA8uDWZIKzGsGP3HlPiLSZzw/Hfdn+u1fIa1DEoduFP0DWKw7Z
GdZuHwZ3dChjl+y5SGxX/eAsxozhJT6kkwcWe9FFUzV5rrEnJc+/wuGVFgFi8KFbdatugwO4tRAJ
rN60gZYwXyOjxMZFEGzNAQbgbQ2TZn4U/IdkIbxq7BqkvU7DaY+HQqkUl0lH806Nb9AU7rP8OcEI
uk+c0rZSVykRfZ98Qx7QK6S/hA7+R7jCzk8zSGDwpsz9+TkZw62hB1zCO9WTFYMeu3mSKifSfY8M
rNl4p3n9KYXGcjCQtaC/tjY+SBKPdy8FE1QqQ4tc/m/Y9qR7xG16xjmBZ3Ponv/OvLj4vb38Jdlb
MB+Ku4AiFWgp98aSVw/5IzGhUTK073r/a2h71AWM0bT96wTeDpGW2ykgegGrfP/EuwoT5yqa3QbZ
mRwmb/kli956m/TcV7pMbQPHv0drJPY45D319jDW/o2Mb/SSuB5a6aS7PZ8NsR0Z01a04/ygUTMx
w2unyDwpcH53g3MSpSXgGe+prXuxIHnoTsEw0omiP4hj3XKn/TcCICxWMtt89hJkW6JQ53FnJ6d+
IZ+8V+7DDoWQ0j1lXlgkSteFoeX3ZT3iZ2IX3DP6WJBnp26sV19OnugTooBjE/S1x4qMMpp0H7A/
bqLcTkBn+hfvY8/mRmCaS2ZnubHZM/4pON9kASXMlZjQIMOBNHja0gNnv23AjTE1j8QM6t2hBlIK
b9VYqVkCkaCF3q1oAuBsn3ZjX3UcgtIgvPUqEybMOOD7h1qlrQZIlw/jTyT/FdCnPrkRQOo/JZpE
NRMeZl1/jogbfeGuchJrNqQavOA5vtGsNqcxC8+sO7c1ak9D2DQ0XVQH94BkASH1s0ZA1qLbuvu7
ZXn6MZk4T49q4LEXI2Gri8eRZVbsduTs3CyPk98j8GEzYiiXv+GQaaeOX00TDIx7c3XC+B8JUKQq
1i2Fthluq45tyN47renm4PhqRAVEQPkX+sICmFQGOvvOunHvFm1r2fmNPeeoLngneI7+3FHbEs2X
HigqPSIZYVyW+cUBXBmNi/NtSApLY7ZNAC2C6ZTGGhD3Zzy+7iJPWaAOtRH+1cqUSLCjCctYIq2T
qiW8owphdK2z5cRo/jnbhjMwyhZz7in7qXjGn55jBtmOzdI4d+djZuAQJazL4h5hmnoFbAwd0JKI
PUojTKRWt9ZI9uyLD7XaJRNgAVpvzgfLVGnuH43YjlTUfEDLnQO9NjPxqTgDwyfAjZsz0zOmhVKB
T06APZOVBO+jax//O/m9nQKUIVLbq02HslVWMj4NRYrEgiruVZELppgueXORocUVFGT1RqHFUaxZ
jwll9rCGmT3DUf8VKEMc5VlF4P1Oz2rKjHRw6Wn+gsLTK/nyLSHkBj3JGI4i2d9gb1dntaG+X0oj
usoB1Cs1qJRGNKdOLTmd3ACq9gWblROHeL40BeDagYV1rdcSr4MpW/p1imYsVMo19k11EgP0K5NV
c5+l0/mfxsPdVPQZvRkgkcipJji0aTkCRrHxDynLWEJvW6XYhs0rcg5VtDaVOKxRn9wYUlhrugpT
hzhHH2P74t/8fi8n77XdmscMeuzsQT6vkVHN/D4l78GxAJRXDcLa7Elx8XdcqGNMe6B3TrX3zIIb
pIAuUoa5QTbb3qyZLbg7Er6xRjzrGGfQ5kZQZt6raw3gw5XODcCpyR/1nfGCZ/Hgb2cHsBC/k5sU
GdV7EDWZ9OaqTvpLeMaOvmN51r5wc6CnCRdH/rXxR/0RdytPlBwgVAbFb8DLae/LmiUZbQ+a0iUy
bhay08qkYKeTmKaGRDJko6IcJd2uIXkPImpDhXLk4f5k2fObLJIFGc6z4cxnjFZRSGkIaML/i46o
IxYKKCdD8zdvguTvnpKBv2W9EuKpogWMo1xVaF7zCmnfQza8Ze7L7LGSYqnG6n6dGvck1Hd3zsUo
zBDVuElOVRtzcBAB+7t30iOEkmX4RS8/KnSJUQ3bSP+wCpXh4EVOU6vMFC07AFbrnfWywGELsOQr
A/HhWd6+ePNGj7z1Tfl04Njod6OKnPqYSPzKeghwLxJQhvioJDBLShprjYxAJjWc9/LB4BHvujjA
4UnGVXl/JOgdudg1xSnXGqBo+lI1ma0L0+BB7VgEr1yUAbc7ZqigdCKUa4Ws2cfJ5Szld/WVWmNg
3KvjEn9/PXFnYsn9xY07SvYsN4BSXVsebIX6qrWXc7O15bNTS3lRGckvMMcwha8Dh46yAsECOYJZ
MAxM0FaDD0cRY7G7dk3iJBtKbk9WpIqeBRBgfOc6u3mZNc2+omGRUzZnPMhCZApKeU1wU5SI/uJE
SP7zVnVovDmTVIepSen7QxxgShoBGlxFZB4SpWRF2kSqqSm8rpF2cSAwfM6jAE9PaQT/d112Yzyb
UN2xo2eZhh00RI/cBXg/bUBiW6W7C1lbDyzbO5ailTXg6k5/gnCLy4pgGhcp1FaedOZ1dSmqXfqp
ixz3algSWBDXhwQcSmaKGAIg3V7r9CLaZ5dC/KC9hI7Tlm00rGfGD3C2lOa7qA4mSRhzSnj8+cOz
mpPQcVIxo359fpBLVOQ7q4ivjJikpmJpHJ26/1VQku8d2KIfsjWWgCSjzYee0P1lC56TRKSEblTO
zJz/2L1XfxN2BGYPTl9BiWUT0LATXlBc3kadMVcTE987rXVN7moTHV6QGJlM4+t+jQksr7H0x/68
AF+r7yaR/Ew+3q3lRCdWNDtEw4MyRGM0OqQ3v2Swo6xKeNJn8YRXtcIarH1Opi23YbrD2QYwqcG8
G25BhxMCkzOWPjggYYX+fb/bd9DgOuK70PoMClYkOqgi6HbVuF3WR3CmHz6IMtO1BHr+YgaZ4F1F
sf9M0kaqbr0rliVqgOuowUzmHsWOszzOhHOPjunGW3kXyQ1A1dp8zCsgW7nJuKvaK3y0R94KtPQX
9E1GtayjMwGrB5buqaw2/FfWnfbq9JixylLXW1fyLP8VaD4cGIgezapHF+K0hCoTepwZgtmmeI0I
jXOLfEAXZbaAPlXIn65IRdN5w8dIZHyR3oOqg1x0XOd/fuYBHkbnErV6PUttKkh92yjJA7kK8+D7
ZLkvlahLhG9LUEyysovU7rm2HvlW1FwXs5n6halprzH6rvAZaeK9LwUA5qQuL/45UDBjJGJppFRb
KLA1Kb8HaJYb1zJRF+7AHv8Oi05Ze4pm3bcRkrLwiMfOXvQiMb7GuZdXwCTCcjPK5w7h+cgU5xEW
/R+9JPaY7aCwBa0qOlFHf0T7rvP9X6ptbbydoSjLFjbPyOxCB4fKuAFbTHsxYJ9udiwpVbIunQlI
4awOMzpcsQ+CzJ3kHpxxQZruIvovYEIMgODyhvZ607DlTMsjRjVml7h0p/XAmTlRXS/6GrWzxzV1
DbwXPlf44eutogSQSI83QwLAjBd4c5OMW9gSz2tjntsbx8aSSE5EMB2ABkIMhKjt7GiFk0JaB+hz
8zNbT3BXmGt/aYH4gMEr/E5kbclqM9Ep63QK5M9+ogiObIwO96k8P6Fw+DMAC8ayloV8hDqzt9Kf
xV0Tipt5T0GdUuVxW8Ftd44qMf/vB3zforhzXME/512CtfqOuj1KIpyZpEjb2Qwu3JeFCwHdZqdv
KMs4vK9Vpc/7WnD5Fd8/y7QYI/Aiq9JI/XN+ZTsU0UGz+dUi4eeg4JItX8i5uzwV8hlGpMCGEdi5
gj4niJPYlB3APt/YJ2Yyo4eKSctLTeZ0tyU+HfnDwtuBjwzYqjb+rEfn4DguKXbCmAxwi8v6VvXR
Aa4nbM+ZY8wzecZp5IijqvlTnKZnKdgMcZ2yzoIWmPrqJ2489LOUX2PqxHlRzua2SBWT8GcwfARv
t51xUYz0C8rD3kpsIWZJTuE26p9Lk3VY2S1XPAyBCsvINtrSempKNtAML169TjNEAO0bGzOKycyL
KkURoxEjoDmFCXx76t7aOxmdWikHFBLsAnxVwLIDXknSa8l1WNxaoXaxCRkFcUd74VbhVQodprMF
ShZNH+HCDjt5gC95Rq9l8XLtSBiv/3DRR42+k9V5YnaCBNO/+16diAhfjUWNJVWkLH7dRl3jn9/W
O6zdGTYYI1yM+E9Bum9rMZJFAaxCSgiQFVaPfXGBzJqc8gKt7pD+7C0Kq2GqoNvMfTpBGf6vPJKl
NClPo89J7wE2QCB90I6isRAlMWFqgzDXUIoEU5oFTNgkFsxe9pZ8ecpLssl/LOZvmAcgd1bpHuHy
BMthkcu4LU4rz98f2Gw9S4Ae8J5wh8lcvL+zGZkZnF6bINumvIGSS80ZCm8X0/wsG64pl/vMA0dK
epEiX2SS8p6giJkoQ1AxZ2BcIkqQBAPmYXcihL3xthsYDMrd1bKgpxLp6zJwi4bCGLw4v+K0PBAu
TxEG7I/S3SXtkiZUBhdGodGUqoa0lS5mln/i1MHPdY2xn9YWZ81kaEgarFv8+1iPqKIkitp4MbZJ
OBmAKuqbXbNBD08SFD/LvsNlw9MSxCsPOM73ESCLLd++3Ws0E6J4ikgEkdXFh2018EdaW+y/xvA6
g+g/UJI68fFt/ARXs00hgeRmoSCJrZU66PyceGfWMpyaHGAr1Nfc5TcJMXbxrvP/1CudoQ9WKRB0
iq+MYjnv3izlyWSsDz5BgbyisyJbDCD7KezyphNlpUWY19qhaH5wfJIiDWyRsJ7zomnwbX04RcZZ
Tvdw49epP+cYNOquVqvRe8jscI2Cr7jl9qUMo9NN+BXeZAgrW2FseEr4Iut/ORPu6nwzkkHg4eQp
CETVV7XS0t5/hzqZ33nBRgthJY5H9OG8m/VHaK32jjvlShc5C5TvaoRFFa/udAJPQJAhUhHfjnzj
H7ncgz9vuj3al6bLWEmSgpWgZL/37BCqVpAeK7fN4uD2S3S+M5q2wnPu5DSINnNc3Z/iXl9gpIjP
muXHqFUdCLtjVFa2/eDFGPSHB9E6HWRdrloA/RWzQckhiO1pJ4IoZq15xfR2a3eiGfRmCBh9dlBx
gZQgBlw3jSzFH4qCMngcsNfK+UeupeYcBXJA9eiamhg+fmC1jo8CZXXEpkuvs2pcrIEXECIEUzR6
FNh+sXA0KVn6aTR57kbs7pkNWFK0cIEgkjiLvukQiy1tzlkxvAiQ0UQdzrhLnWRGanTfwwksMX7M
b5l7XOQuki4seRFXvkrIsDCnq5Nr+1X/gEBZFkq/tDt8V2S2/nBcuAMA49zsCghJIJSFu5uLT0Rt
ktkB07/ufQTn9qzijyvkpmk8CDxRI5brxDUQYCjqqe2H8cxDgBK1yswm8r84vfzFmL9TTY3wNQoz
IccxC4N+f2u/Wj0eyKtxMhoxv718GmBzY4K5p8553cwgPcmWkmnGFJmL7G0acF0PBUhNvKk2P7RY
b8ZlF/+2vE15EqpflPqZ7+9K8ZtIuM40IClwjnj34DbNj1/aSNl4PYa7nsGkuQAEPXzp/+6sm0PO
vNPgaMUaZgzbB14D61zZX4yd5Qbm5NcxE82dADk+L6BcGjH0G0pt8Kbm1MTKvD39p8sE4J8esknI
gbTpIEAoSw09YC29wkSYTZi7bCcBM7/E26npIx7kI2L4jhB9BEF8odhuZjXltIY3F1nFy70iJVu4
Zw82gqCJCeyNNVL9N6KNQ8+aMG8qy6diXI2U9jtCsLRAeHAlBsiJqD0x8P462WAUpWjSdtTUoqMe
dY+pTWw4xPbECSxNeuri9Kon3TkgBnUZpJfmVNqE/inJP1xHKBY8jvWujigIubaSnSaxsE/DBMFu
GAn6jILCAw6sOR5bN5rTL1vognDhma8zEiH/+uQMaXKmBeLDPwlLu6ni6U6T+MDHcPQm/NKK7Llo
pCqrHRHEmAnYUfBhOg4vp/VefDnQSJzkqchXqPdwyx+DlNijfgHow8E6W3mDw2JR2Nl25FNzQJXU
VzIMw0hgjeo3AzKorPsZvmbfGtU07RfTj7vXfJCE7m9q2zfXlWx21AVd6boECY5QsGjN0iM50aD8
JCWjXHWKecQhestrQWo4DjBg/Rdzt5F62yJieOqBl5RtNYmluGV5K4NM276zMlgPq0SKKg4q5vU+
c7sSqplxCto8lo2kA7lsACq7QvZTuIewedsOfE8V0YTTQIevd3RgwQYYo6Wk9RscGVcQXM6NI0IO
3ACCD6rlivJgt3gY1eqDdCOcotoQARcNQ35pZWZYsHnbWUHmTnIpjrTvuZAHsIW1UwbLYrBeUzv+
PO4+P+9uPRIf+I5eohUuKmrsVljXAdpOAD1iJvHBURxB+81vPqHFvN5jOlnLiiH7ckLhlaRJs2qG
0sCtfjpka5bTP8Pf2LOlUTtYuUTHyDx2HbGsqyYcBc3hoz2Wq1AaCqfEHL9R3ggtRG4dmOgjeGS7
pbBxXtR135y9nXOFID9qqipeUbqc9skxgCa9deH0fBfecGY0Alg4ymtz6ZQup5CLYdajfvbNfX4f
D+/zoExwxh43g/I7Y02bp5K82K9kbA5YoJTrmeE9aV7lbvSe9z6dxqYzgf4p+h9sWhxZegxobl6G
n9NXZaa6KwEYkfdObuaghZUbkjAww9LpkGl4Crkb2fAWMGSfkcscKTNYCpTHXHPMwYQ/INW+1Fai
ntaB1YoXXlralwX+/SW7/QCzFY+tFGh+oCs4rTEw283wiFdLc7tnErLuWbDWj3aHDPz1EAfq1J+E
iA6QmmSJwt5FGPEASYRHwYx94Qr4bD6OBGz96Gi7+wrncyVW3Q2AA5BhcV3+WT9AN1d7tAtc1VzA
5BDFJEO1yKh6NTZnYd4ekLIhOg2+WSiMgGCjGHZW/Ez2cVZg79bmHPjFQLuWLq4AvCoqOGcsLYNI
w1cKjn5zHBZ5yZkFbagAMMOXP9R3iHXXrFGNnnJ3ruPmwMbY9MaFpVFaL+yM36Vj7DbVe08vUcd4
tqmERCvkrunwragzPtIzqWY+OVhHmDJgrXn00tWl+NYQ2ep6nL+gR7MdlhaHb4HAtd3TlpCHkVkK
0HIaNvJLCdRPA3a/q/6VAhJa+dNm9hB/Pdv4x3d+Mq6TDyg417r5lcf6QYKVc9c2XdwIMaVJzBcn
2RtZTSH+53Ubxhw5j5EmfCSoKt5ldYqc3+rUpIbE+h70RCYObgF/S1Jp/Ig+pj/XP0sx6K6/oT2r
iGsOJy9cJnn1nND87vOEIUg9igkj4+n3FullRMugzR3MsyqolbGAdYG3HyBooDnh1YhHuIsgAtf7
mZR+5rtv0AwhF8lrjLnqxM9+Iwd+WqwgAK1pq/wIl5OaauHuEuIJb9RGbRiEiSkRF3mTso0YbMwW
Km+gSF5eVeNjhGWFTbiQJ7inud/hJ9yPq1tSekqS+B2vTub3JyKUhaZtB2C8UpXUUvda3WK/ydUZ
Bp8muEsf+F5BxvBFP9jXzQyMelJaAYV+CLYwp0ttAx4Rwb8yfw/YlEshoJanl7EZPym1aITfHGDs
X0aaSe1eAWtKccyDEWMiFEbaz6/KY2YvWtwNtmtzzNd9pE5cgZN5iTIENnGMVh/DRVx7Erp5HNAr
L7Zj7+/zbUrxzZqepU06iK3PlIPiVyGkTBNi5tENBItt5kVJ7a/n9wFr9+EcpA3jpDPqhTLQyLHB
gupdH3SRGQXmgFsZtH9KkQh4SlkoQEpRS1T76wMv24x9AW56yqEjS7pLuuI2hOyvw462aU3VJErq
yVACaEyeoMat4XmIspMDz0eFmB7XC02If/Fir2loQQF9/Z2WVkrS1rmtcxRbkggmwGNhnNrqejEt
rdE0qd8MLUVKKs/ZzTuf1SOI1U4tQDp136vQUE66YqBWGkoIlj1BvMEO0PBpimj2PxJ7JKDuWWl5
6HDrYOQnVZb0U2UvGu4WpRtZsOu2jPVn4Rnbij+2MSOaKLdzzbYoVwX+YLzCq7XWJJbIu64i1AZE
YQ8c+dHkncfZMdoV2KYHbdbyLbL9Qhk/kqZBl1qOJ96sAk4GS9pwDOgRy5zOnhbniZJ4MusEeYr4
xDP9/yy8tVZG2D3zLjWgFKKEirUxL8pKxjRqsM05ydeXEsupO+GMV+1SGkYVSQjRNhChXjjYY/aJ
Gr2lFmTAQartDGvZQamuX13IwsnnvMD2CwNYgJQ0L/53Mx/aU1yE+K5coSuKIlp8jbaQFLpb80lo
gsZZeGNqmd60M2Oid297njxXR944+O9/10XdXh0kZpCcy6cX87dOLyvQeG8/rqNQwI6/XnbVC+Jq
5cjxrAeM+wILvGIvzBI047exNWYgW8QWCO/uXJztNWYpoDuGl1Bcaf8Z3pRm5ye65THANMU1lMhz
rk6ytn8iLD4yxDDwXEl1KCEbmZnOybxlUZALh8oYy/gcydwVjQvLIA4UxA9kixYHruiiUv/Na8S4
7IJLKLldIt1yS8r/d/N/lPQthRi3BLAVdUk5IJOzFhPn9TbvFHRg2TlJVioicjq4cXPLRBuhLx+W
V8vEI+ISowaae/uqi3mfohGs/Ylr5iCYsHDSRDU6E53YEYVW8aSd0CZjI4KP6umDoirx3MBf35fN
D5hT6CEMzzgixTyqAU9elwtlTOps745qSX2JMSLvRHVevHNlvI9MgEuy24fRSkmLvQOif3Tqs9jw
Oxy0U3XOzVtk5JClqFWyaLMs+eV6gQMw46oPE5y/Ey/WSLB4QHwO/N0DbCVNXjVc0poErssM/jI2
DS4dPU79krgv8kMZnL53GiZEskay7HTqZM16eGzUk/Dye9xWXh6dS/uLp0s5teGDBSSFJP6LjTy8
oAp5x1N9RNr/mmsN+5lUgVk/7Qcsg46fmp18E5XCqCYom+sDWy/j5rmxkO1SCHwHkJRUa3ZEsR9f
dcc1DLD9fw1dk3IMtCoFlMlr50P1zYYGtHC/RokYXBRnn0ye/C21nnyooELeCliirbzZ/1uC3fej
66TycJYoNui2nAXr1I6rpvZP0r61+Ge8Aj+3uAXP8tfeD8qu496go9DVpNlRdU4Q/R20Fa+VHsBS
lb17obYu/UBCtH5soJi2y1XOulPBf4TtC1mw+ausqpAaoZNYSDv1U6ITORQgDJ/9Q8zMSxVDlKZm
RO85ohFGe0a1EtlaG05Nq7Bs7z8EE442AgFzpURc6riIHc2J42YL7BJ/vIxuqRqnJHDGA9s7XZmf
ssusmHzO7TH4pn8QGu4+v02VAQC9AEHuu1yGB9TnZLLh0GNrthGfzJixYNzfwOtRj8tjQv6EhWe6
ryGgV4ux6Be3ueAIjcqWCx0qYYFtnnJNUtDRXYxP47I1Ex2r5FwBlvrdDe09Zw6viDlKz396qTW3
jtsnht2LwwCHxwWinW1KnJ5ol9m/sQ1Lj0gR38fCtzFEWyya1hhhROCJhXgrDqdu380OomA3eiQC
BXleK+g2hPgtJtZSUag7ZA4mpKTFK8PnexdzO6TCBk1JvyyhlFcmlgZB0wnkVtT8zP5EKhFfIg/9
Oy2xBD5+bUcucEpmy+sKghkjY8rily8MIOG+3DDfOfyJNuNzN+MoMQ4iZ5wo4BgoVR5tlVNMRC+y
nmkyQ1BcwUGmj4fUR988zE8DEJGu3PGrSNlcEKXe8D+Id39cPnVPia9UUmKG3+fzjFi2M1YNivVO
xa3jPNiOcMpzx3W1roLCkKtzxvcJDd7NBYPAB6WG7ol+r8sgcAcqKNXCuGzTAKi2u/BwjL1KgDnA
bwGGu2aO7IBNk76ocFzzSos4DKGM/4gg3pdC7GeGZCP4C5TwBxb9Wwa91RaOZx4Fh7auJBkhp2SK
2Jh+I4jZEeUeAO3niCDjtvcXG8sWQTANVhSPZQRnJFg6/18gpKbC8H2qDL5B1l7atBJpsYTxSszR
+lXIMsxriFdTeHs2q99gr/oG9WeQhpMKrfI+aqVxgw+puu0TOVz7c4n9IlwF3fgKnIK4eIc5gX8s
MjZH+unSWxahOgqspLTZhWD+hXE4GuNS7fF1efuY2EGZsHRUtveXGfveWNQBSG5OE0jYFgqxSTF4
eMg4Soy0sZsXpp0jw9cd5yyCXADJ0aFHIPRxJb2OoioZLFADdx5cUOeV93uvlPXUDA66NWzEwxnA
nSTOpE9zY5WAhGgowbp4L+VRbOYDVZWHzHOn3ZPDl8RUZ0a4ew1fxfQ2VXzlWny89Khjp0PzCQiW
1DkEP7Qc66cv3DeF0r4/xhdX8Hmhd06Oma8Xuq3LM7bRLals7PJu9gLa81VyZeY2WFWH6IhlsrtW
6hqAaOJvPYFgbfDVotlskZ7vIjJl+b9rC3vkMvoFtYH5JU5chlnL7hYQ40H3VarKi7uDzvWJEg+f
XY5qIU3M1fIA9BQbY0IV9EneVy3PlPJFxMssqnGZv1CpaBje8qs/02L6BRvYjbPJPzix0D3uRMRm
fgHYgLy7Bbjbw8Xe+jY65jkxEt3nkvAAZVJUCCLKOCKMIL7r0d2JZoJ/fhScjRjjkwnbEitfxFp+
ei3IY0kxan/jMo9ugCr0/zY6wrP/3wEqeOg8SH5wUqn6IhsAUk/oWo1iusdhmCW8OaktO0RYmjVE
zgXXet9CBbs8PUZ4TwsA1wbl1kE+AEguXsHq3DPUFV3QmevxfntZgi+hNvggrx1IHILFJljJjMVa
zwWggVkp54dqDMkIE33rpRivQQCrhVGX94UQXjmcAeY/3PfnG9r0noi+SnYrIcNCxk2ynDj1Sa+y
jOoSjs2pyQvwxL0dpMWT6kaEhfbnjA5E42awmTfI6l2QyJAFHoNqxqSlnEqbAD59QIfbwwT7YKmw
PUQulNLl2Q910RiNLbZOGE2onCHjAKdQcjqIkmaCrYPB1OYhIBmvJwRg6CeDp6WzFARXViTc14B/
3f5MEOXIffYjHG64CcILdLzwaRqGlnO3Y24odPXxgp6XxoOrLzfieOydpXalasJ/feyJbqh99xlZ
0lZehsjzb+/7eco+GajtxOJDvXBAKNiCquCSc2rk4ZyyxSqIbzOWW9XZXKBn2I+noUj5JutaV1WA
gkUl2PACx9k8bvl4WsMvWKw854gQqYFNl3AfhJbQysGqg8CROfR1J+Is1ODePBvsGvAiFlxNwgVy
KoOfgRpR3f3yrdxuksfVswoJ4UUSOqBedSosD2ZN8ACbcQvWeDvQGiV2sKcS8nIrudm8sTn4imjJ
EAVmq6fR5ETCbA3Al497ePDDgRZ8cGElTfuG+/y1P+9UwmIqFqnxwk2Mx9JYlz0pc7aY+8S7hJCH
pNbzf+osrO/xf3N3FmNJ3NaryPYj7IJdyRPG+Y188h1xtYWRhYDUbr0YptYGuaGVCTiLP2+xWnCT
pC1BReX8zPIm1p2ghjGZA1jHFEVFQvm3i6J3+FBvGA69MDmfpJOzUcf+ppGaWE7uhIHONzE9F9I6
gJH36O9MNOkTALTaw8U/tQHdHVG/NkbqN9EqubbW9KuFLyR+7kR2wRwgW5bV6ajEcnefFIeqULfK
EhqH2y/br5AAIYl/fjDmhJI6bQmeSVIh3QWjzBVyeR7iBlBZo28GbzKuoOvauMNE+lYwWuTSUJ6t
QICzmoT779ZXGUQLLVlMQYTC2MnW3EqQPa2s21iNk8uW4H86tfMGH7yil7ubcxc9mk6fCEWPBL5A
lUUaPfTbPf4Nl2WIi1J03m75DDBtW5NMd7NrwK2+q1AvP15yx/KU1vRyXj8OUosal48hmqAFJa6q
iLEA8aR7yJvAZ5yyE6qjU0CpeA1Oeu1pSLGraWu5r3SVxixHm39UNos5OY+2VYGsMqnec9gL/cbb
KENT6wHlSq6bE1PyDSc7MFgZnaIuBhUlmYh4ZX97jf7g62xhxhkkwLxyxn3rvn8vbhpoZWdMXHxz
+WPFdbmdR1NyunQRKNT5O+oVwObs2iibAb+dFZuvwyN6rueqJhPxdpVRKcrluBJQ7UgsO64zW4R6
7XvfDcDjVJRDYPbT16ClxZK6ewbYo5pVGRCP5hFmimqX+/zW4abtqlglYAsm86aVkNg1Gk2nMp77
HJYI9mkZORx25zIovLLk29L4huXM691SLAtE3YJq3fq7Gidrrbh0YTM1ABs03pPAq6nBsbm5qtFh
L2ResuqeDyisu4yRtJZsQJbGW8XhyhKbMCdNinXFaRxXb4dqht6l+R+QLIMIZcXW3bENJBp2cHI3
qiydVQK38aFEKDEjQV8BGyOp01dHsHC4EYtLVTEhxMRPmMqYwcdBabyrqtG527eMGJFxT3+Dv6Yi
regOSbT4IFxsqhIGuUA8tXtnzXoXOA8UnRZ/Rn96oG6LTfjmrL8u6yPiTuoV3NJ5MCDMeJSbfyRc
NZrSiPs25IqgTDO7phW5Ey3S6tKQVvIOKXyzbedjeu/4X4ZZrpGC6te9buqZyVmMLyKiNfIzbS1G
yUxgK499GLZZOwAvVCkc4wHh+9gOdYFY8UivyL729kVTqjfIDUg/snxWx1GT68bVu0Uh+s5FJDDv
2pmiekFFF1xDkoAzvElJcvXJlUY99XDsSUGu62VT1lN4Xsc1Hxy/FoLkdOJqgTb8EHGQYFLTgDXg
DGJ1xrXwOwD+EndoTaRd/Kry30aPBICaJpFOIt7NrWu3q/MrdRxXJeUteOKvLwDYSs4+cw6wy2L2
9XLeG6SJirc+zjD4yey/qWHvn5YAPPVbCVTxL8puV4gVE7enNFxsEEL3EUcbyzLJxatrgARy//3y
AndOKARB4XZZngQgyU+ArvLrS/oNMZ2nJFfWPONd4tjBx1uyOUHoIrqSSEMkDTC2L42t9Jng5GtL
TrGY46lYVW8Lq2akEDuyJ9Jd6N9JwWVjZbd18NxcLzqucy5HWj2koyf2263gqbnBbOWwYnmiAflj
gfOBnUKPGMOqMdLwD5C6pu9mWa1+7ljKaoBA+td2t3kyIIjVQUpCDzv/DdKKRDVlj8H7m60vNXfV
OtEuE3uerILMPDsm6dKnqIPnqNaI5lMQyGH43iPynTYAJPT7nipY4S/218aEbb9Sj3iooGRjDF4Y
v++4kWiv7+UmyP32NMOFuDEk2phoHLufwmHo7aryGntD5Cd5qQxXfkIqLAwE4xIRMod1S7kCh8aF
sNhLUpFpIRJ3t19klpOGYMAm/rWA0awo89h28CSaMDDAy0tewHKekE3L2xGRO42qf7jvVGdvaZSs
aVkcjFNgwlNzzQ4Ru3tsT0MBgQ2gXfSyo1P8zO/VdpkkM9U0Yo+fkmwrWCyiobHCQonh+7D2oUU4
ZxiebGqDBFypoDPhO/jgJXMubybdn/ZU2Bryv5Lb+WiXoefaAw9RxdUgjOvC9S4nf/QCxiG4JrP3
bkPf3bk2bb7M5dzviHCq3fBJPzQ/2cHh3MP0AfTz76MrGExrocYqvQHaWhxLFHhbSZeGMCXXjLPo
mr3GkVRzuvNp4xqGAoAIb/Lg9/2LE0WR2+ii0MHZQzBGNcSP7A4bQJNFW3I/jMeMjwMNWnKKww9b
x2YgWKS3DjhUBorxfSsg0Jj42a0vIk/J6ZOdZn1+IaO0RmoCc2MPPb32UeQhZycWAgNcm/w749kK
9vhUmeabycd1RnLI8juvnq+sdu/rNTXJ3TcguuwNS3ao8wag52uCEc6hPKFGBA93gl2zQrMq/EmO
3ieVN4A72QzVYvnBzEZ7A7Zz5vh22dbzROFtykZDlTSPWRLm7QoALGofCEdrc2zmcAndbbpa1U5J
L8wiunhlI9tR6xAGgljZCEyBhWkX4jDKU7NJlbRxyZ6n/gUIOwTAKSH/3isdiFhDkEai9zu/69fS
5ZSdcsxG0DqAN6+J5yUU8lUSkhiSaPnFFMyCOGvqMZmmtQvGqXJ63zSxMG7ocTlEM03aCfNGCy/y
2oajHI/cFwOXGx2OTSNe7rwmTM4/HFGg+emSXr0eV88w0JtbsHu0Wmiq+UK5hnjRcLMtAhSnThZt
MAlerasGeSdBzRKnyfGtTDyLURCYCT6VU35n7kg/xJ6RKD8N3WSdlVwMomyQGw8zmKYfoJRlV4Da
ItAcdpmDvZOdTRED7Jxvd9fBeEt17PsbdgGGG/ikzL+da4zGsSy1s2S85n9gdRpug4dIG+Uq3BeU
+dTuC+WXOpOCA6xX5wEpAQetyl7xfGcdEoMWJqIzREyXAs/0kxTOv+MR4x/PsCWY2aRxTIxDFZRa
2/vf+xwIk02Q0DQ/275PdPcu3SWgiuZmLV+J0vhkaKP8PE2tMUv5vUPDGsjnCslun7Afu4Qv0h+0
iSemhl2xLxYvvAVyYRiU6dU4oRLVHBc0vFfTtM/UBAf1GAyCqjtbJX9C8CHhrO0PIrX56npeoU3L
cxr7dWiC/H60cu12mGI/25Fkwk+ccT//aZWj/liUH5Y/N2Ixa35O/TIJTp15tjGrZ5YWKIgWsFaV
HyuJW1+MGuxt9vpnXQU/J4Y8On379hEBArhzTGOGSmcR/DMn6L5p+jfTPmyqXZUClIWnewrVRCPJ
SnWULhwGFxuUkEJE+Lc32cjxCgzitOnjMGyiCXBSVjFPUC2xVE2fraZXQbt9Qzd6Oe14U65W89rl
gZd40B+pTvaFxIqAx6MyCXNfhs+B0VrUb+G3um7wN5MwNUHPZtAAiRtblRFjCAYSnhMT5VocWV6n
pWYFysVGiyAJQwShVXI641dMzCy+5Rv7XRadC8U+7HbNwUq5C76/MKhxytPV52UKziwfs93mTha3
3/ypTzX44k/d3HpGTHHA7C+qMT/Hb5KAEaMtQhTmF7kY0GA19Qlaxc9ScVBomFfH+f7oj75H5InU
xjTa9ykuqmkllkMyRdf2AKtFMqlV36YfR0Tw32bLSzdukf3EmHrlHpcKkIANHXo/Nlp4tDEYmnXc
zdBPZIE+T+Wtor+b2Q+YLJCvkEDzdb2p021GaYztuBC/pBYi2PFdHfmB4O6uQQorIyftzimbVneU
sggWChpsAb9IUn1LDElFLtaphlHglqawrdSYrhCCuZpQDVhcbjxHWmKo/thzzpr/SVRa0tMbQQa3
/R9f90aa685JM6z1w7o8Zb+i4vmyIz6FouS9l0Pci5ILgOKOcFEqu3JDIt55xSb+q/z9XnWregov
G/6Vat8Dg3H1mEGYTN00c0qWFSyknY873cPG2mH6EiARXo29fBi2K16rZtqHzLWMuFJht5eLcxAc
vL1s99j2ym6GLN05pM89HbkDHFzPgjmly6EwJ3heXv+sEiASEDyFCfVHXF/q/5ZFVQxo9eV4v7Fw
MSPXUZzghYFOERSHTzongpOpjNLxxUcMlFpCYRpab5baLXNGZO0TENAnhE4wQ6mJovsbro9dOuVP
cbuSm2Fi/8xTKyZgrU1WMMg/3BFFqwJx+yzOaQW+fWGkLnU/OTL1lWnD3lRdDO6oOkkEq7VIYbCB
AUpNmNFyROMCuB4uBlrsx8kvEQQrIolMhWQ06jeXmKFQQ7nfiRnVlRLq2/5QjHXuCSQAVaLlD19/
7ZY/rvR2xQHjYbZFAC3YAwoo4rHDcPMq3LqDkpqvB1NeHiYIZ7MpHz1cR2kXIEOAp2sXUPchHs2b
K44zqGo27xdHmc4xB0XXBiBtnwztRMeUwCP/IbwGW866IiOhYuw/FYS3qfhrphGbEYQumwXFtEyk
kdSwMToao6QoCZQyKk2fYseR3sUqnGamEeWtzB6fcUL/12NB4cBzYCPQgZQQzBfutH5FnpuSm5kJ
Kh/iy8tDFI9+XZpfrj9gDRyPe2iV1QG1NZKSfzkXKtf2mwSwtFLbQt1WeLTwL4Wxqbm3jmOxRS1v
PB3isNBZttrokD0ayiVKDsL7XF8Tbvf4q2pFSxNNxDkp+AkQOqqbIC3dswM2hg6VT52CxFzakkvp
k9kWvg8GNDVMHuIDdWUGyxoE7yAp+AyagAfPxM2/mxVtc2nJg9owOS9y8vZq/r++piz4kYHxbvdd
pIldMgNT+fmd99FtHpETTV/UDoaNTvq7agGwv+AYefPu0tHSpPU6Ecxs3ecoaN5o/HrKGre1Ir3o
KjGWSj2IgHi9fhbzzulgchNrQxWathTFKq+tPYgHm6Zsa0ZGQXh/jJJGyTGY0GbzKQYxbwpmlwvt
Sdpz7ek+mscLoNQdIYA84HjmNyz076nOX7R3WlmqS1IwIXrvNT7O4J3OOEkF+Wt9lRwhIQkoqAKm
N+J4c4gsvUGxG/oAuCOsCv2X1l4Ha66N1mGopmXBALYx65rXPMz/Y2tR/Ybq+kkxbnIA+AdxHl1w
3/mIQbfNKU/SmCAYQyx4S9dYgm5GFmat4vFmSR9WQ4FPU/e27zBt1S69vuqH++61Dg9mzpUXU5I9
GFHUJYOTsmgennSxgW66gz7l2waklq9azjEekHYrg7PBrOjiHUHNE0mPGGXaLOa190mHmpIJeDrq
ez3HzLb2FLbIefOqvczZ5uSLpx+3uEUXLur5XuqmCA2OpOESEb/MYFeCNzoaaYmA7nXq31pOpYoU
cJ6HiMasNYW34KJ3u6f86PMfU1x7IG6WYRrCH9/Gd0WS1Ff0boqnEOKYT0H7LNQOJx3a/qlY/CY/
3zGgGbHIiTpLpmAkxEDb1dEfO7IshTcWjyPC4nuLXBw8jqreDTDUVgpnFuE37Pi9h+bYrSl7lY2z
Opww+oisANPngBAdUHiG1rk28/viyspwUbrF2+C0LeT1ebPlEnb2+VR21ceyKzh92tLM5ofrWlSX
SfRpd91bAd7n4PMwVsMlAPuP9mtjMRy2N8qbR6CdwUgFE5uqjzOzSuz1QNdHy3Q1Iu+q9fcsyA9m
GuprXXU5Vo88PUYSIu7GnAYFODxt9lUAOhJDjXyfbMJSQqehyuXYDVWWRa3xMNXZbffMrhmkf4UR
Y5vcnL3HR+3hdDmpEYnPiUfC87TC9AxEr27VFBhz5Cn+cjthRy3eIZHtazlxlHPbii9dFksM9/kr
zr0lPxxkwmET1bN4z2DwaiPTQATecCcPG/bCyLn1Sps0/REfPFkVymJ2TqpRjDvOTeAyjoLmSfMo
/rhvcHKEDO5Q6sWYG96KdsVjuKn82WmqFhC9pQa+HGKDwK+Ehqcf95Lwh/L0IHEBtrevL2YrIeUQ
YpPDwYHhB7DsnJbk4v6A3zVQpD+qLE8BK48Ol08Bsbr28Y7TcxEeZEnMsCFFY6k+jnO5BTUDHcXV
sBF800wwVapidfxy2TwvPKbusH5CiM9akv7OgrThnoOvWqlbbh4L2bW+MfKoX7OsdayTmQSdexF7
hOOFwiKM1jjuL3ysbmoHx9xRcTfgbyOUFWIb4zu07WjqZ28M06zU2/+SDbm5JebnDYFY4nymyELn
ntuVNvkY2ORv6XjYCzB4lmWGJbeR4ZlHkZ1uRCJjIf+GgOsE0z5m4a3qJnxLA7IfgwNS8ETjuAK+
ibjDANBNC8q77JgHzB5yqNVuiwDlz3X/ilgasGaW39AC0QGedxUMtuO5juqIkIPzlIjJaN9ukmma
HlPWxbQVwZHcJWhdbGsPvbcUClQdnHFgBKqx12jP1B4PWzRBDmsQ9rsWVeKiTtVHif1idl8VwZzK
VLL2xDNZrxGheVrMg8P4pLDz/RMzqa+gCwPF3UHSVlBwNAqwt+ex4seYZqd//jCRfPPV24EhEgNy
D7/cJY8EeojvFZ9RRInZAScsLkEtgeEcXh7Y8Ywp1WsAJYcU5SiJzJA+lE4f0hToPEMcVubfzr6n
b91i3m8TPcyfub+hlKVqt/FE5/tfUr4I3ymPgthbIVOjyW0kXLDbroxkXUk/UzdDRVhFJFC/oscR
nZ3jdPu6oK9uaX9xnup/AGytO5/gRqw+GqWsyUZxEIDS88OLJu9+ofbUvqzgseKPaVIdFeceVKxS
e0IN6fXKA2+pneyutRYa2pv5DOMSxAeURdJluyiUnNopyJkGl+oSCWoHK1M7fvzJn6tpFaFEh/3v
UoCsjO4ZaoFqJY0HcNFyA/T407iSAS/ZWxCm0IHxaLK5aIwKmZImsiXTUA9VEkmFbAOXbbilLpEN
DVvvLwO6MZQgldT1j91IQbDTtmTj+7Qj+ZvlyIhQpn5fNiiE/oXDpEWVYvFf0Ml5zOws1+wDJ+Vm
ozj8I4ojCykJ+VN9ELd8nsotvOssWgtlqmfZ+t0q5HNl9EqsZn81thT+KYRC6Z2Kq2twVzeJR8mL
6zexjgIqVW/JV3pVB5LyItqGMjgV/RMMDp4UU5hW3Cg8tMaEMjafz/j5SSbvTzWGGVVlPOrEEa5U
9I1vSv/Da9A7sODNp2qm4iPtSyPZ+vaXTd/0XqwWhM/hZU4mxoeZSo0ZXK44a5clSEVOqCPZCAEh
Cu2S3OVRwEuLh4Sd9DSBzferTKoIf5jqLcgMRdy2Xy8EMyOo9z5Gy25GIkPXnOEKirojMcLJuo0x
69g3IjzTX2rVG2g76w3C4uODKdtxU/boocD26JnP3l57pugVIhrDcNnWFmLMlIp9x4UYdapSpzJT
tc7UsD8b2zOEzzysZ6cd29e4ZHccT1S2dBXVguD5NiqVo5l2JpVeiFfDkpAwUWOMsBrTpK3jDafO
pwBNsOG0vrIAIDylZl8aXg1v8BUwvzrLkWJQKKRvQ+c0n3nz4z7kodfMZDXSfDo71wi7eAkMyRJU
VSDiYnKTEX5rWu3VNzHfjew5QEKesIGCTJX3M8Ml4RZmf2r0g1uh7aYFH6BJ+wgtgao4+cV0rM9B
1UyeC+mPlWn9RDGGv/72Z2flQgeoBl2ZffHRYueSzGTWqxeBG30l2H1K8RbBoe4LMb/b6GNNJXjF
NL+GSWCqrab/XSR3kWFa6tTPrv/g/Pktktw9gvb8sgi5sP9m99ZQSyBqpPtrREIc0K29i0h8IeL6
vSc1Gk/B1IewSTQIZloDaUmx67S5Yv8ub3/IwcghIFiDuRszW9znvfiEcdXAImwMTKcopuQie2dq
VZtaaA+WzYtaYmWPztb07mvEjL6Uv762FrMfzqiW7AnlBxtvoi/JzHPix1miNacR5AhmeA/yfeHT
aIOMjlPSJHJVKGURR2MqQBCkeNR1/wQn20aUKoh7XdQrg+LqDintPeubHnCTHPZVP/16KycY1Aix
duNbTB1ZiLMHN8AQ9xsWmQ/i9lESqSeHdPlYoPu/widJMoktoZVFEQttBm7ll8CstkvXEq4pnsgY
oa32k5dTJefhteQAYEARSMqNqUoypmvNvrRY8h63eOh+t1ya1yNvsfPowvps8oskwOS9nFG8J2my
vxtrE1DMrx8WJdmVLrn2MRnEuBF/h6/RU8O3FJTeLvZomx+ukmFAha0fY4U548NJeBU1Jmvrwf3j
CRyGmsn+NWD5xYdf2aZanW61SFaW7XW0j9rYS42UHGFfSqXcHKRmlZ951fp2NrCaZDOiQ35yaFcP
Yj8VSe8cLGLaffYkpz2LCyYctRvzsozMOA1veZTxhKsDRtVoyIXVzNtFx+6QbQIPWRPvQoaipFEf
dew3RmvYyCPnOzXjsOVOWdpC0hZTHe7OhSqNCQdB3In5R5EWHy4wHIm5u2cDfyMwRR1Ris+tIVg0
SuBHvJwTJtFR28haf8cUmqItWR4IqG8bHeuV/PIdnckCdMDU1R7v0s6edY0fAO2I5I4le5UHAspz
bDZKeCT1rs3KoDEzkUYxspkTTt7EKrmMAjzhyOx/kiZse9grWBlGSexYb4yjy0aOG7ekWlUei0WK
ydkMOCAOn2GQwo/a9RPoUdAZzWJRZxLZYBOeu9MOUWQ0FoB3OfoskVFQj+yKWpB4IbAB9z+jnUsh
Up+qhcLQzPupzIzJczbeI8gCGCmV4IJhG+gYW8A/m9JFTLUMA8yiG43dB/IqdaRrXisJq4yDvb24
mGl3qYiZyNfik6rt/aQkl353iSn9bdBNkh7In1YZ/33vI4OM7ZaVzEgU804EWQAwQMkSJ+1JhcER
GhuSUNpZsV89r0uDq+TBrcTKqNUwV5IY45HmGL68+9yhzqjUcE6IFqTsm6W5NORoohR9HdOcQ+51
xqxjHdFleljaC+H+v7ojuMe6hqkdVFICd++AGmba21YGi4ko2fS7+TGBNG3o1PWOGT8xbQTPy9k5
xXBDE8wo1WyMvu5l6ZEC/lQewiMAI6oBGCBvofIHljhfaZ1vhsWMyYDnP5xm7b5AlRYR9J3Esg4/
+I+JdBiU1+wchNLHCJAOOhIpWAK0YMRLTLAht5UxGpggSTAJAB/QbQOY52rL7mJ38bHWoxScTV3K
y/T5nQ7akZh99Ye98n1MsHt122TRzCnu6AARUoueAU8Xj2eSO8ia9/zROAe81aYo++xVzgGeG8X9
sXY3kx9Ra/kklx36WlRbcDlu3GfSLG8HPSJHTANgI3ltn5BVe/eeaQdZahU0gASokZJRuxh/iQCg
4iQz3RW0y3gt8M1UsqArUBAiGxfQ13LkIUIrk/9yHXnLvNbe5ZXUXP069nsiEyU+0SnYAgPqE48W
Ems5lyUoa22jJ4B6Jf2nGz+7uafGqQ39fHWIZXQgx7eE9+0QF2P4Cz8HSpnnmUUWAsxz/FeZ6YQB
y6LekmVffiHCBmMWd1QKkWebaEDiRdlqf9aaxo5upWSu6vjw8vBKW/xdxeoZdpnh3KpQN9QYu/bN
DAjhZQk8TX09shZlWYxFgXa5xs26rwp32hRfDAJqvY+QRNtwSpdMPP/tBTMxOTnY6zf0FZT69mCv
UVRGsPellc75WazLQkXz/EO8USGcwKPkDppBWNowo1ZFiJHK/szSxaaG22qKozIYwFHNpsaWsX9X
pV+4ayAREQQFwvAa+EjyvSAhPUDRDb0J6oejrAL/tuuv5+7qz/yt/k0n4DQGM8yIpQ9mhtWTffqn
m346bK3LxDqMcrb4kC1QbMkbSjtaKzgn2PxAT8PMPYOm3kJjB94aNtrGXPw7F91GT86R+TBDP0tG
J6UHhyYbdVcv3nHdP6yAtBLRUj5318l+88jX2PDhTBzow8TW3QPkuSG7m+scbFIVxL9ljEEnNvOB
nQGik4cY158DdfY70g6HJ/ljwnQzzf3wenDo81SBrjbGD5qmMKLjlcrQj+MoHyqlyS3pe+cG+TsY
dgCCBVoI7h50YaIaCMeZxA6Z8DKefSR+MVAyIBbno2748WEiarAhHbdWJPftFSrvbZri5ClpNUKq
8S/fRwj4mRmp8PiXwhw75jXokBZ+dHId2cy1bueN3pNJmF9bHaSHMxX11rXz7KB5QtzjpKuk5VXT
u79YiMyGkmYyP7zY7ErzPWdzZqBxSLp1FWnpTMWIOOzCTVY6I5xQIj6thmbsaVreqTBovHqOZ65B
NgN9kfX/jbl28RxqSJCT5MNt3M8xi0qpXepqSP8vpom9A7ChBZYmzULbZIIUUaWUvcCVMehjKaFq
dQZNEtzq4Sx7ue/kmxNMqsPnrp305/Ad3ybWuXPR3sU+5vgFvjF1nxJeSaebKy6kUK7MEKWgrPKZ
O9vRW1xCuqoPZwKlc3js/mVbXdcxxOdPLv2coBcFMV+HZfTAmeTQZn6M7uQHNnA1IDF4qTteDZbq
gCCf/tPsxtFGuQfKemLPu6nSbO9b8ksrXenZc8qbibngWMiM1TCMkWx+uKSYt+uT+s2WUuf+ZAG3
0EEZBgDpFHS38uzeCJncx00n8/xIyMR7xTntK1b8msFHf/d1beykcy6sDYu4tOLgSNGWbl/M3jwS
Y+pAS0y37B1pyujtBOLSI8sfAtGGN2z9MbB9aSzlhFFvX57ZtCvI4Ao7PLSy+NtLx+W7YPVp8FRw
y/A6EZxDfn5NhwEyxMAXJ3rsAyc4knqOaONVCXOvEQ/nU5g79VINJU1iQZzT2nAP7+sWGJH47KRF
tWsol5TgNY6XwcGOMPIF/hsRraefeY8mhC2uJAl4sf39nhz8krv0+vL1uXVmetCyWH2xnPqjKln5
VN8Xnl084qGQq2PCH4VFAc9N4zmOtTgNBGHZOKoJDOOVpCIVtBZSNQUJnydwTekY1epEHhgZlsGr
qhXosuLyDKGAvLdrs+RBLr35qNQ3Gvx+wj8XvA5ObeggoYrH1bYvjp+g0nMr0QGJF2nWfO9yvdaD
6ziSM+BheNcbc4iC2wsx101pzGAd7/Fm4tMfICNo2P51tae24m1kiL1kR0oxOjuSTavZdwvWGRLJ
joxuJd0B5hs2PSTb/kvxXwAjCWFCvUtKcG87BC+mNpB1fyGNRRaz5stV5WhRVmlFkTvHj0vFnSQf
S+Xth6nP9t7NanpfEijPzHndKUvktHhEjbcOVlzKelHp2KLSzTlhfGzageWCmwhe2oCDZ+P1wcMV
Up/jA73tDf2I1ndmlLeBKk5AgXgPAwVWM9QWrIi5woWAb/2mfVKqKJMsJbZHRHbiexh9NOy1Gl8V
2l0h/JdDKcsogdMktZxkOe7+hRIl1wa5qjH94wRAcAft0eCzv40fMkQLh28aAJAX616cE+PStKvd
NsUhZXkS0fnjLh3L8RFeqJyXrOB5fXwHIP9YuTa1I3WEqvkPpsFvBoWtUbgev4GSHPlK/GobjqbG
E3RafssgifOnLxvmc3Yet4+yEuvAb9VnHwjO+jnzoFxDilFi6W9TgfNCmlnBRdYdt5yATUS6T45Z
sYu0kGhzQpGOOeX0mHeNNS7yN9y8l6aXYd/uOYhpqWtdQj5UeNlzCrNyuN+iOQn3zhqJa9AvSQaK
fE6rBQdU+4WzpgDii7l/CKzKwwtZ34AHeRtL3+7KRQo4O1PCJL66F9fksBOiHty0Qm+cC5nLBtBm
3LCeE9SNUl00NHwLelGC4G59nmR60v4gXxbEVLSseSLFDvKAqAxzY7JjkvV3wo7GmkZx22XtQ+6u
DNUJCEbsZTouR/penQVql5gz2CsZi3CLKgADN9KWBrSgRy2O70kweZech9XVd8bnuL86tPhd920D
LX1hrAu0REd0a7/ZQIW24ClrFaINLkjzUuicbUviO4u3XuEz9cbDrVnG2L5TkDoJ5xhUe5VepmNZ
8TKKhkFq1Wr+v70ZyonoKYk+RLtOSnpDgM1iujuUSFpWnasXx/UbBz6OOK+M27bFanR1S7YoIVRK
3l/lB0mr3YgAyXC5+Wk4Q/1zCHfqe/GkUsTbf2lKeeb7SjYP35enVZPoNmOBSAN9etS8ujTHQAh0
CK8IWWp3u3DmwCYKtMqYHKuY1arIH4qFvMniWOqzLokvpx0TalaRawUXdW6GqpYZuKTMIeUE2Qc3
0xsdm4BVCLGAloETlQDaFFjZPFH9gyNDDniBy7KHpjFT1iFfCG2dKUQ/F4M4lwkXUU32UzsfBul3
JEVgLe41SYOfCwaDOuNlDbHI/ywb7H+1prWOs494Lq2ofoM+eoqbv/shldkDhE0NaUdTya5t7q3W
X1ACZA0+iJswn1Y/Xyb4scIrCNrwhGhsEZCnDQoG7lFi1Lhpxu0+q6SR3pfBZGUhZSIZ7yM/fCQs
YZIQ2xLizU/2CE1QP4cZAt3f3aD93f7U5To8YgkzMvRIlW/EmHTI0T8zAbQzizfrI0zOOdaoImmb
yCDZAk9uz8uv2TOI2gtTML/wNKKpAmkdTKwv4ufgXTK/yaBb6LbpYR59YgWLQS03JiQTkA6Y+eGF
piJLyJdX9Ut7eDbnJUDKPLrkQ4XT4s/uMsz8i232ecIX1caQ65fQBn+btijVz/EP0WWoA+MjJHAy
gpPmiWKkFRTj7wA7bZg9raIUIu8c9hp3DbIgYAHL6uVtPaUshTPTLwyTUsWhqfPmcKMCb1AS3vkj
14eqmpHmefGmNa8pi2HNMSqTxxiFDow1oKp2dclUlBqVIgTwoBw+Y5xghOReJfHGILH6evE/H+Gl
NneOI7xImeCh0yXK0U4gsZqwBWsSxwT7mptMnkB4aSjiFTbSR358PZChhCjBVnbAR1SRpylRnRJA
R0lQn5zJ/MOieTGvTPr2D5TfIkLxBmg/lNPo/5l/dwuAmoqanUR2CaloyczxqApBkH1iTBg+hzkJ
CMqyvukozNoDq1uKw+NLIIJKg945NDcrMCV+70cAfM64V1whtUHvUhQzEVp0Z/CcrBH2o80Kt/++
ZNYibgaOHOpR+aVduQqudNHjE4rypvT3EsTXFZKhscUqZSxRutoX5r8mjbHbVxMkB6qrvkztlFcB
8jOPWM36JIHZ3IDO8qZdrYCTewIZx6cYxQ418HVv3YjeDciMVYA1hIoUkY5NmBOvj6Yd7DA0AaOO
7EQVoINwVpwkOrhwzU2BbJdM8m6xhHYjmUESFW8kmNHxFbwiWo7dlnrumunUWG/Ao3OK892zcTVe
msCSw3+sFYcWWjWOI5Z47tVihxS13zBXCh9FbZ70ru1dzDpfKvPhjB6aW0IT6aZZQYnv7Vpip/90
1jedK16ZK4uHJftViBIlW2cUW7FLhUxUz/HCcOWFNz5Av3fx9Oq7NUFl9fnVoJzZh0p/L879BJmn
9wPZzfUqZ0dPG9xzF57zB+70jvKTy26q33QfoUa7CWNIeP+3WQSTQO+NPJwTTUxberWiF/Xg3UEf
eGtE6DFcsOekbsVyMKzP6PE95vnv29zDKCteGV5JrmPCBQ6o7+xq3S/ONeieEcrzOCG6LWddCK/v
TYmOw4E2w1jWGS0CRU65ip0AVc3XrjyfioYUBob6hEqAhigfwXrBtdwuNythjQ9yWzZlJovgjO9W
15webB9/gDGogdTsQ/sxi776NKsDXJH1EQu50V39QkTgSso8EtUm+ydC3D4hIlj8VN5vfKoYI369
KcF9alfzsEeXUWcvPADcBNquCX1yRxznNU3Jyz1egY90bGFZsmIB2u98l0A54SoH5S1UIEUESMR2
+R5Cf9/coztgouFSYGgYbETG97ceBP6xzS8UkBXryvbL7DjWEB2TIHtN18hHsQGP9P+sIPGu86H3
ua7Ak4k57ufwJPOHKMmpsZBhFeoWWWGdITOzMcWe5BROgqWrH0lqdqopp2EJk7ZPELmg8RYA9f8D
ppeYigWx8/6k8XwRwWyKzeyGds1H4Ri5UT7jZZF2Dlfty1zSMhcdllvmUoHZsCZ4reYk85Wz+ESa
FFtVEwdvrXCSDMgV1Qm05NEUN4iUNpj5v6+zjn6iEr7bxpIbE1FUN+QWY2S1NoG/avEO1Aip6Z16
T9LsZsZmR8BzeOIygOo2MSP1MToqUzDPphN1s97Fdjx2cGyYv/pompTkPOigsg3ff1WuJotN3Jti
f4pP3sz6jE8okY5y6VrzVu2FRUA3OuPwZ/RmJg9NAte3M/Xs8d0xFtBRv6GvFg7+c5I2tOdvcyGU
rlVnNB1NT0ryPUc1R5Z8Bxcd3DfzXtJQmWIWNrTzVg0zbDabtn69VQZRJiOGnF8uLsFH4Unjrg+s
gS3xGrPk6mFcqmOCoxwinHxODDJt4QvTELezFWL/V6bhyzkFdw2EOQR6syX0+WKR31jY028oyBeO
BvMfS3pEdzx4hAABVog7lfxlEZ9M895Xy2X/dvJHXEbkjCj7L7K9j7ZtoOJAIwfGzpwTvGMvDrnd
YX8O6V6dKlqcnSDkIPuR5vlzVX5RsGLnywPv37y8Ex7Zknck3P/LSC49CA1P1pRLoBfB+nAZkykc
8KcU1kkqVwZFPGcg3XG2W+TsJiYyCPPHfvBXr0UTDa7iFEJAr2ar6o/v0pr2kjoIGo/Odqc78S6Q
9nQ2YeqMJtkUvuH4ndkQY3igBi+Gmqy750GLjY3+xo31CNc19aNzHRJ/LlQynus8Ixc6d6WQUHVo
NqvSYEl0sy5h6eFMDzSVpmoHE37LQ2eA2HLeHRDUplOpVMMQwBBGAR+KjwWEP4zGWdxQn6ENwRs2
0sst26TOXhNmm/HqBOeXYCvl+sAPkZhbLITJWZMA8aV3n/WTooX94zJxQtWbhSwrLUAHAY3Ir/oy
J8KgZHnjwwTpS8x7McFZxqSKb8FuTc7QcQ9jwDZU/BhWgGfoywaiqSl2GVoNtClZuWuUp0RHAaUp
GOfo9MzAj/6Yfl4h2pm5cEYC0K2rrSs7X10+CR2RZYKg3zEX0Rz6hSThOR5o47Sq0tvWEdFrIf9E
oN8TWk48DDlG/DJZHQY7TbtHcYTlO1NeLfTyiwTKCgGTCZEQrqr6a9NIDtyxhBejh84esX1ZXX/y
MmnTEM3xsE2HaBDLrBGYh8rCx0icphp0bqDrL3+swXHOFzKPOwaqDFm8ubTas9To6g+gqJR4imHS
zHKUZ1p26vcBjqNCKk6kPm3DYNI9Q8uIZpiEAnEbdeG8XCQ0lXVgGP2G6LSDGstCQpb1lIKsNPGK
FT7RSUe+AJFg8e2DVyJoXsZZhMjrXg63qiN80QAND9o8/AstXOqbNT/cjTXbLS8RoT30DQ2l/0Sx
LNK+84oftXuNE7GCfKMhJ+ibQE3uFxycNxvVcDHIfOa+rcP2m1w8fXJgulDXJ0siMHAn+SD+INp2
1q/Wcg2/GO2ynK2G1ymraThlHS3nU7KckGTBm8E+13RpnWe1ZERyjstozsN+4HhPLAy3wu28YjYB
kJBI/FYMxF7FC446/diH9KYc+BCCDxIS201s0It7BvJ+m+pklw5TVjLDkMijC6Wp4VotnJX24ZdR
7s8gpZEDd3wVafDUv1BRQgLwWg2mnpQI/PjuJb9UZmXGi7pfn8uLrIaE/7DbZeA43bV83DNFFZpy
orvIcl/8sScmnoP5vZ4TGfMW60G4LRDy+hjIMeRfB8wjCY+zx/+4OmoC30AuiuQOeCLZOICChCuP
dZNqfK1n0i4ZJnj3gTHu/8jDlxLeS7lWaVPuun6sDOAKVNHJiH7QBXzErGQPFQQ5JP50l+P7o9b7
Z8RC489V+eFPXeR1ASOIArAcVdgUykOOxETSKF2ZffNUwULIIVvEObEU6gPcSfy5uNR6mS0+Fyoo
6AgAAOBCJbr0EnNfl0qt/ZpMJw0HoZN5DMxjdipGOE59yH0MDZagWCy2+hkWEYjauD3bnISNW+a6
xSyVpj9ZH2XxfzyYVc/qGTjaDgM6sgrvrPz1maGk2mllJUXzaIixw5G54nbEFlYni5E8dWqCKp5X
elVxGmb6jQ6L5uQ+DAydcadMdmCG7JMoV78NUEYgRk2vpAdiN001FqataPLqIqg0gpU900YikeiA
hXI4ydv9Vow9usvUGt1uiFHnfJ/UgyrxKNjaaTrjuKNCeEWIBR5HpdvpCPorwKCzZCSgLchxIpYy
1oicEF+DkBVDGHndSbJttPVcu2WKmYxMbHMMQfg+hsOn+j9VCqEF36zRNMy5zVMyZcBpz8ezD1So
+SUAugK8TGnB0GGEiBd9nlyK/YCias7mVc4IwYQRGAb58pinU9TbAC0rR6K9pnK31Atn/0oBeU9l
73s2i/z8IqEb1luM6J6NlvftJVuDeIiZyVP6mqtDOta8j3v0ROqT9sotBW7gn8ZUbo2l+nPKhwv8
sPR28Dj/Wn54ERdi9mZYqvp31Z/m9rnIs4IIbquSKvU7QTCRqM5vb4J8pfx+mtX6D1b/8QbIsuSQ
PbU06I/xZOWvSlhHgfo+uh8UhSOE7ExPgQvCQ1zhJjxtNsoS7HUsmPCCSlN7FCzPXBcKJMOMfx+R
B+kv/0FwBfWb78N1eNTnFQyUWR8WTuhPjIh5Qf1Yo9XUHpubSpkdCmySqeWzMROMzpGOHTUb3u+i
SpsaaZiw0h3o0mnW0z9kouD4ggbadt4U++6TxGS2r1cFDWS/Ti5/NJal7Bxby4oYxl/1HpbcVnzF
FLBew63Edet7R+kvTN6awfLC++Zmlp34nEV+sTvJOBSY7OBQtcgKHankQAOGKFflluw3zKWnSBMB
GPAmUNWxM2/7RD2Kt1sbPdeadeVvEy/EKZuHEVgHK7kEnXsTFl2kGKg9xajsz8fDiPWbMTEwCcvZ
tazJqx353/FdxSqq8m6w596dKvU3fzuHxIiVIlCIZj3z6BhPtavvD0zbfrhLR7SSnNEL/6CSXjeh
jTopiAETHvGUxVvdBONNSieMZGgKnb7pR2MTdUYFiasKp3CD5RIUaMRWdyIzPqQNavpvG2QTkuwi
mjK8xJDCAwrxsBc655czJoE5MKlJQGXkTcCvNXbf7AD/wmcmWBID4gbDK0CoCDKGmgpabAzft4g9
mq5O/4f/fJXLF7YsWyrAboZ94X6X0uSCz2AkB6mAs5/3u9lEiIvB2TpuQ4jZtAk18OCtPHJixHrO
+axbJA4ymScgra8i9gqjmrT1YycgvaJbtMco0n7CqsL0Ztl+yCggGWhWEifX/fyoIpXqUBkrKWfj
M/hbzarJCC4xiNb5ezSugVbJhbyYTKnAR7DK2uH7HwAEYmETWih/npH38t/uaH+/m+9MFSNELqqm
WFl3eY0Cg4VS4hm3TzjvcNI0W0GfdOEu9oRnYscPV3HKX70GNnL7GxGYQYmwyv+R2DO6QZBr3s9n
S84c/T/bDL8ZX2dru7SLDjd/1KRLyxJK16ofALb7m4lX1ocJpCT1+pH3TSJTZ7ysEHoqiszDw+Uq
CYwl4xOXcHCxd2ma85SfoOA1uIyuXGBWC0QA3wWgwCSh8j2VBIuS8lxOpvMwJK7okiDalp6+3I3d
/XL9Gj7eWgM+3UtTIvjHQW0N3Ypcgghb2IRMHZiTUVmaUcgzA4lUaiK4tgV79ItHY/saF2cJn1RB
jLrgxAf0VJp4Df8rCzKsW1OinIgsquOtcguIv8epTAkhUncnTf+w0gbwnHL5kcxAna5BvoGe8B+x
/ew1qHJv1z9YgzrZIei/VODBSNd77tdZMisEO3Gcnx+DTFGfjlPpcMUx9KA/P/cLfs8hLCfrTqrQ
qwpF626+b21mQN3JcpP4m8Z4l4r/AKfaIG+jHvxlvFnEHIEfHcthYWLg1AMw6kOHa0j7MbhHPfq/
G5UWy9EPDOJZVzRHqoEP+7t41wdNZMbUfBX8jAtlh1K1H7CRPmPWBYzIyYT1alewqu8LSJP5I4Si
m9IYWn4xKAcouycliZG43I5V3+mioGphN7ph6TssW39G3Mh+zyvR7Iya3NIcAuNVZT3fkfH14r1O
53toJBWE3NRdB1Ad3DM4SYbpfl+xebSoVQKtoykX8nRQ9iJTLutwe4ljzzqcutdYYFRTJK1UCLMM
Yg8PJbJk/IzLnaO6YWSIzXmGqgY/ERx3YLcILtX5X6pqx4snEJcM55UR6KzK3gcy3K86hwIlcIJP
G1iicCbp13ubZsRdaMeml4M1bgBhY4b9JFHzk5YSVNmdtBlp2VLSgka/y5TYR/g5tk7lnU02lKG+
D0gcmATOm1NWfr5lUuZchiIMpHEbWxCJmBQ2tpTFLw9g5Xhg8Beg5WHXXh/jBK9cvgTREzIDegGa
rT/nWD18dcnle5G/4apwHoEyInRREvwMx735vd4+RRLAYPZ5F/GcQYBycNZ8I3JDzT14uT3oB801
z10NKush4H5x1GTQl4nLNSavrwczvRcj0m7Tjv198TmEG308b6SNl9ZTx/yJDM5SXBiKNLAEz4tm
5OVk8eSWywdMfdw4983QFskeX1wB/2PKzn54BS8fq5OAtAu/JigjbrUNY/RTr8n1apf5EM3JfDuP
05cnXKOf/0zShZGQ07FFDlFBvnqPDlOKH5W90k+fZU5ui3BrmosLVYASu7WllGc83fJb79TEETOt
5CXtdDEyOY0Ey0mO5TVyd8Enh4RteYej6G7vHF1rz829WJaRCozz9fokFrQq5uW4BDgq3Mek+POF
CnCCFfVa/wP5/M9plnC4WQ5s/2CdIf68E/BU6+sJVmRdx1rpbRFZ7JAMUeHHHTzW0DUeue8QRZH/
Pz0jv8Genbs3FsdtvjhRCrLMytucGCo4pG5sKokulo3WPHPwdMAGKNuG427f3/ZQG4/sPYWekkcn
ftsHMtDRFF4APSDEcd//RJK49MN6kiXIQxeE6FkbMS9WfAeqUE6aRzBXpkK2Eb4eDqYRjY818NUN
HNp6afLbMc6BcJUrrT8E4lkAu+b1s9JJBhYHjzYVj8RECbL/7HehyYLxhX6pjcIBrZaSiQWKHQBx
oBOWfVCmGNilsduQVbS3AyhiZsXGmPwfEmlh041pDEUboc1qsX8H9CceFRmtYAdVHrCkmSr1GXli
9tVYA8fnKr8aq+czNufQaF53HJ0FojT01qyHVweNumWBqfeAI5HR7pugcTrJitMQvF1cU6RKn2Ya
F7/1oejdutrYZJh/ikOzXhr9Z+YXb4KPzz+vp7So2ngobAQ6/RFLKfAGSBd4rN6S2Jlqldei+CAu
pdNuoaQ3xVe7sRL1syanAjTiKL5Is5Uz/kc6fWKlF8rhNHbQs7UlyqnfXXc2B51JM7rW/fmGwkdV
p+E5+hqd4Dn9vKS1h1P7F89lOAOSumGHxwdtkiv6VMU+39W6FyPneHb3IkK/BKB7JQzyF4i/rnxu
t0ebnXrHS+9LkWk4MYcwF3+biJ89HbG4UsUWvZxVf4KfINjiNqgc0INOS1u9UkZiAcf/S9DldzWe
azAVt3Sxx1s9Nfyi3zX+lKRhNKYB3ZodxMLGiHqXQm8Dj0Jyn2z7o4ySA8a68u73Z1B7shv5toSd
jcME/SwApI5faQGqj9zr3a+EuA8HYZgbDe0i9zmIwuwMHelx7VRykmvpwJPxDyK3uGGlWnjLOMCR
hsywfJeV1aL2HIM4ZMrBKfyoxIp3T8xsA4lMZCG1X1W3DpCIjcIJi+gd9u+Uvk4pOMNQUCciTnT+
Un5kmKLBh0GgOd0xeLh94MWUMpLA7VELP2seb3rY3aCnEPy8qFYNcNkN5/ZvEcXNliZpwCGP0DnK
XcNbYJpMl2hZXibRSVrr12jUWPtQve0ISia/QMlx+SSUDuEm4SNrY9sH88PyPia/OnMBB7lNxPnq
Fau/CDsQ+ZCAXe9W+PbJ2ZykXek59N0nSqgn9iKkS9nJ2/8dPgy+NFWVVjfIN+dIrZ9FyPve52gR
INeYo6mSr8OySYixICIFmCN3ZgM+o06TJPd+KDQTiMxj0fvftQPCRBqUcfcOOKesCiZRg9mH3sW9
Hfs7SvSpQdeyyZ0q5UJ56NMAmKivTgGB9oAkqfDMBzXaIjH23MYEqbp3HlX5+uoYlA/FjYY2VJ8x
ZNDHQ3RUsDkw3MclMDIfynuys1zBzStgfElCDz+R6kmzQaeC/EbCKfNu0yeJ9Fwmm0Mo7QZP4cnj
8lPw2o5KJhAZewcB2Wreu2TI9fYi2rnzImiVUd2woc4DkQARRKUydoaw+89Wng9ibb6ECmZtVc8T
DliMERNrhhBn0XsPO/By01x6xswR2Dh3p0+I2r9UOhGAf/i+T3q5UO4+71gOaw9ZIDomW7Jd+bX8
17C7U/YhGZKu3n5Pwpfe0yt7zNOHNw3TRXTiu+9XizziO507uLdOXv1EFpJKll/s3koWNWmCVL+h
hpu4QU5bAF3I7UjrMw8k714zdMvcV6bOgA9lMGYWmIK3cLC45Nscb5FrV0RrLFz1QGJBpW2M/Sf/
nEetf3oUcu922mjR+V6ai9tgJub6VTgwNWGB9MTpQ6RyqyKiDuBBGF+aETT0GaFLljLt7h5elP+i
M4Xak1XT6fAylhpsUHnDl9uXOqoT3RVT6mTW7r7nyMfjVtlcWOs+xmt++8ebKVCC+4KbhdpHfGYM
WS34fnQAv00kiz4gG09tdODb5z5skciqxJkpJ1QkVLcr6ulQfYLSPb58L8buiDSPfNgdVPU955Vw
7qKV+BO1V+d4nepnH1rwA2z9Fo5jOLL/S7nw6ceE5/8xqtg50vpPtV1wLFN28I5pjNtPUCesvJxH
/ZkywZpWhSP/b6dZEp36YP0EVcqz1fTBPZKCUjIAZrmhqe3Rdz5gEQX2ZfEJs3wCHNMBaW5pdhbw
i1rV+QZjc2uDnewYP2SjArqgbn6isAprwK8c8S173PkEQlEFfoUt9cUB6A4YydXxCDbbU1Y9Fw8e
qIXd+izConcuPRguelAE2Q77u3k+X58eAW6bqypAbFAdHeKHpsr9UisWzRWy/o1oOvVbC5Al0sEK
A4NwgCCScwKjukE7jq7FchFVkdpubR9r5g7H0og7wepb6YPlYP0mdw1LHWmPiAMUUInyKvNGLis1
ZDOK04oQk252wrrS/9b0+HDwRHeBsrAM8e2cRxmgf36bCTA9BbMLa+A3DXI9FGuy0N+YzH7rIs5+
6omzcoSdAptxoJq6a6DdT6iIKiO5oeagqsnEY8Izk5qL8WU0pc8V3R1MBxm/dLGQwzROS0XzfKeK
JGEYCaMfsjpvTFOc6TfdxvRZ3hrImKgTiKUh1N3oXeHcHPCBAaZ7saapMoGkHe6bD0/o0f8WOoAM
LlMwDWd0dNsizi6LFlbrs/pTL0YuQ3O950K+zL7iyNDOXlXkv5aQ4ntFOJD1kjDE+PexT3lD/JUk
uGOsmb4rZCgwiruIMLNWkx5RCben4U8PqLvyOhpGr5bHlJD+i6XQDhlTETHS1LAj33mUzcj/nLXR
PRVjq5G9oF1pc+xTWexW4RAaGHoh9FqVPZJBvb22cgwRmBXuRHdhq4MzF2oOG0C5ZnaHQBt/6AEX
3WDcpRsCsp4r6iT304Snk14VC3W321jf8QCtV+e3hJ8G8jz1JWIhDj+vlZ4IpIlpqKR8qmCL4jcu
muoKX9oT/vsbqJWgBVgQFGQyK99ZIs2F023NnBEASlCLa1Upzsc4JdksdKs77izou6gn7+FOXDqE
QY40BKq8AsIMliRC1MC3g0NFzGaLXdl8OLg9sDMX3p/OKzxeOuCxwOTimCQKVN1GTz0t97EctMYz
1vtioYN/APV99DLCPRtSn8tNOHwyqaIEORxC8ZK3KVHeaPVU22vtm5B+ASqVZlQXandzWP4z7xQ6
/DiGlJjSKuk4UEdVRV1fMmNpTHlvT0cdYqJycy9eqy6ucBPNxmAiRPjFA3BDzQ3725cdBT7hzAjn
/d7d4PzkHEkTFqzDdano8x5zMNDGt1sE4VSFpgszJmSLNmpzXPKIW8nfccaWejww8XB9fnbAGSG/
OcYtgL3NiMkYXdVda0+rjyOA2oWtPOtpukBofD5AeX5L7YxJ65pHAFJ2VjgWDHjGVW/YsSi3j7JC
DteuHI8XStXv6IvkJ8GJwZjUhBymc+Ea+xEcjDRuXw/0FoiRwYJwnyAvpoccb5X9nt/NJ5byILkC
1Wi+rl1/A01o9hnjgizETAJLRYf5Xx2xMTAUDmlF7Xnf55B1R0WIog3hJbcQklQOOjR2BhLx3R1w
643RT0LXpT/dSxy22hYa97SAdvCNbzbJM2So9DvUs2GcEw2C/dIVkG5Zht1F9J7VyFL1cPRtYOu+
UkduR/NSJu+YSU/delonhc60OtgYgwp8v8ckLasMswsvzje6LTmyGElH9dSx4NTNgeBn8ExDKGDB
SMzOyBAID6bkAimcYp4ttVCiHti4Yi2mjILXwCdmM8ZA7hrKgkasy87/JCVa5NldflGTeXifqk0i
nERf6nst5HEb9JmbwK5C0E3qhxh5lhfp6EJ82LXdGWEX/P4pelrR4aBH27u6Pm+DHLjm8sr6VpT9
biR90rZoVcc6nBEI/6D+4/byImwrpFc613g7bnV9d4HxPSo4YJnYqmBGdOWqu9qJO4zMyFTHgE8M
X7JUGIRlOAXz4iprJVgRMfkc3tUMkwk6HYphXOwfvGQ0V6V6W7nlLH9WXRjolTXXkdTHoMaOw6vZ
4XJMqi2aR18OCoNdzW/1ForyQkZmWzE6HwzwTS3e6KfCOCLmofXcLYg9Q+RtFEXCzpzjQEU6beTj
nbqRtV/EWf8Lt/PA+CVN5qxwPUTi9bfkgrCgkUF3065vPdiPvVa2dWyX2dwnEqR21lRuNTLPbNZN
rloS1gUMUasIK8yrceWAHbG+SP/FoxJPjLsdd2nV84Wu+WJ8gSRecGp77/ZrOWhy9w4JFgSgNo9g
vMedCT1MInvvirJmezCpfySw4CqY6uKlrDC96vE8QoH5xp+Mt7N9Ronr6qa6YJ+RNnaTWEyiEFKs
DWW1il+VkGv7uH+nkybDHXy6IL9knHuWHvmD/KP09kCzuRDvp1yMFp/MRF8TEztxVCinvWGK/YKf
BqBp7D+wcgoWZ51kgiBLjLMdrpyGZYai3F6oXIRIO7m7NyZvOC0PgqBk8Kj/7SmIRUPwbYe9trfY
0Ahhz0XjeMBC+gkxRMwO9KRiKsZjGxP9fqaHQaPnlzV48Tu6dJEpDS4y0OfUxOA6KnGLlEpTHj7v
9rUGVZGG+6GjzJW0GQ1nLW0tZtqGwnUd3ZWq3tU8S4H0Pg49UPDw5iMbtSXGv1LURa/aVYCBP51a
Ozh03ylVxFp+oWWH4tJOgSj5NZkSaqke4a73fjbpNDEDflMZJAP8u5X3TBXTV45U2KwDLqSE8MEf
iQVhmHhWdGyLvRIpB1RlLX99K8i4bsGgkoIT2BkyfSrRwkKClYIlEwfgwneR/k1AMNG3f6K8UbrY
MkxqwJS2R3swk/jlDx0xpTclrJQmZ+zNshee9jcZHLO2ASnI4dI8o3Bbx5qP8bvoE8VBxM1BTlPJ
U1RGdQCdKRDBOj2g5GcUeVfgq/a6V0QDFN/Q6j3C6ZA0B+5dmFZAnR8YP/gOtIz8WzCj7kQMGIm7
GC+NaRJSLZ1sA7vbnEURlKhJ+v4O9hm/pVgZEjzBwP0r+No++jlXdqLemLvnock8rilL7bgzKXKm
/EdqcnrG79HCB3WS9Y1IDwDOIg9VrlrZzpnPVASaJfZh5mRrXaUVFR25KaoSc5fo7d7P0o3+6+tp
rmIUScBdK2YdH9YfKmMjLtMshcIHxPiaCCaECsIXYKUcnqfLUd44QphoQ22NMsMRnqMhojnLQ88x
OB4/Nzz5p5cC3NjMMFwWy9DKX2M+2EH5us76srMvLs8R32qWOPx1mCj5EM+CIXTee6UzzE2RX4dg
41r4l8ytcB1JRULGZ43v+ag57vo/e2rgKHEdkkl7izikbd4/LueQAWq3quHE4Pfi2ajGKJB7adlD
t15YV11yAsrlSitw2yVl0IPnYNjjfZNPRsycszffFUnWdJIqbiKsE7l8GA3a8fL0C/l4lpSiy1hk
NtSq4pdnv0meGbZqCci6AIiWyg/vUHXxps5+z19mf3E5oWr1D0OT7tyZcz44gw3J/iET5PeEpMCq
I7Kcf0q34jSqvzgjRcsgS44Jt8U6GcqMl7gdEv5gGi52xK+vko/KfmlFvI+8YxfRZRF9nn9dNvrJ
OrgLgRYXAVLVEgFerGommuZaqSdVnWYlVDxQBtGw8BBz+7VKgQGPCHfOdIX6ULkhsb9gzd8ZPI1v
yCntthPItWfbFE+t4RAuF5To8iOkBvu53OVRNyeeqtFVJIDQHfbiUjrKjt104kWNxwaCv20yb3RT
42Ke2TBdLYmQkSBqhaLHHImRye7sAlD57vejkJzotSHJ16pb69b+9LOoGbnI8yEISX83354vopLG
AeY7bUzXcpK/IueFcJylyHA9kTbLmVjngNDBjFxIw9Gi2fZBaG8w2lNpq6VveXGuGkxfaL00tL5J
LKrt3k0pIFKVQ2Zd/GfCAqw2DHUmMLDHsOMNXK+3dRu047XkFCDxtTXGXQdHlRZk8JssFshnXj1Z
xF/2soH7XbqwfBwo/RtZBWamnMU3V+wQjRPkKXWVw1CgQSijHXh6mGg4zgXmV8gfYjzTYM1JGIlb
Q0MVVmWC8VexBKUheKdB7Ud0wCCmtTC7LNmuYX+gLer/NnKfhbdYnMr0CNymOXd/sNYJFcGaIWW5
Sb03ZUVr2DyG92z4Oj/U7EEKWBQidOFzPcgtFOKWfxbdoBA7lv8/H5SyT22+EaJJjZKGEGFpATnF
qB9wTTyqyKAslx6ZA5HxSUDtNWOeQ1qhjTV40Ta9J+xwBAZCjflX8bEw7owAFctdGEybzusNvTsX
6JW0gmosNrl916EHgs5BETaXYTp72cC5sA8fWpluZJoEz9JIfmL3kEqFfrQKkTPJxagGY/KYeEgh
+NOLKhHZzrHbvGTRmdGiGrA2AWxaJX0fEB0oP8h3hYp09YJcMOgoh1jgT0XXeWLxhom+9jQHJYgq
Lq5dKVNq0MOIhtQKhnybOukLoIUFJJk82YXQ5x9Toy2PIY1q1f/xfagJ8oBYeTIKEbY6wO6CwGH7
7VjyXPQpZk19K+xnroeKncsy6b753ooLm+3AJWemplrSEMyndk9rPrlWgvdn6fTRKJbaQ7M/Iasc
cja5cMpmSlfjoJ6tmyWTFJ7A0ksAEgHokDRnoRjY5KqrXllZkj+J0XV4k7IogCjfrlG68H7yqny+
G95NPwtieSmuzO2ddlI7A7uxRAMgYN2qsSqMwbNKyzuX6EDnOM4Uzr2igwUDCFBmOiYX6m3yX8dJ
XTWASgcdyA2Vgk4+KsPWi8cqW796mbaE3tf5Jtl7Ey/XXmTouH6lc54qSbj0tmFDVlYHkZSQOpqx
tZQ9ayc3BfF7Yb9yBoLthHCTlVRqQvOk+FdfFiJi3oP03x3AV0clBOfq9l9UoKFODG7iB6DrGrV0
u5YgNseEKHwmxrMsn8lUTC2UkgHy5bKJ1S9CPDVV9QMs/MGDbUJ0g/s64Hu8+gSSyI2Aat8715uu
YZwRQiatjjEhfJA+VirJz9sXoZKxMWsNs1MMO7w9+yAEpYZPe/+8PV1QY9EirjNIpGrhbZ/Ez7fg
awYu9hgyxx7eS/kAwe5bjZhGCi1TneCaNK1koP3SEB3AGOVqvLjJLiQfc3WqH6fyMSAHkXNGDSEy
A8k48rIvlMLaFy81KoD9gTu/D9fEBJnMiMEzUSxZGCt9d4LFZArL5jh+2922QFNqWbXcy41mMgPl
G4VBa4l6N28RUV/2gjnaPWtTmmsgUQS1mZ24rGwmc1MPQTMhLe1b/zBKPofGGu3qHpBtRSyOXlq8
58RVUPg88XX3oe1s3TxbG8gOlSxzUbI19F4EOxUmVLYh678wVC5imY+V07huRxM5x8FsfN1Uahbp
x829WRwn2zJN/3rsGPAbsSuiHz/lkypuUiBy5xIsxrDt8xLkePFPhooQ1BgO47rwFTjp3xK1dTrC
JKYWAlSINNH1zRKbKDVWg1BuLa0Cm96m9edWBItkF4+sEyS/LAEJNQnqIBd6OY79Tu/f/yXAdwpR
UFaFmcUT0rUWrQ1FfNk5ls6oVeHcwToGKmIfYl9TuZrig+rvv2A+Z+xXQ8Db0wBCsLFYFxApAwxv
v5n+jyTwdu6LJP28fUGcP8eJnUr2R+oP3KvlIgXZAiIv2ichikmz75mLh05q1oDSe93H34tEMV03
HQibhYDhDlw4X8s2lyXn/tq1TUbPikVPwRFZP5Xoc3RC2pBdorYR7ntThvv6Skapjkop80vC4oj2
9osvWypqPno8vNRntP1CM3SRqGdJ16IPwN9Kip7eTWsn42B49xmLzuKScwROv1ppdKTNQCSldNCx
hHQhD3Dfuxpo1S2w8B4VfuL9OuXgi36u3a42IvvRrd6cB8oFpmdWfAV7dFFQZvuOwQ5yXHE22WT2
WVk/+NRQQ6GEgugjrg1HKs2U4CATOym7Uon1fsonIm4yjZNKdUWedOcwzekHbLFiQZgQhWC2EVQP
Yto8Iu5N/ChepHLacjlIl81JpynH6KnVadp57FHj2VFRqZw+W7GZsSmaG7go5iEHfRxReGZAS751
Jc9Bzw9uw/OgVdzyh6v6HM5GsOz8Gl8IeZZdCr/k76+U6UYJ/b5T99HZrVm2PjH8HmZVes/cvNUE
PuV6EKyYrUB4lg0dbTbRPX40IvYYcuIJ1Ek4+rzAJztAHxSpIvO+Kt9DwgUrgLStYjaveLV8bajg
VtiJP/Q6EV2SCOFeNBDNAfDI5aqxwL07srU7kJQQDbplAkdGHPBsaQP2UKhYsNmISiT/rY5iYvgP
g+OF3Hdb1m5KHhxGDHdkbq3pdFwz+yuR+sfZwj/848PtH/NZO4rl6BvMvaP/O4xtMQ9S3o+S5ScI
6M+D+Ab06iIhQxh2N7gJSdZbDCYOzbniYk2T9vl7icRrTJJM9AERd/63za/0oPST9qSKU5iSfkqp
rWznqqGBIO3ZzFYLHPfkNCpYdsXB0/SrPCwwUxKlO7L7qKqIwZ8Xo9CXdkZjT3rqoFLS3EnvNtqN
pKj8dpXbTUCQI4APfZPmUVG2An7yH26ToCfuqG/Ac33pkPH6hCd8YL6/bhoohe+nb/GKNsQyjYPG
PP45NXW0LFHv4M4MjqFxtZAov9I4xi5iAnztIXqruotcs1+i+Dv3paxCN2si3j7IauHYG2hwFMA3
VIXZSDNo83GKCLlfeFYEuXugytrh110CBGCFqNOxvf0ijLK2gd+0TYALMhGItHAyaDF89zCRc6zl
K3acAlJwWZ8I9ga3QaGW2XOFZkm7tf0nWlv4sDbZJiNhzy+AZcIik9uD6ML//tLeYzQltafAsqb6
YT9r3U/AvgZGosaGHQIPzl4N/RX4HfzT/uXbMelmz3LcqZslxVZMcA/SDv7ZUqQjlEOkwIY6bnQW
Ff+fCPvy+QtLw1EkOB0k797QZiMy45RLGYSUX9iV8N0p4u/oOI8zlwcN00dD201M0LB2lMN7LWAi
mDAyIkPNz38l0jrxXiQxwA7QFe3J29m2ArdZJmGD1jwJOYfR4XnDPvLd/Miw2PFSAGgHqCMXtUN/
X39Mb9esJPdXKc+VGbdAFCEWjcrRZG31sK2JWiHQ2Tcn849yXFiQHRqC/hUuGpKFv4gtCl/2k9Ev
TVvRlHi9exqnvVRfFF21xxi68fvkJs796wpZINc7dU7xE4sJfCTnz/5J/m3jcEwytRKjeIwDp4Cw
6zzSdSmP4CY750UK5a7I1zdgsYBVH8Lv4s5KVeTLcBMc/QOiPXZKqTPaqXc2jQHuW8YiZI2QI1GQ
YOLO+50SIrgrLUSKS+o9GL3WMQxCgeh5RmirGPlkgWLBgYPUYwyl4zZY0xL21xpVbQYWOIdm1g8P
3qQkLEmxxOnvQeg8jONAq34XdRwGNaBzDiNhLcxHYNCNWNgkWVR8qG4rn3X2SnkltZPUCC9YWapR
ujyzX+2w9k5tODhIrpUFr3w0IGQK2jnkoJjV7AGBF1ZZ/N3r1YMbhf+0a/IwPc4seBypadQHameU
mZhTJU/gTYlhT+Ld2CqThUMfhtPLU2qKxQXakDW2W9C/LCxl+4W57a0pYt+8qWZId9KaihpWNmLf
E37WmITAJ7xjO/iX1SCDMPVAi1o7olaPjSb/ZD7aiwQqFZSoH6wN6g3yucBsWJ20X9p2LQomkDqk
HRISvMKN/66soJ+XHasbr6CwvouNW7fl6iCLoSGOA2zVIGwLp4rpDZxHQ5NRRtxbKzNCvgPQJ8Q8
6ONQ0WyxDm/JwO75sLw/G5SRXhfv2c6326pMlhpEpwaNHRo4FW13AjopYsnGsQ3p4rNi16N6FZBJ
gELjoRg0crfyWtE75y5GP76otldI9CHH2AfZ0xWWZ2mlEYCQNVJb4CFjgUfIDfstY2XN+LENxg9H
4zxIvbCi7O03pV80eSdrIjI1OhzdqbSHmowC7SadXX/sPtRArF9V7V9NUyxJr5M+T11P4r5D2RAi
2a2IU1SSW257Bm7KM5pMPMnudcfZkrPFNM2zcn8x0pobIkhPNQAZWPsQHr5h6PS61WA4+3xqexRb
aXYvwNspbzOaMKathfdMY/Fni1JloFEyLg0Q2GgMRet/CbNEnUOBI9nrQXGSbgnh/1cuQOxY6v7z
yuhNAiX8DT7Pt5q3UQUWZaPMOVIak7TkEUzxAPU4I8W7Sh16vh/ArVa79xKfLe9Csc3yCOB1mXHe
lzYC31st2g0i/a2hf1O+I3jUEF3d9r93OOd5F0AC0QTSl5zMkK80YTGEUjkqONlzsDx2rW2jo/rB
flwD4cMGR2TDjD3zo2Ds6UuwlRzBKv/ml8bAo5pkTHcujBQvZINv/1UQcndeYPnuv/cDhixl9bLA
aI041ye2GucAFGMzTu53SO+0TbXLeh5ZrEvFGzsVCQPHXfMpVFlfaZ7ADOANHTmwJeTly4HtvhWU
yqyeL0vRSqyyJgEXj+F5oFdsWXZY9KAlpT2UT8Te8qfishx6x35TMRtS10iLyHlGTq2sVnCmCYgF
jE0IvxkapMq1Ku2HzRagJCRCqUqf/cnwUGks45kQ3Xyx6ShF3ed/MBsis22jwrhjFngJWpFvMovJ
Sj80R7Am1124XCV9aBt3UfJWsMqqTheKeKR2QuTmA1icHbjZW0FcnIi0TSbDTl4Fa/aeSS55QiOh
twXaYFbu6kFldRVM2NInkRS0mGLXZ2veO+kqWVf30NSlH8V9rq6fwNIy6D1aeVg/Ebif2vFuN5Fy
fgzZG6B7CQj6CIzM6op7wIfaEKvbKd2fMBBqgv/ybAi2yNzJnbQgNviBe8nNOZQYY47mEmfaWdCi
TRqrixQnFUP603arYZ+ikeSWOvUqhiiwk3HZyxU3O5o4BOw7vVpYL+Rz+zpnrKqFYqR4o5omVKHK
XHqiC61ovextY5xJ+0yiP6NUDNfLmDuVkJWLej/fhfVxUiVtUhC2i7sKcr1LDOBMFQByc92bvls2
fZaMWm/PBbuJfi5XUjgAAuCGYeIGt6XY+6x20IvEjNvKCsBQsKPGzHE5gsjwp34ywhG543KWAFIT
pUDuRxbBiQ2KwhPIJRZP+H6VAD4ZGBY9llcuo7DDTkckRv2nifBALm4FIquyQ1rzulg0jIP/70SZ
AM3sAXkooscGczAZEggEKqBJn23fXsjsYY7hq7P/P7CqAsPPI3JHSsHjsY4EJWZRUP+nKFDY285x
b4ShbD5YIMa5Apw9yC3FLNYoXOtzqxF/r9OSM10Xn+20s9vrwzAR1DROZWla4JtsXZEb5UeCSrUd
mzA8caCtK9LniPNAEJ47vSyzmChAEAe4v2pNRZXYksfs4mOIakGcp2d141yeDIfTgFjgDnLtaiWJ
wjR6NtSpLj0EsxRCAmIV0XWdzSzg9umbvY8EhdqMiw8ZsJhfD6RrGaFlNt+xR2+pS0o7c6MN+JzG
v5Gns0mK7tkZZdTQnDhSBnBU0wX4Y3tlhw0Pp4EZz8Wdzk/UQSRiGuevvnBgYmE2Zmo10ECwor+4
5Z+oe5m94U6ijR+Jq3WZDWTXSSfCTBHwrUE4f9494ikFGxqx0urbi2fP+LBFfRXFQT6zFmQMYHVa
F8XjDDE+8b36BkMBTQ5QxfD00i/4nAoH+6dcX6mIddNZOuv3ZEaeWDm5Z2LW3LB6bRAzzIMtRgCc
HSeVCidw679uVQWetIqoXC598ISa29lqdp5IWjjh1gw46H5H4q5CdvIfqXUh0lNuFt7C1xIR7q64
XJWExLucN0MDMq3RBocWxFQVPdI7pFN+n0cHnOPBDYozeEi8u5t1aKZjB8tvn3+zGfbaE9sAkWvY
/+YpSEsIIVz/1jOzcG4G/mwy23P6jS3YMcY8Y1Gw8ldmZ9nFLJiXSWqk/MqBUUydCiQ/rwRwuUiU
GibKl6rXY54MMT2OY5R8LvpX+VYKrfL48/rSwVw+LAC+2MzdojAyNrVczCK2BbYFoF7R5RbCbUQv
Gd8y/Xc6Draddl2ZrsG/i82jUwa6U4x5bmN121JK4BkjDqsVHazAjMesX6KfpqaEA5r9F4xPtLjS
qgbb0JdhvSbi+6R2KB2Ao4gl9WerjcmNg5NmRieI9s3Ufv4JVT0Lle6suDRvtuZzDFGOLPIWtXq4
HKDr1bCSqP/4i3t7Tpwq01ipbFkxs1YQ9Gbkq29k46eidhaXnDK5Klku3qOXkwo0ZALiZxexECQv
6rh17Rjp+OYFwTyUp3hhsGLrixBuOtaaTCc7RYUAVL5Neqeu7iI0UVe93+Zr1mvc/5FfaYgMajYQ
zMugHB8KalEuLuZ/iIfSvlWHDjqwfeSgOlE4IrQRjovPvavDJcc+9HdQGZCjULlZeNpFfUeTXETk
9Dy62dV4fj49nntBGN5XMPh06MyDlOeR8/xg83wrbQwTHrMTTEfUEgx9UwdrnAX7pniwGBxdgEgH
zYdtgipdEU3JL/yOmdJpTj/MB+yanjObTFwoKGfbvBPj42FqJPNp/J3jvHkndrGF3gylN4Axv7lU
W5meNqMvnewySLzGFMwChAXvVbDYEe6ZUvvd33zxcRJaM8pRGBhGPv67XksqWj4usc2dIJo7obFL
vRQ+dgfWybKscoHMrtE5aDDRbbnbHE+wcV8YAcYw5imwNGrcwDEgoUr0ale73kKgEMdN9pXHi6TK
SeWbwdmrqclA4xWWobYNvN2otLZpVXIL12VIDgq23tuECWGhJzW9/o+L1zgpRvQzreucNB+tx3Hr
+M4HimmeP/aN0QWJf4NWCQYzs1HTkg3TWBioHXnhqeZAlytSY44u/TtpdWqWJe79b+49ny/Bbkhq
Bt7mflExCV7e7oFsg+HoMkgoJe9S1nYlb0eAPXz4HEQWBGIQPmQyH/c8Qr2iaO9EvlR7F5UzUJUZ
hM6s1Y7QjH9mNTz8657gApvH0iBMU7qwH3QmMp631Bo2xlDGSVDOH08WKqEYmUZ6mbP94RIE/OXY
gXuxI+Rkt0H6+lqgO1V4LeuC0XJ/ociLLco2BCbXwupwvgpNGGIjs5CZA35njqQAmK53u3ASUpCk
uTpgEQ7wGL8FBgDN7P2tzU3LI6SOBPnHgvwO8JBF94PLzmeq8vG1Tks3Ms9uLX4ObPYOXms4Xjgm
C6OAqepOUrLlBC6yk9sE3o/Vcv+zbwMa47ta53U1tXm+u+zTtkWnhMMH1Awb1zWu5F54sKC7ACX0
JYakgIwUQZ5H0X1u1axth2s52IfBe3ZzX5xxutkthUb8OzDQwvCGqFcmc3AxUrAGZ1KDxR/I4SAt
kZ1WDeKWQiZqCcVVK8vdeWvMoesGUeUFbuD3l0x4jwvlKWLLPsSNlT7XOxpCJGZRleADcCF/5J7G
PPKg4ocZYpRIR2EoBLscsO8Icshr8cy2cwjXUeoU60xTrK6EWrYr3vLYWaw3hxoiMYeln1VK/C1O
OCwPGn75s7oNBd5lIboTPYlESHeyCykjZ/YH5GbLqhPvGq9xy2M18X5IV1XcVxKNDoWIq4pwsx6w
PdsIJk+0g/LbzHGf2kSPcdLvM9FgX0KelapAxv8uYup2v2H0T39JeSsmRHs8TGP45j+IFPXknYxO
7aad2bv1u0qcKGm9yJfBf3pYOsR5U3FqGcC+MgpWtHAnPLjDUkb+HuT3eZvqjOUHi7vxvOMrkN1U
dh2UTk0X/QLxAsdPWDitHbhAiYH4vpZvxyqTUh3+TnpHrysJPIdayKXyDHoBP1Szofzco+GWrG5W
WdBB35sh8xvj8iMFQ9rBsHRDS1noyphTeYPN00Y1rkj+6c44mBxPBqbT7gNt+YCXbe8X2G4HjYil
oaf6tKrdNP/rZpHrsa24lpt5JDoU1RFME3lgaPf/wSJWChvboFylNCBFOtQSqgJ9FtzKGTM1oYjv
DpG1sk1kRY/LBEV+ERTijUdPQOl/tLvQlSq0Wqr1C6Sq5NyzmBegLgTHZZhQrBZIlMp6J0lZXyzI
8UazNj8780oP2CkXNH08573TXRVcPQkpTsiuzOC028eopznfXmWVcO1tmj6VZdw4H+vhmDRLPLKc
y4t4fXde67R9dy7UaFxVHxNG0ivYcx/QjwnfrShTjL8x4eoxmdnIwyFgc+J30IoPfyEM9GicdjJ+
yuBGvT5Od1t4v/whxNH0iMXP0jFptNcYKXSAc0lu1AXpggd8zTLrpAzc6uViyfrbnLEwwa1sseHZ
ZNGcXZDEccd/fYNxUj8VLxWTXQrcyvfMeW0NT3tFVPOqRBNY0JwHBHbbez2n/iQdJDDdqa4DPZJO
f4FdTeWVP8ge364BgYBYA46tOkSp6erCZXu6TvUkl6G9MsdLPOByqiFo0FIyJukaq3tiwWBzHsDA
QiacYpQXsoxHNzn/lH9Xrvbdv/HVY9WS0PPW0nQ3NmY82kNIiH6g9YeRGth1oIY/vWFzmfcSv948
EDjhHUjimzsigNiVoFz0LBCmukeVEFRyqi7ffqRwe+NmED8OQsATbz4I15TSoc1D498QgY9bx4gc
X3UcVFyRetwiDxXYdYUkXuSz0yzdWnByTBaFn47TjUWBhrNx0sWI/yGm97SbNDf5h8PhJVqrRmrr
GPm0C4y23Z6qLMzeHeIRZSpeTcgbqYrqcG6vgESsPi2kMKJDFxShH1Q5Oyg64M7ok244E+pQy2nn
29AyT5e2XGK92abcNphNe+Ad+niMc1pkRz/hmqV+hnWQ+1cSBshOxa/QIywTfIB3Ljvi4YrIDjsc
ClFME99DawPx7wH1yqr+IQhXYiv+8kCPCQ5dBW7DLR3dXMhUBk4bTsOaBvD28Mh7MBCXTQRWXn7c
rj2oUCFPnGIh65gqxQeU0NsTe1g5lRJJd9SsZg0E8V9BDSXIIcaQ/g7Fx1PH3lpvs8prCYZg53D4
sFBzl+83g/mlEqxODv+LpgwVToS+BkAPMq8q+g3ZCiWLoVAyIv/Im9jxRhwTI0PLScx7rTXuyJJH
lytgDpqFRzCAN1qdeGMpssY0I1PQ53l2xgEsqQees0cjEYRmh9ErBz0p659sH1cDRlEW5gokp9dF
4iclPj/r8WiMmo6bcXTBxYMl7sHDv9+HoBdKsHfBinBY9F/W+EU+swEsWl+QsZWFbbbr9nLIXON1
tGRcNO07RchntzYgijqLKeZf+CaFQkrKJJ8XpYfzk/4iVIoF63bSLWKHeHpyp20YxsjEnLqmU261
wUe/on6cU2trsHyeCiAFngpU75hKYyteH6P93Cnwk8teDciGXxDovt5NaEXCJAgOvZqu6wXxpE+G
1ncqX/ZSrKvGYAsV5UGdaqUSlUc80S74GeajYBftoBRoS50wweNB7VIvjqjGlL5tXZHqJhB7DFp1
7DucXqOEYAmEGW4JL/YZrMvnQJ7FK5qefNJLV+U8omBpa3H2QcT8Y0Bm0q8ojAHafdS31v+IQfvv
MylEDbyifKpD/YAAz0X7AfD7lHUAHuKTuJYhycP6JnKfBCQymuTSYMa9aVbwPZ1RXeCrOBdYCD1M
jfzN+EdaE6ZOp2WaJGrpKXOWFOeiWTQ5jxZpkqZG0OZ/haR2WBrOIxaPR4beFiCY3U8a80Wee63+
n0atnUsnASJJ9lonirS8dXNCQpcCQ0MPANyDgbMNwiYfUUSvYr1rR3rss+VL9va8w7xOE46QekoI
HU+CzQ8awzCKJ43xFHd39uGM85D3pIXQr6p7hTZA6mcNQcJ5+f9V03Tx02a7PXemX6X9pRd3R60t
AZJAGxVr0C2S6Hsh0VmBDP9RqVCJvVIcYEI/ZF4XnqfLeyZnxycsVfoDyxZ63PFVgVUQt8Hd/Jb0
/ao6gHMftLqESqsimxH44cBgf8Ro/aPgZ+pw4hVhlEFXXV9oGure5kc4wKk9zllGJSfLpjwAO2NJ
4zMkgmEYQSg2IRjsnyS71cv8RL9wuN6dN65wCDDyINZAeNsELrxQAzzHoB9ENLMUWWJAHhusd6fQ
qXyA4P2l2ko6H1ng84M67g4CXOcbKDXGz20qjicRgKyRb3fyupgVfkLd+4MqtsxxPXWXp/7b2yL8
M616qaKVaAFOJrvW7tF3khlxNsZV1PObMdjnuitoWpWz8pCctfPIjVvPDO6304Hl1+4ZWqPoMgY6
2d1kzEJpoiAu4qdEQue5i2xhjq/z7pLcL2/R4NCPf8HzQQaN0ira6HPdnG0nNeO2PR+bSkWjDnJ3
BX8OZJFpJ+opRZHbXZNHXodsYCOua6pZPPrAAIbpOfH6Vd2MEsttgtPmYc/fu1ViJ5CIsvtohtVy
OvaX0oh/M87A/flr8ILnT61O01SsyJ02Unh4S9nfqhIzeL4xesf9IffFwD2MMszvxZekfrobT+jV
NhvM/uZ0AcgP0x76/d2YwDXIn5Il7RG87lcSVADMICB0zHcfvf0GfWxVV7/BFzdssmLYmFCRmogo
EOIiR0ttoXkj0DUbYxs9ac5MIh3nt/fYQbDXJV/2SaMg9cehOIhg+U7Urf0lyWwuXR6vbdszzEpY
cvLB9h6k0qH1YWgIncXwhIBGkofVZIGlSSzDPfG1OfC6+5agoyMyK8lsULrxEj59yJSQjZGC6Pat
+8ny7QsU04S3OvWKiYj/Z2OMtxprnQCEi6OxmmlskFcJAOPwrcx7IGVyCywb+O0BkY8wr/60aQn3
/QWa/EP7cUexqYhkd8cM+4Kp4DpxUZdjAjhn/Maeh/rLTM4LKXKdU1nGgW/d9+Rt2Ve2ON+BBMGE
7n2hEy66iBAkNGPu9/3kg5ICadiYaT7u0ombC580T4CbRojFbqmJQxj9U29LeARQoHkpqGPgW7JT
nCoDiRDStTADnLXYV6hQbg6NJM54trrRuitG4fcIEm+KlWRtcM/rf2c0HFHkGhdppZL/Q/cxl+55
2R3YJXEMYSuHPl+J0xQdv08LqxQYVpccqxnhy/6bNnxpBavybqPoTeyjMI2bmuWdG0ZD45Rdl8I4
3e3hARx/ILGK6x/k+bLIjL59J8NXHimuVyWW3UKYmMpH7utpm5TQKxFcHs3ZBOe1DAWwnqJao74j
Tzw+/6cd+MGaRqmjgBDoDPVEJx0Dj0l65tpyhfmMEEMexUeYQZh40FLScbzwrnvP5lJeou1WMTxm
qk0SDA1iAGt7GtzZkBzqOhPfzz4kRk3SgSs2OAdL2Eqr2Sh9WWYMg/O9B2yBxl1R8hYpciZa5Q8F
AeOprjC8KFvoL6lHR+YQV5IHiagpKAI7rftwOO527YKEkGEGPmmKKsXJVNnHxRQbEuvFkNlSOjtH
lwj2do4aoxuRU9hO5DrDLap9ehETwMcei9OyaYMXfsEh6d6E1yb9cgGBV4lNm7JdaASJCRtd8YGD
9NIbBd8KJ8ExKvuuskUZkf21stNacoozO3sL3mjMaAxPd3X5ZCWt5mXrg+R9a1CykRUClLy2dYpN
YbeVkLW74oIFI7gHYEzAxu52pKyju/ISFVccpZjkW7OGkQVpP3ZtyiXaJs4EpIqwWDS3K1v9D/bI
KwNoEZ0WpOQs7vvHGq6y4SfJuIYAA/RZ8B9Dj4WdDJS2bckN3sdP6aIX7DAqxnFX3CT2U+maIiUq
9/KLDwAQbgrdHRcDKfz92xvFDZMkoQjrg5uLzqbfFSP98nNj0Jq/JeSv9HsHKEDHW4rQw59dTezM
im9MrM2+afrQjJaBym1/RIn3M/65011kKLgl+aQsQ9GeVRYHIzy76oxkwqyoRs3e6OHSoXGYy+j2
L/LSG4AXm+A2iGgbt26GahOM/5ZysJ1Zht+me6Gfm8bZlYLOz8cvkLMEka4kKwodLZeDcbSlf8XE
OSQ1X3u0nCipGgbDEUM5Lv+vyk2N4gP5k/zp5niL1z7tyOhRVORVN2S5JuTm7/aowpiCLAK0acAx
0RSCvl3kCswldaJEThfQAyAWV/BOxy/TcGIC4FnBDAqG1ufuywEzeUcsU5nPTnRTJmZaHe1QhJXW
J3p2JCYw4VGCVkgCx8iPmii9hAAlWZ1JLkEpHpYxjhzduRs+oC4WQ0vDdG9FkgYWRq1LvbJd037E
Cx5lDcfSHi42zYttbMNVC0nVxxkMlDM7oJ0G1pRbZOkYCa4U3+coppBY7mY0NCrsqgP7Z2TaGPSn
3e3IpiTIjOrXEit1h/FBX9Wy7/dVZ/+pfYJiXLqzH5NyY7efzejEmHVD/UljkJdrgPhkOMW9+2C0
5Qv27T8PfvIhWnBDQDywG+HXM/lMjCSx6DC9wk2BnAPS5RZZ+IwBkzH9x+oIkSReZQ1z96l7tWU8
OxT/+RGN1daA4mbV2h2TH7V/YKWqGrO90A9N/cneTrwZwNV+cUQVBzqblgdvAWMdnni2/wHQ3C8Q
UR5265NKEXlr2s3GTQsR7Es3zId2Y5XpHuvn9cTRfhwwY6l8slruJWamfOGmFbpuKfntmkmUQ3Uf
fXoSoPNH9hG2WpS40kOPpf4cz9OG5DOVhVbqgYeyoUnmM0JyrHQ+vbBNji+F5ioS3oT/uCiyPRoa
Btmwp8sP+3y29MWjPaYBsvMFlPtVIkMmdMAKDwWnwQGM4/5ADJDm+IslClRqaT7p+LLUj+zpV02x
T0AvNcSeymN8X3eLDtlsXVwG8qiVdSjuqUb3egX/rfYg/HMzWPjhyZg7eIhWvepsNIXEJJ7vlftq
DrHvzxL8jFS+GWscTqS2oDvq6WNnORA4s9j68gatAhoT5/GCq5fHe9snxaRtpj6/1xKb3QKxifv5
fzDjosnwraHpodXbZoGDnLz+rP1Y7NLF7yMRdXAJV+i7WBRzHfyHkQ9jXGhqTI3rSR4NMlk+UkQd
hVOBwRXK38UsEo5UHT9DdikLN0h9SmD1455iVriv5HRb6MDwiX9ttSZ47TNdtckVHIXQMOrHfjWO
ghTp8gmIcgRm/9rwi5VIyo7G0LoJGJXxtpOaJNfehL8tfaf3rFJVUrOTCU0kqAh/wgak3aTDXvpt
bOSZ+o71WazxhoO2kACKpG8aYx6Qs8f8G3MzKPLRYJx7Kd1ZMZKbaCVq64NsN3m+hje4Q4zoCrOZ
BraOR1HqGzLJtNrmCTo0Acq7jPRcLKpX1TdKi8x4ZJ24UFb3jFNYWbB/b3tE+8lZmCTNsqx6wTYN
LdmvQB0fmTL9Ur07S4EB49uGTUiAzXrBysSR57gUSW8bIqkw1MsaRn7lc/KzNXAGgCdSNYebbEPY
Yvheou58RfxxKC/A/RnlhjTFtwhUW7GBWXZdRUB+NWEr0Jdt/Dpnst++EsKDoLdmH1v8YoVPoTH4
3c8fKPJu2es+fYyDqXd5iUWKzuVWdT9vZoA+wYVxbMdNQjmz4ZWkqfUYEx1WA/JAZs+iTSh+y+1Q
5oLNCFrHDEAo5U0Vr/LJf0raplIF5Bub70vT4AvazOEVq1597f85stSMHgP4s9FaXcOlvbhoD0rh
zJpzdUCLI8gmOn9kMGJSjrbkGqxh9oPiQPGefWTUtKRSoaQ/FAXMt8wMpF1poQVEwUEZAGX0kshn
5fT+lIuIQyr1qKQu9LfEB0zfXh2k3aUJtPyqmS071Qh6cITOV7VcoCqtF+tpbt1K0K72ozo/3aAw
WEdbdQix1EJgAevbK1NEo1yXrIdv/wBSwxFQtS0gS0SI2FLiO0VxXvbhFrxA9ec1ala8PIufcqJi
39dzEq2EGP7sbTn0DHuT/rhqpB9TyfOX3paSeAuhxxZIZ52fuWqhJcFP6vTNkr4SG//ezvI0uFDZ
uY7mneMKdRk67X6MPj26JQqYRKuwbYkGkWnD5NA0SPWX2Zy9mETrBWYfjpbIFW+OBlUpEZg2pQOM
MtGJgkUg1EaFKB4423CBSmhbCYUMkzzubPhNQ44QZlNr4uWH1J2M8BzEDGzVejW9Hbo1LWgMKfc5
+gqRmFqk2POcqrdLu7riXySOkwfT+QYEoX9oot8Pmls3QZrHj7BwsMONuRV9T1LnTRqg6adwMJ13
ycoT92/akaAs60BgqjDTYny+tyvJ44L0NXQsVUSDaK+SzD8Nx5TFa0OhAwNzCTeD0lbovnZohW1W
8pVA5vtvMVYCtmvVcX1yT6M7MA7EGjwYtkRGl08+cM1rsk7Jdbng97uh6KJLWffk3zHTatb4fRRa
1idlF1zXRcZYBdPMBqHheCL+BMpLuit+A2hh3is1Ms+yqpkv2yPXLCjBlvMqUjDtgITvZzmGB+Ks
XqCXv7qp6dByNE2asAiAaVfxXEjxwsCMeZzTJ8aNGpF8RQTKFguxiEMxT4h/6bbQY0C6Gk6RSuGx
bmO748YoOLfvzCtCd4R7ODPc1pk4Ac/1OBSj3HlyiLTXFEzjJ7bKKEUWF5TpZ/FpOIhHnHloFZY2
nz/pkv3siELgCQha4Cv6scqqMpsUsjF0Rgfu9dFrWiAtbEeGgXfqVFMVV5kUk2Vc2xlD6sxKk/rj
qvg/l0Sz1Bp/gxKBYIC/xuxbpx2qJjp9pGDD4KPfFSXd7mW66PxaPxIozP+td2MUYODsFOoNV/hG
h6qaJoc5uJE1CAzzqKQSZZ5R2l48xFhZKFXGoo+o30cX5XiVVxMwhzWOQf8nimhlW5CqqclZhwTT
nZRlGCdzTJGc//Kky/25rzpU8E1t+ccRm55xjGvWoE7RKQlZjizUnegOjP70qO3INB0zh3W3xhut
ir+wWNuk51eQz7Fwvc4Txf9rtQNYYNY1KKnGXj42p7rUnZrfudd1QfjGPBwGzVrKb3Hqx4/vvptW
XuLSBWADxJClu2E7lcVelCELqKicQ2UZa2YbG9ArQo9cjl/pPBsVIbRwIp+j76yKXnn6K+ha6Aut
FIps2bPPAj5V/oanKDQpDW8uSqjfFUHf3fZXFsyFbSltYC81abrF/BbLe3GPyGJ360wfeEVraD4K
SZbL0UmvE7pddJ0MfNL6T8cM75ZSbwlQU9jbscDjwW7AJG6kjifMovQdx2rR93kZ1JHIBPvEzNES
1LrQHpyIS+A/yEk95MvTyssFr9CoHsYwvY9Gct6wWgbz8lgCVWyyUSEOXhRChll22TEIvlThsMxA
22s4wQynb0PgeNnG9spaHocPryUj3VhFm7oKeV2yr6ZAQvNGONTcAkAhWOEdE4OdYiK3wszi4ssc
8Cf+5eyUPY2H85wp/90Ci2++J5aJPtNBRGUPhqDlvGuuZdfhAiN5qEW96ZBYGQaT0RR01lns8Exl
+XclcLd1oC38MV4zdruwWp1/ndN1ytz54AIcfzhnP71oNS1QfWOf6wUvdCLcHEck9fCMdR6yv20y
Krusa7gdgj3V8BdAnDxgtTd+B/J1W+jdkLcRWdtWvzk5d6WImxEqeIuaJFtV9wbMjJSHec/P2WOP
mHSsFRqPLfGUNfzfKE+c/Z1zO/aZjbff11ncsxTjqE4klGYj1VLwY9Jtje9z6ugTyg6gRKkGsg9v
PNJgh9An3Zblun0iISim/bvagC0cGHxjpMsbUheL1TIRyH7m+v40/FVuv5fyrZcTx2P4LuRQah/a
h+zpKjnJuJBQ56zFvIiWUwrfqQafaSAe2+zDjUI3Dstsi2Ez+nXyxYitcohXHsdVP0FD5479D/uk
62Dso8uzCC7etXrZ99ziNplruyTy/qIRyXJe8bQYhYR86vN+OTnmez5AoAAzZHFcMdQUi6HFiWMe
onOi9lGJiKjSFqYXESg6UOneVLlAvxbK/d7mpGRlOo/NcWAjvb57uy5P9h9W172FTE2M1hsUyV64
j2ao1YayBK5lz9n5s9LrZ+J7FEF7m2HfVvXLEzICqQ0zgvl42icKkbv5t18iLdRc68bepE4HwM7j
V0KCguX7oZg9bPvLtFGWvaiP4uPrQOaRggZdPIA8zKi4hNJd1mkJypG2Dbcc0tPb5b1oaa6ODmap
qkRHp4INfgZ2XSyGqFlzUiTkamG1yGqR3lDFzyg54VOjikz3pnrDXJ57wbF9HlM0e9kuTHyU4O6u
9bI9BRRTt1dyLTaDgjMn5/IjVdOv4IXhjH0FydJpI2fx4nSwrrW6uIv98OaQ3uCP94ye3HNZushx
Aidruhj6SlB0q0Cr/mOcEnzRV04XX6tyemmhCUBMXJxFrNx1OjSc7HYvD1Dvgz9iJFk5aylZSvSV
e8j48UtJgZNNqenxAv5GM7M81jnUpXoqpI69jZ6e18gVmTIjPu0v/jl/SazZ/3ltmey2q2A56BrI
ILR2hm4Bq0dRkTcHUa/duo5XcYO+I29U1YWvNfOtRJqtkQXXInRJeqVOlsUXvzx48CQSIofFhL59
bvDnJJkU+CxGmX6NrUbQE84sPbFWhjpwTlkwQgYcLv6qdrBvBPLslmfzWOa9ZzAVU9h4GwoDOxES
hzgKZwAh3Q/1lgSsZ+C1tytac0FgGEE4NVnsNKgA4727Q045PfAvXAMX3JHwq+IwcNhO2mMGzzxO
rOuf5Gb8dbli6a4AfUeSjmdnECk0W6Hcg78lO5wM/+TnftTOCmBRXRsAaAOqgAcxp8NiC2cqvQ8Z
ydoaxIfzStpbzYKGFmKp8//e/eYL+g0g18ruolSQLF40048lUAMiCzyvFudcgK36V27FV/+WJoX1
nGdaQwFMpPZD2rYOcUH3XBqCo0DD2jCdp/vnh+m0Nl0DNRJz8J+pY1lvtj0JG5+56JH+qhf3qe5Y
mCbH4MOdyOBy6BJFrZFcpEffXUasBp0saiavALYawLE85GKhWfkvnRFUuRGuYtSThx6yGBoR54gG
mxM+Ybp3F+DhPtKXaBRqOFE3Yqa5cH3kLvHuCwQJhH7HvFYPk5UJX9t1mtA7kYCe4AIOhPrShJGX
kfu3kahvmixjqSqmz2MRgGoM26xrNneu/sA0kilc8l5NLzCPZY3NLcB/JBhz1wG7gc+NjRVR9lff
KWRX/dfkr4/4HsextMx8H1JXcn1eVue7ne1H8c5m17JzBYCDv9cloibfm33NWP9lsDpTmfWX0btD
vjsxLUPciPnNRJLOtS0PMvqqMcB0B5dVUw5KsQM/X/2YPNBAW4e7eERVYJe07jX0hhg44F4PpcTs
O9cQuAnH90Nx32En3sasJUMcNd8n9ep9kbQQE4D4tTKprAIlKABQ13kMVwLTf072O2fvPmyijLTj
LY0A64UUDvU5eSRzvbmQVn9LSVZAH/duccCr462yAiPgMWJhtvs2JaiNpx2Bc+319vwggmnrVR87
8zTnOolWSigvueotJLm9i4NcSiSX/5hDMDi3ZeO/T/vNorDITAiil6TyBFlGm3N2O+8/qrQz4x++
3Rpway+HsjNWjdZXlV0jFTSB5Q1cx0psrfH8yyLJLnfWT1xhikikOI4l2WXzbTouVRwLojqlgaUl
YW/ijqr4CC25lPH4FiU0XatazeOBbWnyysQ04ZD+DIUjrZPxA5YnuJ3Md9+LLvDRZ5tAP7i4y6wi
V2TmHVDH7McVulcmQFLaTPwzYRkL3C079YQ02/2pv4lud4GL4Db0VP1ueb2kjDfzO5OzvZ3L8s9H
7lV6O6pmcbxlgTtw6rIEAlMrHmmm5r6E9XTjB2qRUW5yKjpWhzMNB4Y1x5spqicaIo6L3sUjI3wB
qWEAHACA6aYmKPhqK0Pfu9H5NRAaf9RoHER8v9x6OXCBTBRnfBanCmHYcQU8HZv+GmiZvfZaBgJt
S7+BYl3Up8vpnca4TtQ8uC728xffFqUtam4D65HyH6opMDQWDjlP/5bCmwqcx9lqPc5OAtyf8ZfP
xlpvAsxIHkQCr65c3/0QKApfjE86Z1995p5hzFQQlR/okSTDdBMrS73XHGXpsk+AyWWneHHPaDD/
jhVIVjK9LalJckOWmYv0IOoVk2zaOXisSeeFV4zGd+c2ngoOru/whVQZfFHt64uxQilLN5fD2FEN
ByQFB8hBNSjMPdzr8G1xcFyDuD7BkpZZmjdFIk86y2kQpQxk3gAv6G+Z7QmjWul2gTlujy1kAGIg
Ha+aNc2J9UWj0np/b36V9zRWL1IfGJftFGUjJCFBxTQ75pfHwJx+knKpb2tL6Bq4DJ4wL7MQPysK
UKGoc1ZJK5Qplvy0MFiLbWChaSewtb5jx5v1YxRQhPoryZ1K2KrrSU6wJB52XFoqTUlu/r64dkVa
FpVOpmVz2ZKpNcPl+mj3j9JGCI8ZtNdViMDYJcvVttlDI985gICkUma0z3YP0tLgfJOcrxGFpa/D
19fjdMYd/agG1/F9AwRt4bLkgmn1uDfHI9ZcjKWHw5Txgw0aw0WBVSMQZQx72rkDNPvfmfFCMjBP
BmO5J/HJNqkNDR3g/My1+1tUpaQ44SLcs+qCigl8ybYwsFIjIc7ymNo99esgtIBFjfOSYTkmVL7p
QusEe04/3iuGevAtmruDdu83gRZUTQ5dEvy1UU+2jT42NHRY8Kg3126MIufKx7o3qt7SUX6Rw1xM
CkrjjaTkVbGkKA0/0DnXlmKKFeCfJAcM9vD1irqb3c2V+vsDj0TOTtkKhRQ/va0EtBICZp5FpJe8
W7LhrBBVFeW7ah0rHu2myltx/WHp4tvgTr2dGdY73FlOIehzxMUtR2QPx7+PmzN5Wj+UPsyRkJ1I
PrW3VqRLN/esjhvaoowTwtYGialTvgYqCd3MLn1ANzwKuOFJGxn9owU8qRElrzFhgyGytqmpGm1Z
GUMvM2wCTpgNNcYFOHc1pJMCU+FzXhWkiVP3iGS9UPeyTBLnuw2K/TEWo298ZWwj8YvCHeh4GLJg
3M3cgWynlH3qPGw/EHoyta9OGdMZLzt4BqXnJgHQ12stQzQz+Y2KLZ/mfgs9qe6CIAqsJ3RFNE9v
Eq+KDd/BEeNfdk+EXS2di1bGgRldX2TMReZMhnXxBJfb+WJTASOQJuz7CnK2AEttO6vgjXHjpzm/
Kezy6DUcSPvaZP3dPXnQioCEgyC3XDlBaUaPBwsnJDcjA1erO9i31jsvatb76xPH/hjUJJONi/gU
m77RQCwJxzn7Al7egOMteiwuNhYYT9zJBBYuHD+5J3ToWkKrF6H1JjfMS8BgfIPUU0ftthnugjc5
1gevqClKdM7mCmtNWA50PHW4hwc0jvwarj0F+n5etd1CDKJFiNorySfp7GRQwUEeC1VilNlWCOoJ
NYuOjD7mzoYdzw8Hi8GKN9wiTAPCTFWlWumo7BfQDN2p3op/Drg6pkvO6bgGOdFda4fFaSaUUpsD
rVqDoEhSNqR3qiw5mBM5t0krbKn75jhNSVjPBsruk8iUSBb2/1kJrxBV6NDm9wbLdXZwa06D2C0W
vg9fWgCtXKbg+avzWqISSo28/Jr/slK73OkX9yyK68hSJxzj1iyHcDo5WtywZM0Yv3bHzGUcK9IK
C/1+w9Yqizsra2QzAf4201u6wnkB6vqShG5y2Ce+DCZSqpzQwW2z3RgkzrscYZGaTJJ/qNQuTAWK
j8qbJ0m9usf2dJAAQkhgUAJnbNRCjt520HSGrck6oaEhpsyPSJoY6grbH00LWxKG/MPGbe9iwjT2
6xYHsN2POHmXboSfimbggtRAjYzXgx4sDFCcEqmAIx6BvqWNMtgDSl+/xcCf0Vr+34Lthj7Of/lb
ioEShm/24uK4L82LLfS2HqC0JvoS3Lm6dSgF7945WL1AI6PPugOHq+Kd8Cx3EufcquuaO5F/1nJ6
erUmaku81JIwSwo+vlTiJfnw1ICRr+341VF5oXz76e7F/mFVFVW8+u2NP7ELfErbHqXjjSu442cX
pk5j9r8a2XcZCUHa6l2PWoJYR0bEXm52pyps/iokuDEJidZY9jJ3Ew9ua2PAiuIEhBKNx3sfMBGO
m/pKg0NGqW1AgfC8qkfnjGhjkw2hGtXBhU12GYzbAZ44zdiEqP5PVqgxOIbuioW3PdtYLk7l6MWt
2CpuJ5jwgC+X8xs6SIDsSn1DuGn6/LEgTYEJuPZj8B0AzmOhi5rSoPgLQ6Vl7AVx4TeXf/ASOU/G
ZvnX0Qu+Z1e6x3Ttgto4fkaJ632FkaHRDstw51muFPogrQc63F6mMCH3BeK9r7OI80ral2Q1WGlf
Ro5p40ve4+X2xzqDMgJqdi7gg/hIxs/ViHmAkGBKpcf1EXQNKINv1JecMDYoH0BXOywvUTfDgY4U
RuudqIeKiGG1SxAj2+ymDM8H+8bHfmn0YHN3bzVi9iXRBBD0Gq9roxaICmNf5BvcZSP3NdLSJolL
SXYV0imjylZyS3lZ/poCheOZI6k6KvjOj6SmZoSSLhRVuhKTgi1rPX3lROZfGiCp4lirnQxiLZdF
AOwuekMbqGIbJT1sdnLttCl4cCpcgYGvogmJgou+zZYSb5hlBBRKD8dDKzWgJb48DtOuHGeCP9Rx
4T2OZa+WW0LS2dcwAvfW6xLOk7sfWrAAdE6rJGWIFVWvS66lAEsuBiYOVqDwhHQTJJnevS7kNozl
lDfDpB2bExvXmTaudM1s3DWu32lwEWR1WqAMGW0xdL1tg2qf8PPdU++iwtoddHuCn2Bxw2Iy7nCy
mcJC6OpCiehU1HspwzfiNlYx6jYqmAlPVMEWpeAIi0hm2VB55umvJR5PMlYL6141VEcqYUDysujI
35LEW1dQlRh3CZNAhKAG+uy5HTqxz2CGXvHZ941v/FN4O7La51BkQ6wgVS8DRkvZqlUVLwk8Rc7i
7dUW995hD709gRJB4UWNZxdHjmddy8dII571zxxDDxHqISB1TYSkQppy4qKoTlmG3VlL+/O43mOs
CYSVZsu2jYkaszUsvMDeQtzvAbwuOez0zA/6HcW29KSOlXiVIUqKtTlhVuQXl2OeY15ULQywM1j4
GT7sM+JsSAqyJyiZT/6nLoKvu3NovAuVOmAPyJKGotYbRuH2VcZIT5nAwMjGcg4JkB9NqaUBTK4D
hRR2AESRWUFO/JDetLfTGyIOKC3k2bekB3aqRdxT5bPOc0ZMwa88i/DEYhVT1V0Ih9MvBqphg0u5
F3o9DGFRZ4+aJMgOAwbXfKA3Bb+Lp6KO0GR61ijqBYfgZyiTy2rttigrxFHhyKlWtJFQEGo+byk3
f04j+EuQhLrboz2xaPJLzfiWtzxLTsTkTE8Q0a7dZDEG7EFnuzM1SjY1pEiKyUygp/fJ8T49BSiC
3n0EGSIHjXmU7CpU8mDWTqP4k81xqTAlYuFZncRj/FOYjgLSOo5OPxAKIzoiOwrfsUlECg6zznl9
MEta3xKW7TAoXF+CalCTJgdX+s5oQN22oNgprNYbu6V+sLFuf01fM2FdNAD/HihCZZvUCoyp9xzB
4XwjGMhMdWtMmE3t1Jf1GrKqNPXqVHFSOrdA5qeSzW50XccZ2oO6wHAZ/ar/TboEKlwaZlihrw1U
Xj6AIajCbC1x7cVDsb+i7z3Gv70SNuPNZbKdfJBajBRQmcz8ZBXxP63v5jiYieUotMuZwrfF9duu
HKq4l4Osi1MFyzDHLS07MZ+6RjKTFnCyGuKD86K75b4ND0kkDTkbn9+tis1OTAtULx6WufqUR4mR
e5Y52dXOogkEtK5fKQE5/0KLryM8QiPTej4tlxvdeuJiRPjy359flNLufvDq5H8ZGzesOAzW+CPw
ZHLw/aExRNyAVvikdpAqMgFdqyztc7WZyt66ltPojFL4KigT7Bfmggbb32HRrI/5geNkVO0H4IeI
0LfTBf01tX5IqUypvgAUUMteCQos7AkhJ3pm+274ub1VDX1jLFt8yRK23fiVigxHLrkZDRZ2lMco
NT3hrprhuCG5nD/DKTAzOXYe8QQ1ukMPdO/EsIo1+aJw4CnI0tYKdecDgdsIIcZXhUXprL1ZZonZ
o1L8h9/YfrieRvjnid2uDNEioVbwp5+BZATDwK8IpGOsoCvQkZUCaY0/x2g6gGzA76zFWPQPax43
qaoIgwc8sSItWbWD0efES3SNqVPJ9K88aJ13cMBrtXrLulKI3X+kM384jnm4x5WSFHhm+KfOBCWT
SjFcYLPiXKrIYz/FApei51Ks4c8k3o4Jrxzy4OO7fjss12Kg3KdvleRB06LFivDLuY/b1ExONjJh
pDx41E3cX4mExGeQ1K/Z0gKDLETBSXSeQr60W5IkVpPtbT1hmk5fyHa64gnP6eG36Wm0yoloShyu
HqNXxrv/mvoh9HxBasHKujyhfgqHnB2DvUTHLffygJiTtxwzjZpY48jLBYfXtWvDAVz/KKWkIfji
mvqCYyBdrTFhJ+AI4olzMkeX2SHF2P2FZECZmoA2eeaXoxxuKpoWeezeoB0JR6VgqhkVrdIhBiJH
PxbLaj+b7LzktcXa+ITiXxdXiMrDOWvT2V2AbyMCPhrdTAMPsrWl/MSGCVzPXL8xmdXbtneWhy4B
6OauIk0mr4UggQIsSy84ED+xvaBH1/x4/DD6dIJkfIUX1Uy8LcprGXW65ODe5BJyU+iQkywVmwr7
nVOSJuMOKC0X6KplpXpZIwc1An01zCjX//0HWZPg6UX7r6u94mQpk1QYpWUrXCMr22JvzRO9YKEn
TJpp1o5y0l9TTpK+DbHfGu54IqgwVt4iQvg9ssZZs/770eqWiK17VPQIQA1Er/+Zyx7pv6Rzn5eI
2w6SSrC95Fi6bshQ1gUMQ78ffZQtpn20TeH+BtQof4TmymYPd5fWOgnDEftwfkleubA7Akvnsl5s
zTzmnj+jvb10kQNMnHBrJLbAkpRXbU81c+PmywvyOvffZOA7Ay4kcwp1OrADpp20u14UfXvy2MTd
srsaNbL/nvihzzuj1+Pqq8K90MmD2zeh2hCit56UWZWh7Cyb0UYCz3LzIZSLg6keEB7mGmBl0LTe
QUxEbhTLSwKDUOe/WglyJ42cMkSZEM0HUCn8HKeTOueNTy5LppPgbtwSTF5+ew+Cf/z46ysPq+KL
ZE6PSpvX1avodsoh4G3DTTt2kldV03Ov8ftRS0CZK1LFTWIQGpeGpGIBDx27VX0pKAqMxRyKJgJf
eB6UyxR5CfijZOT2dC1LrCdn3XDsTqsO8queos3KNXuhodmVgrIPq+azVVXH8Xl7QlA4+UiD4+w2
0maTlh2enBuIE1/PPUEa3js/Pm3mq9zurIDWJdIZkJTu0Lkf6r3MFj58xTdKo7M55VAOa7Um1IKQ
e8Nv0Idc7hVX+wqA7OsePL4hSXg/SSaKL+PCt/d9pp+uD8SRFoCEtKsaOQ3xLkaULROnR43RIVqG
Y6mCmM1ePt61Q4/xw5DlEyQeeXELMSRcsuBJiaS0rB2ByFwuDj+sionIApUAu6T8dIwgIpmPIYmt
igUMKG2N5hWqFZLO0G+c21+LMyq0cC0i0ovE+oRD4RryS4RI7sC6W5bdrQ0XEQA/+MIWuHU0at6/
dkpAdFd1Or8xhAPi3fySMpNM6+IwEdjT+FaUh7qDOKOAK0qa7ID6Udt/d8pY+0FhwxjjdFJqW9hA
8zg4hYYEI4JFli3SRzSPbPk2ZSSzzf6HDmL83bZcWE9woBPwU18r2GWRgI4//X5jszBxqNtx+Xne
sWVE5FVg7NJgUCtF/kiI43BmPNa8Eihzrj5OXyWXKWzPSd7cxPEiGl5NzvP2/e6mrGhOn6DYsLuR
dpJglamF88tMpI6Z8ZO4zfrmcvgBb9lyyIZ3XOqJ2XlJ6kNZT01jZDG/ARw+DuqP7y7Jux0q8lVT
z7gQbDpUCMWe2uGLMY6cJF7U79/f8m3xnz9g291ZKRqDxDj9UusQ1pAaffJQGkAGhEDCqrtLqdp1
MskjkHfXqI0elPPK89+i37ef57PRFI6+FyjccqXI46Y58Nz+lIRmHYl3JXMAfelaZG5vfxyIRsSr
Pr5/doNrkyTi3oYKDvgeXZfUQsMuoDmXBKUId9Gz8nFofilePEnt4giPjjPpbi2pW1Ej1HwuHiOk
NQhsnuku/bH4UdX7279mEsocyKVRvBowEwa0/t3t9Gk2TPgRVMynVH34TsU6mRQjg0A1OAgl82if
FZfglfQhmlQJY9e7IQQTtqlpRl5SQ7md4ru38xM06LSK9Yk49IrwxD6xW3fA/AwvYS3K5vzGhw40
iIxuZhKCyM6T6F21sodfvw9qAd8hlLZtm9RDlatxv8KvoJI5FOSdJAMmVk75w1OvVSseY6K8snSd
ffFsKy4wUUy29g+61DCc06gH4XZZgq1S03BshCrmHvp6FhudN1nrAhdOEgHiSf9kxUJ+mNzDybxs
ttzURXIUNZXddrKl47WXNYwTiO9qM9lCA8uJ3C4Ss1BlwfLkGlL0JbRcVpaINcxooAotL8XsYZ5u
FMEbMmQCms/9ZiDWOh+7opzFGJAnRUnrYFmoLYJ1iFW2pTlzren3OsvzEVGE/d7T1/2iTcyCwGx6
U3fm1N9PuONXijlcM+piOsOZAjG2FELnrT151pAqHbZiXYWVZgKozhSB79XJf6ZA4b3NHZY2NROn
sfopPWXGDOrJt3KdO6M4nOKsXQ/P7/7xdPi5MiqJU9ODxVo0YIZ0zbRbPEMSXY/jmkwVwE9F5AqO
ywc0lgjT/VAIq3TFEGXPG2QaVOg9vKdb2dUqoTzzD7+2KuJP4WIwDpSie0IIHumKEo6MwuWbtqFo
p579Zp0spmzwUz0SquMGlwpFoQJ5OOgbD26r3guqjLl77BOs9brkeOzkSzTALbYUGi2sEOZGtuTl
8e7ylNdY0wvKKU0ZhEgbf11fOBZNRx/p2ScbR6cAAMn/lOEnT5gpVRyXvg5v62xGKNh9cOywsQ2I
gMxHO8iQarDsy50htDTyUTMdiuuFpG9rrNjGs2cY71cwxIu+X8Sw1oqxUYr/B0P684Mu33/nbLjX
pXspPOnl507VRlUfKSsKYYa3O+HJ2TzRXG1SyuNkvoo6WHztFE7NZPEutzc6dhTjD4MINGbdsuQv
c84NCOgcZ/B5pFRPLXd0X76NzVRCVEKprjhCabRIAUOW09C3cPMtOpd4zHMPjNyrqawVKsRtLF9A
8M5kkXw+qv7X1gHJRQCZkTDgUqD/SZheZgGniwbknD6ij0myIT675Dx9lswSL2gMsOHNsfuwrE4L
DSBNDqCpbTh93xbUnOfVYsDe/DZHNpWwsNKlD9U50q/2cORPTis7QdpTHOsSk+IKpupi9nrT4WGB
lNBL8XHkW9l3gyk8AwZzmjRgWwhCaqYYAp0JxdpcaiAAipAdcHMKIPzTvDLXqIBwg5QK/NZ/Ra1m
vw5IXRvNnQnnueAC/5M0lm7NWsYuQbvQKr4TA4lbnwLRe8MQV8r4ZbV6MVFXpLer02WfmyfxOWB4
MQJVuxwDeLtopYwCxfMMI4uehG+HH2rs3eKE0s1S6SJTuOzAMq8tQRwfMkQejIvCp6WcC9K+ovj/
0QN27G32/Vtv75PdP/RWaM0bBoIA8lEVwqfpbBCfQ273w3FBXVgubX6EGSyYqaFOFmBhEKcdGIPq
ju9UyuBJsiM53Pe3NtaA+CEEz949HzzLlwYSi3cG97PpL2mGsRQBYPKtcKaYVMMHGEU/7/DRa57w
tsbU4ZUHd0l/8lOHSIljr8UaKNBliiMgWVgJV49K/zg0b1dDHxyMjdAXuWWtHTsM8p73fUHCFrZO
5C0H+1cDYGvs9p3Q5F7G95T/ZPKYv3dl2ms7HJahYj09+VyAZMNY65bno0T4HdxyO8DHE2voXGdi
/57lV4qbGuq2Z3ZsCOK0C8Ey3xIaRG+ewM0Lc+JdzGsjBUZhYCe6adQq84f+uiWdGeGZ8CVXFbRn
fhjYMsucrTBcjA/EHnBqoJRI7i1o9PkQxBqsO9Axpn5uOt91X7/B/7VVzhQjisqNmXr8FZVaNjPW
D4eBEqUKlphQYD8ypDrdlkRgWFPlcCxAc69wpREttxAIOklR3pEUQp8XXMLGJPBLG2LjhPBDq/gJ
i5n1uafBjUSL3dqG3v+sHqtDjJDWGKft9igY3LBKyGU7NUETHYfmw+kwUrjKemLrlqWMnAOCgoDs
X69KCcjxs0AIYjrTHGcHFV7DGcxzlViENT/Rhel78YsD3Pc8rutk/3qHjuJoFDwzXnLh8m4CrHH+
CWHWINLVbfZRVFcLJvdhk4bz3AYLEJD+SZIpI8Ftmm2cemJy5iLGbzVY2qUI2oiy+ZZIvHfvh9dG
RsP1kZSJzpXyYpWVtI250Kn7rKLCy5YMVRsYPPFLEuH9VJXQcMJp9Rqo+xoUqnuyLYpxf6ZX3Izc
9/b8SiKFkHyd6DyssVoIh8v38ra3Inal2Y5P9TOj3aYiqpmY/mP90ITnXtIX6sfTazNuy4gXU1t9
FmhxyPAoXLrDmTdk5JRiq5DUYm2vSwJ3d2Dunmk2T42ky00M38yDQ8YYIRtgnpl38PU78F24kRL6
Scd/eAyMeza/FzZoOEhi4LHgFK8BOTkU559EP0fsUsSVgcBUOIf+9uy4fngnrdSowPLGJDXtdfzN
qr44fhi9W+uW9K4QWndC1zKRnBRN5TpRSHdD6suYQyX9QHVgCk3tLq3MPKzui4IUJWzys/upXqjF
ufK2PmHmvlebThVIudo3T0evDSKYOvzWJjASV4eW8/U2Xh/wF7GoLV8nBIo73zrqAD+BulfQA1AI
ZhC8kPXLf7qvaVtbxOKckjdFfGRYOCuQMfLGlMdpYmPlsYAbsXjrElfVodNPu18yDBS8lAXlAzl/
C4LOeYRf3uYMDcLIT2u5DvVQWkaZkb6TmgJ4EUPayLuqPRWjbK2G//3SvW2RoT3RkZ7MGfjSO1Pk
yvKC9lff0YbcKzR3IDrqTH5vs6Vws9sCACXxsYPZN5YniHgMFh6MAmzVfJPcHBLI+/87FGTzbnYJ
9PgmmsF51Ndv1gVioDjbJmKtdIn7Mt/lNLi/dGxiIu+V5/GzpDWhcuIx38kchB1H9v5dZE/pn12+
8/B51cCIzfcJZLwUr8ZirgKv7dW//XPvTCanjLlx78XA4UTKerDHH87EIAbQcvBXq7QmO2YmcvQi
04u8VVSVouuaGrFBiztHyx+gUc0WQi6gVP46/nLLy99w7RdT3oq7JsPTFTSqmKtzRxMT/3q2GY/e
FIVCXrQwj2IvPNroFvsbRGJgui7XRSiIBFjU0AEPsQT5etQz9rkN/oz3f4Vy5gX3Qmjw+UB+I9x7
WrvreuEvFC9DAnS6AbgTNtStWq4kTvNWbg6tuvgd5OrWIjgIAVcUoaYB0xD1JhMtM563P2X6HJ75
v5vtj0I29WaAepUVRqXYo8Ti9JxuEHHuN9G8gLQsYsGrshhInOHnB5tGgEj98ft/qCkum3DbsCYy
sNIxKiDBD1uTMfKSZpspq+QAQg5LAxx2sIYn3whuaw9+n+My0ow9AsBUFr9h6FML0PTjiZV6t/qb
iwscK9FIJlO9PCyPMSIcBBMsy/SgE9I4aoPlKhT0eKYcdKbW6gAZDCWd0qSFiggd82JdCah5iQ+0
bGmxLV050U5lhAxvVY+D7Y/U8T2fSibGD9A9b5D5rnQvo+M7Mp6lONGTzRs0FBsY4w0+/tZprjXo
B5kDANLdJjJyDnlMB7JDJELGnXEiA2gqb5AbJTbktmqK9WEJ2zlVmRSHm+zik/BRttR7frK9qGKH
nrKRnOnXyUeXxA4wjKrhTWBvyJLiFLWny4TYu1od6k/F3YlM75HZwRhT2QItRYJupxIG9ydWZVqH
b+dy4wb4XIasRJ+SRQSfXSvWXj7NgY4E6MGCOliqJnQwJ+vUsssV9EPRkpaCqe39Ly7kdgU+kP//
xnGlvvuCht7bls6Cvdt2uKDahijLK6iWeZqAom55IrVU8rtJIVmCnp6Z0D2GjfCMoaoKgTujKOc+
RQI8CDPKzGpNkuSupVNuP7YKr+JMN9mfSOhDUY1jnieUC9E8CRDPyNiEunzeFLtdV3pA/OkWP5d2
oX+jWiHoif1EhuNu9CNy0nNKYaNc7rB0TsKBjW2lMVJ0DowU+Qjh9dyuJI70MbJPtyDOyPFY4j1J
5EZMAZ889vVjFPHd0DmWj8SQVKhio6LpXF6uxEkl+ywlXl1+jOP+qbyXKlj9staSiNcHq7q4vR1X
53/oiV1z+rsVo94jDLToZkXyh+nkoodN+Icqxyc/Npg4M3jw1dEcJk3aI0yhyYZeRdchTlEGG/Mu
9RkPjOG/APuYmHvK2h472TbVxolmlTwi6qVVW9bxA8QZrtVJpanO8YYbGJAtLq/cSVPq1kVfQ2mJ
KhFcQ4JVdiet0/1zrGyL+9phmL9jOV3xlRjtN/C4Icy38cN01xg2sGi4dkUQHqoj9khPK/s3VYas
6XOFTep8/r+tArQ6X1c9N6gMs3Rbh6Q2mEoNqsZ4vPgO40gzyTNMiAsh8T7r8boXIC4/ZfLVy10V
52GuXrhmEWvgb51kFXUk9XK6FPzyiYTIZZX5GS9thK+ZpI8eiIWv+GSWbdq73mQzXM7rw+HF3yD1
gntu/+WKfHffDpQyToKxDIvBfhev9L43x7GD6PHGzv+zI8h8S/qxYtLuM5kvO84Wc4CBB0Q8meZg
YCTNCgEfbV1137KvWtQbgFHA3a1ZhRoRQpWlnuOq6F8W3ZIUr2oOuq+mrWKntWm05doS6JCTYR3H
99oToSoqnu78HgT39NaH2lzFJFXvHASmowXaObP2+YP/kxY2D18qJbicYPdyWdqZR3mJTUiKgJ84
1KGo5rAqXpGRo/d3YxeXgb9njWZtMo9DxFQ2mNrcJsQpqLpMK4DklMZBwaEPFodF9ZTIg6ZXsEdE
z4DdmjH+2c5plnslA21LjVUoSEu8WZkiHO9fAyb6TJ3nRT847lPv3hPBO7rbSyQf8AznDcpeGaTi
PVZJN8+qgJlVnMJ8f7tzqkC6swIV3+lF9u8aI5XmG7H/P++zMopkB+Ywl2oNuVhE/lWmlqL1EcuA
M55zAWxYWL8RD8AllR/f7wO524mNl+I4Rh3qo4H1jqy2fhzCK9GwHcGv2/Bj3PnHbhk/RtDrrKHy
NnrHC8AL/vTgdCin9qqwZc6Y7wKJ0m4GkWKKDJf4iSXXKjkdgBuyx+i7IHtk754FnAnqXC4cmNGp
ZIULT6+NtqKBPCrw82LATqU39CiBTdBkYvB09UVI3qQXSb3uCMAiVgEo/B0DkMdEDaFv5lZdzTK3
Q6EKEwz/K4ms6U3csOJSTbxLMuE1tADpoz9VC/2LxmngHks+difDFt48I6ADCMyAiuePEJZrHqMg
1DLsBBGEjqU0rS4GPd80CBaC1vzjN6/c66bVp88NZBe8ifGZbvjkJFAMCMt+hfjIaimmmji48pot
GIHMy1tL1jMm5HxACR1vrOVId0g61tBiTWlVmSDYTSPYXX47A1DN4nMLN3+UT0EuH4WTw3LRJRnM
gjugCgcRpaUmMlmIvMEazEuAh/o1QilBcuNE1slYbVMSU4KxqTsTAwWnoQphzkFKFrJ52yUJcGYc
18LnWWKFmlJOFzpua1shfyPzZq1oeFBeM6+n2IK+O99DrPs4Kk/fUUgJl3QqzsE/SMpDoLQJoh0d
FZTafXtv+/ApQDrkhUPcY16pw0c+P3VnJRIy/QzaNjCOg9nKurT9wT5viqsV5WgnjInZIqHFfwWO
z/Y1bd/Oir/PNFiFajILyeG8vIH9qrQu70Xwm+wn3r4+J4dACItJp6Sv4bfws5V4LjmQtJ++/GM2
Ow8Rt0uwh/2JK4dVC5jwJP8jgc7ddOgk2+fURG1xYcMjVpReuylzPq4bPyhbWJBVNBSGkQgP3l1c
+riqBBRJ2ksqBwOd5DyyzGkrR9ovSDCbq3IP1USVyCmcyXXgNfsW0OvkugBkYj7gojccRd1Wf8qj
viISDPkwGAcdXrqX02wcWFqA4/gIKtnLDklUAVnSmiEDkTLr2QrkW+d6AKfXTrfooJe65K7ZXnPZ
3UeQ8PTKSEi4TakWN45fmQktyHzfCJnsZaldNh7Y6b0OeQRp3JGK65Q0vAqbzPs7zRNSqkVH0BeF
fX1tzJw11csmGHWhus+FgIfzuMxuHGHyaIsMW/PqjuB2U1QV/SYlDf2lN8+6o7rP8DW+3ceKzmtv
wrIdcoSc96qHQ9uBUaLDQ2csnApflS54AqeShh8ok90mnw3AaZXFl+hfaDGbjkji/jOLZalr4bnD
MWNgRB4tfrEpLhUAsVmuyZM5ciuq+GEVh9W3b6Cc/zaFiL3OA9yhXcmVvIw1sZIAoGEsZpO1ACNI
63uW+9AfmcJQ2n7LCQ/aI+HOgFxUDAwFXfSDMqMZ68Ti02Q4PDxaD/C0fNyUqAnc58LNJ4RlVXdV
SNq4HCIgffal6D2E7vQ8vR8WvXbcYVwDMd9p+/WSml4ZrhLrqQcK2S1bjqeN0yD2NESSOG+9Qs9w
w2w573p/Bzupuj95GeQ440C0XYVP4LNvGXB2vGDXcbVHbOea9YiaL2CULgZ7dnE8s89uSQPI/aDs
bIM4817bouQR1GbSpgDoyH8Cy6MJZjTDo3WopkFKqmOjJtbvmr3UaY0jySfe7u+MxV22jH2uBvCp
8ew9C9a/wksBtxEdFMGwgDVZggrLQ07ogK8lW9TJnmlSqDcBC10Tv/oAKTtoKPWeAciROyA8rmHG
uaKhNPe5INZcaypg4AKiZ1EjiwxYxGbx45cq1M7X/Rh4rLprXbgCYE63Wnxfdxa9ZNNsgTWpPwDt
PSAkWOA8NUd+ZGnFUzcaxHpEsrD/PqUecEUm0I0PGJS98t/jM9CbjlBBOF9Pi/s+ygKIoQBAFDxS
IOFDdu34rwPKlrtvHlAzLzyDLoMor9HlhU0GYifqfuiFaRiMGxCMQ4FLDPd+HpP/jDk/X95kiUGh
WlxuLRj4vxyRbIZkYJgljj3qVn9iUPblSTdPGMVFvED9pOPmOuQUOmUE7lXlIJ7/5w2KapYZRBgm
YsMfd5RSqhgqgGIKc9vhRZubzaC7quAAFSgn4JkhBXTmBhWv6z6L7GnmqabnJqE8iz0p6AVYi/GO
p/KOLNA4GpuW2ggrdLovn5kSfYPm6sXvDgUvZFsoyGYDro54QFCDISBfBYvb/CcZRVOqdoPpq2A2
sx5Y93SPOSVAs/8u4KmQnsIBzkGJZxREh/QOWkm2CVVHmTNPoTYREqZqSeAeVB0AqUBdzwV2VPpe
ppCM65MVPz1Nn3sJKhlE7fCEiLrwKFiSdf1jlRsddXPe1FaTTXRud6XSS59kXfUIlX1fp6E62ROj
Fewn+ld6HWs3dJTiuTv4p0R2StqCJ7V1vNeEaNOeE51KHH23MmFtk5e5na2PCQdN/g+GGlcps8Xr
4psCfc2PQlMIrY5xClgHZ6/xauvg/3Sn4mGsi2/F30feKFL+gtunvcOWbbiGr8tItR2r8GgzhlS6
TFH9UWXIYwTBMuVieS3MwterbDWAAL8/37i4InJmGS8tw1gtCX3/U/dNF0fti7aK3gfn+mCu+BfW
kW4zIUh42Aa1NlQhlCOs9Vneisms1mWLi+iio2eodvvmCqAJIyWFwQQx4KqhfKShqcRvRVF7nhqM
e1p2O8yhDj/9BJzCAH9JHAcXHSPTUptBmnmKBKGJ3eoZzK2Nhhh/PVbl4bkAwg5B98y3qLF/VACn
A1S/F/REY4/0crXqu5DbqzeiCh4aQavJ5MXNkm7GTkn1sOpG58EVYkmyW1gO98wf/sJlQwk/yzwC
HGioKzbdKRXdvacppiHl9P/1H28H8GTfCRtuvEvdMTdRCfOKspgU7WRAabJ1S1gUWigxUJ1EgmLb
8TXVBUANFKveIxmfCKpRxdjS77JT68U3F8mzbtnY9byuRm/N4DAr8G6jRZ0HtLFkiArqjJkeywvR
cbV99/OU4Kd1wHK0QNhlybWEkXvQbpe1TQ4DzebmdmcOiaSdhXdqYZjPbqsgGeQgCEy/ctOeP0sa
IsMN9C+DnyiAbTxeGHFGT/zLKqctZSxBfRXPwI7OXg2D4nRFAGHfJj7ovTKLa8TIpsHmD1ibx3Td
Qfq8Fh3hThijFXrXUhPq0+cQvvwwvMjihwqGm84WTb90E3+1yiI/sk0GEVMSUmc5MZIoOTiuJnFn
Oy9IR7Km2JelsRxdVFDCcP/3xrJtSxp1iwxueQA/BtQ+8bS07CmVctjiXu14lVoX0cHA+EE+TOcY
pN5j6LsipPxhzDcKghvSzP1j9GzWrKHXrg558oR7QAV4WOgJdC8fmYxGTVmO8b64/Isl7sg2vE9P
ZMLKTt5wS8FoB53+XmgvcZiI6W9TMGS9fLj/oM9FR871xkB3O4qrTFbTbjVYI7bgtPFCmig1x+W3
TpEq2DhB10/QHhK5OUT764IfJ/CL92BrOFtqXAWmRX44MifcKEjmxV3Iq8pqibQzACUuHOQdwk6V
E0ZFUWv0zDO2q3gwZQ6urGiL20HJUCucqqgS2l+s4k8kjhtkw0cj9ozhBKo3SO3ofsSLNcoa4cjI
8LIa+69rDMiqXUcz/8KZenJwzgO9YfxX47Y3YKYepmCWfyaaAwcdNcm+zd9aINUUNcidE0jwPRHd
Z6B8dHwCClisioGv9ZPsTcn/qqg0/2bLgR677aSd1711DD05c3+wdrB4F0IjoTp5ntYVVEdWSg+/
krofCTmocF2IpcIy+J+4Qw3eutQArhXseFSlRH0rTkjWRF6cBfL0nGo1JyZYpi/gh0Ul1nDwf6gU
qX009nRMq3CMHIzXXSFq5ET6BZlCBkAuXjGRekhLpFVfJSftFhXgv9NxUM8UsfEvnrLzKZaL74Vv
X6KfglY7xg+KURiJcMe0fTd+cDke1XVRDsx2iiiSzFlUSqkQqcS81LxfhMvjqOliREtss+5DE67j
w3SRfeSXuruZTNkFNQDP3SyU4Zronbw21oFYn6s3SmcK5k76rC6hb4lU1jaYLhSiKPafv/oxMHh7
s0dANIcMunRVNdtUDITCKOJmOtoBS88ctYkhiH6eMNw39Hiqzhl+ygdoE0QiehYxvQYfIhWUyibu
X5wqs5i0QoWVBUtQWyhFtqYLUUWr/ofMSzDbw8Xhsn8BxoW9L7a7c4tqtU02UPf7Ouo3dXjDFVwz
tR+vXRDiGQ4EfYwx6FGrgpB2AH61CguPg9fLyr83xsYQEsa++wagb12wwCxc7m13i9a6jy1pmWhC
a4ru3v1vbifOl5ljoyiNW+tTYRUvvDWz15PxF6AKA8HpkaectPYq2LMeaU1xKqI5FzRDPr6bRA6p
WeXh2Z8kC93TBbcdrTGSiMCT9bQfsWr0KxJXdS9rVeONCEYSpZwI89IjMIU02ko6oTYwUUDB0TZa
tVJyYzm6u75fTci1S2RtPSBa1jhogC5R/uqG3qKAsouDWLppPr1RVcuz7GE/Y+9h7o1Ms+O1XOpQ
K24hyqSUFyfPM1kFea2kR1n6DqyW/Hb7rZU9UoyUGrQiKvBuU517yeVgFSbbX0JXsQXRQ1A7ExNU
fKy98FYNdtYdJomqIwFkv+ela8MxGDgAU+y+FnS6osLtGYitznr19sZSVrm44sjr2jrO7Wglapsi
KyotoThPHeHah2oPClAIyRdQSdkSlCagHHYS4RtwCeMQDdJkfW6z1cIYGtzH8fML96JzV5MBCdVo
HI7TuHQCIWh5PYOVuLFMVXTkHlzZJuhwzr7P4NHGyFZXz6MlijjOFw0gcx34UPn4g1k3VNA4k/a0
lC5l6b/OCHOC4XrllxAnaxaCXT1DukjUmbEddD0R3OS2H6j8+ecCafruiGG5UCE+HsoKqVXJAlgi
uO5fiS/Xf1AHSJXsQJlZy9X4Gr7Cpv6x81jr94vSZYjxxkgXqL99J+HxlmM53gcoRUG8sz71XjwC
5Qv7lc54ZQ5AkCFOOwWEmMCe2sHfDVJURnbdaF0H+hmWYx/dK70vRro/87SqNx4zaavtjSqs6RSv
ZSIEZb+H2GLUdI2IUig9HaAJJvfjt+DZYEb+wmO5kBPeiE/uPZFfIN+3e4bZERqnnjdCBt7Ysnjo
mSXwig7yZJFbINtlQfD0KtRWhsK82xBxKqSFhXgvhCiFgeTqG6QcDHxeqTWgcZPN23DtI34xCJvx
n8YmAr8NTPI0tGyP1torGEA74WTOJ64K38CLnQM7hRmRHA7jMXR6ird4ZO5jHy5SEBbJG39Z9BXL
rzA5GEaxhaX9Nk99Y4vrEVVjjrYA2YFr1JvMWkbBsUM94Ly2fqNQNwQ0XQtZzMtXwUI7GQ4IZq6O
ieYtkZuzNcudG07HXm0E9aV2p9WLRwRlKZNLnOkYcAtsjHU4GkBG+o9PU/rQMiSJY3QTH+INLVkG
U5KANMDObnCAX/3zT2wy9K/77FDbIJ2Ye7ytOsP/oVDuyEoqpYknxxYtWiDUz4xqgCLf24krdymM
cn6pt5zhhiKQzNoe/lTp0V4H2E8uFHST/cvMmRb+UL5jMOq0G+2JHQ1iCqg7HttFAyUT4Ek3SAHn
Y56ESItZE/aq6kDhlhBjGW3G5J1qFQh3jNsZ/3QuaPOJD3qZHqx/mEqu1xZ+Nv1CPtItl89Yu+zV
bLzqh/Nqgq4SgYJR5fXkHzOJCjQHCWdYdRcf2eSVPg/aqpKvwg2KoxXDX+/gPgIiUNxukg4V1o0K
CclIqhs+HIoFdyyKszAXSdkMyaXEgzPhHTFz6GSvIyTp9qCt2W758FQj0PiXUHB4qCj0np421Rq7
OZ3fBFqwE8EBGsAdb/+kVTcW73/d1RQ6p6Y7cM0tpmXKzmDU2WRc9k7tgl5+wvqKN1fsWC8xihea
CbdElS+J1hp8frF6KJRV0Qd4deZsotNJAWybbC8UQYk4OPi3P5VZYe6fAO3C58YaSsdaCSbVp6gS
y2X6CFMX+fuGBqC9AUYQTd36Ae0FcZNcd4heQbjiAitk3nWMI5X8ZMHyHYGel0jUSdQc0ixSs9EM
INlpYkMrC52x5vuT9/6rGrOToxdWZjVt2Vul7BFdKZdBhME3vq5KrGGAhbNImu5+h9JQwTRHlCVA
oQGTg9ksa4P/91m4nwN8ZTireR0L4Fn7eT9l+b4+oUc0BlqkITazhxb2gWmDS3PsQOX5aubofFeZ
vAPjOP7CWarb2Pdy3T3uWtiUvUPpeMOnsULyxmdfY1JyqpNIF86+noW/bibYjszYQgb/hENo2085
13lCGGjHinyrnSu2inFQJMq9pgNKf+EqUQDY0+7TdxtgnYp2Hgmm34julfUhCzOmw31nYqyQ3SVw
XrwgDCw4frd8SnZf4bn6TvAtuoGu4+g3oANfpJoVJ9zab0ly/seb3AnTL6Nb15a4djZ6OaAk7fms
BkuQT5E5DszKY7w0fXIgKQyuFP4n+7FT/hQ+YxeBIH83w6pQw2Slrpxt00yVbM1AYucus8F3NxoQ
bASF6PQc9t6FCtqgNFqPaWFX/ULyHQKGALVQrevfUXfQKMAj/r6Gnq/lfE/7mC672T28mpDxvQug
qZEwiphcd8TpCJPQ8uaELrD/pwM12f6aanL3p8ZC7LROUCJx+DvAiJWmxE6iM5FTxqpJQzaWMk7t
fN9QxvcQ1YfDKbHPhlUP/Gw/YTyy8iq49+Xdl50u/nazmZwd+nrmwh1fv5UsQomg6It/rPWtPopY
QS2cK37V8NMTyyytZcUkLqQTZVMOlorVaLEv3eMmIh70e3DCq3QLBDBxQLqR+xf2FZ5oRB36aKyN
dtGKqznv8kBJCPgmK5oVtLxTn/Hk5Tw7/nHAlDF+EC302QPJCY7MZbX4SjwRtyX6VMcwSlNvW5fg
yNnxBDuW5E0xdgYr2+ysE1JPmLC3CcTET3i7t2wGJNEzHckRS5M20sO9pZKPEQk/+44gj2y/54RO
3AdVDsB43/HZEB0F/JL2tITlIS1MaUtr6RDgqqOroeq7PuI0Jssr50kkv3n9ae+Q40keljV3SvHi
yJnAEm8djv+H9nK14228mtXoRctjb+H0guZSp3lOcV943hWQrmaaaKvV5M1LnqxC+7FzVY04Zcm/
BEMIKJArl2kMZsDLVnoldnDGZP80dTsJZPnglAU5V4qg03wJLSbakE6DNOpQ0Gfv++qwXxXDICVx
NNKj5CAcnNffbOEOXcemiLNMqNR/DqQiApjsUoEUd5y7w8URF6WuHhOIns4+WQ2AcBKrSOIIRSYz
bkY86D6SFS/XArpeBWRDmxKAGxcbJGsEqXp4tQhI3xaMuiIteGvyF3SrSP1mljKWmzLP88WvmXgt
lXDXjhJg1OJA25mE8WJy37LevBkqsfrMICV9woIELRCjhUY8c3CU+KSrNybC59YOOFJ6MOKCGTDh
v+YcqdE0VK29x43rWg49kxM6GXc+Cx5ov0+yEfkcJVCCK7A0QKc++rFqNHGYimgfNDi1UQF4QKt7
xQI7haQGXuIvBXtsjfvawPvXjSsdpLxDEdlwoP073540Bd59x7s1ISWOyRh1uJu2OEnn6HU0UQC/
w13jZPb2fe8vToZYYfyz6rc/pMYqP3Hm0/KAm2+DQv1a2KdkzPzl55igryixjgccw0by4BVZpBFZ
C12KVUcrmKGmJDr1sq9nJg3DHx1PwUjWY3Suk4fJZ1CIfxxOBagCt4fQ7RdcS6q/ZjzSq/0K9o9D
v71vemPZW5eIDAvJH6oQ9a7GmeQi0GqJmPEOhs+De977UapX+m0Z7Iu06ubH7bEkXczkX+PEoaNf
QKLs32UpOydnoZamjzPhMbKg9sIwA12tjP9Z1TkRnw/BIim6uq1/FArgg+lCP02nM4O/lfXT+Ncu
6mBRy/I2V9yKAtK06pQ/cd+UKexIKb6NkADutV190HzAfMqCfXkMy1yBWmG/H42GKdALlGt8Hq6X
ZcCcUb/xivCHrpKUQ06Q2ru7siflvuC8+B99KQC33FdgPBwF9LvO4A/N/0XoiqfntsCjjNWTSEot
SGzd7zOVeIi83VIATsDAVfFG+YsGkb5nNE7K8ce+iXydzdF0dWZlDi1ReifkCjrV9FlXvct11MZd
1SpR1ebUVNvNEeh68g77Q/hFxjJBtaK0Jwr6H5kAcB9nMbCUxlS645hof7TgpbJasAl3q/3Ahj8f
VdW+s9FC/6R4oXlkvFS7cSmob8OejgYlN/ZPbS/+zwuIZBl/FYbGsKb2Wp5cnBSFYgGZT4wxa5g3
Ajxb3KEmtnpLdxKw6qn5kFAzQqpVxFF9C3nHBLmZqorDA6p6iNc5vCgxMimynYQWFgj+nvNxjmPi
mqgdsnWt2aKJRcN/HO3QfBNkiwngmfMKnanha10z0NuvuOM0H+fSYdOON35awa4Cdjb6w6FrItRg
jtu49Ss0177nMr/iUllD1u4WcbprlRkDmbqyBKpyzaWS5Kg8Lczldeg/ToC1rb6to3Nzij1fQsjY
GHSmOZtdridc/Uk8K93jXDAJPLthwIvvPt4v26ipHZ5X0tLMee4V08AulWuUIIwehqgvY9+2z0lm
X/ToqREu4hdsLQBb5td2fIrnSGxxzw4ml0gvTUrdUcQ82VmhAVU1nojb+Qbq1cUaenKrH4wEncBm
aNyxdQHc+KKDTEjQrW/iYAiVO41qVsvrC3PNmB7p3d8hPfJ+4zQcO3XzEari6SN1SLTGAxrdpgBG
r8tSIvAIRcY73kPEZR3fwOUaRVc4+K+sF7XnuCDO9y8epjlms3GTaQSoSV07+L1o3XHzO78fdixx
Vvx7OphaJZtzRJ8swmIMsGmnTB6m3ZMw2UtJrXaPMGNvRSBWTNmq0jY9MmdGQ7N20KM5qmNHwXPs
V2zfaMRdVmpjiianOUxIVNdCWIcaFhXhwL+4U8xYtkRdvC+1pxOXRXqsabFMWcaisnv3MNvZuaZU
lVQv8VdIzzNlmQRLnRLXBJkXlQsIkohR3WEHIe2YxUwncvLU13fhciTVGpg/lFU0kngbF/gltgKN
PZWtshW8r+tGteXAPNpRQvbQ7Lfqfxql8xyHggQZ1PFUCttjwS9r0j9l5zck/32Hqc02Xxn8ptaA
DKCGhZFamB7vPN2om2G6Techd/9GTWxzP9nN4T4vscKVpai+Iv9uqOKy30aWk955Vkc1shOtUjHI
/LSNYrL1dGBIlIcqU56haLQ84IamuWLBnWkpj22QLGbMn1WCn5phMR8ICMpUbbBzuLmpgXJrBY+k
l9nppFaC3JfSmD0vRGcIGgPqK+2SVleBgeDh0XKmnVTlgVrtnyWJALAT/wtRrvamCJnzum+0d9zb
SLRd1WbkZU4Q0IBvtdWfy9WLSy+LzvP2XUa1K3DVx+baMRuHYfGtu7ukf6V7fOuTAQ6oXAITHXKr
ajZ5VqTBag360ICF67jJThA2jIJ1QC4o2ZkQF3SSprskqfut0Cc0vjcpKdhLBlDGuMabKLoGEkXp
dusKHnZfb7M2cIezYD68yAYiEzHY29l4YHkulLicCWN/cJDx852kJ8TNM04iCg5P7/faNVAe16rZ
q950fVSF8ABsHyZENTZMt4+W5/lV80mqGtwhK+N1BN2bHhbIeTF9PjdV5QWBWtSeo0V7SnTzhgrq
nTGSwLol1vdRV5l0FBXh158JI+fQJMJAppK/I4DulutxxCIUTjr6WYBgzo1iBVpodkhR7uEgt1JN
932jsSO8MIJbTWiKEg8uEzNawC/aRDkjDbc+alu2btBlRYnlqqvWyakiR1ew9Mw7YWu01IDoTDLo
LL3+Bmlkq9A4+MozA8VfH9xa9/HgV1RyDvToJQtindZcCig0qccTtfQe4JrLTZ1nIgaP746thhJ2
ulH6nWhhwwj/gEbcbLaB94bA0HnXzsljt2wuZVATwJdJFvCRBHm+b5Zce12axFBv4L89IaD2bLPm
Io5UDUufhiM79XXl0iQRsB7OJwApxfVEA+Kvh54CE2A8Ob1n2stMPwWwOAjfAzCUA6RczIhpXG5D
enxuhDjI2vWq8vONBpawrPMhMwZyuMLFAf0ve9ZQiJZ4XXbFy0ilzEAJQrOUJ7YndPxugMQssFWH
USq+xh6RtptDsISZ2HxjHlI6xrSzea2D9unOUy6Z5XcfoO8FeHU7bNaWf7RIClJoS0XPYtx61NZT
hSaPaTVb/ZzWyLqTgeGfupvJqWIlZVGT3iczWuRdUv+kvyQyqDve2CLHVMJmwdnizKiGw3Z47uvL
mB/DQ3tcrCyIMWpAbu3AFk0mhnvdbn5u3XNZjvXrMlIttlmhrxK7hR7YawQUDrLSWC3TlUNhqSfY
+EjhGrVsKzCa7S7zgNJcJLK9238JgbtO0AE1cwtQqgGOZ7uVLEbmPWP9saQaKAqU/6ub2hB+YNAk
/B4X0kxL8LUwDdI3AtwT6U0CEiNqzXo0IUtH8Jt2p1FAvGP9xVD2XPdyamc1B52hD1IRZCL6TOQo
jz9q5ySqljsNuo0c+ukR6cLeMFaiU1AZQULknty4UH0U9C+lkOFrWtfMQ7xe0XKcndHJbPNHbERD
i0RA6HWFcQxgkD7pF6sW3E9BXxJaDy+QJzZyhY/fctJqpzTueHOXeBheZ8i8jDWEzBGiStOkQWAo
bNzGg05I9P37sIuPPFdo8h1sVI7u4oN/oML1J75+XzUQCJzu7BQCYVvA3W9JYZ/xsw/DQbYTH3tG
XDtrTihStp2DRR0RTP1RJdeiDIOqrWQSZy8DyaK1KDNJqUxoayAqwTWApl27AiBkLH6S5HidCfF1
fdFTyPNmE+NSaHWBwrcgW/h/PCcMlRQZT0MsI5MFt16o1f38jtUo+QOJmGoTIxueRw46oAORIkbM
WEHByolklRCRXNR3xTGnjjHm3lDQGKTGaEbDVh+5lf8p3P/hPYi67An6SjnzH94twXQrmbBtf8Ea
OV9sB457BjgIJ1zlQSRrk88pbVklGm+1oZ5RVhN6y0RRbHBib5jv5pGUafVQSYUH59RQZUPo1jgC
5DIm1Zj2d/9Ph3zjvPXMV+H6VNmoBS3kgxLfxA8aCg6q7LH0h3o2iZZBfrPIMWxI7BJQDHHRCS+y
UVVO7pdqRMgsWoQf3gYLsQfxONRjLPxEQ1tjwVbzxUo6CQdZmN/l0USfkKQYe91AcE8I8Lq6hhdy
CAMNmewg04cqg2aKLvks8eArjr3JdFQnjthFGbRU5Hxj+YA79AhnhGDe5d3EFfbomph0l68105s4
Fwzt7Q6YvqTfEZakVDxQxfP2DVbQp4e+kAkxf1shJjX0AiCPOsBl8vTfCpxtuxMleGwGRGu1kY3L
z8AegpuKJW2WgPN+eQffreH8OS2sGF9mk/1Vhc8Vl5KnG+dMEkwSXzgAGbyJ8iqFUymnc8LMu/rn
LvdbgxCDvoLcDKQ4XyZQqIM3WUvqk460CJ3YptZiKPZ2VtGzeSVHK+fSdTNi0hIhZ68Pwh1eX8T4
7CT/+cfB9tYyWC1lAOL0DIIOgXWEShb37UrYg91/ULpxRZWK3q5mv0GYwC8zxq1WkJG9a7TKzvli
pKF+aqhCLp4hBm4zoVEeWCJJHvviSnB+VqZuDu5uYo+0yNXOAd9iLFRUTzIvjIWC6ErjGn1S12rq
FsmcuGfJqm+nXogArl1ue90xXDf1/wKeV7DSogufKijrVTr2NPyZ36FpyLdyjK3lhmkCfrufD3op
l7hdmWw6AfoR04BZ1t4MTKWfh/BnjI1jalWNawTbQDekkCaL5mT2RNM2mUubJNm5uhjIN+qE7HfW
rwDz+oWlUV9YgTWvPjDINgy8PmG3ow7U8x4FRWiZ/OzQ239qndlpDBC0Hfx4XXK4MyyyyG7aswes
9e1tJtZKwUVFK8dgsJW9Cp0j499Zr6mrfSM1d3Cy21ApwmRT0pXKTMizJ8WTmv1j9mMJIM8+wEZD
+cGGida7c485e7WB3ZlIiLltckLmFh1uWbQrgW+UhfRfk1dHgAaewsi/ji6OH+3XxwjHG0YS2TLZ
e+wEZIDCrbNLF7Y3GswH6D/rhiD06N17+VHg0Yu2Q2gtHd91mH87Sbx+3A2Ktue66ktrkPd5oGlV
oJT0omzF6A4mE3CR4btjlSnlzqDGRE0iI2a7wHSxnidhVyRKC7b2jq2jfnYiDuFjcDs/yUZpyppQ
fg+g66nUm9YqfZ2Hyg/H9dYRDURKIaUygdS36pt21rVHlm5GqLHuK/BZHIBwHhkDqduQONSDNgT6
EiXLrfNNYLICl9VvY5EwwLtbK1dDetpL1m2/U0SlxGTskS/FNXvhiIMshH9SQvXCnpAKFIFe0tNw
bDYkpdxcx1002NxuB2gkBO5fDElYQVtjcdAPLt1+E93XKOTA3e+nOlzQf8RUVxfCWEd41wqmb9eu
juY/BUGYBOpHEVYa0fFI72kF4gSOJU4xgoJZfn18Vd/reWR88yiaqVpnmyOw65xlPSGuzKfjftFL
bNvQAJG4HyvyJHpaG9YVXDJqQ2ySJsFknjuhAgqpBDzcUtovwDONdzKzPes/CiesaxgohN6vYKXb
60/1664MUnyg79wxGZ9TosuMGeavggkFXca76fAU2oMTqAyN22TMJ4QXltKnwLzmv4w/Na1niYAD
S+5pDaTbOziNEQH4mBrIGfYJqDS0H2WVHOR2lXeGUMwGXm3S386SviP0pDyvn2nFJ7OdWKwWutNv
6IFsuIulStqhX6pFO6Xzj4ii64ce+jnH7nkEk1uyMa37L16GyeeZNIJqEmwouYNLw8CCxBgUyY4O
12bTHFiXnWAQNmMYIYzX+RuTymDNVNCHxw9nhuRE2CmA+jPwq/d6Zty8JCiJ6ZRKyjfKB/kIoSf2
pIMp0W87S+KM9S7DlRKwU8pSlT2QHvLShz049RJic1LeYkNlDaJtl9ZbyIkBYdgELo8wYZMDJgdK
s9yIYCw5mVeqSo0evccITCl3YTfkX50dZxJuhhcgJJREF/fDP1kpxsh21E9DDF9Z+2b7ftLS4b5p
KlywUleKMjrFDJ24ue3dZuOc4GTsRVS0sRU2YjhbCHSj0/9f5BAdi+bmos/3EdQkP/6K3C5uLkuD
5U2Z1YX8IIsH75HhtStVX92FiKr3tpjIax31w1Vig2tz138algGcg+OUkYUxLzmCz9rZP3/BnjOR
qeas5i89+3GKOtNxBO5nEQIMo93lRy4ALV9fBsfEZnDqD1hWyMqMOwQA08jezeuVsQXPRCQg9304
/5/2rNfz+b2lwnLfptBVjkLA4iQhE0Gyh3XSNjoLKbW+0QJiXaq8g4+xSedhwRe6XyYMWElIXMS5
p/uuVlo1vF6IzzCdZeH6sexlFQsX1BtUNrElm92qXZ0ZlKTr2GM4yZlQO/mOOm6LoJ7FTZbv6Ndd
/lRwqDAcG7dBHNI2Oitg0hL6GVJcH4/3wrSCSdRXnK6WgWLdOrqVvSs5LcuAX4epytHPyH+J0KBg
8T37BQH/hmL+I2eWjBFDYSeNrPhZkWtD9NolwY+JEswiU/u9fAZL9mtnnC9wbSajE//t6HkGZVdu
YV7zhWiSfiqK79aMwrG0R/q7+hkvbU24HTelnoZ0KRERQsditr8OlhYy91itLa1VOF2/ie7btcZ2
e2eJIcDGLHZ30cCOvN5RdbI4SOo5j8y/WTsvaaNAZde+0loWHUOUjGlCE1KLSEgOP72qWS3NPd8V
rMIINOsyMcLfr6OXyKrbKsRS9p3xpC2iAArwkauzYfKWaLJW/TnPfU+0FRgEIqaQ4EKpkbWsdYYi
S8SIFuUdm6VV00oYAp4THK01VXUdEploqG3/ki5wn7YfgCLAiDQYT4CvYP79UkDq/ArfgZfxwb2o
Hl7PMhEVJjkwbAkVambAD4QyUrY2fdgoK/kpa4SXDgTNeog623W2DOUo1yU65C1dTLXVENaORrIu
7UOAKi66vI7b9ahkSHlWlpOLOJOJFCKctG7apHILhXvvx5ITHTQ9nOOG2Dur4OBSpzoEzKKBqhgo
PsR3Ui5WXzmvGqjpX3Jg9EznlXJa2ke7dKpKmWAR2jwsR7T0kYVUmSfyEE4TY8tw7DRg3as25GaN
oDWYJH/rcaJ8ZTo1N1j4hfJ3RVBYxh8Av7BhKiGKJUl8OsMoT7etn9KoK/IAaTxGrvlmWykebIPp
qTU5ZGGH8AqVHFRGv1WEMHhF1ViVR5bVkDRXnFI6jZdqnt359Nu1ygG5mza32ci/VMa19RgDrDEO
KgSBksiiVEwkE0eI0j5QK27y0JfrfgM2Czpl7OMUzsTbahZvcSzS+/XQ+3uuJ9sO96s0JJRkAtdB
0q7kqTJzlUC58GPGwDGSpwtqPOwwMzN08nPD6qSPWmZR9WFemPF+HaF7noKk4e/nxczlAXU1B69+
cm7Yn/syareTx7QFChTCvG/U/KFRlGfZzc7IJnouCZHQCA2JfLXtT0/IS6tJS/FveMNUkE3X7qtQ
2z9aSDP9KYjZS70cOW0MSZYeR/YFC1iiFbIuhmSHbuj7cJmmKac90hCzO6PKRz6ogJbZa0BEIKV4
IhugDPUXlUkjiVXSqtaxSLCVjHGGdMcl4FlVg8k0EXDpdNcrWhmD+vUViEZ/glAlQnkRBULoMqkG
dijOo1/Y5qFvz1CA4VXq4gLJTFfQerj3iAOm8gtehVwPXifZ9Ln258WDIrgQ28fMz8e/SrVZBm8Y
HCKGASYIvom3xaVEa/XxddoTivKeSi+B3LmulLPVmWYwkrilyc34uvJ6MvyL7ODkyvGsmg8psx+5
HTByspQApd4Jz3B59BVExM6xQZ79U0E+oxS+X1UIFJ10LACNSDRa7FhwlJCrdQzwi1S1JEggSRuc
CsBehuvK2oqnR3itw/sPQ4ApVOWltuR/GtpP/SdEh9IiTo7DtMOkRjmQLZHvHL8WA/HLE8yxpDCy
acxLpTFxy9YfpA7FXd5TZoaN7jBwaZBjZQDxi+rg4fvqAc8DdtW4qxX+1UDYC9CN7AXHyFYG8PlT
eRzlzIOjtm4ocpoW0FrvfVheOq2gNEwaLTaqnhhtGtVTKq5HDD8j00ITy4jdZ4azDKfsOrzDrFuE
9VnSwW+/fAF940HJVWOeVDyVtxvm0px2i++SiEm+lTK6TP1jTz4IF5SvbdmYg8tQOQUIqKyy1kth
NM39xAUUZPKu7EJeuuB6xEt6h2W8az9o5yyWpGLizpKYM85r2wtfXbPEnik0YkeKYs4qHpa3c61Z
tl8k/+mvJuIZAwQxDl8aXm2eQHQiukdqRJ1nOr5oxKLCh6CrK6NaGBU5s/00KUZhbu69yPc7G5nm
Nsog7r3qL7fxdqNyo2LsGbZh7181fKEEOb/padHp9zH9E6/ZeuBg2TIEr00IDCDACWmas181zW1t
R/JFF06gOmLAxiizuxfwzyFUuTsmg3z5178IUr/4HBefqgpTx3/uJVa0c2tkDCw3BKcdCQ6wjwsH
LiPNFaWXwynyj+9guUclh5Xyap2XJ6aeowxpqT7IXahWol6M8dNVrg9xRJ52pf2OH4G3pZLKUCfC
mw7doorJTYEU/q4BpmiGCFhfqRPLDBcBTdYN/TBkjWQa9hn7qf+G0p7gpD0Qt1dfH/V5wgja3n3W
Y2IVuc4dpDAtT49qGVhVNqYFsb+qNHXar8rvSnHmrGWWnRwZ5kQW3kS9bGQThPfjGSS7Fo9p+bhJ
hV1K+uuYrMhsgXUKFgTM2aWORagBw1lget4+umWNfq2cmK1WF2fP8xjfsVXHwulQqAsBwvrPx4O1
QddOYTqLo3dBgqhV70B3J9QS447j1v5siuYJgprPMZ5vmeESHKZ1AbYCMRoqCpTiyETW6uDPPDL3
ei2qh2nGqR6/lIrnLWW6zxUK928zljI6LVIndTeh8iiyhJLDkJhuNCLMX1wtud+QKe5YjqS2UqfV
V9mFxeykN/SBspVN+cjcXO0lrW/R/0nZqU6OsrpfetJqXFtu6lYmgA3M2rYele0vXimFbpA/wT0s
iHfS2Nk5nFI4lVIqu4kHAzwgR4IuhgYjHT4lnNNdtkMqsVueBDjeX3x/9BaU+k/97HbmlEZRj9wS
SSRVjtGCVUD253ggAd/rbboK5yJncOQU1ok1S9vKf8dFNQpUV8CsAt7szfYz+x+MHPDxJhlDfHJD
3Uul7mX8/dMWQm0CXAn1cPnV3Z9BEpoEV/RSR49LstF61HrLCOdCTnvbYwc6eUtIWXJiEpX8f2Lu
gncstIK5Hll+esTswcAbUlagdMyDavseZfEOhpqyyBEDKbkQAyYH/EFd1dKbr0h6PZKx7PqUNeGv
X1C8dD1F+A/EVvklTsoQfnmP5MwQc98rW/6jU7eZNfPu6qGAp8F0YhKmYGsYUggr0z1gXOr1INZ0
95SkNt5JxKxst3vvxdKL19ocZGShRgj9OaHUX8yJVpK/PTTSeNoZLuXg81Wb+z+VIcGl/+Z7gr4v
+UEEzJ4Xjo9IIYP0i/b8ceh1Q+qAxIsHcbLQugyZ7fuaiD5hrfqqdebT5gjkyx1ANmQjy0gqzaam
uyBPDXF5SLfVzjccyKu2tXUuInVszGyarg3d310dmmbHYdXfDNMk62fTY6mL6ZDZN8FPYQVOUfeK
lKFyna2s5Om5xvkqspOx1q9pDgJILV3AKhnBtpTtoFu9Dfu8aSL12JtzJo3LtfztwnY/8E5oodKP
lH3ngP0XPGyINH5o646JW3WOgbwjp5ufJgebg459kH+WxFwe4jqFEi2wGtTwx5SqxV6SIElJE+Nl
csBwVyGzKUTN5XcIKrrxgqAgSEdfdBQnq77H0qhon3F7dfH6/AkszssJwkWl7FNIbvyemEv0p3Lh
x5HMqznCRVUHDG6A16UgCDobXcQMLThu0wdEhOS0pLZz6IULkZRF2fzCxLGwhqpM6Dq0h6Q5DW8+
/NDI7kJhrFlHj/QlxbrpBXrS+Lju/nP5Xr++O8VggLSuSKAUn0G5ly9kfRoa2reEvtHvHCK3naCe
d3iSi+I4vbY6t86W2NzIIH+/vaObyx84ieZNBxlyjmnmjO4QCXMRep/l/3l5PgSOdC0y2ugUBVh6
OnS8jtZHCm0kHLKGz+xL/LlCYgftPUFaIweKBcxopvxFgljA2+FuWZX6+a+WYWbjz78B+HpAjr+L
dcviP1iCXbA5xH8F6jmuG7zPyf2OoMCKgDVw7fG9TI/mwWQsiLkcGLw4/3Lqa21uNxPX6k0ke8HQ
+NjiGZLKeQQdGJUMJws2UKeSTgvMxrQdHciBGfZv/UxjAzAqBKuf697nJI9c1CUYM0ghkODzA2mf
WH8nb2Xstt16s1broH6nvjsphtAJ3PIhJSjZZw4v0HKxUiAaBX+/9v7iailq277Fl+o9KPtrDpkY
f5m0KtxarzCAPX6dy5oXVyOF1kNQrJpYVY7wjHGPVB4W2IdWL/R2uVb+gIznvsffjGh7CPDdlLDG
IanPMt7efx4oTJ9J6ZGqoe4c32rmh1FY7d6GeYU1AwTWwd8hc9S3CM2u6b0uMUXjwCeg/2YChuQm
XmYVWZ6NTuRvsdzrF8QJKTFMnDcOyTMqC8TZ6gouwXnWp0JEMBxaaZxxUxhOUSQtXdf7JkxlP+ag
uJn4yfBB6ZvXpDAc4PdKmLXrBS+sjaxjyKL5umuPj3rAbxj3t1QqMcCHrBu5aRxj4HtDcBHMRAj4
qRAtCeoUR03AMN0fv1TUZKl4WpW337D2LnpIif3K0MnG2zvduWGkSYVheMyC23mprWZE6yAGwapo
1td1d3/3y/ROCzYSsmUOKLrgG7Hv1mf5C3R1S9+lo/B/VjOJ0vkhhn2Ovq12NBLgzOQ/ubPi/VUz
nU/z1L/ORT7jpykIZ9KuI0/CveUZCyGN1GcJjbJTXO0tn58oOyf9+eLolRgE/iAq8TgplzjDm6MK
1WgpsckF7UzCwVn1ckuKpX/Q4nk6GIhP9bxtbz6aLEuUYk2sf1EXOeJ+aGXEb7Rj52eT9BhMGTve
K9FXNY0vMQ867n4H2hc+ZVpZMDZynubk6QsWmoAnKkGHd/8g5J219RjobiMIruzVYDXA0A6Nh6Bl
zZ5vwEydoEtJHbI3ynOm1u8VMWQ0YgI53vo05ZDzUkrTvUl8AHZ+U1KV/sSEc7i40Y+XeYkcM0J4
910CouqdPdhEV0tTIiI5DdWeyXUBhwqW3Rp/hExg8n4o+gaS7PH8Of4Y0K+06feLUY80MO8FiDqb
sq8P/bb9f0oMQrmmZ0wSq2uTo7cdDtd8mraEiFCztQDBuXDQaywOnCoqNOltrJPKg4xW2R2p6ylw
xR05QzQrgMgfOIxwcH6xVFfo0iGvKagGIYyhy1Wx26Go08DzRdoo+ASfq85fZzBeewEURMvlToL1
09m1Buc1R3zRkN7X4jdGuM9TD7gc+i6cgY0PwtLvwJKZF6jVoQ+3TSQe3qpnhXmtlzL5dIumVC89
k6GfW78RtGjUND9I9FblaFqIhCmc8rEEB6W5ramIc59XqElkIwUQZKYMWo44TZ4xEdTovQcIIhb7
Z5DFVHDzV1V1LdvabaBR2upjevfJGySKoNHcUxE/kqESpU0J2Wy29mlexZDVwxzUiHBsyBRKk24l
5f/xBaJoMhpbasZ6+DSgh/DxFvgmjxjugCzmi8fC9QtsFFMjqIth0jvmR7dTkP7kKc3MePOnuIfg
kYxs3tsTgoHNnHSXe4iztol0ijIWycQSvYJU6WpE+Sv8tGlMj7zwlkMUQp7wJJd6xFycgtBbt9we
+/6NCC6FN0NQXaZzyGPjxnNdRhhsmXuQEPCNHT48Ko3+wy6oHWOTUKeI+8GokO3IeJ+TvCO7+iuY
hLEvmgckiqIltIrKhzkLmr3PrtG3lu2dplHCHjJESiUsFuR7SVpv31I+tXm2HJGQ5b4J/oHNm/qO
11O6SBHZ7eirvfKlYVxKsemL32qnuxnJafKx5n2tdEntJYT17D2TPfo5fLZ8NcEFpFGrH5hbL0A8
iioMm77XFl7zVyQFKRTgRoH0XpQnjfS05y0GWc6xtyO7OeUWiGtgBT4C4RX5YIpsAsb8muh867S5
l6TzpMhLLzGqn4M9qLPx42cR17YnGs8QGkaRa0wmuYEKw3QlbYQ/dZEeVI8EecccpuhO4/kqrmp+
d9IkF8/13Rg5t6Z4cKkHVDaW6RPjrlMBM6GFSqhOzKgw+zRCnRl8/m1kMdeJjt4nPOmyuXwT7fCM
2JZoyNbC9bsj7frkEMxkIHg++HexbvcvMq4U+BOO464kywXqoTBQfp27MPIP+KsEIh+bozGrNsk+
cPTHgdWD+Ofh8vjpm/ebeD1GbPXErFoYyIQLNDgTokoUKmZ79lqJ/wBJHdfgtqMfPe+B+SnVr9Kw
2FRd/F8gvCSD1/lcEL1Tg11l00QWsPLhER9wczQlKYOzM7n54xf19eBwM5tNFgQ2t1lmKICZoVxb
XEpknRfec/028U50QHQzDLTCmV09XRuoo3wX5XK9KJ25LHz2eS5Y8l/uYflUcn//7rkGV1qF+4AJ
nxTiygctBTMuy7NVEkpqpi0/BkbXgcuDsAlvUOGQebxVunFWqfoZlR9LPVaFqLy9jJldo4G9maYD
TZDbY7lCFU9WCp/y3zrwnLQyc2iFBJZUmMQEtaGECWUwLjeFaAVlUYo8xODDkbuf4VVDGgxMQn3g
+Q89nytAniFP9RdwkGZxNvobjTMP0fMpucPTkWJl9qlV4yuSAGIUfbF6euHpvgY/rqZAGwBEGsU5
oOmfDqAMU9xZLhBHl53hWRXof+hotblQ971+4aK3GHXZKyZap2f4E7q9Z+M0318eQAVGjTM2+zC+
81WmIJzkVfJa2ydziFvh6NEJuanSp6n0dRcRFN4V3kxszAahpdoKMfdt9I3sNF3e/5v2UVQq3XCp
r3pXrvH33PGTBIkXJHiF1DH4fHTy98afiBkDBkknu9iHJLqNvxlTUKGvs058UDkUw1TrleJC7ZI5
g3bBPzxsmCZvEwlgEx+QlA1hIt6b+CEMgXjMdhyplxY2uG9N6EqT/FMcsDs01ucepzmYwfcJTBBh
44Ub9WZfKOZ17RwEA7y8vfc5FcrnJHkNIqkLAHHsxPQYovg2SP+TJVWd39JlYwC3es2RVy5kb2SK
6WBIbTezf55XU8A0xOcncSGdUpczs4x2zuZNwmEirZmqR566pcdpCi3OmwrR56UFat5tIX1nDmtU
Gx1NUw+H0LNWwL/pwtXeKK7EW0Ncc+N1ObfRQvw7J3YXkKSoB10hcRE8TexhF86icOFRjtYWQfZL
4nPkte/A5SlE57e9pF5aPS7tXBl3BCZto8fNWtn8poauHECQaeojJMx1y4oJPQe60LTQeQ4wgmcz
NjYDo2nakJfsR+kfY2ryqxI9Rw9eOBkHDX9V6Qwicu6ctKqKz7YPG8uw4hxu+eIjble/KD3dz+Qc
zvDnPSsx2FJ8pJ8EBu7CxFA+eIdOtoPS39GNuMAGHVk7jaNazSY5sFA0USu50Cd5MRu43TfS4OVe
Nr09hZffvGiJOkLG7QUsvvlnkKOILdpIYbhyH8E9Xb9Tyu0OrKqLD2xC+9fC9o7nzfh8/1PNRZ9O
eb+hELQZn3UtdWk/v96DLZ0zWos4/QJfLAsaUXxKXq2AnntnEwGp2BarL4a55PU4o453Z2tYD5zB
o9d1JdEL2qH3LMEFZUZnL0MI0SPZBRyJ51P1aHCYA3w1qzyo0UGmwYdRrXeQNcOhwX1pIruY+nXZ
TcXXg2Jwrb9CocIc5XyBKJi8867RClPyJcVHXTtUvjxftZmvxef3H3De2zoC9VCrQTDekugHHMOq
Y/Tfpt/5VFvKtOlDLccCBbclC3dl2aEn95amoZ6rzt6q4ocLArgJlTbCSubP4pK/1dDvv89SovcW
omUlxlfLR4HAqVcftQlYMBc4ezxDAXABdfvJyEeIeMArxeeXLd3taANPKjNCb24wdUJIVlfkSGFg
4Z97dP81JGH7tB74IWQadX9Hvu8YcT6YHCS1iRdGHQQDNkALw5LiC5+HymCQqg9/5fezr1kdaoiq
tCcNv/HdtCwUl8nzs1HwETWzTtNJB1kvSWJhGybDS2wZBD8MlNXNNXEkOusq6ofHX6woquAk8eU1
6v8AYWkn2ms8czsBCFhE7irMafcqI0ZBpfRd9XF0aG2qsTJJdwe7+y8XCayN/F+2qbpIiu1VgtnC
Vr94Bdyzs3+hUEodZsH9Mo2cLsCT/hDyZirJEx4ls2vHJi4SuPIcURCD7Hi0pj/qasz7YAq84/rY
ze+/iO1NdcitYOgsi4Xb+JYOmiMl3hUTFY+OjaF/xWLNxC3zQ1DLY2ukkCmzh0EqByLAA1RcennY
qDb1J80t6KHN8rzx+/KKwEewKUbiviUtEVWTxZgMG0jXlXIH/TKU0TAMfWdHY2YRozDDtlk7iNgo
dkPUR72ovM4/encB5eVzk4GCsUeeCbx5Wxl2IujvneQ4/AVRxswmJvEmeeMACjYetOzjII8mtxFn
7qr5/RRc5d26nTLbZfl1q6Lwzoh4JN/Bm9LYFsS3ZrQY4AUYWkeqdTb/y/hRHDt7XN9ZVU7hs+Ma
D/Tqwo/0IsIv2nFD820LGfGaQiH5AFxW9b2tNO0LLTsS364/x7+sNXGkAsHFXHNKT6KK9si9WNHY
3FghCtIGUEHlwNL/ypUpRUk5Ad8N2ZXctBLJGzQhSFFNrr7JBP3T5YlHcMEy3mnq0U09V66PqYAp
o5UrYzDf7h08UKW450z0t4+DPjY3ocT6+N++rfxRinqtcbVlBGd8XvGNhz2vsSuvpXWcAVlllI12
2CVio2Up6C+aZ7SxrE0OKwpsTu+iJLWx5kBR9NHxVnQ2ENIZNUfHLe+gXW/gKVVLFoQrPgxOrwpa
+JY58bjx9dwze7l8nmIMWleXDGr+Y3VZucuauvABc4I6afXOE65d178Ynr+ffBagMMnm/xh8QEgS
sUwyIlTveUKqn+YkbDX6dIXWEEMdLj3kj7e/X4cDv9PlNnBbMQXbzmvYe73PECqTmL4YKS7NW9xW
nnIv0Wd7aKLj5zgvEw1Dj34r7jR3U9yDRbIXMiAncUw7LdL8ijMtM09uRVyQSAYNGJ0SPYjOT16K
iT+nS42WRs410KCCZfZvf2kvXmQvxU5cZsyF4Du3zpemfAV4kCW0lfrnkdd+sbqYN8KUi0aLqqGC
Q6EwQLkxAIpAnFMQ/FVFuLKhMW4pO4STC/Blrh8PBTHmVk3JTZ0EeSvpJPsYcc0IbsZRanq2ga0A
KjLWi+G1Ik7GVqn4w4s1j2KJ8qwexGcaVutOGASTOX3GwZa8Z0DcJ/sn/18Pdbbs+Tj9cuoe2Jc6
PCYRflr7JfrTx5pTLWPnqXF/L9DX0MMbW7MoGYt/5z3pIxFvdUD1sUejToWoBJjJxcl9zdCBAs/i
GH0SvgURY54KENJL9EsSyj7icTwoPLHfTl/v7O4cOd5yvewZWXmB9QO33OzDOk1nbxmEgzxTkpOn
N5LQGlhhvej1Ti/WdWUtsLeSs2Urib+hW1tK2rBfGMeeN7BiFBi0fdTcz/h/6SRqNLfLlQ3tBV14
mci1EHBXGEyrFU9JjtNzZoUNSummukOIbb4h6RBrRm+T+VwbedW7+sjSYmF9Oqg9ulgnD31w3/7X
EvQlEnBBS6qNh1AO4eSf1PHlUxScVI+8RZ4S6B2/FHaXYojsZZeGL7g0Q6rW96EabSjkNzWd18j9
vPBmurB95KzwK+ZyOh2MmqYxGkonhV1rtS54J9XhRAMO8lmswRd/bLiaAvJXntSrkuVOn/15YjQP
EMA+sqvlaZGAmEOIVYJTfkxUhwGumrkPJIYUhQCABZK07vFR/3ZwVY4YCF/8/L8zfW54aQSLl3D1
ggp/uoxwt9u3ZzAQSEssmeczK+7jlCugX8St+MhxfDP9zVrKyhJmBjgDTjvbiMrCk0aciyFghRXd
ax1jlxXhYhlKsQe1duaB/49usSJ5efNoVHMK2K5tZNKlOxZzaxkNEFOUQ9MiUlw/JVacdJdvtHG3
wldriJiPZjXjKa+uXzs4jnRwnTCQDnFPmO1RkcxwT7kgnubqjJv1335MYbYFOSytFibXhLXT0WUH
YX5F5d7ST3kHBokdb6HAqx9v/TIt53hF+UvZWy2LBVBQChHEBDsE9w9u2jnhJOcAMarCHc7zbAbn
IBxK5rXACFA0/CzlLM7r7XvQ3Hn08n59MlRAzSS14v5l+9ZsH+XlSytHGvI2sT7YqMs5WvJDGKtJ
9+Pa1GoffjnQSz8kktZ+WQGh71qhzpgJn7wyye+Q1YP4QWETneJ/sjMrjFEvrexpkz1Mvgakgpxi
eFtCigrThyWDYj4gC/xNairE4nE13a26F3UjNHn+TAkxT2VybA/8SQMl/J8Vpu1mUAHRH0kFqu65
gWzs8VE8uA3D1blRl8T7jAcwcZIvkJo7C2kFW5FSoA5XPlsUaQv6Z52gmpBGUvOVPqDP9oQRgQnl
nH4n4Li4JCdudUg/l9/0Pd/MP7Y8oTMKqfqeVez2bBiCQIh2a+rZToabS9cNcp9QP4S9e3CGZ5nP
aD/T5XaOPRT4S5nrGjNWqW3D2gIk3QM+DFsfXVSZsK5hnCSNzP7CKI3eA/3ZGg4jwXvDTbyEL8SP
S9Xw2LZOv6Pb2Ydu2NKa/PShABgJ76esSsWgcPf9riiAzkxeimy03Fn2qvIhSy+w59Kp32QIcKDv
mqNb4TdanHtddLwWdb1wwPtraAYNb5yPwe0KyjfTV6AUu99yhGwxL89L3axAmitPLfX5q3YqeHf6
3GHMpHFLRSt9SC9HEMR2wDD5HyqR92Rv/xXp7H5xeR+/w1CWdnF46zuz5xQk0in9xGc/K0Qop3Oj
qTkrMztPGkKPA7blk8GRQmkrTG3FSSmEnXkKcN3Uu9+GFQQrLDxL5AJCSWPx5+yGybWGEzCX0yqU
xeijptYXmbqeths3UA8UzmF2x+BIZpwevd8BeV7N4rZ4+4+gn2U/c21+kiOK/os+ltXj3IKOwySS
s8pAFopYDcwbH8loKrvDIu2YHNK4r3MuDBwYk1bWfEzz3LmBO3Wknb5TsqXpp7eNia2wywdrstq5
KxYAf9HSwwVq69FQYY5jfTMgtEsD62kMVnxAqaDoygQhRv9Xw/VCly292hL66/Cf4rMnS+UoH3OO
bIdARB5AfIdYlAmHS05603pFQ3JXrnY9WN0SrEP+7fndKnoZFtv+a3297dKgjJDljVJzbJX0U78R
drPN86hsqaSSUHQkor/FwnHfp0ftUuPTlgBTtjmN5K/R/5mj2Es4SRCXjCFuD5/6XVcy1HryJkG7
/cs8VdPYBsoNqzWjSWSj5HGGxxYHntVHf4FQ4rETk3FGLKCwDDIe4aRpsYFsoYNwwbjYkyqtzN9p
VPuOUXRenk9kpOJyHBhsVY9WoKi6sqU7QVs6/UVYodpti2jOx+O0fMXjZXAENjgEt/ocE7pbUfg2
QfPx1Gzlyu1r1MErSVWVorvkbGGemuydt/87K8JRV3UQCyAfmUPz/dr4FS1EJC7zcHWJmIJJaezT
SqnF5LvVmmB8XBSq2g/PijTEn+IxYUkRJSUkdqnzOiJaf1WlkdPj71WLuNKQimMa59j6oJ6KwHAz
fBXN3wnuiKcO7v5ZFJ/BegM3BkVr1wqDba9i49cGeSQH6+iqyNPxMcEB1SxuJaQ9jP65EsWVDIrD
js7OQPY0FK/iK6PiZOBJr8SB+hd2PG3PHAuupNlb0U2RGGWZyiKqAvK+voQzXRsMAMIV4rvPFIIs
2lPP71whaO0dHufr4miwKvT9q+hLfbeLGSHE2/EFdDThiZfpy2Y347SseTEfKlp1ktho51WmkpYL
FLSsp16LA/8T+6ueV8g4hY8exU240/+LSl3bwhHC4wToMpjzjQShcrc5GKMtWzWn9+gM9O/6VvnX
So/7Jm9asBVufzJi6S7EYnKLgJ2skAiTLk4vC8WUFeSCyTMos7UMzKfisChMfdA2o1yoxFrJKLlz
6d34NEvqhabrKMSvJMQiIDSDoY/S7E7YECOG3yFTLhWL0rWYaYWi5CDxGZ49SXVzMlAL8R2xJeCR
XQ8qqY+EXWGqID8ip0Q5AT75XWEppuTwSNOyDQNOSW8IwMyLb/SfCXAL1HjhI88r/WRUuQujC9oV
Mie0joiMlawF0r8axIpM/oWXfAut7pB3+LKJzqaRjpdNDVyx9+ZX8mHjplf4/I94obwFgPZ9Nf4o
7qt8V9PnsQ4DaLpr5I7ahkFTJixr2kV4cSDtCWs+/c42sRumx3PBgaENtgOH94YW3Qf3u0kQaq+P
lcdWETP050sri7xsWBO8b1xlLqycqaTrsK7lR0mpcuD7d3ypVRWKQaWkwGV/yAcDtc9+XhVtBOPy
TVZFOIuBt5loLNWfHzSBMsVBJZrXYT0xzVFgY1ekeqTLm0aQa1s38Y0rTIQ/382pHNHAkI4pGyP9
ak1L5Dzbnq9k6GiI7BBpO3bLw2qKFuWKN6QVrk1eU6IxnuyemGraxiAYfwsyB8JL3w46KcEoOzRI
CBTdllt80L4gSpnuPhbdAyVOwj7hzmOdhMdvbi4EJj7Xki/ox6y0DwyKOQj6I1ihySdFtXLWnYhM
7spUz+Eir33Jtr8qAw6BfawywQxwxsk7Qgti4aW8pJOIyMcbe28dJmTSvHbZ4VrL5CXPnwZWdQsh
thE9qntQ1S7xoKMKlcYtfdT26Vf2mzggAmtFQTdR7T35+Ny0TBUgSqjaDM94oM39DNyJ72jCeuJ8
aUUq+RDyVbsrXGfV7u7G+ayhvJ3GPy+isDGGzsTvYLP4+RAXT/n3prvSvAH52non3Nuw7H/DATxn
hyVsW0ouVC/T5AOL5ce7KoyU8SpeHmc+xlGbU9Hp7MZ07GDj4Tpl5pesILPuTv5g6yRtkXU+H2oo
H+lm07PaM2SuCrPafV07Ltya12RwYWjG1yMVB/KeChbS80qkzTttqsapBD0N1jxMamEJrGdPnqsK
G8laJgdpp044mmRB6z+yU14LePlNk3Kaoe9ehXlGTc5R4phWNRGcCTgLg/5Fn5pkevPnPBTcjyfQ
sdghYonmO2w4DJneLV5qPyp0dUqvPnl+V8nYJb4qI9FqdRJ7r5oLT06GOnbtT45YBSyqFqdDKu0X
p1VwbGQpuPv1SwY+cuYA5RVq0F+QnvXJemb29rBZzV/NugpxBAJgWH44vxP2zyfyLbgf5yE2CZLc
Fd/6P0nUJGLvbbi5L5vG9Tn7wAhaPH0VO+R46ucaMPq2h54MR/hNfDEF/SjQMZXkj7lITMcqmL5B
MrcgmQKUmeTIvZph5oq7ALyX3SH7CEsB5/5fsaWnCAvpeDwVnXcSqrAL1uwjIayX7kZwzT59tGmz
1dZbTlNyGSpj5dwvotUEJdzlwQH9MduVoGAMWlT85CGpKUjuLVJqKLo5Xdsvs0hgLjmsPeiLP0jG
UIx5fOrMyD2Vn0HTUnjYb74p7eMNH7YQS7T/xaulWrjJC/knfHyNsf/UOrOw89hhXlSMVTWWO3Ro
3az8emuy7gMpHpchmtXvwT/Xf2DFKvEcqY/Exw/pn7zqVdNDaxc5aWyEnypWaHTUDLNAcIofVvC3
XgK7PRQANKXfeGxYdqI9WXb/dfN7pD1p/tGbRiwX2vrW8LP0vKfSVX/b/dV8atFmd5v/S4LN6tLu
rcupRRFLn5bTEXG8xfVVRfK3DW71pRQdLkie5k3ncDlh6eJKi+Z1OP9Otiw2d3ZV4scw841LlYdc
AufnzkPqZtXD1aBHXKLqgCqX0ndFqJq8KGNYR3uBrEF5Yvw//qlgQXevyyGDkUCP2JKQAVxd4Pd9
czuXaZ2bozikcEs7GPTtoXmu/nc+dewTbA686OvB3yo0QhlpIvs+TkpLDskldddd4EgNV1YUgolH
msUvg/RhU2JBmn4Jm5GIrVepfKfnnhXhWE3BB1v82B8nUO1sbEwV34qU2ElgZiKefBtDhSyQ+rQc
/4Kt2Vfho0woe2r+jYsKrCPvqUYmn9zT1RaUXHd/ROXQW2jUOV9LMAIuvVTcFPEGh+nIKpImsbNE
Qgq9Fvm/Kz6YhEmSVX1AnB9r/APLZM09qjtBLYOWiB/d/qc/gYuiqdFVKaHziqWyYwWnphDUpRpd
4jJgeb3F4ZaOICiGXveYtRulnxsKnwIQkBUQPJHvJmYGrCacgDEMiqN247yDQDSTCMgrfDYNvU7y
kY7ABWdNR4PUQfJS61EDQoV1f03utQbOd8Fh8y6XFMpTuffsen0ZxliD6EGXY2MdQezNKJ/z8iWH
KoTgy30XiFVaIaEvzuPzNH6JGT+OjIaAoBaU8NtAuALCOFoKUACpigJ/aEQ31Fi6kfeYr5tRrhCk
qsNISCiN0ysAP6TCmTNDKXt5GnEYUxDroFiEddfOp5Vg27w2X56KgTZsCr2gpNryL+Ra+kKNZOQp
JyiW/21KDMmyZ0+jld4cFRB1iZU9wMAQ2VekcEr6gb9BykOliB810Djzl7b4K4LZp3MgFB4B20Dg
PB2b2L3FoMVZby5VYn9LNalU/wb061q9GHBhXvDEj+veuBjet8CNR9tfR9sI5IznaGny3djTBc3C
u2ZaQUhVkUpDY8TAd+Pgv5edqrV4RD/kL8ACVPnb/dW/5SIlvXe+DVoxkdF9mArDZw3yjXeck1Io
YyuNiAnefluLSeCXT8QJk6JXSv743GASyHbAtRlFeTsdg0To9VCjCf0TM4g8ozdSEDMNFJPN1196
T3zR2plm1lCHtu3VLBZut0a/4gQmRPtUvXqhhecFbDWj9xF8AHkeW659IuotUkSiPNRDvCKCvcLU
tLz63IoRpe0GkdtG4F90uhYwVPn/z97WbuMHT+UtihCgQPozB2RJAm9y203TwR2kBDod+C2nyyoO
bs7ydbm08FTL0A83GLjO7Ph+qp+6ju5Wdk9LS7LBpjQXPjpS3Rh052u8XLyyp4mzbtczVYxQxaGK
kvOrcOcQAg8FfSAmNJwKL5LzpG0Xr413dPNHRgC2EpeVN7MsFb5y2l1e5BYxqSGeySHB1F7LMer9
EC1SS2yGiu+i0GhAobVe1Jg5duU0NyRPb0AbjiQHHNwm2HAsjXxGeqKZ1AY25wpyZ8Zl57HjCjd7
wKFc0DuknS4OZt+nz+ysdMKCTDhTlPS+nr3bYuln5Sl+vu2La74LHarCdx8jKKGvbVYGxA6jvw68
ekniyWFOFDkLeLusRYmqGAmXjHDxPDF3Ca+gE9/a5A5DlyuvAtu1YA9gLq2icq2S+Xybw29ub4X5
JtqAPmAmFfG8nuTAKb1KhoNLSNfIPFcaU0pVlMRofybvnaPzg+SHnj7CZQRRhOWJJEwyXWqN1Xm8
bTOY00PZK6j0sclCpI6M2D4idyfs7NaRpEDmBPQj3+HmgD+qu+ql+oeqcj0XZgFj+rWfnlMBHTsR
ORY7r8vsORUS1ukIHtoX4EGgjZuopWbrobCcDtw1FOzw0DYGzrlULH/71Q+weMvY0UhzEfqUsw8w
MPfb7Fnp9H8bviF9cQ/V4heD+AE7oBmeUFonF8s2hz/T5Ioj78HCNNIfHJgBxLzhYpx4uppAehct
FjyvpWzihKz4nQXY6dpu15R5HtJBDYQO26u8HU/XMK2dnBmJGCkX2k2zQ6CdSjhf6A+8oIZvO9Ih
61lV0Zct0MvVL1Frl6AfuvKRE0m7DjX5MciXzbw87lqkWHsxFP26dYodlilW/ZqL6eZlFMBOuBiu
vQEuoSPxgDxtX+8+3bXjXDHr70tgtu0x6IgflTFsEpxqgqTo6EotugaNgFpMgrPxY6VJYlgPy+X5
HUjsIZ1eQBTq6rAq+6ZGRT6DnMiCc+z/3u+7NY7d14XauvWnfzclWDTdv010+usOdq65K8VAI0YV
SEee8HGbq/Liu2mkZcOKdVit6C/bKQw9WhMH2GMkdVHKLEIvYh8NcHkrTrwJ+JLHzdwfS5mOxp3T
Ltdmv3dhu5FzjAvRLuHWJq4G8b6xyvaQYDL3H9y2YLNIULJQLlw0vtOOPq8WE7/zSfzmrSoOL25C
RgLBKkISpY7OIsCg/Ahx9L5ugYfvQnf5VSGLdYVdGpF7jZ5TRQ4tkRe9xcZftROWQ2/PhfEjhR2S
wkaf57tPNstjCLc+0oxFL/H4GTgtNp+VQ5UUkknVvx+OfsLtLgw6XQv+jOmbMxVRLMfzMFML6hZM
Q7V+cRgBwBuVj0VszVFhLiAbu/HAlY4sYXsqeyh1FNuF5K3UFbiR2CbWLhnocTjxI7IHRBgxSepo
P6beeCP+2DcVYXNwLliYCuy842HUlCQbvxFPdckoAd4rETvNQtixwrynCd/VCvsUkqdw/tnIPbl4
MoFRpUjP3+OfmuGn6c0u7lDIOKFVvB2TtiVl1vhX1MigZVSrO2Rf4PqkjD108llac8rQRRkT/Dk/
c+xNaDW/qoLaNlRsww13YHyS8yMxFF3ghEOJPatQufJckkJ3uigvPvoOJdmvRrvfSbPCuaRcPbgw
sFzx/sFMLGcOoEzCejzRk3SQkzl04JGmeq/DVHQIG1Ck/ktMCcuBwkZvrgMNuQyKVx6k0mpNix1b
C3ru6Fjgl4KERMNHNprWOLaFxXu+onnompItVtzPEKo07JDvDjZKOh2JQVCz7IpuKHFudon5E0My
Fi9LSQI47Ur+0B8/jrIpiAXnMwvrE7/R3+ifI+brWF/09GAl7ANqkRr+H7C+2kCNxNkfGF6WG3ke
RnIYuNh8bhvlyTDMlFTTOOA2N61RTTtEmb8UZ6RDjmI3/TN5jPaobB+iTAg+zCZoxY0GUKoCnAuK
lvVbSrvzz9Fgv97Gik+wz4hfWYuyrPF1aCPSPpzSkNnX4x+DFdAppu5GZRJ6PXHhMTHa67g7G8yH
rdAOBN8mNHrRnbk8/Oy0JE9IJHgM5tOz3UDIWU2/Sd5a4+wY8kcoPCn33BkN7v8XPDPRMVlws/+p
aDABco5c9w5DQ1yUeO5eIzmhN8JTv+ctB4fx1fkfjHHJkBBWjNQfrlYLSAu2yMEGWlrMQ6uWK5HE
QT1U2G6E0pTbVtF4/mA3wGuxS4X1gFJkYnz/ep0IpLus3y7Gaio8lirR7TCqqlV3Mw6ViPZUwoSU
neTxuz82O9ezRgUQQ9llLPFwQnslAHSnkPPeTczxJPFu3pliQxtji4HoH/qMHOmosrHxLqVlmDy1
MQm4gzCWds5YbPgC+kHSvEtRPyfRlX4Ncucf/tVb0+jpUGU0JEo67Yn3fSHjS2qUJSjHgrZJsWB6
Jxw3GMbeMPpAuQvoMGQbU/6tQsjeqsqdFwxd4wO3/34Lc4JN0531pH6c5F2XIwa6zFc8qMDNv9gX
ojhuVZ2XvSM03F4IFlYtbVZGplZyZd3Hts2K0KBGcgvioxMFEx5r70OxkcE7CfgpGBA7FXdZx2XS
uJzKq1pQFZ9cxkX4SiAs+H6OPVsAK3A6yby8bg+MIOmn+tBaCKdIH4Am4uEQNiXpK67Vh5hmdIlj
Dx50UI9BJMIq124qOVZsad2Bcw6eKl5wJeNzPMMTSpkkr0TdX9idAylcdnF15qpg06dsIW9Ub3PF
H3z+XYeA3td+GtGWi+4H+Adz/VhgSyfzEtrDkv96VmOrm1ymMVYeUpO+TKcB8w9j7c0lBwH9/rP0
eS1i5gFS4jtHssQATG3phsRxnXgjRKm7KSWIbyJSDExX95164NnamUl6fHkvy0+nslzo1SQNruW1
VmXVVsibnek0tQ2Gs7jDSn7Ph1eeAg/HB3hswfVoXxNsPf/cDPSXkJYIJPZHtYHZPsRuXtiIkURW
qetv0MmrQZd5wbvu+lksjvrLiFtSrNAW9BcZbhUHvy4cP01VqN9hXbncQTvJm99AeGRI05HLfzwD
Ac5SK8zMXw0/1uMS8jezbwQQeQTr6iBaA9DG4/2FOYYUo9NeVK/BNmbk4Dxpel2OTOLmxCsE9A4h
jtHvNcd6qD3bgWuAZ1fTgeoGAubhA9JNXnvkQDcLex/sQD4KhLctAzboOLLn58/kZk5T157HKUqF
OumiAWkIdN5goaBnzdtPUcQ36VbetP/3HV3A47aAllEI9WFkVFWuNk8aMbZDj6A/agqQhSXL9v36
wBgjnYwZZruqDG8RlovbJvDjWsAT2pSs84C8ky/vKfUPZLv82In7s85RyYJkhBAJUekcbqzolNRW
u+gCG0OKX90vNP99s1EWOrt8Dz5nL4//oXJJ1B2djcdYZDERXwSRoLKz0c3gfyHRC7dsy1C1/Umd
g5hMKcZsoHYf5tK4KciqlABDvUcjfaly8AEP1p6ObgYjEQLeCFU3jvXkd4f1ITwAqW84IY28Ntal
p8W1mjWgkiGs8dhtPn6XtMCfT+ljHzS1oMTq1hflkWjBs2IpuR94hVjWpx3qMmeWQMGr0L9VOKPo
OtI41dRux0c1u0EuB3dnooIknmYezkC3RiEvd4PgWFW/sIxDtwfyCsGT8FonrvmrsA7AT1SpYrod
usNFx0Et2vKQC0MD3AIKNxL/zF82EjYUCHxGOC8hM8cXrbgGLTWacbc4fa7tEkdf/jMN7DNzmwAZ
KcUHDtP7pDH+i41TbkE0duMSqEwznmwX6prXSJ6Ov+WKNi3R/v2/1ONjme+0BEEnb3PYR3/RPcEG
nvwEYdp/fi0PvUCqKPqalUVmHnI+WRuG+X42Knm+Hsga1HnHXUD5tVGFxI7aBp1Fs3oilrAy/qwO
e5gA/xoA9YHm2uec6Rw9yy6KCEx5QBxNeRTWaj4uyDDoXU6EUFrJ0w7uIZ7Vp6wTACmlL1iqgCAd
5ug/KvsTzOaVbhiY4yFNvlYZkzn0ZA3lJbQOogyKT0CqrbFyY3d++seK4i/2jX/0PIerqQ8YB2pn
G59AGGn0BN6wW56gCf6ljnSXNTlwdjb9mw4CHGwqhSdkAcI0A5o+tzfPM1nxCRtp8JLIBTmdGyVR
xvn3IAXNGToPFSgc0/Mj3JXtbkLr6LjLICQJsLFccp9HyUlRhDP7SmFHp/Z5SAEpF8jj6LNMqKR4
RRE+2caO7wH9Jw1y/4yuGQj99ZIg7AfIvyjIGwoykzTrWYjew1xFI3K2zTOlazG1WU7vjIA8C8Sd
AjpHxHsmymSFtnF8pryOP1lv0N1bS523Nlzb6FErabqCgifF97/5Q+hm2eQh9Su2+Ng3EOqzmhUa
1IxEmYkkPQC4JKRhY/zUy+2Yziqd9wL0GkuycmXzM1zZ8h16+caQyC871s4B1swj06FyUegynX+Y
qyYk6aT5Qg0NYc4CsUjIZhP8p/Ox4eThJDmCB4jvQ+3I9QwjA52BxxoAi2FfE3URVCxLrKFvQR5b
OGfg3JqppzFF2hMEfuDr9SGAJtOnyH67++W2+nDasR/gIxyEXSu0YRRXVqS3omJoj2FAiRw4VSUY
oeTR0HH5NjEK5idxhjuUcBky1yw1xFNntX7Qhk8qWCXWaumqAHZW+BLICMve2pr/ajdZ4g1pqyQl
z82lDCTBY+EtF+6wg9jbHEesx+W2pk2mVaBOal0OwceQTddOeyqvFDRLudE7mQN1DbMMeWgH0JFy
xAF4AGBRzECdOFugyMq1+6gRad4Q7l/f44TDk2xPmQMzJc/UJZbZdTsv3mAlcf3AJqKLwAMsKnk2
z0gwhdMdU2im5nDOf2HmWzNZcB2CR/A/gIGlGmq14RzJ7g4PxX7boaArcCSzo1ul49D8oxgibecl
aom/7HHVFvnyJIbUsRLVQaU1OqvSP3af/bnUFFcztnHu2YaRMcBcayF4tuFLBwsM1y8KiJsplwgo
DYG8Tz8yKNExHmj6q2iO5fZFb7jtiZIeNJytykJsZBx7Sh8fYzy6ATekKJZLvh37dIr/NdRtiyTv
RixXu/tBHZ3HySfNUe03prR7GGhPkIzXiAzC+1kyiStRvC/V++ZI7OQ5O65KeS034XL+JwbqXIsn
X5xtNX1GuYmS5muBUc+49/h/UqNwEsfaRt+K8pI9l/KX3/5REFgAJS3h+eFSZ1kSd/IQcmkvxWlD
i/iw3R+yFUjG5pL5fqCYPsroGBmsqtH54oLrrr7duZATUkxsKWKYDRopAGuEXqF3pESthhRC1rJ7
Tolc9qwu4peTyL0tACdXkEHQI6b5ZUPhjroTKoC/vkfvL+DsNPzsQd4/oQB4FieN2qFpgDChqpH3
JMraC/mmlTNEou+GucNhGMNRKpI1yxJJhw1XU0KrQzssjXNwaLKdPlkQQrHCYCgpASt6eG/UqGWU
ZmIEtxC6vlXMytLRWjcKJd1IvsMUL/byRXimK7SMF6hIQpIL7En6XE/Zb9Pxl76wfHuq8zAZIk9V
nT8XRGBuO+BB9wAtZ2ZjeVlzmESI263wXQbpy9x2oRKqfgJBF9n/y7HZwVgz/LB5m2xm7HBq0Tns
jowknge5MBy2ZKnjZxEJtUA7pxDZZ0xqrLWnLicqwK5bXua84ZAnZ4WxSbrCMOp6Ky1M911GUwZE
V8INqzgVoG2SnNYL5sEcvPyDNpuXzcytg932zeMvqefpDcOwYJRLMUVgVRht0YC18euEWLoGreM7
cyl3hxBBcOvHAbTEfY0aHpLK7N/Dyu6CYatU5Ao2pSpoyu8wD2UqUkQTS4Ck5bvWJducrx/Wc0PS
ODlv+MZDJdl8r1dGeko+U+yCrD66n3MAppMbTNLfevv1fixl/fLJth+i/BLCGNW4HeKHgPuR1IRx
JZ6TI3HRRIaysmnb2atTt+sP8f/HJXbb4nPDzxv84FTKAhpjIEg/yBGabBYqwfKvfV/uMoeVzc0P
D71XM7X1ScXRU9HWXVQTsIGQhglgWfczL/QfR/f9SDD6q/pI3bvO76RPRGELbwsuvs/UexDeDexc
k/xVeHcmzohgVPa3YHwMUL5cRvl9xKuM4JB/U8+eTlaNn1S/AzxKKTQxrfSCnuT9edfBepPLAac1
h2nUMZIUJVeemldcIkRmTBuazd6BYI1LlLCXNMABWOz87WdK0Knkpfwqe1IcMDAxPMnWoVM89s7l
yQTOnQKy+z5phF9/jAsxjh7+S3JdXmqwjAFM7WfD35CDpcE82LjbW6M1gmq5eEVe7NMSQUZ9k2fS
U5i0EPyUyc06Tx0oVrAs+DyrYC+vuOMcKiNaH/fzr9duXaD4jXAXR5pOyrPswdZAdCg0Eh6d7ezl
/6LMPuCszRWDLDu7Mtrxs89khWm2xIPIsJJEpELZRIwnzR0AD67WUDPsJtiFPTkS1LCVbD4jtsGj
V0A2jj76GPmD+IZrwVeJVC/8F5A333ec2BjH6sUb+fAqZ5Y8nPD8VpMRXGb2a/KXGzEbTp0ind7Y
uGqardHhKjrtUdPZHEMWOMYAdGiw3CskmWyl6CzIDcFD1EXCz9S6vtcfic0Kof/8r8haj5nXHnBh
a+QxFCGe8GKvgu4oENXORF3N+BYRVNcfwWjSse4njQyB5pSjhfZGL/VNuDn7U70VUMFAVx7KG99P
ux4QbaoAl3ItlMQm0hi3XW2gMlzy2cMtd1FmJqYaFKQChNDmaTuudXa56BHOw7QxnnWW+Gffrjfz
yGxnAayOEL8TkTxu3rz/6/+kcW+ozvzP3DBL6An4ubz3zkXxcf8gz7nga6n4DPHldp10Miw6FZvC
l1r8smGPQZ8cwQXPAMbT+vxh4auAdlrxnsbVNGpfPVY3BNBCWuEHAD4LvBZDweFSKOd7fs6YlNwk
AG3Z0ZQLyQ4Dq/XweypKYCZ12THGzuY23TyUlSjAjC+zmVdbB40BVqV4UcJRoMe2NmFnyl5RR898
3jNKl/8S9p9i3Op4hU58xGQLYAXxVQ4rCwkqdyqE5eNo37omMmOw2eNRUGeTdOeKVZ70WC7DSA/4
nmPlNLcaVniZ2R6FaBr8ITVS9KK01O21Dh2ceQ8heK7hnaoR/2Y56y7li7/EACgr9mTO8PU8nog4
9A5CXfp4YiyIkTTrah+DaFqxEU+nZSya1MSe9NgE/xCBRnIv+vlo+K19u/xoimak/5uKEnJYn6Q9
9+FcC8OJjHTCL39O35/WPQj8G4ybCH9CxiQGpFfrTPkJclhKPYu1TD79v82Wgjf3dLkBsBP5wODP
NomeyvLWDfB+orra68Nha3cNrf+7DdcD87BPveb+klUAOnQEWDuYVr2oLe8YnRc6WheCo6S1RzIU
4gZB3+rHPqBKmKX1zjR5zY+knFfpg86uV2rgfQErfZ0F0zFJP1gPjsgjtGs8qZ5GJxrc/kdm8m7c
E8PVwI2Zs12/TM+NhjHnNYUvDbOr4JWkLmNJnYybORhZcK+hfuxYo7p688SYvC+WcAcylQyFlFA0
iVZER3MOGuLZlvG4gjH/c5yfn/DUtuI8WIOCLBU0ewqj8vK9o8RkQMfMuUUg/sW+FAKBSaSWlHw3
X13/CjhNJHcKwT/d5GQkFFRs7ajYqAmHLyhAg14Ry8UoUZmHizWKTQ+BEFjOFzjR+yQo3E7QGGkN
HJWbSMkzvrgiPeUsF8/rOW2U9FI/oDZOIFoAOlu+TmTti+2+Hm4CqClLuTM9RMMLuetaX2IX02tm
A46gsy/Depn6A3MdVfFpXIRQcBf0btijGWamSdvm3oxyyOPuceBs/gQ+BKqNgp+CI44jE7LqNOIH
p7R06kMeCIFuLaKds0qdj8t7HyiGjTX051iAZj9GSi/1SP4WXJx9Upb9KHpIoxMODc5B/1e46sF/
HUaDKVRsGArtlTIjIHisbmfMsduqa/EseWpLCfosyFY2MooHJKaNg/ZAw9itG8uW3D8oSmGvjErE
JKxKEV5n3AfTJuHyEDV0l+WGdsN/1wmBpxCjkcowgsm2WbeFp9P92wAitn7bHT5kPZVtQH/6fE39
oExAi4EfqUmjFAeB4We6mdqaMPMK2LhNrTK9u+1X41uywOZG0qmWQMwU/ZyQi/UBJc+DCHN2gQ9T
YNNWLD+8mqi0R+jRXNi8lq4GdLeX+hg/l/o0bBC7I4jr4uTnSkVvdHnT/yvvP4BOju8+eqy0mD+g
iy+/p+HgSPk73f5t8M3634s7eDMg8zJ4gj3Kzu9z0JnnpE3J3OX5nq3LwMPTqBrhQ7U2G4cm5jdM
xLVntOfgJ0L48bUI5bC4Y9pIy4J18VjQWaCeSqGo3zoZh6OXqLqTCQSyjZwsSTWM8KvoUkVXfTvv
Bu5BE6G69/53aOA6rkxU1DBIyMY5iCG2qo6QJQsIXz3Hgf6OB8mLEJGZLqPUg6f9PAQa0LnYvmad
IcHMM8tAruLqCC5KzCIIr+hMUWoWoAnxDmYtVICZx1rTHLymohI7ku6ANb8XC2ma7KHVEvtVm19m
lN2vpGsuQMmiAQM2WswNwC4IEeqf9TBrqWKW8FoayrEYmbBvxtq27LnjXFC8vN6jVymFVO9YMhGY
jpOLDQxgMaZiDDqBqBGdIAhPvdDuo8k5oqsCTDH8OkTsEkJbWvYmfD69u5/HATh6Ahg2JLPq/2LO
po+6tC81eteiJQVH+/0yubzO2Mj7m70Wm1nQ2fKcgOgFoDVL31VF0IGgK6DVt5xF0rZQxugEF9oS
wx8DhAMMF/p9wBZ1OhfHF3MSmWf8ssUTOR7pq9UgFSBewFmNGWyWQ91s8IhtuazV8B4hu71TAve9
oEVBpfx6fPbJ+4amvYdVxev74IOp42vP5RO3nWuc1gstqSevpp6R9ZFbFKaSFx0nW7ppZDJqcOmw
KW0Lp9o+fzsZpHwM0dX/0tuT32q4T7iuPM6Ubs0TOPVFZW5XNsKC7Z5ocGB3OT7WirSwN3UhEsJA
FljniF/L3FC4LxhuO4i0noZnKMO41xrlXwjtz3T0ZD4CVl75QMxLbTIz9NWjbvk0zUsWfmqQfP8x
RdRctkhs/8yuWeAOBv8dL9vJQFvrmSTunsYEhq9EQAVBKmDdroaDknRpmJKYVnvjySanqVAD/Ojd
G4xfBNhWiq2Ah+EeVVMn7W7lcQ9ZZgP78H5T751rbItUObsJT0wklRnhYKYyyB+N5VH9i9vu/LZE
TjVZxKLFmdTsp/6WX3CVrP3TV2gGCNXd3v4RIE3H5Z11AwTV370ffDjjz56OPCb19iiqkAG7Ytqn
39VyC7G/CbZYEkmAZhoD0CXTQq3y9l9non6lMDq9uGlKIInCtgWu+7+lNzw3piUrof683tNgW6os
KXAoctUtrPPHvMmzXdSwWooOf/gokfYXLbUqSf8oad0PVFPdPntp4TC51sQ8eDRIumAIPn510qyb
r8cdxfL9mqsJdGUdin6Q9Np+d6eaiTMixjoj3+YRrsBI+VZAJM8LVDdU6CCU670IwngAUybt+Iuo
LjOPchopKyq4J0GQCASjRXsLeIJ+Ajic3K7RPxuC0YIzaQnrtBHza91vKT5uUBPbe9YyshpZqHQa
oxkP+2IswUfR0tWMjpftimmAhYaYaFPPqEp+Mg080FWGkHA5PCDsK1ZbUbg1NSaoSbdcXAikJc5I
H+2ETfIB+Fkm02ZSCXlE500aADcLOS51bM56XbIIpo92ji9Df4KbiyCpRFIvzQaSy/LUHUwfWhHA
lHtgZEuLhBQ6gFW89K6JttwdOG3Nr/p2z8oMy7/Gal/5q85zdNmySH62aYiY/vjUNl5Q8gDbIgSV
2NLgQD8mqxjn/LZtabpodX5y6SO7BpX/Pf2qq4GozW+RSClSPBrUiHfW4ZdOmTMsQ7OdfK1a7iAP
x5FmbpRKnOWG5GwWz3NrHwxRGEcgmOb9og25EF/WMMZFGgdIzCPft/CbJTh85A08pMI5+lGlDcPP
fBF8cGQ5D7US9SXzuBNn2xYDkktHT8VYi879VR7WWaVzM8D9r69Ri//o40LMWfkiW+5fZ+pBibKb
o3bPNet8m44fKSIgtBVhvP09iiMybxRmqjTXHt1JOpQZCJON8+xMMpGDKdF0/9wk0JJImH/R4GGn
McdkFoK7ym2EvTJUqquJBIdsRcUE2zch0SQNcEocWIBjoVmQU94sXlyWATdc+WdswKGtGvKIm3+A
wcK50vMgJXa3juC6820U4+fZdwN/jYlYTrbl6Nj+/pffzcnFu4cD15TQrCrhjrBcPGucSWRZ0CpQ
t5wl7btbnj3x/fcKGRG0maIgtFNDeYzz2sm/TrTbAoMCjTMGUywZ8t8tO1qpY3lTSRYYuhVa1yJy
khPwakjHuEbezTDVpA2FiMEZpdw+dJlLEnI7owzbQMGDgKAWRLd7Q6Yt7i9dNaWfR4OJ3C6f+5tq
b8KjJoOFKApJd9CY76XIbq+LdbFuwLenMWnK8wjcqYDGHHZXDWt58MSCgM1lRU+gfvfV4WiV7zJZ
+umj5hqp5XTKM5eP2IAlVg4sKnfB9PYDj1wEW9Rj+G0bRO0J3ZSYxtY3u+gNU1ajeF8lNBTD6Uio
vlkPHONUdRZzCeA1Lpc8UwxDuX3XdezZLgqL/55RkG5cEIr9krLHNvnuKNZ5bCnxIR5GH6ukM/Bc
jh88NZCjsNR+weLfp8QentuSafdZeZ+WK8S9afr+sRxT04fvOrFy5XeH+EiPww2h+idcWNrz1+BC
EIu+OLc9JTgADzONaiM45GK1QVQvMoIOVqy4gkzIIEmVOMwEWHwMk8PMkNv5NVMbQlPeQX+1Jt32
UWE29q64K5KqyarxL9nAtcNSsOzRK1F+IZetyHEWF6NzCAWxaHEwOrIxtgpNhACZUL3ZbdA90Z40
AtmHAA3hsmQUAyRashOnMGeX6cIYK09QYIo1s9cVYDWAd9/trljBgDX0XjEnWDnVjP636D2nakTS
owho2kpUzV/bc1WeldYgSX6xunb3YXNy/mbd9zLNHvaCW9uWWiv9R5W/pCkyYN5apPAjAf1hD1AH
5kn5OcD6D5DYRfLPKnxIf6S+CFzW2A9BBgVAG+6mEeD4wUlq2QshlZ0qJvdQsKX2gTXPpcF5JDar
ty2Gp/qfwoUywBbsJj92sAGhhE7I3oqSEa5hUxLX32fgUDfRGy3rLOt5fv7Dhyz7NmMNc4kOObwE
39qN38PpD7L7KmjBhKHPxPsbUuJOqn+R5dlBN/Cfv/mZPK32HcEd5ce/zdWcp7nnR+4buMvVG0a5
iJiv8jyyG2JpE06+hfWKkR9taC+JMN9nHe/CiMJ26n2DcTKGB0sQJW5PCTswQDI9a33kJpFUNBOG
nlEM2RfChoZXa4pWND6dwdmq+ZNbWezB56I9PvuzSW2vcuG3BjyQpY3dbE3kHJevyrN0Ittaclfw
xpsQS1lyYepW0K4JxVcgawgQ9qHEbzlGzlNpFd/ICigIk9jdMih32bCiMNUnT3SDZD5wYx2+OU7u
NCSfkEnpmW2PElY/C9l2qRVkOwu8c9OBRfSdzDCgVAnzsXFxQvUGkGh1byqvE+r3IsScIArhpV0k
hlzA5slQQ2bRRLG6OYTFSRDdio4iRlJS7vRY5G0BbgKZiRIMM5DmoMs0Uwvp6p/2xl2dLcOISRrR
JOMwDCoohoiNmGbhQYFoKTXTzIdmcv3p6FUlwmJMsPFKJC5QddwIy0PX/rBzVkvTW7VlogGwGm0J
0WrjRwLyI1O9foRSFscRrJkW06Nqtz4nvpZDXb4Dnd2nV66q9hZ8+U2wz/qHmo8MIEMVRUWIlkZP
rTcpi5dxw1o5JF1pG2cP0sITOjarltLcyu5A4EFgTcUolWlWf6RRxb+bBvg6j8jKRmxwSYre0Ctp
4W9mxZElvPjQF6r9R3wjTmHf+82Tb8AKSehUyHJWfvu7SAYzX3b2gteIj4CVNvAGVx2EM97N9P9T
bB9pALiCO8s4SR41XOBU0ndyYcoVLafTfOgx/7CrN24Z1p5yCZCTwg6f4v3yZggy7c5Rm5dZ3YFG
41G9A9tyxuhjI5p0LxeqnKB0V0N7aVKmcB9t9xduFWJrPzpOTc3nWPufHUUoExkQZAR06++ymvZS
4Qr5vxyhtcipBvtd40lMfN2R3nts9f5ZjM8ROxRBvBbOBYeguJOAwjgB8tccIiUxiSr2CVvvACei
5hqRU8d+dqBudycHwE96Ix+xKxt7deRmaJ98/UKlT9sGnCKmF77BWZGwzdwtG0m37iavJMS+baxx
Wt2c/36J38Cna8X8zQCpch/xoPi44wl3HT1ql2muR5e0Az4U9MWPoa7XkbrrZZGlY32spxuHcGeC
35hR2PrYTkvaoFVdty8AYNapvrHM6RRh3oC4b3U3K6qy931+WowIUSquSQOKzC8ps4uq8IEKgrlz
y7h+rI+mEjQysYFR6S8dh/hcKhtFKu4heq9edKYj879/fPfIXV7dRk2oEAW4kHu1ocx2xPTAUkrl
J7XhXoohXv094k91IgBa79fYoKZwYX9GNC7r3wBT1xpXR8BuauuoYUO3qerQcB+7K/NC3aPxvQJ8
vVb2HDsjjJTCY7sEsvi4M6zUxvRZhj8W7YeEuhPkkwOMbZTbXpgNHyvasbX1WxEqxAI08sJNpqjH
1tn1FS68391IhfSAy+hrm0tp7egGwCmZVHbcYGL4n2YQhXe9Jjoq+7Uand9bTdnJ0JNI5lb05Txq
4wDS877PwkK77d+1hsy0zxGDQpgGF3lXvodfFtm/9gXCwBEyD8b4Pu6DA/VO54p0wcDERYBjGW0W
IppZ/P8woStg28a9PqsucQQxjaoDn+PrhIY/L9clcRgc72DmW4iIHe5YJfJUtEhMxjnCRCuEZEar
pvzw/RZ6ARKqvVSJzSu30xsGU8zgFgmfOYQjayqlZprrMVNY0moq+bB/Ng4plKAUvQKDfQx3KBMM
aTlVsckesQgDtBMCIIevQvaroaHePR2vzAG4oDTFMr4SIIiE9T7fpE1bKbXb+YRdelxNinTsAAej
HpZNWY/t+FB+Tm2gl964ntfsMIsSwNM39SjlGnDEH2KlkO0/zBYVR0lV+YChGh7/4bCjRCAlqdSB
wg1X+J+ztvnUwYnV1xEx/yq8ESJ8WuB/Oj11tkUeoba4ZSdwxe+IVHqEKaevDX3werMXiGLBYRaL
5kflmaoTE9PgoCSI/Kj7GVkFbbHkZUyS/W53Xf4ZSyeW9sBJLjwJsNsXyustKd/g2SEJNmW2ayvh
IgyImnoGx+lkHI6lNfDFA1VG1QIP2qenysJ6k60Jo/8SwDoLOoJvACs+WwHBwp/NpSEy2UnSX29N
cpTFcHP+/osgeW0C9fQysMGMFTeo+ZI2UzcAmhx07KVa8StS7vl6vdeUwwjVIAkccjGmsb5I1yyt
W467YykmCFHM/mB/zygbmI0SWCFhI5DPrCHR38nZkLl1wagIQvBOqs8f5uJG9cUviTv7eWqioWdc
nVWuwhhLQTOYFoEtMTbuc52kCMLlfngUutqwZ3+mxcdG5DvLumE6o/vrGk3S7+DGvk5JgRi/jxBe
OZUuk/ejVUhK4NTaP3ExYezcyN2j02GJarRTXLIjRG6X3CaE97ug5VOA04V8M4L7fNfalh4IoL0v
OK6v4ctCDNQcPfTxMEOS3tMzqKm5X2UJTCgfYssVV1bEApe3QAZR4tAPaUO1Qpo4vi3J7Le70YKS
G0N7ydma5gFCh4dQA0xKB6Po8F5IwUsGeLYCzG6/mrSTSOE6OjwujW473FoNnBE9okGLrltn+6H5
VuthqrcDmW+A/CCwRYloZuromVTlIiHHQQQodvE7KdGSw7atyvAjPmpOvOtInwnoKUAe9Kk75PwF
OWjCi/bdA/EZ+OzW1Zcy2qpTqTLfsnkGLxtJYTAMpH1v0j+uDm3dcdTalQY7WVQ+dVJu2jafSNrR
kThzndXYckAFwGITqbToI6ktAtHid1C3RrypE1nZLS10ZImeGO/1F5mF6f87UDffGPPvNPEFg2ZK
FESEIbbwgvkJ4/KNdzcRGeEtzcbO62pGm1PhdvCOW4qhd5Wuu6xpm3eBaRFZRvvi9bEgYzZWugq5
QEypbG0a7Mcb1Px10oY2roWOIM+dl3tNsEGv7pfJwAUxGaReDfeovr9D4hfSJlBXho1bBzNF+7VD
TWGatrYcw7MW0K7EA40v5aqgWS443jOL/OsMVI/JSzh2wcUvspPIBh1Axu6uQQRE1GynP0unYeOQ
C02Xjw8NSPQdHaqOKosjztY9jhfSHvxBBM3OOUOVFK6ej5XYJokeysdD2AIVxbMb8ol0h0lDmohX
Vz0U4+Hlo6yI+4wxsmH/5Nu5G/tMBYhyZTWjzthNFMqPuuUNyKUeBGzpgPhXTD//iS2q6+VCK2ac
5qx/Iv4wgQMTIDT0l0lW4Uzr1WnS1sni3hWmfMm0Wx5pFDel93le4QHkTwUgxpxA1zoa3MR4Vy7H
c+iNMsl71YrMrPhVxEiVT34w7diF/p4demRIaIBZSYD2M7VobV85PrDwTRPpYRlrWEO2SWvyAXWB
okLhExm+t47t8JdnCBkQ64ZfgsxZ6mQIxCW+3YZdsCyokyvZegOgXwpeCLdcgGdUCvvZqJvkEzVn
BQ3euPKwKJMTPZTVKtQlVUnPe6xnI2iCG4insZCZgGS2iLKw+05bR/6NTnPCUldHyrB95MevmZo8
sqMzexwZFQeauZFMgSiyOsrwBujRfQcI1RyHuMXuif1jtcRiC40bXh0DiRdlHxMP2bX0Z1lC72Zz
eSd1QyNr91WakP02OUJLcWT06JbgrNaarrFWq0sTc8sA/oTeO9KxAamPB7I+NdOLm2g6k0xDy7Cw
hd8h2GeIuw9yfoSyRIP/2jhXpCJdmvmZi1Cw9oAa8OYLvAKgV/w4q+lRo6MTfX0e0UwrIpH8J/gL
+FajvZCv694ANj4chh+2MdAdbFhGPxWRlWNFsacOck6vS9/RqRWFv7/DB3KkQ5fZyPokDCIU8Kfm
FObRavVdgq205ice1HfNXbh4FcbEdLF6um443Sv0sYglssujE/aQ3NFQtyEvvvvDoukKKPRZnDl/
SdpDflyrbFR2WM88PbcPQoLjI/3pzR8kOuU7wEM6VwjeYvgk7MaSYlq9bKWpIGzI3l7bydPpUaT3
y+gFcMZSLOGfZUOgFJO0PFGwL0LVw8AnDTYdPyqrqiPhvJvfCyZ2+tbn3Vgu0dlLETSCe3UkJxST
gixctNEtjwM/Glop8zmev/YhRcbUD/BvZSAW3AuaJz6lOv/o0RsjVQUHFvlHLhFgMMzKMr6q4H+h
cofrLTdEkcavotK7oo9ZgH862WZ3jy6MtMcj/23LkYAzj7d3hFB/IyWzCEYgZG+LX1YMNZduNh1a
8vREqP3vktfCcu9O41o4GgAVpZZOJ86QiZl/lwOMxX7JUlG+QWjcDMsIf+HwK1YeqSqKO9yIgEFM
Yqi5FhH2MusWKrupOZ7jikYmmhMI0A4+Ue5vbbw6jlaOUOxxRbt4Ck3I5wgFDm4LdgtY4tFMFEQk
UbIs8FHo2NQz9+7/xGfqjhtvSQu0ifkRYkdk0AAdE0tumkNMcUqre/mKU8aFHNViTA6Qp2KgiPxk
6pMWph+B8iq7Rj6+FAr8XO4lgmhvp6LVQfN7eYmEEaBNbBp7l/1Jkv1t/m0B22HSqKKtnnAqeaaT
IXZ+7vfhPWUacqol/c4NMwGYmkgsWlvuJNoHLAsiMZranbP9Ly9wLq/GCWsi5HREreWSiQ69F9Gk
1JE0dcGegtMQ2w+cj+A0YfVyctj27vghyb80fOHK2MVgO7u14a4kF7f3FH8R2+a1Zb436RVJWYyj
1lwJHQjsShR7tJYvMuxV/rxUsZljCPHEsF5nWC5ysOw/yLIDT6D0zROJkvVn9Ez5huNf5CLjwN02
YW53b403AJ/buSRvGFNgVIlcr3OG0NYyYrNn1gTfyk0q5Tl5UONtYw0z7n1Qh2vmwgm9mwT/xDQt
lm9uNfu7o7+yzFcYKVEWeK1BhHcuJEngFOWBt95bFNRT1n+F91DULqt25c6HOKoFaYPa63yTV+jW
clLVgRMT/8b5G1GJi2k+e745kUk6Bo15uWBFdFz9AgE2BwVtHTBNJ2IQ74DxJM1+xk4JXJu0LkGH
kHGRoHcC63sdBxj67fEYLAlI+uYGaGFZwuLrqWm1hI+il6J6K06YSWOC62S5brlDHhl2wEHcP8SW
fZqYSbJJLClGFX+3KK9hicTMy0snh9DiLfyLNh2h9ZAjIZdlHvkiMtjUNHsTsm0pHZcxz5ALT7U0
pjXdQfacOW1vFxbhMvv6NP/uR24mCinjZK2NmwiHyOVzl6gkSYmRVIJDhSmtaCP6iE/D3SPofINt
SvJ603lGm884cDJzVYLxihfFg0tQLTb6D3qPzak1GxgCeITu+lhU0nKQXip0ijdsTbEK9Hq67p2E
MJ1qDjy9JN2uzIoOoBRleECXO7idPVWS9VkZnmNjlyVoAEVY0UX+rFnAwul3OAnaoj16C4Wm9AcG
G+NVnnhlCtF70FxMB5piqpI/vHb4TSQ0uWVTZIQ5158L6gDQQQeFZNcv2nJ3vAUiKLrIKSPC2Uwh
XI2+RFeJAa5gCH3mXRnpRl/9ikfaPutlKj6p3lV5TBAYR2YMPyv6CpJ2FggVaj0pd8VqMfGs/Ws9
ipx2BUSQu30RQ7VuHEI8dv6Qx9aIMH2zbJ4uFVR+ftM86DE1FVEAnvNmPx615wsV8OstspByl0Fg
/RVGUnrVfInCJw5kbRTB0AA5nPxot8AZ6uuKnT2cF88AA2NgH5R2eoRWhr2w1TP/+k+nECz2Y6E4
fSAMRUt9M0huEPYgRTSTNvpzd4P146pfGG3uo7kHks68Hfiz+AIWrUzCGoKV2f0+p1DRGQq8I36m
MEcMQB2KAHpRowIhOMPLbBLxOftTUMLJGdDxzAeZTSriT1YjcYvqJrqHGKLmvxtKMC852d5nhxMg
V5r4PMfVTR9neGh/ymnhvQuRNIld6Mj1tDAl1i43ho9IFP4iZbtqb3R6peCTvMuBnt6f9n36wyXl
Q3hUuTI12hfbWM5A84t9JDv8+aIPJvi9+L6slOQ/lSHnxls+Qd3lQw5C544/SsKxaGFRDxDse5Tv
2mztId3GHTri2cR67QkdSJxn+eNR5JYUTBIsFYybF5zhOu/tnH1cjdJUiBAR+A/1U6JTrpP/Oyso
t8netarsUp9as2DZaMjUn9ajXeK5seq/71kfQkuDpbqnHdTCaHHSDe+JKnVmMLc6vxWXhQg88Mal
cUJ1zzusaWEwfeBe7JO4x4rOw1j61iScBsyQ3dN6epDMco/VTl9V1OpSeNzwNbdWlFjtIJqfuJHc
5mETfOyGlgar1XSXUi/ocT7O9+ZAjTZQdfqG/TgdVT5ExHH/hBQQHJ4o07avNTBExD4sTTZX/OmB
9Xx4FB/EbPSmJ2zl3O7oBeknPpdHELmuvg3BZ3cliux3NObjjrKhEginUKrmInGUXFPR+sIXcANu
iUbkNfER/PfGtKOg94Q5hlPSN9zrVgiv1ZmgEkGlRCnwJZqBMsyoBFbr2BOD90Du8MkuSnJ1xoFb
h9oOk2GGg5ZYiCOucmRTmT+OB64nuwZVUta/MH14iRW128PJqLxN1FWJSTaV3MkFLUF3A6q8J3ka
KFqXVlpcR+7kj4a+LfaB92dD2zKBKBeQP9vzHByQFzpXM5fUOf9DYh5BCaOMvl4bAtb9on7FW+TK
V9X00BJBJujnIfQdxCgUzdR99CtjJO/eZd94n6jiSejvfE/zaNvBDgQiWQtL/pgvjwJ8VlT75/e6
DXQfX7CFboPIs6U0sdn04PrlJpsTqNw1wqpWdoYmD5uEmtFNfYgRKAuC3k3+ZLE2AqoyGwF61kfx
q2keBfPHMk0ETrji92ft+Y2Y781NyYET85o3UGK7MhyfCWDhDCDtuNMSp6QPXg2UMFSKMcvh9L4s
tjo6mhLCxTaj7WObTFzVsTy+99GuibzZzjmf3cJ/Ij3KkQ23u9clm8w/PPHEUry325UWD+qOtvDb
eGERWj4eUiPa70qNL0fzv5V+Wd8t222ANPb8+wCjMaItYEcHympDs1LDXFVRIVYNltKgOlrpOP3U
Op87XIettys/dcsx8ecvr2kK3aruHC9uuohc2zCOYlkV+tzffx8XP3mN2XTPD0nSKdm6SriZlLGv
S2FEobje7UDIV7ol9PvMAE5YyCXMeV14MFQ5yTDje87AQBnJvgia9mU64R0Ds6FauPgfHzN4rVT3
9cLhcEDTdR0F4DU6ZEnLmtDTxTUbAWhbeDLWqq1/TwcArS+81c8NCjCA/fC3k1mwCm9Yt6E16wdG
HM3ZUQf+CT6C/YkCYZCyzHFdT7atDFLwE+wMgyllGMiSlRQ2sW+MusoE8i+2Oax9YAUZucBJj1y9
NnwktIFk5zv8h389T9y17iaeeHpGFWky87rBsJDibwtBV3do1BYu3vb+KSqXf+9mxf3lirdM6ofJ
mWjer0pDX6uIFNVQog2Zq5FbxOQEdwtvvcpngBeVZRbV59WGMZknW+1NGQEajISUEQ6Hp1JOYKL0
xiHvidFchjmLm+R7ylKX81b1cfCniuuu3eoMBi71nwt79xWjESFOTvkllcj9kCjzOcBzpQpmHMvy
YheRzpmGnGMWomFNnMcPmLd8pI5+lGaUMKqLvtdeOld6ee2wfJEx8fPRwCuHKULcGFylZZN6k1U2
XFClpcnqD1lBOw25/iF21j1Zpr4LDc/uFr6fASm98xWIga09u9mrGnuKiTlLictuog89zY+hXSWt
PEj+7JP5s9DwH/tNSRBlDcP+1BqxpeT0B2wTbc6eSCW3uM+5WEDc/j6c9sgayKo2AFbFt3uz+KLy
+dLnMjGxkp2mDMIkOSGG/EM7cB58ov0fcfFoD4wp0MD4TmDFQ2M+4kQZyrsaoNC3dJYgAmLZ+XBA
a7IygaDeIkTGHzGgjL++dyu3lYswmQAY365XfuwuJxuemPFAoQT+gFLflCI83aW1PGC1VE9UsDQv
RHZPo7Q7IQAcvbWM9ONL32Kq96s9h76P9DsEJqjgzA/lz5jjFPNSyC3a04JrfSGkhinJr/GVsuB4
/uNyoXZ5aTo1yYyd4bmCg5615KBzc5p95ybiZYIXZNqP0CZd2brbQUkpYb6insDr/g31b6Tir2kX
qEn4JsQchTMATklozU15yD+4CIwQzqoluWExxNC5FQYuL0+b8si/jMblz6ZNg6ZOCijNqHk9dtHH
xBcB5F7jbRqK4PUENtw0op8J/QINWoztyZHs9gWzZMKEfL+2CRpy1Mc9ZbJ8zmJmlOKme46upynR
R61GFH8v7rX3l4Bv0Xz2dQYeMBmFBC1vSaqihOpRdTAuy4DBi9ao+ahYdQbyieJGNRdDhHis6Xt4
d1uc508QW76lL1BvsCJP2FSzmJBC9rBz5aVbhgxJ/xEbCHRhAPF440wxu3HurqdJkhZIAs5Gkx6H
MfQfzP9uI1sY+phiJkMvq0W7I6NxDjQwA8ITpK2r75ytjhxusD3iphUQJr+ffYtTyrohRmTJjDSm
7PXuWiDBGK99koSjZVz9nRzXMM5TO4h8C1rPpoDgxWESw3qWN1Ilnq6OilBdaevF094VdRzC8wdQ
+qwKkxGkKQkldzEnV/isUX6aKsNU0oma5n3ERvT7onYq9j4kwh6t59wF8Yzl3IvrLnw0vRucq9ev
bKmH1i4+rIvQ0n/CkuzkIYMeM3w8ppXazrW+r2Y8s04TnK/WZl1XkQ3if/NeZgUP178qFk0y4FWc
CKJ3sQsholfmsMif2Ota2rFSsww9CfAMpvUxlelMDIvGPPwq4FxpAyPoCMeXpIqAMon83Jolh4Gx
0jM1mqcHwPJd7ZQ+v9D+FqPI1aE4EM94SQS47QNT3wms2kWWuEaWF6Ks8/kcjU9BWsg7T8MXzsYB
erHJHMxQ1h2ZA6DoKGDK7OhCnbS1CbES/cPAOYWPp1Ljd7cRFeVbPAOiIAI8jh5UYSWD/IP+xsYV
z3uQTUHNH+Pj9t2joTXeAChqBWe+g4bU5Pd8ZaDpROrXV4yh4n+nzmfz501YOMjAZc20ebCAYEya
Y8eKzP9DZCvmgGjGNc/nCBvMNwW4Y8d6drPzwu7soDRkqS4WAKUk+RgBAmksC/reF5zpCx72K79u
LMJNdwkWnj1hqBSy4YntW8yBvGd89dYbKBake0hRGOCdIsQ4l7IP4LKyBM2axS953Ikl17pG3CRo
tvsvet7TqPePkvbQ/kgRzD2IQYwr80p4f0Rfcl/jSZiRqs3JWFFbNhqdsBsDYymQZtQOAd4069LT
8wQSzFibfHz59cUkOjRym+T5crL09t+RZTNG0iQ6bGEsftUxZVpyT4ccsIS8ncr3tDGtR2b6bE5b
CyYwkkCJLMumks8OxuN3WNnP1M3EcwSwW0LapLFctiI9t98rHMXIk1/WSDWFErxLi3EK/bcqO4IB
0htrUyyNu3Bii06WSOQwo2l8A31hL3nej7VHwTmLiuUCL6UkfQyBoWzksp3DLWSwzfgRpEJd+fd2
i2SA1V9eSoDjL56ZAQ0H6ZhRN7VUBVHzrWAQhBMusgIF+98tzieyvfXCfxblKfc4r6pwhc1MYTO7
zocf8MAz+iuhLv0cD/w34DSr2YGt1aSDZzMuwEkQlZQHnk5gRdVxEt8GEj+6APqZ+K6daBZoanmm
N3l880ro96r34SC5NFst/xs2jBGnm8Gj664NGTebJnFj+Lk9Iwk5SNHTFwVUzkFu2sVYs93MkF9S
4x1lF6DM67kY9vEBp9Y6E/7SUmGWt4LQn+NbbKOynUuaEUqHUVehHVQw42n818hVvWtC4MDAPELL
H1XI49l3Ap7hecDgNwAj2JWPhTD/zLh+fJ45JgrTYr6qfhqOOyN+AgMCsW8zp/heAWZqeZQMj7Fe
kCExvpzB5wy3SrQao9c6170uM+0pHEMbJ4gAROxafyzQp0UXhfRm24Lz1DdfPw8gsKCrpvpY6VpG
24TKL81388qtzg8ZFH29XpMe/6eHpXwMTksTu1cfv75SpsOkPiXFl7OBHM7uROruxuqn+0QAOf9Z
jztYtHkYUjEhxDO7vWFl5Yswbp3KT/LWAw3kCqAf5RomD11h/AQh+Jwa15t5E182yx1b+SDTU6RP
ddxwWD75N3IQGdheEXKiqT85hE52aVjfwfdMvLAxeqAwdhPk7zZTRGy9s0CFWNy9CZAFr1Uz83Hz
nSl/Ly2KN3ec8f6kUclcLOMIswVG7lWpSpMthlxiqu2SIhQYOAs4SWUR0M4NbYtiHg2V/DUt1p8O
aK2lDeH0uhgr/erLRhnDxs72XySEPxnGIy6nwiWD8HMX5/RpeR4Q3IwfKKaRq23ed3CcpFCNHW17
GWNyy+BHP42CLT/X32w3aJNPWBUL2fT9axYIixSyfQdCwbDVaz2YbnNJ9rQ1wZyhE+YGpkINGwuz
WZOL4KuxKDn+VWqLAkQuC8hIG/T3QwuX5iIfmRFUtmXctJ3a0/H8gIP4bh0Y/Z8bMk6Tt94JmPq6
3QWMuOv4UXZf/b4i+z7/QpuXlA3TcPJpWs80FdkDgA6G9ZcEjQheXGZBbw+S2ciefOnm/4XdCNge
BOCh+JP7bWK3vO86X3oUivS6GFbWUpSEHZeXVyNU8GkwvA8oMPyPeI3als9XRDlpjIxJA3UOKPz/
5aKXIflU1rWtDv3NTm7A0bBuBtEmrZceHpx6/Xk6kZh/IkDpil9sa9dhR/NoM8taPcbLW5y4yhvE
NqAMeramSiG28bSpFO1V3uFFGyd+d0C50ojbxvRuMdHVwRSQ0cJxq43h7kG0uCOkp8KC7WaIhtfj
YlCSWVWR+PiW15chQ/dTBjHIX4XrQt+u5MnwxTY3qUnSfokocxZ8LGENf4n+b4QrELpWY7GBj36E
TlSiJsAhXrDFMt161BknBRo+PjN+v3p5DcG6n9D2FtfBO+UeraDimFqZcNnAJuD+SC4RwdsgUrR0
Ek1c3VUj1MZUwZvGwI6A2GsmFxZNtgO4kiynK9fYCNYgAJwML1gaiJAj2ncEmmhr01q/dLvSEOCo
wWwwaZEEnXmMU0BvOzO4bRWCbWF7CjzxmsjzfDntkEZH7aXJrHCDpRbgfgforuc5piiORtr/tXHy
hmUhCoASPseuYzK2XU2AWWZxX2iWxpD0MWCnMnsJzRAv69SvH8KA+LxJN2xy2aco45PeaRDCdVnz
w/xaGqA25CwLc9kmcVY7VHOGRVPqFlYpJQl6lEdiiGNPR2fpIRZeXqWaY4RoVrgvZFEAZ/mA1m1d
Hh9MA6Gl51y49AjUYDK5LSAOy6behV0OhkixMXonXC6vPqaNa891fdfcUh3Oe1scN2UrctFVB2jj
t+uWi1G7DWCFnr3icCJrdKia1Aiv4m1SIKOySGGINZzjkz3DS2Fngj7wUO+/mG8QnPlkUJS58Gl0
a6wJCDs0iQeTsDWv64PPzhz8H07F5HxZcVp7gT/Z8S+CDfN7irgCQ5rIH4DL2/L+aR1MeXYf8HX4
FsNrWbFgQCn51akknfribaaP0I7RzdlFJEW8loYFy21O9NT5dSSh5/fEhARFh4JYJZb0v3Cfkjpm
EnKnL2kuH7kBC4rxHQO8mGRaXYGsBimV6iEkpkjmXkiUqLjkn8UdEtZ6c/4Z0Ie4UqaR4BMqdfDW
KXe2pMQa5kATN5qME/FPRwkDy3luHXtZvcG3sasV/iWlsv/Dz7KFMJCbAzMz13hEpxouu9DTk8BN
lucDmRVDnJHEj8EzwMJri7Cpur7MATVHL/PzmGFi8NedP6oRmgLHqILopGnyZHY56zAB0ythaNgi
DxbXBMUejxpmcvBaoc4ZvihGoOI0R7LzpN0WQ/SO3bQ9AomtH9sRQtYWZKPYjsUvsawL4VeG1o+c
7Xgmq5/0/90/sioiB/SZVnneI+5ZcRn6bmtLRgyqfjFX3OFzehYkdlpKIdEeYfCbwODTcWDNhODC
sRik1EyfX9ia+cRFLgIMn5BlHiPTvhXENKQzsCZ+FxnuhjP7E82R3MiQSoa3SuwQdlYqH3L/toY4
cQw06uy8ohGjUPMwZK/grj9MrFoyQravBc96MICyj+ybbsF8wbwVfvyV5eNWhY5XbLX1N2zbWY+n
VIVBOq+DnbWSOBON2cjOOJ+LNs9bt6rkOFiGZbDinnVzk+5E1UFxCcljRHdugmC/fZLW96OcVvZS
bmK0S+KWv/OMghXNeUW9LS8M8yeUPSZWOsOF+Rjttl4WoSHRBiKTuw6POlByXhZKlPKl7BopJQec
+eX455jXcK1BG8l1e0jW0sandGAWQbQZR7nboLiYhIUp9eRFk47FarKeQmjwgTBCk4n0FIlW49N5
+uptNY8SUrf7ownZgyRow36bi8KaQMyT6IctuSJwavlvwctniCX2BabwMJcp5z/tt89NJMTGlhRu
hEOw9V2uFzkSGcPUOkotfT2Fg2aDXo7lpDENLM3H5ZLBKAgsNyXdaU2exZxSKWvtn2X0cQt8wyE3
tddJl8XPbE2CHZYU/ndj2smVWSpBr5CPssSCz1Z7dRx68O93GYwhFDwmYqgTkjfd9VFhgRS8mSpy
waCAj5R6emCGDd/1QHrOJAItjVAy7Y/dmu3eLp0/NIiGb5J0swvJTYWwecOScQ9EkHi9B5dQ2J/U
WU5IxIR/eY8GZHo9EsiHOVtleIF1OJjCe1oNmLgazJlQXFqTiKalG8SBgO2nLVQ7UJadJfVu+I/M
7GRIAFTXHX5PZ5Lt73VWDz+zhD43rQ9J96dIxn/s3PhnMn2stQTOQSZlZaXRWXN9QvhJBqJqAUaO
TQtjogYbOG8H4Vnf9CfJ31S/bH4i3wgQdKGAZJ9y4T/FXzzhxv66e8HgbyAcOSM741DBfkUle8dJ
YvbMEoQLnlDiq9LpmRxXo8YjHxWmkqDP260w3l2ff+xL1n49aPMVB82JqIocM/dl3qnemeXetMA+
Q0j3cdrDXW17J0DbzzVVrW2eXTew0z3WfrLmS/8FWMb7MP47h37o8xr2tS53nUjKcBsIvN+ud3j1
5i5Um++6ZIfUVJMKQ8dYRfuE7H3FZGha1Q9Q9YuOzg26NNhOMDJr6Z4GthrWvQ0g6OXFgzH/FrA+
9h+LZ1+4XkDKuVk17tSSvHWY/ub50EwyWFCOddKt+d0DMujz4ytMThaN5ReWX/qyYWtK6HMHNIbV
ijRg+y6mpi01dtvinr7Dz1D0WtHHAXdCaRn8+xwqY0TKDO9BMgk0kZW5xgskDnPybVcLomBeElx2
Y03Zl03nytaR2bq0We46CZxS4H08HLwHMPDkVRXDDKxMnNy9DLQMqwHlFfxkSzm/FEXNSbFiik0D
suQAdNkzjG6a3AwfgwDdyMc25KNmS1NG7PMuV+I9DlAc7mpeb4o6+hJWKnoIN+QfXGCnu7aJg/Vq
nB9l/jDss2jnnMW2hJfBZuS9fuMErgzqWuu7tWp2TX5asDfh5ozOgjwYV09r2+AWQcrxhH194wQV
dV/6m1BqMV4efVm7rIUosxx4yogJG1bUDvr+9pWEvc168x1PQzrdGy+yM3GOrfXmy3KHbGX7/Dfz
tumydCBiGA1RKjXj4cEDh5UeKWELGPPCKeUd5qjeCumjvnect87pTZCwWOvXs5XJPk8nONaXF3EO
9kt1rNY08555E9I3U+wkewzIXs2yf6iWoYSmVBL1w/7zQ/U3Ax/8Y1NWSRaWIivngL4DlD+EfThK
uVmvQ/ll3BDfHO5La1YI0VTJg/kQhrxdou/pXgt/MdtVB5oVBP0pLz5eBqhzCNX17qJSyXeIPRLW
3dfM1cB4Is20AtgRr5COTnihFCvLLvrzp8ruAFmFTl/HRxj7fp83ZOYCKpduw4HHlwyAOvwDaWy+
0MvyWhFfbwbAFdkSp7yAJGiDpCcqIMM1mYDM8rLHScFTubQqEl4/7KtNDYZfFCTPLYKkqn+JL8Rt
ZKqEN+hAozKCpE1/AlNCON99fc2T6PJufseDNaAwMwNVtq5dif1ZWPa+BMA1PYK315S5Q/2NWCS5
fWuI0PKW1k7rHFGyKbFb1e9yvC8nl2RuTaV0j+/MsxLoSjSUOdwUk2YMz83XtAn/52KVB5DYOTWH
qrX5E02YHAbMet/Wm8vXO7MP7+dsKywfoMTHLVLqfesXU/pxtU4sS+A52Ln3sPYaHxHj/UkaCzTt
h4K6+RZVA4PQkOBsLZEcrUdnU/dpIw/lk3HwRhGPTXmMuk6OYwta/yLnJzTNklXzBQR2ndmYh1RI
KeVrNxQvzwS7Gdqe/GafzlO9dPov+7aSP2XtV3a8e29PHb7BlWt+RDSiAqocaps0P0p0qNBIVDSi
Cqyp0wmc9YUPM2LLIkeTiDUrejpjozShTGT3dViQhH/jvE8qEPMJbR08LuZpBx1EQb3tlon06wDR
OxSUGxube8qC5o+EGpR6iN0FSxKBfD0g4vez0fMSdq58EE17G1tZtrCXEsexKDMLDyJ507d+qkjX
iDHe5Cn6RUoo0Gumkp5nOAzXqqDGCIl4fqlsO+Td34lh96Oj/Na34Lx5X+fQKHNX8qk3Qo4uft00
bGPSD/0X0v6pE1IbtCx/TdFY4hhbMaYLB+TqsPzvH4Jl6Mg3ShmxeyyntcogteGFv3URSKVmHwFR
Ib4/wEN9JaVpwCh6cphQUg7Ly1tRqzS/azB0tPB5a0XHhA+0JW4RiiSLmnjZaqpfEtN4aeV241oA
ZQOUT2EhPARnKWx2tfIA4mRZpATyXb79pBf2aKRP7yURP4ABOrDauRB5U2Ua6U5rxsH2XJIL6Wwt
Bka4JpOaVGf7evfVVCsHaKxObIH4dmHqMHRH5NT6LJcaRQZ5QIZ35Thd523mKB9v1CGhX1yXKmRe
cRayCmAsAyaAPr/24x/Yy5Qhcv35OgoSyhtqUdRvagnfYzGQ42VG6aiQFTsxyKEJRnmkOryMk6yp
ZEo0tR1z/b6iQlaJ3Fl5ln8nUVc6kC5/6839j1odLnD34P+ifIntumazzeARWYgQJkLT3iOleNfm
7iVd2/G5GWm9x12ziQD+YVAqiZGDi9HU721AVLCpJ7yd9dNcsUYEamQBLYLKGusYV/OZy3fMFhKD
c7jJHrDpr4cXecOTkVKhkYP0d9wWngvTzxxtrvDljQ6KvOwOqbpqJS4uxnNVKpEJdWSeofeEjMkW
OrQ3fSrlbiZOvv1HOehI64fLNCif5bwWCPfnU9wHwBJiRXdtVZ1Ij+g5LCy7OnLSw3froXQTVx+f
wjHrFUoX2q/NaFLWtVSRJPJULWVHC7+LTmxjdTkozmCwO0JXwUYxemNNwblfSNXfiw28vw1ixwJp
zUqF/OnNx+BcwjiG/PuvNgd2Ez0Ho1RKYH+wzJwBMUEfGZMJgHkxRfMH1FeL0B7f9IuyQmo+9oFy
IJ8eaS8hfyDWdXpsJLoHWyoeExPbyS3rtHpBN/9FQFzdVcLaY7Z5v7i6JVF8i7PlAI2JmCmdr2lx
m41Bt9koPcZYMNYWe5OM6lcqzuOKFCgM2OnayCtAgNw9eOf7iXeP8L9CcXnCSCEE/dJEQtsgSLR9
LnaEnbnFnxrKQ6sqqnZsireVFvEAZFqAdxI4uz7+n1rVPsSPs5CwyjGIvkYp6VPAsLulFdhdg1Sc
FXHDrk8wGEPLn9yMKlVjxK/6q0mYwJHbGpFqJ+fJCNYdbz0sURibQu2hslocRtNL4tCY6tjb99zi
lQcKGeNUfGK+iZ2KhjAtElrsl2x+6Ihs3J4AO410mFw+LO+CkqD7hU1uD/FzeHWqpgMtgwVWgHXx
2UxqzHLWT/ZeXP0N9UQu4aDCKbxGDXBzXKL5+cJuyHFLJoW8qOkRvU7CIfmfF2DV8MMx0/ODG3+b
5sKNLExW7hUl7MbEPrT/2TgwotuZP7yrg6VMcH6ZfDmQXi5rjccQrypVBsc88WGAkQTmJdcfRLsB
phS+RUOc+flUXNtTgsmufbM9SyQP/2PYkkYDjLtw0EIhPnp9FRKeKTdx9FjeuA/95RnF7PeT8rBZ
cv6OjnXSueHv/jtmap6sOOi5OH035i0PX1g+HqfW8c+8wqnA+WLeDBGb+POyjugGS+uL2gwRvRxe
IAigu/ppuettf5CIq7irctf4v1r2Kteq3mTx4wccx7I6gAMVOU5pa8gDNeoKicjhs37QKlbvTFWN
+0U95PKpaDRMSKPvhWuIA3T/ewxD7dikUtFi1E6yTzQG3BkrX3V0e8pMHNKjyZ1n5Sensa+uLybH
WWAFT+ibWeaLKlWnahWb1b4IsXzJY7XW1Cmjo/U3WzGq6yIRMTicFGrkl5GLmNXNHE/lzXSBfDuR
eL3Xvuama0pv8QHSFURlbpWp65dnsRYpH5WCU3nrAQx/NPNnSVEjTcCO0hBMvIXrzVHURGoWLsse
fSV2X4pmxr85GZq7jP9P69Ral6sSySx6achsTtl/YjlTDkjEZSHfNQ8o7MLrGt8ydO0rhpEhMgkw
SrhQX9VhrkKdUERoFjKDq0eJTxaz0B14RyAwoXcic2/e+gSWe+mATPq0l74MZTIlc8uT2/o6M2e8
YBWqbw/RyuZwHIxps6WfnnZ0rzqbrbMbFTOD0uOpc4cfi8gfTpwEyWc80XILtLhkn2ZzQI70C4an
nkk1Da4+TPrUcdV7YBAwTFs2PJ2mXq6NbQ8T9DHiot5LFgf7ag0JXl8Xo1qYY7W+BtjoLJKdv684
UfPQNtjCCwOYJNkANwXxN3JOdUXAq6pyprGjP/L73Fn0u5Fx5SrgutIV97BIYCDeu3SaNgga7c+m
mmWnOyNDI8kGcpoZNtpGuXRLcp1e94NddyDat9VYkFkvXqhYbPwcp7IGNttxVbg97Bog2e9wGHSP
Ag1XePvBwYAs4RJcwRLQrHPFs3Z/LFwBqJVBCbEWk+oZSsptLHdUlXlZlPXwj7nUyg7lgvz8K5VF
XEMH70R84UEvZBfoIbL6sySit90XY3pRYIX6G/m+0gvcV12JGYNJmStoWSpgZFpUMAaB6Pyjn1u5
Hom5vBMJOhjSxGhT2clD7oKuU74FJ8jT+/HpzvgqHhVaZK/KqyImNj1rOKR4vP2Q2aIu2mbI9H/7
PkEO6jXbn8lb9XxOJaJJzs8WU8H5YpGqXNZniEYR7QcevntEagXBr0abnBiUo0DJZTfhd0EDVvut
A1kMxhyyxCK8auyuv61fVlF83SR3X/zV0XjQzbP+6o6dMZUAGsxR/wJqmgvJGWwHLE1VlAUR+sk/
AxLdv/+HxwNUtLPXvSwb/hDC/br9m+hKzVJfl3gGCJD+Vsit92KL2l34hCOIgjL41misfV0KOJ1z
pFnQTqhaFCvYqL4hUFVZjzR6Qa1QGlOOkX74lhu8hJOzCBRTy145x49Y5/H56/FqWe6fAB2n7Ki2
X82S//5MKDtLrQasRdWPhecefcSqDdxWRpnnqYo9AC7wpvPsSkf/v21PrvVqFq8CGiO+77IFbIGm
K5ABoNl6A+5/qwvzq3sgpuxL4fuNeHij5i2a9eSA+5aWh4qQcPyje35oOEE8WA0qJ3aItBMHrt/0
CscNSX7z+U8B+rUuysoBW23eqFN2TQL605bdA8FLS0s6C948swZ7X+vkjlXbwAwheFVvLmxYFuNE
zBdULbNGKQJaXSGvhC3F7UJCGUzwIaWNckX4o0zXow/hWaM2tUm9MOp+WIECEy5y1pDNvv1mJFFI
fYv9/RSu+ITKOuAuzeRPlfJuc9x1zQcCgkOyFbrshOx4e7T1EzuluG/DZZM347Mrinu20TMilhve
4Tg/EpHYM5dWFhmBjeLnbVYviNKaOq/inUimfGP+APBa97tiIQZoZLCAe5Ruv0yKxcBBcginm3S8
ftrgrvCHTERDj3MZfNOU1NZA9I3wo6T/gPAkVmm5aVagACT7O7V5XGZTA8c+nOvOjfS40O3GLSkw
UXSDS1iYf3ex5jbg4dYbdMsFuWpl4+dugGeco+B95RiHamFcnW2N2epOJoCEIDWeX1SbFTh5A/b1
CVQWZyU1tDPQsyCv9mEewsmgA/NYw25Ht8R0SB4fRujMqXPN8DdOssytLcdUOt8GM68nYzsQn52b
eDLI1uzujDxLA0n7riqFT4U+oQDf2JWBqGxNGH4qV7QxAMkjDIkWJ9I1D3cXzckaTOJwGgd+B8KO
Z3OfwImAiIOiOFs2yDO3h+h+7b5byxWoz4q1fH9fHwFdF+DQvnTerboEIFuC2a8qkSfY/b99zJAL
2tqUSi2zO+0U1IRhiIDpbGbdSzGL4rDyFN/3M0EC1YsLo2OBUp8/vBaDZRxbwU4wE3cdQ0MmYJ+n
Cy0aPqpkB7TvcDwzfaN8iIlntObdDMf+aJDEoi25eyLwSeO3FSfdBCrI4pYGcBof5rV+AjWCprkh
9l/IiNlpNhOATktRXRXYTmb8AzfGqUg+476tEBYhIFQ58dl5JPNUPn4lhrwplrfzut0tDCvK2fKB
CWsAvpAa+/fK+EEd2kjfIsldixPHg6OjD0+oogTfg3vwnkRnADRc2lAGVGHF5UfPJ5wZC10ohYoP
tZXJZf11vblDBG/aRyMZ/VT9AQnDlVc/Rk70vpBdgkT6mTeqrwTVyeIphu/Q0d0oZghgySqT/3k9
83FbmAN9Z8kUUEAc7CjzJzhTqkQAzYf9otc7vanz11ycUuoHlE0AwPYbnkZeCIPVdvl/mQH+WBzf
XRK0mPnibD6N/0bSeOCi0BZ73hIB9DfL3iI3qjTtG7fNo3nqrD+QIo/RasTQzmVZoSwzcBRwyJhR
/sddPVfKxRcZRMUjHJa1GcrT55HAZy/3yMiK+CuiBEUqpMDFph80JnE0mMdcRD/yPhrHlyhg1oOc
KZmF3ecBy68rn2Hu0Hrx8YQ5iTVVb3VGZWANbleF+NtnfETEj1GrlG40ICyKZQfh49sjHIG8GUhE
e1jL/r2pClFTAM794tJB+qKPSVRfyyaqVC311D/X3c23duSzAfFEHVlECGSbg/iE07tDERIyD5xT
CSzBuP/6FLkJDrxeYL6MsMcS8Qbh0dOKhPIgFMkQtWLOpz17CtchIIsb5if27U2rw8LMFWKAtrj4
uC7Ri9+f+sVxFCn456SdSFkOdXt8QukK9YjN1yK4xSGLO5VPkalV3Fa4ywG3lY8stgtxjfCy0J+Q
AEbCA/GQDzLWrKzPZH7VtYHHOZuBWWWpr8sxlSu/9ALgOgtJqJHI6675Y2hImurTuEKtaHDW4PXM
xcW7xA2Px+RCQwoGF9r2AcF28AHSMeV2ux6yNmd0zJhl6afvqpwGPtfe1xZwwPTt/RdZhZA2gD7o
AjbAlCLHdNvYNyBcGRtaM75AF+KcPAQHKApMhzLfxj0CibKDwGwa0VLpOrTxm06I0YP8rOSiBVdT
EpkbBG91e8ClrSIfAAggZYpmN5Grd93ezQOxBufEMUKqWHnVEU/nhiDC3Kswi9zbJHfkyVqd35hN
7cmC45oDGbUu9Z2jiINfui/UdFm/6471CrOOEwITVpogVojwOBktSzLvcv74Ui5Cv53T5NnjrrUv
qhsQ1HRdkQHzCQTVp9rOEwPjwnPIKy0q0YlCfvi+7sS4osJGyxbLPyDOaCa/bHmEu+9fVfF87TVl
Nwm9vi4YmUnTwn89XgYWpqpFmtMqsycJ1AtMkR6lQK6X17BgP2Qp0aX3CSsZliePx3b9VxocAMmA
b+aIiWTqyWGlxBhkH0q//2LI+RYrBIftSIDibrJFIRITHSoH93sIhssxsafiaZdpQwriU7eroN8J
HVkLD39sX6aZ/yiX8sqV0e6EpHNj6X+ZAuoSuC68VkTKD4tpW7KkmQqXxbBov8CI6Erpp7DT5TPP
Jmd/mmp3rN1WFSEFHppS/gxRdgCNhiaM63FT9LPSDFar25HHzawLZW1Nw1n00q1jhCWgzQs8iE1d
Y23C8lKUmvHTs8t9mCwM+D0gdE8HS6tfDUXwpkMQyhok2Ck51l7ua/SISzo56EGBv0LoqFc/ir9J
uPrXXWiDzFa5QKt7vPN2JCX3TJ9yMdVR5holE9jqswVZRvKVbuwbRgRFliBaYIuGFRxchV4HOBXn
qcWkTUbir/fnayKfVvvBPws9cqn9RDuiTjZZKEVsb7YHDJv220h6tVPG9C6C0RoHqHGmyvQJA0mR
xKu07irt6aswZkHJFKrSGZTbqwXEjlHpODa1ykA3z7J3mJOVHQyMlsQGp/tsrCFt99CfoxRzXLl/
RBjXrCtq1INk0guhNXe1sSO/M4+MUe30rrmO7HKAZVFaTQoMvYbC490hzf+RHsUMcQVlGTOrLm9B
m1ZXdWM1BTg/BPDP/NNwrApRwwCnns2Q6HD/BefVPxbGUR6wGjFl8Wqc0CauNzrunfvw1931jUJG
UXzbgLHtBpdZZwjwK+WeYZtyHgv+yTXtogILvxYShVatXSc99b26BbRISCtW80Z7Gfqav1FBlchL
fe/4z1dZbeWF5hpTo9EIDkG7JJ833pZ0/gePckFW7ZvtLtl0L6cW0TwPGW3pvO/jeqmMbiBmBgUV
nnfl2EkkK7rQ0TK2bk9QZ4oCJoCZHh5633vxWflaZiqF3+j9lHwKPWdl4Glyfm2Mlzz8OaiTnY9c
0ezTgEFbTKT7XKwKucQvRKtICwWtyUBgx389yN9lPRA1w4Q3ktBn2MHAkYpElLYdhWX1CIM7duDG
N2E16Bf2q3eqqX4XyE/Qpum1ZNvTDXWaT8XuEp135LI7tA02uR70nFMAcINMs9roWCPWIQC3y0ls
7IffBB/G6R73+ej3+/QnqvqwSz25RtNSXMfW23JLsSJ8AsIoZ5crbOv8tA32LFYZML0K/kIm58Pd
Z1ST8aI2r9d6CXH/mmXl2tAx8TeXZ04poqle1DWTQ7H4bhRiD3E82rEzUqBCPg6x+tCyfDiUAUA0
om7Bs/SVuczu+O0KMf+Tha4+PwcD+xP9BwulpZQCUNtsI7LuzbNQ4+4XmeSwgybXeift4PjvGbAV
zsexqyufXWGNrfrd49t4iFeHaoktH2RWSe/3vlLqIEL9otQhz9Y0op+Bz2Lmlgr6NsEMKYjQONc+
dHl19s1xowAkW6WOpLQpy6s3Vxcqx5K0aKxIEThupgBe0D4Cr0KzM4jXDvNPkPzECXQO740V+8ib
Wwk8pxjW5NHyVoO3vcnM6iRM7QmohNbZiIRAH73i9fvIWzFTcgc3VaSztjDi/o9KvMlue+OZi6N3
kU1SsHYSciV/RHnXPoAASrue4NEbeh5ZI4gP3XyrGAKebhfgHH7vy+s1GL8TWAlicORiaprJ+RSa
SyYdmXF/26E+yxQTU/nOQqmypojNzVsfcNDYI0A2D550TGjt6U3HX/BiUrIvKMyANPzOjuhmXo4B
Dk99tdftUEdUJxk5cR5i2mlaXEG4goLZCpDVMTC+LldUe5wuEY9EkVkHfGy7fSCl1z4bi4aA2tqA
XmO6HAcywv5/tVWrJF4TvcBMTJsbcMVk3vNUXbcJGEGckm3qV0j1yZSm8sQc997s0XcZpkTbIcir
D3bQRww+znp5G4hSNxX9VeJJ2+twX73FnD7zaKBEDarggZFLS1Vgo6rZ1A/yXoMTOlcpFWr9elDN
AZzLqjAVJNWa5Vnj8tXpnYfWylzQ1mtDk7JOcX+tVLKSWrfeRfrjetANwI6YhMakZ0+yT7/ZpyyA
s0YuRqsdDWWFLDGZDfQDHLsu4y/M0vRW/1+MidBHTgTewbhFasOrMsXmGUbqGpAk3ZMdYWeLlLwm
V58bfEvuwPN/BnvAbruAoaYN/BcJYVzaRtr4tjm0ycP4C0AglFDMbPDknZWxNWvP2eXwVhWqsUYJ
h6pyaapcBWn5zskPty6CoeyoN8iBGNf5gVP4rzoiybBV8Zixk7BG7CkYiKPHx4F4BB7OUqyg837x
ZoMq2bX49c8j14SepNoG/WhAoL2kNUSgV/qfgBg7B9680KkgQUhpVVaDHSNCF7fvq2GV1fdAAbt/
Nne9TOOL1AmpNUWhJRtIXwrfEoYC+uyR2jzzoOL/xEpYOjPGH7+oVGaFMNAIk4o/XYwWEpR8TjS1
Vxz1vB+BTMXTccfCT5jGIxGo3hR/RjHTlolWbFUsh+xgbRw+uDIyxaJN++UKEO057K65fskaHMFR
lAOewSQnSZlnPp6wDjfLyfLAFo5dcwRRAMTdrDqg+TKJFppNX/1NxCqo46S8/P3LWMok/x2gRz09
d34pE3GpFHHcFfFcVJ2WdWfkaKILMdCyWKprGNRhNMSQW4bRblsPruAnI7vq4UGDhwaiEwJKXNLH
FGFWpx7sdvBPPerMXMhEnaFtDVR6nKM0Kh+5J88zcgWZS0rw96Yogd18ugvrus4j3QsmHV8DlRyx
dNrhV9i5JumYGObghdpo37cE5gYjfJ9A0Yo6cq5IVt3mZabfwN5SupnHT7lqERy0teSFnfEeLSsG
dGi8hEd1uGe1KMM9vXgNE9ERju3WzrvQDswZs+6LyOkOHiVTMTiSJdfOCPwrXbhrC4byY2k4UDNk
UeLEccmPP0yMfI7K0OtdKh3nNKBTfjELIOAqBkICaaCqU7AreuRwHMLbv2NOv2i2P9sPud8atQLN
zfq+yes7L6NJ6dOme/OYRsxzNnPnOFvulWja+VPi0Ue2iH99THrFursDSfUF6nIvwAhaES/Csoha
vYr0N8CuKax0Fb9qLI8OnjMTJkncLJZfrki41gVs2a50FNW1QB/Pz5mGEZSdq9nc0XeIpwubYDl6
dg1wFMO0z3GFcOFIQY23A0IE6+2aHXz53SJLM46F1r+qtxKJksGk49Alwi2uKACv9/+y8wocroWf
9fknkIW93Aiy7V/2/85EXZkfN0J2fkXnOEDP+Hl/JV214SXDvEe8t7s90vyqqSB9Ioo6eP8ns5r6
XLl1PqjaLNaqgvPZgeNcbT4l+VPiGDhZr60tDf7x38KeWygm9mMFTgTAjwa+eUnNx6VwDnwMHEaR
gMbtG/QeH4d8f8R1dRjBTQfhts5WqpSG53bEtAPGvyM5iL6/CeP910pcxPjm4GHgqZypy/D0UIkW
BJfYmmSzM8fCB4i0XimBL0h1iqyjHHsZ7XNNuRberZM+WddtbnFOmWnQKsTkw68YTZdRzK8pz10x
+fyAjHt9DPgLZoQEJkoacEBcCaM1mVg/UX+lmdLt79M9dW20KnJjqp3MsBIW2uNC+z3erEP6jBBZ
CqPwvUwxmjgcGQvVifrmftCIiQ3jITixWiFVXOq4rUaKLNJQPwV404HSzxqlv0IFi5I8du8xL8FC
4g7Z0Gbn7k7U8ZDhO9+7HumncRUISXoTMhAY8cojhFxEhwdBjhpQnOVW3RQZJu3VDpTO/FVpuQQF
IVhX/c36Wsw94FFy/G6X35cjcdOXec6bysCoovXKRCOtKIjwhpkYfyCLPU+3sjueKwSc4+tYLaAJ
KKDkV8w1xLfWyaqQvqCGRrCtKNtqsT0bFD1mhh3VGEszdk/C0r1I2d5xTthgJpzmFrwzgjGJm0me
GqH9hIw9RhwmfoymosDSIq+RdV2Y2r2B96oDbwXBYvq2EcjojQrDy4uR8jc2vESZjxl2gN3+yTuk
LIpQN9Gj+1QF+Q96bvhY+6j+nVXOOFWYYogYcnGcv4i9Pq9EDuXr2QQtKOL/LfpKxXfD+oOUOIHF
5UYf4sezaSLN8xUxUAmjJkKL+L60fXlXm0zRSwPRdoHaLiUiTq1PaRXbFPFFmVr3yf0cKdV9xQHn
wkb1jadZsUDYJNpWVXl4XLTcWBkfXD0K/NR5YfGSCsC6XiL6LjGrJjCSbKBQse2w+wW3i/DL5GsK
zS9+5wM/o3E/9msI4z2xXyCmFrSrhxA+XJc/qq5wfmPZmIM6rzQvFSB5HrC6Z2RiMJ2pUxYLIgFm
xSqYN0Vnljra7mz10B4nWhYTSiii5woF01sfBbOwX9vqLBhOr1igDFlLmfPEpwE9DXxEOP8WVGEH
NuygK/ScT4RSa17aPwfrSKUqzuctalFer1a1O5Mf9MKyERp9MYBlHd9Ve1uaOGZkzf2nvVA+O0ja
LnoyG4PzHn7BgL1jx8Qs1+Q6mg3zKzZKHq5OEoyDxoJklnQ32Qzyr9ZLk+YZfYR0aOE5ZmlvUkSX
NXGF9Vc9x0AGuDWm/DCws4PG7jyDP7pJhNrdRq2ZRb8hIaqe7SAvFS8tTTXC56jGjYtosQxLFGtB
FwYbvl9OXnkdvrPzjXYpaTr/TAkFlSLX5kOM4wDe6RRSZ1xOzQt04RGSVkgM9L2mYfzpOQs4HpuN
rom+bpTGxDyUThxM7G3ZzT7OdQiSvJtIl68h9ehVnp3uTrv4Pf6YIhXQvTxy77/8giJd9ZoNSne+
0uxrT0z62FHxxQRQqG2GWD/gvYkc16K718zxvEJBIBjJxJ+0QxPA3jLbNZF2eSsMRi3VGe8rIhkZ
kcaxxknZXk4NwWoZZGnTLs+VfDJFFl2SeJptr9doiwfmmJdDRb9q5dt4KPk19uDogG19GcYXgdNN
g5Bp5qbLsWDAiD5VcaAPGqhiV0Q2rbwzeThEEuuhHlu3xuw+wN3pa98nvJDRLHtJ7a2uf1ysJ72V
0yayn2s6MeiSrk2xARLddgEA4Vi13e7g5K+JEUf1/nD18BJl4W/b1KlOxUqf5kA8eOi6psZ6aBp0
fX6nxdA6j454BwJ45yCKSiCA18OMtgXJPFkAWuBOJCR/9BCeRX6QY2aGqtazXLoJ16TTUVPt8NNS
rYh/5J1NPTkBm8ux0RUqu7UZHHYYQPVPYqxaPoxRaAzYuDGElmcCca5a7Ay8u4VgrYQibDS8pLrG
OJD1WJ3qD/V9KrD00BQWp8auzBiA6f3Fixg/QsKItn75P27y/1dBw0+JbCw9viSdaWi2jG3eOpdU
J3m/TdTYatbbgL/BBZykGMNKNr29N39OADPOJbyf+UJfqcNKKIGrF8Ps4ME7MvUYg2N0fy03uLD+
KCvPIl1GCLCfQfBKfmHyrNXRWc5HJvjR903Rg8gjs7y90QhWjXHgYWqXjBOBtyGVTmmepX2Ow1Yb
b+5VNiNpXYohgHA3UT1Mh6LchJw4TVGLjAcrVaeIb+SIsgH+NuItY3G5D9IxKUViGsGSRa1F/RsF
bf7OvCwq8N3c58qDVliVmKyg8zdtCU69FeazwVq5ZrnMs2ff0Ylckh5yqzWOsaRv5ufgA5DkdX+Q
PkKmsvphjHBFZYSYtMnuASF/XER3yW8sAUEJl2uBb2N2TslMpSiTsa4sVfsGXOdhQiijnlvq3b5X
0CfTVeBUD8Yf1yOsfEED8HM4oSdTeegfClnP4aK+9LO3mzcHj8bKrzGNXY2yUb/UWRLGkUeDaZUt
PTE5MWTwFpF6Hi0r2FfQm+yD5/kGOGFg25VCmFj+qJ6hmfgDz0M78feHRCkHaL1QNvG6k6txG8Rn
1CEygl4h9NWmqjltYAYJRSiwvDKrNqA+bpRMGhA0TOvIwD8zrlBEGLTNKiU1lTbqEtPTzAZC7VFY
t3CAhxg/cj09lFmUfIH7ddxuGYhZsDQef2f/QHPxrdeqwUjmaxCbjWi2PNNj2E4qIATR+iDmupzH
ZET8V5rCAHmqohtO/nRY2BFdTz6pdDRd9ObvS67oVAkJgExTqGYQGe7IFGq4yndToBbr5eDXqFWX
I1WUTCHbhaih4zKVt9NLawFE2asir4CVfR+GnOcdw9CneLDWZgrX2ZLGCLPMsvEJnZKzrsLiyN/0
GWSw4rlJ7G7YMZimM5yG1XhlXa9nPaBs447L7Tt6Mv0km36u+8VGxbCy9JyWYQv7G0w/1NsUhjg0
tYkB0e+JXRyUUlVZTX+ibCxanBHq/gQkEkfVq6+X0LnfIjNCPjBq5Vcxa55Am6HGCpL6K83laDa9
/rLB6kLrluJL/ZY8vOYeUG65EmuXQkuaXAOOX41KmPt0hoAfCr9gxtDHakaMwYtXYwAEjXkoN3w0
mljwTPDAj0TsGNTscpDi5OYjVa46r4SeUU8nlkfSbMfC5o8X4nzjrep5nd38VaYXGIhHmijZLe1h
dJY4S7w5bXGTz0ntNIxFKXiwLQJ91YNk4RxP3Ti05wlfcF8FUhYXJIaWTX9dDdgjn6fEczN0flaY
WkIjl+5ktBYW0V4pWJAJy+wHnBHNqJQREt9iUNe8IvzqrDBs7+IabIv1Co24tFjcVVLcWmPfuuQs
Jb9oW2aD0RsfSCLMRbGaZU52cHdogvZubomphWTxGilEaGVQ+Tn8Zz0Acp8d9LAaJCoyvS6HRIZK
PYwP79z7tM74B6+PVIjy6G2dQBGLXM7l3rWlvDLXpgXH4kRzQwFJO5hjvI24OVDcFNmx0RjGmb2k
7tQA/fh7pEqUmWcMzxqPk9kg/gV30wIFQ6eP86XmV29n6vmhExma2NL+hEHHFS7ypHOhISX9eNqW
vtll+nScL5h8P1x1H6c6LDkXa5q17absXOQVIGwWhiHaeCU97uQYVfggYMmfy3vPzQKUBd2hbeFo
U5yhw5TJSvcybfYWM/8tJ8cZ4rd3acoozTz0z+6x1gDMH2sZHueaTmOka0uo53YQWIJwFgE3MnNL
Gg0tVqskFtkN0YpRI/mBkAQ+EK2FMp4I6ALhLSBWC64Oc6nrxgdiufoQv9GWE1HlZ5cvUjmFCrI8
xJm0lxnZGPHpDUAL2Adp15B41MuWEqbKK4g4MBXULAEpGLDkRJckmTaicWku+Z1BAnMQCxxI4ooF
PHhAzplpo4t4Kpp2P14Hs9BFBhRWZ9kWb9Do7rdhdWIrj/guGmaOByPzEo5MGoCtohrHbtuHy8PF
WhuSJUCvNeoJVe9YAlF2JY3pGviUwaHMeTCDQvh+WAwyPsbg9eOzIknm72x66+GbvflzBUR8qq0v
4g9Vf4F9tOJvYoNGcORkc7eLiakqh4JSTMRzznNWIH4LYzYrdmTUz8WZ9GNSDNcNaVd16ZCWOtSU
xE9ObFtI65yMn9Vq+CNC0qRyqVBChhQ9CB671dggOAtDMrzJsk2DyhJgvRe+Y96l8mbohLtwr11k
bXtbqAnqOIge6QpXw4SBfUOmlpFMBytI4kRjcpTCaG5BgyjxFmspaFpTKVq+9tba/6P+dQ5pFLYZ
3PZUDlFp3Ly/ShMcmCZBVxuZ4bPeQnLsL4xpJtylft8zg3WaDyyg7vMPMKEFty6gWaWDNrd0CELc
RfBVhk7/I/WLnBXEVitN/+h4Zit5IVQRdDl+au7aZ+5OLlJdKstI6CEwmUCYH2AAvQv9gD7+TQeC
wiwYQgr2+FbM3QtNbUHfoIPvs06+9j63VhDLqDiSrKCAnCSNA6urAqdBw/7UyznlQaGaz5s1gQ8/
2RoIJuRZLm4S2DxxvTQH5rBgPaws2q1q4dxHb7IJbpnn+yzp6dnphE5ULLwY5Lh9YE4RfWyFYSTx
Vg0k/iavPBWTm0b5iqXmp64phkjI/bhyWHUnjXCIAs7kb+Q80kLR3eYP5q0PejosyYYyFpW7smwK
6b9K9Wozl/phwYS4hfRh+a7/+hWtrc9LAYduHTCzBDfDLjThNcmhAgicEppWCoJY06UQ6d/xmk+f
OPG6EHoXdHjG+/4Zj2ycGHkBZJdu8py5jJnJ0ND09NyARk0un/eWGZXd17pyGRWjSFBtVKmNUBmk
koZHgo+eVH4dlQchYn/zUDNhiNN7Yj8nt/ruZeHr3avLnD3ULPakVuauJoR7Xa9g3giga4OKfD/q
y9SX1UMkqagtkW5ZrHh4BUu+hzOkjcdV2IapnzCWlOWOYJ1doANEcAJvsfYQhVXpjNV8XHKVYY3G
r+plMBTj+nlRuic9/l05RX+bIYkc3RWJCE1pvg8jJutnlhbDrHBS7g/JaYObh4EOoI9JGbV8THGz
oNARBkgAzKgVzPD8NQQ4Ci3hG5fUkIBrhg8l4dpXhpJJ6sPyPtdOZTGUYhs8Diaq4aE2pVGYR746
US/+VJPdLMnxeRJNI3/GEC6x0LJvB8n3teXaraUIgc8bQ4/lIihzuD3yORuLR0IxJX/o8srQg4mQ
lLzEM6RzjcxbsphClxyj/R/FoHJUELhU5/KNSpIEVRKy8Fc3t/D3nM0g6NHUNOaitmpYIVKRyhI1
F0ehiJ+lj45UMkEWjGlDOc5UCPaGgpypZMB60QtmIlF8V0oxb2z3tT4DhAy38G0jJ5tFSPlWoAbj
Ml8aDHrQVIiCHXsnPFNN7w+X2A5TtvQoaD/KbyUvJEl7FnOJyxp7+GlAxUep8ewHj/ETLxhckJOs
ekhLtupNCE1YhUF8aC/VMZqr/vULwVEDNLwA3RgZsdTPIrXs9XPzczfgMwvPAugF0NL7q8BVhuHb
yWDovQAs4VaIWa1O/PYL5+aCHpEOIB8sHP/nn1vxP3PaGSIyEpkKxA+xMPGY2yIG3puqnjR8rKHo
38KH7Mhhg4yhqsqnmrAWKDHOAf0UhHY0N8+469jwcJ4W16ydjViQRcpn2/bJKT2WjIGf9QU+BlC/
KT0m1EUR95RQaArrHwESb9CuTra7xz45Fhr4eEsfuuQGFxOOc6EsJPPjpzNngRoRquSOBAG/z6Ne
fbIYXZpdQvY2qKYHYDG3+QLJaOrquOORpKgpnEnaOvskRUY+jTtwTtUSZ43cd7U4hRnzMq+9kJnk
NambXmF2yAxv69kXhRS1z+Lk5oRo+DtNUArRLRENhO51A/9txhD/YWpu2z4l+H3KuEy3kP6Qg+WU
1vV0mxp6VDLhNbBKK6oKW7rrGDR/mmPTYGeztRsfp6cLKaAlcuSyaiyfMO6Wj4FaL7ePH+7X1fIk
vESLZZdxISwLF/VzznF0pZxPl3x1p+49wKKGE8dgVI3PNrhSdSyxJnAfMVvwAlct0PsSQ9xoWoV3
h/l/LT8P0P1xqXvReV9GGDqtn1jq59YOBx3cE9PGPgHMO2zPA1beOhfWyxgbvLikBlg8b0JTNneb
PE6JnomdkpSxpjt72Gq9rGWqvJYRjIzCBAzkb4KXaDWqZjy0XVceatonkRN3XptfMltydWnap52t
hjsKWCkzbmFTcUQefpLbX8Tu0o36U1S2wiWS5arFZLevs63x+dg6HDuLrmrP27cXxlu3v2k/6Wa2
/iVWPIChYJwhEtIk2EO1OOnuBkru5nMfK9MKv7R6rXP2rjQIQWyJ1CotSuEs+NtMnX5vPTkupYFW
AAnMLYR7NybzyjMwMkOkGf+ZyNEQn6MSlUPS7WDwk2UNhffXXqNRQxGlBpnqfGQUXEy0+iAWKIil
bx2yTmfiDO8Uctc6axdNU0UNNSZQT0aWXBcqfJtF4mDPZJsxZ/OBlul3E0yofuzalPgit/RtKdvw
kEc0yhBCnzV8mDkDvIcyzLuthx1kpgbY6LDIcBB43CtmmS122deXnhmOkTxMKJxNSmi+PJ+WpxlZ
eN7Zv0YvaGVigsdUhkmZrH59jq3qq3FErGXT85QosMAgBm6Dop0lKBupQCO2wHBpWhFGBmHifNe2
xait8JiWuVhIgM0QDY5N4ILkb6eiA7GM2OYj0J4hlKo2FoD7qFITdbYtUo1ArtRz92IA9ae4Eufo
yz8E3PZ59dCPdy/0ZFSyHNm8QSf9V4ufuCrebNU7LfMgFmOyJfuQGV+Y8PJH/yo41EdIrJFHhmGz
yrLQ8uqWp4CUgXTxnsl0p3JI1YpNzGKUMsELbzarRRFHkCIJKg1wZeqVXFIUr1zW5QFBj0d/vGfV
+LftsEcBjHXzq+Ky78DLKNa8rsn81YBnkqjtT5CPnzPDr2T4cjve+Kt+sfiQNKp5W1cdw7Y8NKHC
AkzeQxVWujbmn9H/1d8BqESa0sU0zGHWRwfCHkwgb+jgLc8BC6AuAQLM78DCIVZKRmI+d1Nf6+pr
Ebes8DqgMFQQnxtz4YU696ijan5XBZyyiNSh2azPJnujlfR44iNjptatcfXLDuKKSjy8DfesesAe
GnqPUcgswQhSWrz+594++cy9A9vR10ixLtJkeJW3BxymZtYVXo85hbwuS9eRqz58fKAQDsIVasa3
8qz9XcjJq+rtViGjCxn9RP049GC8nQiEb+RZex2XdIfvSfg6f2UcnEwXUuAuUeofxKXQypXHSQjz
K93KP6QSYD/ByCZ7aJ17F66jbpq2PiiFuW29W7aaXe8GzkyN/IgD+1Q47JYA5NBvekTHsIzjqE03
Uxn8QYUheAewumlJJVJyEzhHvImKUyU266+0vXjOyLEmQqvy+1I1p1VPahkv4J0jROPhR1KwE5Eo
Ue3DKTmzO0cGGdhYDzf2D2Nep3tGfbNlxBrF3RrSzJoG7TYTtEPyU0hNPaBNf2BsEV53GRI+0Mmc
y9R8ixu95WUl1qX1q45wVDuCHkDSpADx8DItinDIso3CPp8frYFbnUTdXX7cYPT0s4l4H6/dxxjF
dmtt/NMx/BDD2viWeZxQ+PKtPGcxdCewquWlcisYpP+F5oHZIVsX07ZSPiZtIYvtzZiaFynQPX1i
BfNYG6/BXNO+1U6Q3J1/aNiHk8zlMTe/6Q507p5EpPbzQW7/xDwy32oH/ysCOAN0HQuCUh7QN2JW
vqyp9acZIFrT5TVUn1OnDOUfZ/XkornM/b9jwSDEwlim1sx8iMwG7kmVQuoK2J2C9TQWVz/YNOaY
PUsteHp2Y0pjlKLbXvM7PNBf+RENVEE/pikcbWfTqK1CN7aNFeWEmA3ExJvKDKTr45co3q/aCTri
qjI88enmarmGdZoKCs6UVC7Ght/7OkPR8SPIPL++i61RlrtybiPygGVmr+qTeEYV9N+lI78huUzd
zaPJ5EYUCEcZ/DciAcnJqjQXvGn043qcgDLABgyNj46l8zsK+1ZcVi7XkJRC6sp/m7zbj7cZGrqv
bY9Lk6unPX1Hpb8pneGDgqrZOgQ0vklULTEzCaBFwlWAiSaT7CfWduerhYTzpEr+bKNJm0OHXiHR
O3zXnipHUab+sc6udH6TUI9m1igYvilb0NH7ySD0B7G0ZwCgo4Rqlm1attoNVFDDjQhRJOAzoNp3
0HESEL/Yz41TtfE+Uva6mAmtqVN+do2SEFLBVjoil3Krr413wi8bcpmlYCcOP+4x27CYBe+slhaS
SKfRQG9Fiox3/+ZHJf10PtCDxLbmys0C1f9t8up10Tv3I+43+A5wW8Za/5sHFHqlUminZmLeO2So
D5xKa/4aTC+rpMAoRmHArRDdfx84stdAFWqA65K0InVPHz2QR2A1zBlrdSbu2G6yOLM6cU9zJeVw
5AdN/3syFOBpMqMuqjpuslZ369zmtEQ9f2Rx2RJCGCmqpHERK8InZ5/QF7m8iwOOxDx07FCyGnLo
Nx77sTotzq2YzEWmhxuW1TcAteUkwuzQIgEYRZl1XBxnNPZwWdg3DhV7N1r5tGELkb1pW5LpGPDI
WzATbxnuT7Buq13HaW+qocyorxe/72VhyUSyANCCtUM3zPH7mnArXlITRosje6Q2x9NB8dYvf5E4
m35b8gc3BIR0JSwu9MBCUPwTpzPA3fa0g5tYAEg5tH4UtjTshl4TjT/WjmUDrZRSruvJmO0k0pAW
sqfPP7xMouaTKwdtNhjeiqnW7TpINJRwM3Qs02HWOcJT4c35QgVVpcOl+EfcajTtu+eArZfek2gH
cmRGl2smxFyfYYKEAQeY2y2gBd5waCgqG06enCM+VnsOnPremC9V1kLx6tI2GY80LGlp4lXErLbk
NwBY5WSNUnHTKHRN/2Mflpb2KJ8xPLYfpMbdoeS8wb2sLy1rJ9eQ+dqmAyejoZ9U1iJZ8lDHXgK6
DJjGvRjPaL8UW3hI9s0RkY7KKr237qBs5uXHUuB4aTCyQdTLZzatLgOP7/5Y/RryLXc01M2ZX8fH
/jv9mfU1QPaZKK0XDkCZf7aG0+I8jfHl00/pFTokv2n+av9WDnhFh9RR/y8Ivg9fnIdHUSLKwiw1
N0UFzejJ758Ab/qzIsuxZ38WgNhxxJScPyojkOkDv5XWltim8nMrmc6oWDhhfup9GCtknUD/PuEE
6p/Fl04PQDwaSTvextyXFcYR66mKmw7ubSMzlocW10J5FVl68v3MslWN04zEqtSlDPZif2W79wKG
chNNHeHeqDv3uidsYCqT27dTARM4Z63XTdtvd38Px0Fs3y9w/pBKkNfd1Z7Ekiuf6NZWDQ9TOp7U
Mu9ayKYOnK5vmkj1KrUYpykS1xl+umSENAEXSLyC3KXuDT6c5MFA4zJPM4NJJPFxiM2i4cbPoxJL
6LjWZWLFaYaLCEJGSCDNOnL0tsr93CZdL9XCLVVDYh9qsWIR/JCVxd5Jd538lgiGWE/MTVePIUA6
5Rroy5yWo0gFR0tpS9PQARYFyr850cUTdqalPnifTSKPt12ZFkp90AEGHNMZjhwZ8itfzEYoVQzk
518koXhRmetoJ34fFqs+vT3ZpOehLZWMuKLyS54ysoHbPUPoxyqVe8qtVYLHVjroF5OWOxkRNWgg
VmyF2ZNC+c7BakYs4chfsUis/kuCGbdtkXnNKyHs2jQQaDC14ym49+ZL0gGaWAcpNp57Ufy9MEQa
crlOrAIKDVIBog+VaJEQrkWT0Pf5OuxQNPTV2EGY/RfWKOmI4bg2oW85hncAa5xdmRHS6W8NPhOh
HUBWCSXz2WSzOUFeyxKywn38YukbJzIME9BoZWGnsnEhfSTC3a5w1ZT0q5qr+A4p4T5oR3n2cBaP
3knsNBFJfVVScnJ6PSmvdqTQLwLTeR4RqPRZRIz/4Pd/OFDj9VgFRS64kRXMvqRAgT/eSX7J2PD9
vyA6n0Ve0mZpQ1Wj5E7oyOir8YGhdr4D/TUpO7yKSf5kemQJTDdWubb7V9hxB7qrLfR6vEBeqGoQ
2IuS/cpLsph/sWNBEEavhaKWe8KfFvYrSa2/sjzMq75N6GFVW3OF5cIYvfzH9K/1PZ3yqK2UjDGR
Y2UecJVxqVlqy2HJqDEu8JvbekncUmyTdzXi76Gybg3x1YIwBDLFa4kJimgNC8ptfSirWIp/qlW3
+75jaJZsj4zYLVHnQ1rTm5iqLXe3svW0/1X9Yg3uyl6ZQ2eqjFtvzdYFKUJixfZ4HibrToxy8MRj
xCu/p41ykdq/e5d5EKt2qmNJ3pCKD1RDKRc8RSjy2XGLCCVZTR6J0AIPZe7TT3d+n/MUbxY0sU25
THwcFT1X/357e4KGUcn2PLTPmU+OO2C9JH1dbBUhR8K4c/ygnLq5BP22atmJvXPONUu7VxamTDQ1
8pB159O0qNnLNNTRaDvZO+CgtXOeKsorTSQ+HDFJpVKbMOxvjmwjjSEHJh58f8x11mZZ4G3w4mf+
BZsMq7zIf4KHF8hhJNG17K71G2kc1HipDnI4HUcd/NV+T9HoQNgW96dguPSg+oqn6bg2I+o/qJeC
SZK2NimraEW6M2XnkAnPpTxJLDhlfQIWGah1TRfAcSr1niq5inhRnYWAQ5UYJIgBj36xwn6Ll0qw
XIiHtAFqM9oOThUVjH0Oy6fgV3uMxgvtqhKt2KYbiquhGxVRkrtNzDkStxEzklFQ7pw5bC8SPWyf
8dFFLSl4Sjwvrui7/tIKbij7x+MSsQA7oasaumI64GhiWE9iPjzU3NkJLrh/we0f1/BijMAQrVZQ
gV+hH3Eh76rls7QRHjveUbdaRcxtnNNGav1MtQUxkrFbri0hfTVIzKSUEGJFcaFrOeXnWH/dMd9d
KgqhPsIYsVNRZR3MHsMVgSWk97bp9xShGj63BT5ZxuCjH0RaSP4aal6HSDFb3fE4+VdzwiayR9B5
MSTRV5lm6AmhDgwChAJjpJvWfkXOl5iJ36OcS98I7aAGlkaLoquxuqLrV/eNpKNTDP45eDDwCHKC
Cc0T3i2tB9D94cupBoXfUTWeCBUiJEbN6pbfeXl6edLTMoUmlfmKLJG4YIkJS7Ssc81vjvZ6KC/0
1Lla0fzAOeS9Q3FqOuSmImBwevN+3+I7L30gPPobwGR26TTdt6OJ1CGZi0YefpyOFDXun9eSxt9b
Rl2YE1ZMwZBJY/Nt9Rpvb0fQJ5Nexy4FajA6SCt6QbM6dha+6/yx41gRLMRD1i059RHiRwCpxe0h
zK8owpWSfh89lBvMYt+OlSrtC4amDbG6s60LVdYW5rf7HF1LMdXYlp7iRQdcLy/sJGGg7i1T5x9X
2BvhKjyp25lBc5z66h0s5Yltwjk1oPqM3xlTjroDg30taTWVyiBsIx+UeF7la/nmkcT40Hg2Wup/
5buis/wHzGNmdqUymFYCqgZhi78ghz8DNX640nghPeaGNegxqZkGeWarch4msVluLqTgZdL233+U
YnXLvTKHzxYrfNuhp79bTosW6lj2L+D+JeeIihBM0Ww2TsZ7EnuerpqCfHFGKJ2Cr5aX3xWAAqL6
ANB5iFV63w7SvVW10lHvP8u976hk72VLXE5MMOJ3RtYHksjHt3VXTqIUYQQ29QjBXYmuBFreP52t
CjtmrdfSb/GCtMwb7gVKWXl3WhNkHU1aWq12uoVjBoHrHfXD27vbC7gtXragiku9DYX7m2oZkrL9
t+PxG7UlP+WXI8tyd1N2TelmbLeHHF3+e9WZbhmxfThzP4cOyAl1bWxh95UgqPo05DBaP4cLbw7/
ZljV8a1Gd8zTSaAM5Qvrm66KIFMkuhh6WKjTFjvCj6z/VQ/2uIY9lVIJAqd6s20G3OriBfRkdZ+i
DESwSN7xDislGewLeZPFqwJMeWFF8BV7rFLflFRQCgnS+GT1MMcKd731+Q0b2Jtr4VlsPxoqQPoX
Ev/fYh/Nc4ngMlO/6z/QS2Gjv1BYNY8xKwHuFcbHpqF4mY8ve0GDOqGBFhSkC+ZYc3pK1IhQdON/
Gz7k7HczYS3auvNuTntOjXBi24GatsW67gtAgZc0Xh0pqHqKhequUYAGFSINyhmPYlZSv7oUWoz4
gx/fhicDwU9npajju/yQvy4/0EfNrDHg3Z0t97lOmMk25l5oX4F9fJEx0o4EHhs8xw1jGZl6JSo9
SmuzdCxDbYdUod1EEhWCtfjzgj19VoizAyGpWzyqQ/cW9tucHGn1TGWaOF53hmf9CHcoQ3Ix3cD5
2oMJGGTiLRhxF0mwtXsqoWh0+kmUvwbGGupTA+3xvA6hBXjwJK8TwBqIkafdBGIt0aTsFZg489nG
i6ujU2FaIOvDJFu/PUSh1RuASTQXph+E1CciTYBmwczOTXQXbxIQ37uyAoJvjS9CCsRL3y0dG9aU
UkSUNznuS8cbblQnv9u4nDXVHXt+ENXkf7Xa7wMIDPAoiF8DtloNpR+1t3YIGp7abvydxjzb3neK
BySgfr4Kkf9Q1NYgdBHxjnNieJBOF1VD+kw30jQbyZcjuU+Ua/8e/ppuB/Q1jBzG1THGh6obU0Az
s8H/qjJRtvJsr3a7aS9+r6NNcJTaNdCahywPWz/Hebg6pclHAQgizbu1VDXOlHBuomrF1ea79GTV
ePTgz44T4C6ll4dSxPFqRBprCoGG9/y/Hw9sw3dRxHLWCBmjZMVv6fbfgueCkxsFwvcpeDw167kH
N7QxqB+tLHgqp1naBTmrQ5Z92q4swLs+lisvUh/CWO5GzCYHmiX5E/U9163sg1h1QhEsHt58K4V1
cxHciTuQsE8ofBji45eRyJHRlkLduyhzgnv1uhPFQCN3kenJc24kh+uKv+Gr9rYkvGPOxgCYBifg
Vea2u6m+34lwjSUfE1ZcxED/Vk6UHUjgFdVykkW5zjd/YJLg2vWyxelNm54tE4ZNVsO453EIFYwR
UJNPURQ2aq6KjQ+julSbsZwzjtX2GrVV972FKQUcuuLGGhJE8MOB1iuVpGXr6qKU6eIBgeU6eLjS
llU9NiFkBrI7DuZTIohZd1Bo42VUE+zmxRHAxQ5MC0anOkjhkd6iCqxED4QsP4VeNq8O0mGGQ7C5
AY8OtTjej8nT5IWqSA29lH5a1c5m9dn3fcziAjhBUpW2RWD8FnmnqMMzAhwxpaIRRNsxMBqV/BmK
wZ+y79FSVX+8lGw3TbG65bQIp5o7QirHX/vXM7K4iomFjAi/9DODT6mU9EIMjCVXrBSdxVQ08rY/
yl5V7smo+05EBu3mMKMQekeynDS0oxaICCn589+iSsTKv/6jwIqmER7Ofs5UTP9JKEHIxu/uKdtX
n1CP46MM4PMyOYfQ55Kz3p+NFN/QJBzgdxUw/CCqmRiGJ3moVR+sQKxmiJiyQftlEqJU4lkLNUfI
RcgSpoEv1F8Crpy3xXbvjrrZsoFVYuivlY+XbnfqWa+yGk2rBLU2Bf39wXn0iOIizSwz/XzQohU3
sPdNVt07hWjYwkf2fXfbSkCRcnJCaQwPv7RlMMbWum9diCZrhGhRmac+fk/gsBq8QiTCzMTm5lNv
WKhDf379EwrQ7UrtUjUrh3ZRBHQaUsdB63thVBk5KW5qOZz0zPh/7CxUf8XQr2JEKr8dpTI9XKMv
NHhT5z430kYTubv7AsgTZFJybR1WCeUmAnKdFtkv0RhMiUowmD2uN8SFcRIL3hnElnISehdn+LOT
dS9vN3EW1QjH0xZdM4Th1tmFg1tqlYpn+8xqBGYzZbbK2IoaVx3xH+Hz5tCjFEqFVfmVCQJElqKI
tb5cY2II7ESUbhP4bFIT8Xo+RX+ncr68WnMd6otCmM4y5vmHuhem9yUJd5m8p8NmNUj36YgpiqAw
g6fng6nU3dy7iWZvby4YJAwOFOV3slySRwd2rBFPa8fQieLHdMpRMsvVEQqZYm5u4X2iHtXKR1qD
o3JG7Vy3m18zOke8EEmtvHFyFlbYHnHFVWXKdgcJU/86gj2IQ5UBfchXT03sXW7VFZHER4g0o+xP
rU21BJw1kMhbrr9GqCmGv7TE+gUPTu9NsUpk8JanDvNk+ESuudOkzTiN7tyKvIz/M0Y7PdqbGZSI
5YLsg9uaYh3EZzzysfA7tfxC30AYXtEa2R7tuJyfMXvnCFYEcFCHF2nYjG7CIgmZ267XbLMQWAQb
GsEIzpLqWpK3Mbc9XcEvSkny+fvrd6Qv1tKnmkFOQ8r4nUYy/jnBPrlp7TC44Ohv7FBfaGs3eSc1
BNQSpIe13E3W3LgxACY2pfmeWCr/KaWiPKSUyKoQGwXWtTQ62tITAN2oy3JY25wljIJUyXwMcziK
m7lkbq3R89zOwPmQCuaCQxZuZ/NAQyUispifTZYSWX+2Zn4i3TjBmpD+FR6wNwX/FkulVHF59eqL
wxxlm8ECdPhUxXwEkAFArpQCGZYsT9n6i5w3uAmETyh688hrQQ3DY/j1VDy2FZ8qRAHqYlQ2A15I
AF+sZgJcL7YQ/LJKA6mtUfJjGNNzqAKuL748XQjFFgcf6kOznEcXVuWmcxMD2vLd1pUU36q/0p8K
i22+k+KN6/Qbm3PAoLdemvc1AEuZFzbUa+M6N+u5w9r2Ve1lSx0aPDWHzVrOzo7GOoY2bbU3Pt5v
EUX7ofqPrNIuDlb5WtOwKehM2LDjwvbjr6dEfli0WO4ZSnJpWbQrKEpgZBlSi75Fp0T1eal3YJYG
Uz84dufIGtCNJagbJKqtpeSQFMmvYjcJOnR4ZHFBUycLSqALLOlKeB5gPud4MQJxIFKYfOhCCa7E
MqZ1/0mo/4UM74WxDllf8OwEp3BGP77ZqbnJrkfqNUp6NgV1+mfq/oPfopBZhuobLECqFyPcfTxw
PXPcAoppgtuoqp8ProSFa5B5TiLI/FMhxcZGskgku0xJtKkByo3BRSAG/qxI4xkc8UljVz4gdx/D
+PyF8MBoLDJi2gAnCyNCINBLN6+43mRiu/+DlBZeOBTeNhI1kPbFDnF1TP2yteW1p8l1TLP+dIDr
Wt1yEeZRMk0FTzaHUQfQibD3g5HCujfbmYKh2As9xBiMGCNlTm9W1taMVXXxdPBAd40zSokmi2TI
oGXlBsElop/Nhk5/KT0KGHrA4fulxGKSfhtMbmcJcQ76jgaOigCMJUIqKsmY6vSK7Lp+sfgfce+3
RxcPCxUszj/1wLO1+OUhAsuGIj+YCcKH3nBILgn7D/0C48zHGv0pC/SEUNjQ2itBxv9iyv0iRv2p
NiEpZzkkMxbHfZp3wsFDxF5lUg9SOso4FhU43CIjzA9MXv2CCFJIhe+uqMmT6KnwfzSDPDIOgcuf
qIe+2Po26GxvuhfKKqflJMWVdrezBZL0Qr2CYUct5CVKE5fHMbaYF0BShN6Kj/KyEe3WFmRh8pZ4
4TmAdBWLKqqvh+oP/xuHk7Hdur8sKfPY5hiwFL2UmRmXT3jOvfq/VPSnGr9LZhx6sEKpeuUeryBo
awSL2xI378P3XVMsaIW+aTaWhQcYSso3RAyJ6aRwok+Qbg/LZFqDBJzaTfCGp0tav+i6tlYI7GFJ
g2qBVh/IEJsoB/4PMaaqD2eOhdYyDA5m1T1xFSD48ZEW+VVTxNalt+cBY36km5VBlViKSGz+y6LJ
2E5gUz5pnceCTLl5GpPDT8IpcRpDbNMkAd4i/NQveLnxT++5FPah9oGBAQFwrElL51nFJ1YaTakg
KSi6n9gb5KpbuY7Xbdd50amkLOE2o5tEMEt6U84aenYX1AOS2ed682j9XzF7932snd1/H/01wGNm
ZOlmEj9FSu/leBdHfIak4n9PDxAo5gjutv0PtrcwjT0+VR95LwgcKpXk50Eb9cX7FVMhGAZEvTGM
P1Pzaz5T6DZjZxv5QAt69DrDARnHJuX3dEK43BowNixKFjeMITqBstiQzBxvL4lPUeH+o4nUBw6c
4f+RVEUawLcUTytVo4NYyHIkV64I4ehljP3xIIDWfSes2aXYx+wF/wuxe2SvsdV6GphX0HlUfZ2B
lYs60gKzmkZlGP85Hc+ASY/2prPzkb7pF0leENH0+/Cc2rGxCRKBv20qTBPLn4sICIzidmkmOzZB
qai9AL4lskh99Qc7bDlPcyiYR5TwhH6SDGXe+zxw1pnwDrY2dzLSan7Hc9wYfp8COi076FYv3pmJ
l+dLEzkgjTiDEnPzLBH5532ou6hetbhn0z0t8v108XvCT+G2V4zsN4GoOUn7alTQoRvQuTZEO8o9
aOKvjcTPzS2Cd/kp5pXgXkKfVdY5fkQCTHrj5QEdL5Htnk3JYamkI9idDeS2bZV/vTIVUC4Btr8o
k6A01B3XudkyJkw2Bas51CVmbEKQYAiK3eurVaL/J3njaURD0CUDr3CUWxzr2DmFB467UQCCzWn6
VKP3apl3izxXHV5R/RMP+Y4G9JrDjFVRZe+3gk1WC73hccEdu5W8zUqypOQwYkG0wCZm5ZcmWZI6
q7CEfXTG33y8Ih4ack+kk+qHZh9bD9HfHUV+SpYkRyPW7en1L53jIItQtQ+0EOSwhU7bmoy3xJW8
Fnbvm5c2fsb++lhyyb8pumcNekezZ4flqbCPyAI5ev3q6t2IYOvQU7GlpR0NwzwKCQb2ldc53e7Q
/mIuWfPkBMOynWV5oKfjJ1qtzyBAaLRWxUok5ubO/M0zEacmOnlt0gs5xZknozZpWzJuz3qXf4RY
JlLIIXraWt4RyrAISOjuq8mJnmQ6IFic85HZPvSPUdgKVJFbTmM3anURgk4IDma1yh+8ezxOJ+vF
OrciCp0tqYDu64pyaKZLxdP8ENs0Jgf2aHTS6Y3BTBZjbPXzUVFnMT/Yke5AqGo9rQucLU7YglnS
9bLZlnkPKl5V8t1YznjxWGFtp20LELPMupPal7Jpk2acz0GSGRVjqdRMwX1rB/k7ETvZpooUC1sO
P88eQa5Im3midneWG0ucjLqWvXsvwJn2g48ClRGVVBfjfd2UE0MRrbREz+rMB1ZGRCgFrLaQqtnG
d3rNFoLGBwjbbkQrdm15fxblFgbSn45F4+caY1NqVog2P0eY/7crvOtE27yEFMJxBlydwaq/3Aqi
EsdbfZgTn6ngWGuCnT0JSx6qgqTUx4l2PA3CFM0hQ6YDuj/6bDNC/YS/1fMGxbB9hEPkp4DB4brk
VTx9A7a0jDwE6ZUDwQBDIi55aQhetVJPUHIBIC2mTjruhoW172WlV1qtG7OQ9q+5zX6Z3Tet7qmT
08cH+sp8g8mepFhRHF8W6TK+cYZ4bDOVwGtuhIFXsD2ZzLWr61IdE3/ZoLn4WovQzxFb75nwIvav
FDMI2HRHoyVUvzY2Spz9s/2W83W4idTAcMcAcDieUSeiXRITENTEF/jLHe6NTkbwKWxSimst72DS
sM+Hw6+vlHzBR+Km1YgTBjdiwyeDD3qTJCntdVdHX9Q/S39+cU6cyomLC+7lu/IqMZpKJUyHd4bV
mnYvrOo+6XDEMJVdJnXQfIF90uvVNHdcYcMTBlnmQbGoHZJ2izazhs3Hf1wKKviC6YNAMFm5S94h
6oG/4BBys5N3meXt8wNFoRn/7EyIZzsuYGCX4UOCw2CpTe5EvrExe73ml4asXVKmLM79lYJMveCU
xKh+mqBTHu6HDJy4rjaUsl9XwNOV8sAWLeGn0VpAQQoxjvVeDpUSJVbkbL9vSFMCiMSM5Kufqyim
ocbC1X6PT9sUQYACTxlGAHDA3gGhJ5wZwLpz3yfsAWNuFmI2LIOp7cNRJhiyrB7HS07CFMnDZwc5
MNGk6kRTA/rMHeF785L1f8AuvA9KFn0Iyx/8Y0FCv7OTfceKOiRzMiNKOWcioKS6FHvIA0qoPgzH
cC5EaKVZl9v94Om6cZlKnAQlMFALN3O97IZl6rNwFcwInbnc6iRFwOaFLByylvwAtoRukerE9yJL
WTlUvRNoJ9KZwzgCJna+A9sH8Ew8Sn1wA2UqKMMVZScDvqocOg9VqyWMR6qQYhehfju3DKnscjmX
QpmDAH4BkEL86yvxKR2VpZclGdexiEIY5gZsoLIUfGnkj4k1b3M+z9dKFhN/FNzyD0GHk+TMCNcG
zoXXCidcyl4SYM7QVHTDRibhqI9yB3XJeVNzsr+d+1xnqiT55Pgg2G3q4zsY2Fq62AsX+n7zBOPz
tETNbaoJK4TeJnFGwrwDp0fgQiPs8QYQQtPI6H2HCFbm1u048Id/m8TIzRApFUMvx7nJUEAjjDIn
HWySx3laeQQDWypxUgWxRAEvMISlqG4xdJB+hFC1cHpJWqtPRNzJVjU18syQhYWBLRlolHuMXVlV
PxkhYTo68mZGrPeB/wJbSxOHGkzORkt01AGOntGVHIalpYI4Ot59T9IYos72LRLNaOFTM9Zt02k4
WVdKOZICdOyh71oB7MY63QLOzP0knm15Pba8Z34RqXtc60FHVYNxnPXIOHWHswL0yFmV0FxYZKn3
rV6J+ZIHqmVyJ0uUNJGmbVTNA5zMETF1+erz/9LFmh6BVepvBKFufCoFmgRt3DfbOadYsa22iRPP
cGYV1Gsvorob/G/+3tPPPppTcmXDJx8YWoJ/ABaCad6zn4y4bEm6QA34hkuZGLkPkavCRa6LyNA9
pS8MsQm81wF3EEnA6AfDDTrM/K1WUF2aC4Se8rCM5Jq+vnjjfwELzGHdsgyWzUj/C8TwTlRWv1Yh
i/h4TA7H8Yo48EeR16ePA/ck/iCM74HeFAjNmc+uqX0Du59z2LIR0aejqrba3UN8nDVWIW8JDkLB
buZblEIIwQXmLZb9hGXVHcauDIdTVaYST6BCgvcwSjn4K0lRVS1weJ8IqjApzVDsUhwfn+WQ3rCw
DyEnxmvai9Zq9/M4gcKo8cJ3UTSRkvLiOPIn+hGk+tVjakq1hWQGhT+Y7BWhYXuJoo599elQDaCM
eOofdi2l5UOhZywxxqhGRHmQQP3nlHUNMXzir9YEOwd8Bh6YruTq0G3tW5QRB16BoaWS0dCPL3Fb
kwX1kOWCO1z8berT/WSomrusEPqUfm3L6L6zLffqLTuWmGUZgLcxCa4skBG/AE1TagkDxg95SYVV
eOaTVPx4gLgn0DiFEUIv2lQ/EqvzJ7WVgP2VX1LAc6gi6tTHoCHIrTkjFP+4cPDvLu4/0JnjnX1q
HFQWKIzgqBoIs6V+cTmJ1wCIGSvxTPYjZBbzqtHHz8YHxCijQWshmJ74rpvNfzjv9wexMSGCw/ox
oojrO4J48hqCCdyTEKybQBwAbVKCDKjt48tLC6nD/PkZnJ7u3SGv3tKpsaxxkwifrF1zmQTMARAa
tZqGDQyI9rZ3wZkqX7jrUc0d1n0hxItm1+Taf9EvgGrAXxmk/u4sgPnBSh2s5OJgYInXhKHOEKnM
KMjryTnZJ/2sr6Gb388lXvzzD/1ZbQl8dXEGIj15MXEJLPnz2dtBQc3syvHQ9VQM/m0PoEe5NkyP
7mV1OQxlTpgejxGn6kcz+qCY83Pe5OLWg116fM+sMtkRcH4l/jLAgHju5qqQLcIEGwxNFdat+ckh
WZAiJ+kNoX06m9ZqPJBjaWy236dchwDE5u2V7++wWleyb7whOy/aPAjJ38OuxoLMxPam1aHtYuWZ
cjSbgOr3xspC10UbojOM8atwvwingWfizsffqmWt8VR+ioPv2n9mlNPaUL7Q3zLfmNTIFkiQm1cK
f96RpRUU0Mth/8TidoRanLSxWydg7AM/3/R3ucVLsrKlNvD9sK32uq223l4Rs5+aDmnD/G/RdQkv
Fdl6ycyjBniNoq6SsP4zb3s1kKLVvGSBjhq1hASAP6H3Nm/qNQ34LG0U76N50Un0sRtDQ/WC8X8Z
SlvkqAUvTri94PrmyyxNvv5/heCZ3PB8a7SyYU2VRO2QoIJtXQJUe06ydNYbgYSxjGwrTje1PlMc
Y/p1OLVTeYi8w9qKbbxefyw/3wR0axmww2BWi510ahtLUi3X++6YOFPZpmmOfud9YSuLPaPvhDJQ
08Vx2DWyQqvu62t3YsCl1ugbE+NXhOH+CNice/GciUcF30O0kubQfCjFRf7PikvlVZrFhYUH1gQO
PUxM+bYR4cRzpUU6FwdY7ogcwcRp+F+TBEtjH+ZdPejaXB34dLvOQoq1aTyvmEyQTUv9UJwHDTpb
mOb5Odbj4AKiCwi8TVm/t+r+H/06T5K0PE+9U7p/s0tX1Zty3iaQdUVNQc7Mpb7Gl2cmH5Gxq1pe
sj4vE2N3PwBH6jD7hgJZmOezpZzwsBwVLYEXEdSetjxAocEqxHDLKyw+jcXug1gqpFoz8p+UteV5
jDBlKCsd+Pno5pyfvS4NTnBRtOdmGn1a+LRNDv64BQIqfM3/geTMUlcuoqXA8q5MjuOxeSYrXjIs
Kbb77vIATM/U7OP89kEaxVUeZS0pKuIySXYhNazGRnJZgRhCW+hagfa771cc7sRRfcRzxrtZfPLW
rAYO/HeZpF+t6gsCphIgqawsapEL5QBKMZ/XGGmVfywjgEtd9RbgDRndTgKROm4a3kDykRBD03xc
ymvJTT0Q4annKwEpb/UJ51xitfzC1lGBsxzhu4nKm0yrJM7Xi5KNpc2sQUAlgJielJWzLVOEuKts
/ZpWpJB/Y43Xn99fBs9TEWFRfPKx0UCOagpyfLECbWC8G6+fK7P6dLpDTFIgeLi0WsQdJqzbOhmC
WZJij2JL/70hm19vzdAnBSC+DVImhfQWh68P/krR1xUyMkzhWg4xAkobrqF+UCoe/HL1DIgdwtt1
4DVEyhUkgIWXwSQpeuapqlR9Jv7kj5zAFrHH70zCINjOhi8VuxILSAuslI7XCj5fx+WJ6+FTltQl
9PkGhLOVP9Tw4Kn+PiwVinJULLp+i1qGZ20R6ag9zElM4f2r1IJUMKgqniJqTa6n7OvJVB+uAfcx
Kbl4hwZsHj7l3jBgc+h5uQK5sEjg7TKUDd9wqDc2H1Xf1n7kS03jRJiRm3k5aOm0ZTjZ8FOkIgzP
OmzTMx3HJTmi37NTvXhlJHPbcAEtl7I8ekFhRS56YUIPA3OgKL/I4HU/PmJrK6dfVJAugK56/I0+
54lAQBcgcHqbyIisEkEP9M0pzGvbyIMk1W35UfsQyJmgwJB9Mr8dMta6DpRGHU9XjngQg6IvU6Uj
1ZDvjpN6F0sGLOzTkySXVPHf+dtKsd8gjOO9KH8AFugQIsw5XkbpgJ0/Wi3fOST9ELq7z4JtQob1
yLcFcngIx+gVq07cBphW5vHTVQ6wGJpoOte9mXms+7RJorrdCQTGPkNa3BlKqxqJ4vrrlHgIdAe+
T9GUSwfCHTfOgyxhCwysF+JEfkP3SKURgfCEQmGMEjmsDRDnpL+S0CeHFG5A2LFbPf5qsn+NyCve
TWJDXFJ0SJ7Jf3vuArCEpHAKcKtQ8H38CRDR5T2KVHzBQ+3+5XTgqw/gS/hg4ULZtOt2tyZ5xd5x
iSbgcySmaH/t7NHiUHK6JjxDYvFEL33TswS883xMV4gJUrxrLkqT5o/NV68gbUBjkmlrAPTPTw56
lxHXltnNCmtGuEaLYVdmaGRvV5uYU8e95OC4H43F2OJ+Klw/4z7zDpkAeYEK1AnZf26oT7pC8FtP
TRhtdqZMrfBaN230gk4IvlhC9Dq+ejNRjxcMFYYBRe2/EAlkog/DCf32vd+VV3I8DcHwpZNAwr44
+ssGiEVUcsiDW0QJZnK4KPsOJT/rz7UxBuPQZ4mwmNS3Xfe6YqG6Xqxgw8YDyD7NP4VNOb2Vp8qg
rcnjtiVUPtydlpkCWFg6jQkxD6ibeR/ejmEaZ3FRHq5rxJRY7Ub6EcvN0RXbIEM/C3yNBidw9bjP
2aXf20mwG8pnmLK0KuS4Usil4UfDjEQcd9tug0csDLiXWj/0wIASL5TmT4klQfInqk8UcYwQ3FvJ
lKD+gWsOC5hS6/nCcob8Pt8Hr2uYi+NiSwMtJ2KW/xuDMxDAbKssneKIVAIHUF2Smf9X2S4nJcta
yeahT9tcXTRkyeP2Haiq1qQ/wN17GiplmY0kZCKcMm0ZW+RCai/Mei0WPu8C/3dl6WHO+6FPhT+b
ry5A4g9ScLdTDsbnXA08rGs1WU9OHfOyXx7Z2I3qV8s/6q+nr2E5YAIJsW1kTBwke6NbTZhWBqLY
C3t2n0UrTpX7uL2maNCfI2myhQgFGB7yrEf5pCHN3Na3j/v2HWlnYZZE1HU1Wqre7BGgCguV0Ys6
N7PKBhpmGUWUqO+wYeD4IZP1PrI8boDBnJRPMeg/pFK0J4apNRHT0HmdFckGThIodXspHqmQNUmU
h8TF2vSgNIvPXQCZu6XJCWcrezVRAq2OzJ8c2d3cTGXsUTDC8SEpqXS8Q1dSo9Ra8SW+/jy7qRHx
E9TVXlVQGujKuireLlB5hxY58gmo/E8FkDJZpyrtxTf+zxOmNbcsacQBvbxigX5CKkPnejwzWPXa
mKuTzS9jnblDCCNuduBkEQo/rK/aNp9QklhMMPtr4bXIenL4mdPssPHfYUf17vCrA8lxCulE/b6p
QxNdUP5WAV7icmm1BmoEmQIc9ppTxC1nqCqbOjOg+MlD82QiG2NCKqZYdZLwsRBAG5UjTev5+uMM
Uv6P8ddJh1h56HlH5d3IG7QxY3cAtVWC5/NL2pHBthViewhAjDoxeHAX1rQzI+MmS06gyOraNNk9
4xKhhnHxNPF/5iP8ZQ6VUGpQyIY0imE2GfFq7z3KjdWh96YEJoNAtpaGzQTNklZeztq9jrAYA+F9
XjFNvsKNGTcag+QUiLwIe/D2sGcX9H99u0LMh5SMh7lyi5AZgUtyZYaWv2SVF5fb9XYWWZXJeSj4
0qDsNvPpzIUwPBTRifH104lI9mxwa7DlN6T+CDJd5fpuWJqOsWLaVz7vZDcQ6yEwEsWfRTIGgAWJ
YANAVNRrwbLvjnDzvD0XOoPSpXb98+5cmw/W4UbR+DL450sBWFqYfGFfUgU7L+0GY5ED2bSYwJb5
BJtWJKBdZ2WlipLNK2G9QnRzbT1eZENUVAIwLMFhfT6xMImHJ3kcLRFF3mRwt7dNE4CcBFjdeC/P
Bmgt+niTZeK6sF9+AJlZxx1IGvD8jqygcGfYlSLun7dY3Tq0qPv33PJOcKQ5/UYfCJCOR30fXgtX
DtLBxrdk0JCBzo/YM3UBv9f5GES952J+R/4eXvL7xoPdxyalTHxbPy/m8MFSUBFO/EXWbq+mFCNg
ptyqRqhIIh+ijblrX5lu36CbfhmTT7y/vnM0DuJG9F3ptckkZeptFa8am292Rc+KH5Jb1GhHG/ti
163HGs3RrUiqAbTmfoVZrOBbWy+f1YqPAcDzoz3/0cXizxue+1/I23rS0KQ3No1p/oIvoQ8506Yc
MNdUmYf5RS1OoI9+tPEajLWUAuWj1x91SZ4ExGonM9aEoAOyYi6lTY27FvulCmBNUwkbnLs6/bYm
hRIFRwEm8bOITX8PRv7jyTX13djE12aptTey5hEjgFI+rnVgNweDsakp11EQZR1s16naDfCIniLR
v0sUMvbgvCVWnGIPrMl5WhVZ5ByaTMtpE2p6RgfwCSnQHdaD2Ffd4+42iIRW0vdThAgOUOIbna9g
jadY3OMe1gnrYA7HnRvcCVuRGA/awMCp3G1MAJ1Vp9ejzZkc5jw7vwGNk1vA8RV/SVy48Jp0LKVR
3Fzduu3F+XYIWFmFI9OO8JnqzDBjlJTQtqn/33aztzdEQnm/NdXhq178SyJbCTXe+Fa9m3vhE+qw
7ZTSC/TilrGiytr0mhjxOqY8iJ6i+GIynTq1urJARJSOR+UFfDDJYcccU1lTNmLoPFay240g/qm0
+GcCzm/EK/tpKPanMpgMkI/upvyUhW2+dEZuWni6BWpIcPaUg6tanilNpuW8A/TFuXNIvCvKGbf/
WqxX5SgOmNaLvwyksMaP3OsLI/NULFULDD33ApFr35FIjqqE18LdtLqVFRyWE0j9B8IYiGq71QyJ
fwS5nCT10R3gXEmXR1508D7rkT0KA/srgeyjLK5CzapEna4oiu5Ymc4TrIOe+tYaiOvxdVlfIejY
A5cgILIiOqNz4rY8op5C4WvvzlKQZfhfI/gXNZuSguFIWGR+5R8fM4bicUreQfalDec1LYptRxVl
Le+rCxCdnjm6ibmz6AQKp6+8xCzoOqJ6dVaJfOjP9+90rcFrmVgGWJhwyut/5Yo3UkAKmnMDImy6
x2mdZT2ecP/2F74rjuJ8dqUzjrZVwG9Uz0udA2reMrJRgQ4Dvn5RUf3euYVcm3q4UPEtIBI2yvxE
Vf0Ycf1Y5cY+3HsWeC9YiwtxszMwn+8iilJEk+AAzGMSoT3+LMH2/cMI+D06STQ5EXAk+5T1OplK
Wo0zCZA8YeB2nX40VwhGk0METXMsjl3CKMauGePR8futjbf6CXBoG3w6nCYjdTkBITpW8CZA+E+m
10hNFy4uh7/2axzso+QWG3vG6UnRzfvgS6TDiJ8aY/OlaZdGnBDjNfivadsLrchRNwR/pGKd/NY/
GN9/vnU7FV6O7axkRY7H65jKevAzisvPu7XGN15wI7L813eWzz3Q+lIo7++kkiUCadq2rEPx6kYl
SIcqh+qKahXXD9uvYlsS5AJLr18dAa1fctIlOWAxou7c6tn3pUUO6xQnyFc7W2EJhAJurSxx4OIh
i7242vFCHqO18Cpd2ZxC/RVp6x8+6tqqLX0j6WU64weNUNgy8qyey6IYvthnexEYYESZiNZhRWdB
JCX7kZ0SredcS1kxqxDq4U9wghcdbmvBPNgv/BKNpeqwGWObx4LsS8OhON6dewHmrtXm/g4zb7LI
A1tWDLFlHkmzrhLdqU+oSYXiKI9KkYy7GzEr7+naa9BkQjMUbN1ZgmSUcQ//Olp7RtuD6DaCvt21
gWBYgAjCvkhjtzgz/sWoFs3sIS8uSnT0QYf29wAuQmq/riOiXBIM/vXU+4R0bmkELCuUmgCwWLed
Bk3AMvg63I+HfzhpRc5T+TDKlpRmFobK+99ojlTAvILX4WhJ7/sOtxsqn0FLwmq07gnTJYpNf5dw
Ocnb6uwCKu1is3G7Ou3rBTqTq0+pzcR+iIN2hSxnWuwvRPtx0H0M+sdmzVOFga1XZdjbwMLkGl7X
GKYdPY95rpLmlMfm5IcfstVdXkO/cx7g9nQTGA8wPVcKDhaXSyZuGBzUCjMgitQnv6n6FESFwU2L
diuYGRF4jcDsp+XgakScZVmMjeDu/i0ZQhhPQcKaTIVQOKwDL/mMBseWxUvld/bhocxX808ZRhAg
b2YFZrvwwVzs6i1iGaJtdLNctXqvWf66JLmHJn72VS5t4vWahY/6CjJLggSEceW/9+uIhQH91u/N
gwBTafhblmiIsfYRdt/6qJPG+LLsEMbQ71uniBp0Z44nCGUh6+wnADA49zgg0kq6E5DWtc7r5vZp
geHkAGJRDAhCO6tYX2klXiqUFe5KzHjtoScrOC/Mb3n6aMlQTKaMr9J5wWxuasqakhjyZNMp8VKN
j9mJhDyqz/D6fseYeF2+ZynWUrswBpw3VHRXo12aNAnb3GfGeUv9cRUmWcdkclV29zAmO5+rzVUE
KPY/E4R4EVcvZuNphlrlqu8JZ0vVSY/UuehcaGZK2eKvTSvItTJ8Ix32FBeX4/4ow4eFjwWVRCqU
u/2mX/5kz8k3f7hUO51ZFbUyjJ0hLZJczxgmD+nnnzGlgTXS1PWciFjw/5oxg7T6SRx+kx+/xWca
LBSGfAn4U4MmCU3UFxTGswvrNksBK1+I2YiOENY1NNlldUCAvXsoG6ONf1b6ll5kGd6k4iECYVSw
hFKc61IaS22+7tGfoDDgNtcPzpJFQ3eNDvNIrQIX8BcqaJNEd/Kmc0UuVcUafuE8p59Xx620kFzB
xmMjM2ly3agiiH7zQoHukVnsyFEnCYASoYpzAhnOswuL9rjVCthWrastTZegm0DUjNX/sDHJVKvk
nwKXFZfPhYWCm0sIYz2HOCjysR1qHLYWb4NdpCHrFEIuLbJl3SqHg23php577SYhtLf2v5XdzY7E
gfN5EfcTCZBYrmjCvXkTG/bdZ4jyGAExg4H2USMQBH8H5bDlaq9ELyTo96pG7ZOxwbve//Eqyg8c
dDCH+ovLSr7FgekA1fyOn2qnG/93mtjPgjHnF9NGa/k40emHf/s/pyXKdSMb3jhy2VK1CummUHRc
p4vL6njhEZkBfNJ1ENGjUcPEkCJN1dlqNG9bm9DHRtNGPApRV3Wyd27eZTVO3Z02Td6/gWKVvBOH
Jhpfw28LHGiXSE8cv7Cz0fzuaRczg4uWql05P9+5BHYGuQNJi5vYvqc9/J2iTWHaDS99wC2smet6
HAs/zgwaJqnepqUavAwz9rsjIi4LMub4I1EL2r8Nibai0Mf+mjfZlbmDNztC0KtDkRXxHmjHv151
lYGIeAdaeFoHANCTd3jJX+cr2r/Go//9/IlUAl0ljV6mN6e7foEnG9AkiRrHX8y5laVTFc8mFrQk
eK9cKVoWETDGC8BKzeMVgc2FMuirEl71wrQ4LxHElmI/HuBsIdXVCZ5qbeCJGrO3EsP6jKVeFShh
atnPX8xWGStfSHZmwvsrKMfG+nVcUgqJrw2sKt4PigYKA/yUI1tHEkVhmecAfCpD/DkeJYRoXSQC
TPngzqIHRChkpYBZ7ApMndxUZLe2My+Z70cBUwv9JVsqrTbyruIKyC1ZeIUHaxttYUu2OPZu3ZNK
jsDnpiLvnJTycXYeA4BOKL98vZcZ1iB8h/O9xDTKP9r0UIDE7GmxqYe/Kg1ND3LsYjWtErVJJ4E4
3ERBdyrt8nnzElECXyPylE4eba2HYiJZkX9+I+jsMYJxhDWMKZh46CwYYvkn/j4LHDF7qL90WYlk
+l012dbOMWpm/4smwWS8qzyb0weEyrP8s+7OtxT3N8OgVLOkhMuEWz/WdqrqrfJoJwGeZAPNS0HJ
upYTBSqsMs/MWA0d+6q1Jwo85gbOklYKA+cAMacEiFBtkwQEVGxzPsAAK1g25ERtUJMm+JFXZujN
Ow0c6/UF0FkkWMmJ5e3Qr0gm7fKCRidfo0wZdgPqtup8tDySy4sX+vK9Bl0OFoApfeKOPCwr2j0k
bg4afxnSSs8JIORqDN1feDB1HBu6UfTmyjHF4Uu2+eZnH3WTYXcOmZ1U8nld02cB1QJosXgL6bQn
PRe0vbSoAQVF4kvI8g9psdWaVasgAvLpz2lDE9pAWaDKjqPERHsegRH8QMg/EglAzVsfGbNRWSRi
9QtJWd2JPQblmv7J5Ypv1WPOkkcwNeGmCP75qMlylWafQNIY4i2Lc+WgzueWrklJfC4f8CfEawtj
hnJB4IZn2mlReZtsfdp3lilYxntXM5R8zKauizUYEpcpnHXl4KGe8EGIKIXMTIrnrvYoHPX/bwHP
sWIG21zxeG9Cu8NqQ3xnr1sYUgpw9kwuOA0ATyrC8fvo81apshO9srjoaqP4RW9Y9QdUNoI3xqZj
XJZ/dR0HjjAuCMGkYFbEAxrWKOjwQ/fbpywWWylzXDSp7Qr6xEsDLrIx5O7vCKGaOJoz1LY12Uwk
9ALGcNml2MCo5fjpTWBLtJFRVziUINXvimMuI2p6m3U2CJMQYtZM0QHykY4D86dCWKFcVG/ondEq
fMFJAVlDhAC9KxG/sAYNoxpETNTyd865e37l/a1xwqbY2DhQ/QKH568gGvyJo5xU57fLXW2I40gm
TadUroPICI5QoeZMhKWAnFM6JPvOktgq4XjSFl3mU3N+yHHUQQ93akHAwDT0F5x88kevRjPhnZSl
SriaDpF1zTDMhZv1ppiOA1YJBlFAgmPdiIzuvoKYhRNVTLoSFxUKrD3PvrUxKCKcdw0/2PcR+yc8
P1ajyBFXp9zt5z7T1Lul1jFWOTnzlwPqH+IN0oYgf7Xsdlyc5w+JvqAL3f/yHnxACGgkMLgirVih
f3C4aR1pLHgFIy6xBjvGpGlnEHyagXwVYM05fuXpiVGDK6wP6wqdZpQL5B5GzPxZAKOkHkHQGbFH
cEspBeQsdU0ESD2gGPVC0rfBRNlJNKwJ9SJmgz/ImudwxlrERHgdNAq9rjFLI7VPaipERuAp1SG3
cAiLEUoV8myDhLRH1f8pUUH17cWBxF0KT4kXW5JvjocIUjeirb7VMjwvEzkGHJ+ei4wbQeGjge+S
ztRNYFskqcLTWuG9puZGoTbG2QLjNLPkxSgBfizZlcsYT+ddkZ2sYWPdFY72PBorfYCxbQ4wwFW0
UuJi9W7/95c2/SsUoaeDcUvOfND31QhVap8n/bnqppp6WN8iF3lHdGBwoMwJq2Zh65cI0KXhXnIz
QhrMqcgM+A0osoqWMcso166OoluBwGsxJJnHVGEH095ePssi0NNR0YYVHb+HmHX+ON5ALjmCRvSS
7yermljh1/Uv4XL7PMXwGVp7q+zoUAGIjtnlZCajoj+Maagl1M8UFl9pc/+QsAnr032k8o8LC9+M
848SdqpmILSHIvsgxKqFk/ztFsTe430r3OesrmFJMEhn1OjBbJ26Y4ilIYtysQBSbwoarIA00ySI
kDcIzJOM2mRTPjQh/ghIP6KUHXsdGLnK2qraivt0zj7GavaCn+Qop4Vj+Xi8KQsarLTwqiNOfpPG
I3lZLbE6HH0bZUNGjz7pkGmdbECsh1dqZTv1ObR+LcOzcSjxykdR7sm6s8wC4Ztwzt4FoHIYw9k/
STlcHvCwpTTUJWCldi5M9tlRmBThpxzw5xw5xA1GIJ+sN/I79lcbAPibm59m8oBSs/UDJrsv26IK
Lxnh2MB3TcnLAYb3XOUjfsSPZwGgjTf5s6ol/bgHzt3R7I2/XE3UFlXoRNun/Cl1V0jSnWEnDjlI
iQOP7yRc96k5NeY/yTW3ZEVD8CdrsjadwHcjoqNmQWHepiUvJOvl2X9TM11gppr/SSRZVK19agOB
rNk2hBp3AzBrRHzb+jaAM0qDmAEojeUeMvAMpeMg1qBn1XdwsebhaYK6ap98IoT2eNVCyf1d4uJH
sbpHZsUPWtRe1KXKujraxsBqezkhhmvmkH0G6w7gp5NvLuZeRm6pLdd33V4WMmZuRHtIiAAz1xnZ
R1Rf97/O7z4TPWbo0P3oAEJVmIhh44IteB+AKTIX/pSH2ESffqd5iPqcW1RgzxZKataPP3TYOB1f
byBVqJJI6k7jwSCr/xAc9Eng0VU2xzVi7kcYMpQVcJTIE5ytAjBOBr264YoOy0U2Mli7zFgC56+5
2iZo+FIYlXPWvx5w9/H6DNBiiSWF7MV05XjOoXfPNXLvgs36bJhWfbqWSRCQJ/g6xsPhEjUNWP3k
l6W3bxa5jEU47NJbPkFR8BF0juqSuNaDfkNjvwfYZydL7AByRa3/oEi5UosBjIhAcGSdLUoGI0sQ
9jZ7YELINvXFZt429rnQ37gK8oUJ4d+HAMTbEIC3S0zPb1W7r37S3hC9LAbuOzAjuw1ReU0ydggZ
JFyHRNTCumg45IceLBDXySqeg6BDJE0UOPg2ca8qCgY1CiRPwaY63j3zNErD7KiWCCPDIUhlWPkt
glAhRstibIjjOiiMf5fTV7Ft2KqbxxPKT+lTRFhCNRABIudTF78SOmc+ddd+4KWGLxHDe1yJFM+V
+rvxK8Pn9AkwStkEaOAHrfzTGjc6OVXbc8hhqkDj6hAdgnDdEmlhv60HA15KEjvBgaC3QtHomXfh
+8hIp1ANBdP6eFJFmWp4KzMOB0t5fL5gGojD5SLyigvku8SpRudIKxm1xMKUavR8uc0qkxAzIDJM
In2+9Oqcyln76g5LKDbXb2hCOUyEeq2+UY8W980QH7GtRobZz1SHUZGeKJF2paKUI60otNDk38mn
WO2/C+pAcuLiFeZfP6PjO8hsE2YET3nYVwCh6pwu1sgrDV7rFWWWVRge3kIBLv4JTNnp53SJqCgq
iS/x3K2P82cyZ69MpNe+xECEl9kHqAaYqNhCcuGfeV4DbOM2V2lP5sU/rk6RCqwk99Fs9zhmuIk1
oNTy83CRIp9FLjxsgVAcQZ1xBLOrIwtxuUaWLOjdvx7tCA4av/yJZ0nNAYi7ia6tdB6vo6ijPT33
sWuOaz5Wtm0ChHAwTBsotGNpeXh49YiiE0nhaFYrgbUdsONswP+hP/vPBj6edIub2zTLhSWCTQZ9
MWOlo2bXKgSbydzZpqqBEgR9zoSOY5Rq1KYqxtJ8V8EkjoL1LHWdF55Lb3m3ivvw79QcriBZXXn9
w1/yepSBVRiEzP0ny/GiTBO6v+UDc5iEoaRDpqP6D5J+544GvPmVleoizvSdR1TvmO455D8/fYsP
Q/47170HBa7F9Wage4xlroE9HIOij0IRFJBFecurizX5TVMyYmMIZZbM53V5M/7/X26McWsMtKsx
EUHjvcgUJWrLMlHeVoSmxcl529GX1p9lIzjzDM4TKEvnr8S/wxf6dVzAWe42QB1zo8xWI0PD1ZF3
KwwEgxsscWLCv422As1RJYpjkewaUjQbZF8K8KsGdHXoKOph9RK8pXdffJ1iVY0qZs9PnXoFkzk4
i9yLFcQJNM5xjWRnT5athUxIpjF5mwUdTkUPkuNsZav8lE0gs/lZv1QtgADgBEVTuhseeRi+TZUU
6RzGBIFsOJumANJAzcRdsUBEZpNzkusOnjIahdhiWiEYp4HI4X30MV9wfcKDlNLhdfi3MhsPbPXM
x7n4WAnuGniABCtWkzdC1ReVgKFfEiwbdZEiTZ4sh8h5bYMid/z7zwy/vok+D8in3YRDQWIXDhLu
xdjHVRZS1QagD/nimuQ0C3UxPmRKSvWUV0TagnwfFE7cQ9zLUVyfa0HUZibIvZyXCb3CqD25idSn
RXmvvqVnzSLkSDymxut19WCmmwaOsrJMdEUfP9Ze2nffIRj82aoYaHnhE229AKFdAw9pMZlwYU48
3hf3L3f1w66RuZUqSDZsOHlmZbbpT/JUYJa/1l4uUCRV6s/p5J45+vfQV2ra0JU1EMROD53PyfCd
0920x6lBv6LMKX9eh714vUv4UihX7KGwslE0U2cT7pZDGNs8KTgMA6leDe8CESKZ5eusSXqv8ard
Vn2jCovcIvXAQTgHukU3BzMipzQLp0fyaLBG9EZEEEq0bMCT/7wZJYh6BRIAV1gwrJ4Wfq64ass4
npgDg4zMwOiLisI5Wo12/+jtC/k9Q2G68GYgiToJA7IPj0HJyoY8FL87BOjCJ/24haDx533GKtgP
cxlbgeITqld2S0Aq1G1+8Xk30hm7dppfem258J6Ka7ywVVxPsQqJi3LkiysocfxhGrakB8mIQPxM
Rmo8Nsb9pPMVYddf19HZTm1LyHJQ1nXzPrj9WvJSOJDT8FIL5av6JmP4QXKnK7JrPtXzIAQoqga1
YJ92snjo1pRmSFXbFDTeIaD4Hb6SOQNlsP+e85C+cZKzH1egG9yXoGhM9y9Qs2o+O2eO671vIpGI
v7A/EzWT7rgK7/vh+SoAHsliiOilZOIdnpVwmwqf3YmjsDxY8hWc+TdS/DH3MtqB+O1tylNSELD+
6i/J+b7121H7urzkEALnwPRZ0biZuK0dnlJmoCDP6rAT1LzEDJiWpyYKgRUBtr85U0ARjSaZOljR
4UHMedF4n85HhD1wRs3OTTm7lDlE/0ozJifjBkL77Oru7sDGBic23j6yIavzMfQ4pYcj8b7XVxWD
JRp5UNU/TSfm+ZQht2P8Zf0n/UcxdX0WHVr63re5wPdyOjO1afl95CQta9gIaw0oFY8rAOrlpAV7
1nyD/Q5KmVbslOo9x32342dq72r+fmo2iDeMwVA/0inxv+BBIHxx2Tac/D426zRAEkgIAk3DaPFT
fxN+16/SbptWzj34kjgTIlnba4UOUgkYWngwmzaa2DM8GGxV7ZcEGPD417cKE5I80RdgVp9+NJvw
4UxpD5YCOy5kIG0Syf+2zYi9RD3tuDlDPPsRxjQp+dXxMgKUKupMn/ZJvZwg5Q1Mhrvoc/75M2qu
UUG0Xn7ZZgO33x/T9aMVWECU/COMrwhgTvwE7dNP5ACpIAy//zsI+KxzY6u3n1bbxXaSXvKisXkw
1Y0swBSfPj2+jrW7E07SBe3mnSU8LqVOExuszu4dunVqmKtUn9u/CpCZhMzPXPmzR2fb2y4XSp41
STFr9ii8OeTmEkIg5fXV2fmPKMjBkq9K8vY0SVNnSq6eAXKs7akdy/q3rk9s4kxTpPE8k1StYXm0
C4zvrqpIRmIBAP4W0ga5eeba0+unYoUwnx8sraVLiyjAqRs0QY+YIa0fzcVmw2tpUhKWGAvu81wE
wV2ydwPEctFODfCrqOrNlpE7i2UnxCsbLwmWyiA4BDLyg8Rt548HBmeQTYbTV/J+Nm3VvxUfQycV
kM1tgSmyOTZz7Bdin0TBb955UXuZsHFoFiw6w2TteV0NiwhVTs8/PARu+FZyNWHDAQGSrwzc2B7q
92Rb32qCsqNy2xh+QXKdrG3CpiGB4gmZW5+9Oc1N7vXiHjW8o+xvNpB8q/pCw0/7RMiXV2nKi016
0RoT2jPecvPfj/VXvN8jkh+PPM+XRilsPvOl0qObUp+wBGHMGeeu1HDL5ZoJR8rUZQsFDTIY1QnS
Cg1+Z0Ylv946VzS05MWooVOAQX0ArepWHpHuPHL1HSUPMU3mcZKi8QTZ1oLBozO4sfOj5oVlbElQ
cxqkpZVYWP01nFy//uLPgtr4MulgS8zWBAwltZLi/Kqa7gboBVOacEaLM2oPys28v8xPN1vN/NKa
N7FVhQ9hhLeGgsJGpWpHp0lN1s+lAVHkUZsJjrbRb4ljLSx6YCqLZ6tRGBfT+kP5QUcUfN30PKqd
ztMlylka6hh2TsMC1lSv2BE+PFDQZojdjZNoPlxpCvMzJUS7smLMvqHN944bpQuATdsIsDiy3r48
Rn2NLkFhwmankIs1lo/G3gDZriSpSLTCRZeoJAR/BF9syw5lV4qqqiUMKsBTCnRpvE7VreOtucxb
YMehZxOnXEbnJ9neOxOy4Qe+96oMOY0wriB+phxCXqSAddMi7CWpAb1ufJhs1WSpKvrrbznU/1lC
GMiEwMv9kPLiMDKXVdNko0X88URCN9+4zyeeC80PCaDGv/LkCiYhSEafSkkcTu7SwH5WfjDPlpwE
AneIvFYHwP4WU/nDphRQlEN80lpt0m54yWbVf3ZmnqjYU3oyr4+JkjenCuOvFb92zZPjuX21srbx
x4yl6aBUZptLN1uuOpopPh+AItqCUdrKp+gajGy2gJvjLT6JBXLfH85WDFKsjxc3J4lLvNzkRt9h
iho/+7s8gQa3Nubf+k4X977K1LPvFaNM2OQCsKlUaNmZzPC9FGfmKlBwFMo7hYHiRUxuz4FswKMy
ZSZIWUQSvp6BTYFEVIQWU+L9DCoUxpwHXLpAmBdTKz5VVZBkpDbowuel1m+9gykkx4zDfOYYqecX
rdJMrSMUFSrkldqyqJx8wY5GC0CnDchc5EQZgvd9EQlQGSY5QW6DgiI2WVRNi9JCNMPxWVnFzHOG
oXStJOMAt7rQZ+pTO5cVGxPfG6Kt8DaMsbPxb9jX/Uq8vDlSzIk9BAtxTfXLIUKsCwpsx6vFXw8T
a2D/SuHWiXY7jUrGi73h+OWWrZRbU4IPY/Qomab9i2pIi2vrpGBmeWtrFQXuDqZTfvd0KnGLsmAq
kXnDFNpkehyToodw7zNgqd64JkaoRv+CRBNGgPHkChX6D7oznlp5qEP0gp9KtDQmznIV3whXq1W0
5nsLN+n4uLkWC79EGEqpViZ1oNyndZD0l84tLOp9Fc5ZEe5Sp7DV3BD36q5QGhk0kZ+e7GFy22uC
gsjNYfewoGvVTzhASZ3epNBiPICSJvzO4EK6jnXagWqAPsYOv7Vr+HWvTIpz7FJddtOc3Td0cxPO
m4OLmskUfPl1kCHCr5dHr9qIFb9++IFjPN67eX0GihbqJ1JjtDdBwhfz4LULG39Ub7mYVnPM7qsy
Awwtg8z+CLOb5oVd9MiSHab0cPMptmRhFdprXUmU0w2UdaJWlIqKg+9wXzEUaZeKPkKVp9X4uzZQ
tRrIuaS5hZB/Z5FreGT6CkAMrHT4GxSE4dodPNl8gVX8xpaJVy3/nH4JEGMzeKWuMufAYw6VOgiO
4W6hF4Q/DQ5dObIEVwatUGssx4e+rLzBOn2JKOzfG3AKz1Jsv6VHrxWjeL7+SDGIfkyBp9QwkUdU
c4Rof+5aKo/3N+l4KlGyENUsRKi9KMoTWfHq2AA04wLa2HPb9nG8n3JcP/M7mjdifyedUHBlFES+
1PjOefhYybHJcPej0zgt7Kbo0FuDeYLFko4RGhrz/dHU9bpNwsdNt3lhtrQd5oZ7n9PnllowbkZu
aoNQz+t+ETvgUEvF2OGvXI9jzxiQK24ObqUp4S2vilp00Mj90ANDLtX6JBbPpPH+ZetoNrbYPtZo
e7DFab4UoI1qrqB8jIx89fbMutjay4Bq/XfrhHKWhlP6iOpqwPL8L9CElopLhwyq2kfDy/BRIge2
jU18C6BAIiq0a4qahNHei3LmHYet4//CHvLyILjxON0MvuGtx+OxbYAmEVpYJJCk/hAXxy8NecTA
eTIiuuXdBv091jW5wARRRjpesYrDzU7VjW8atUy332p3NBedwxZMFpm5XR5UFRLLrqVQ1+bzTPM1
lLkMHOuGwS0JMqVhKb5ia9Mrruk0IR3Cqav4ZVC1T8m4H7NC47Y2isZXi0V7JxGkG30M6EKYM88e
N6MPaIFX/8c1sMhVCU/nhz0DTJq9Mry+Y0fTajhWrQZ684kAPe9QqMC4fFtH2YIoCSbmFzVnglKK
g2FlNof16iuyb5D8Sg7AbpaEH244XG3+eh04/csuA6RL1XMELb3xXlT3Iz0gFT6oYteveem2rl+q
wD9TNTcgyE2aSJNwyGMrWEhbWWU6j3vDt0ay8X4GSWGKP6DrrkY4FJWM8n33ERkqDEOHEBOI7xmg
bxgrOXwFc+dvUXyFkCMQQXW85fSaHx4nhJVT8RAybgOolzbSBzhYz5gANpHruQakRhKgwiZ0PQAx
szq0pFQIObVQc3VJLp6OaGNC1rnW76tpIz0ivXhpBxIlXfYnAlC8N3h10btDuBwb0hO7c7Azixyj
0dulzoC4Io2H+OgReASu7nTLGawBUKMY8C67/JSAFjQc+5PtKHSzvcktUoDKntiVBtfNOvDHD10w
a5oKE/AtEsxXP1jIMCNG983+0qjJ5w7M1TbMTXZveVskzSXC1BoLnaKNwYjzpka3+Tw4VeCSOOG2
oJIgXkgE6WU3aXP23Lu+qBzeGLJU/RZlFME6PPegVWXTuQiXW53CJjVz4XRf1XHpR2n0iawfcfWu
dsR9dvmNhotItEfIqXbu2cZXOTuxAoKlNUVk9USB9jJn57Boxd/GBVZS9v8NwgzmngJ/VPlAcQ4+
0A+Hoc4kqjThwGOzHqGSmUuQXMlfYFHyiH0zzlH5ezMIh9pKNKmlhKBBxkfL99aXw2fYBu6qoV4C
3KazlKsZ/dxyq2lWujpo+enW8d02932rEhnVwvEwVCdcNNVnHnrldxU4xCJ10nUDo1qS6JfNExnV
VUCE6BbJ8wt1dQz4dFwTbGnNrYAPwVQ7NK/6CrQAw5s6yj9tXRWcZCH2R1cBmrpJfrcL4kk9QEbv
kHxDIjs+NnRA3wDIM5Q0nmRlfeTR/hXmOM4eSsEE82Kz+dXMYtDDaAzTAkgqL2clrlQrzAN4K36D
tXih8TUl7+2Bed4xRywjmeB89cDU0ggHnvwyzLR0OW2lTWjR2cpWOgMfAxmNLHrwgaZYXXEOFjJm
Q9tnSDFPlaKUsrSvFlW0OHBcWGgUZbwxym1F4vbrUvmIzKtbakdQhs0GokCyDogr3CXhtKy8LWI8
zr7XXe/dPmEdZpvZwksKmbGWBEunVdUOy5mx+tzsoUuaOUJE2ddncoDnMu00ltk1e4jzPCyFQ/sc
4aPY/eLT/z7X31UXgbwYXw8HoIgYaO8WVC03wZoQht6q6noDYggqwp7EbeH1MaAIRReddPdQY9m4
kqcZ6kgwx9jmL0FmIaE7mF725c6usG9CfAGM8UcGE1NiWEtokz0c5mBzBgLBoE0FSxq+CLLw16O/
GiSFeXuAwm9HJyzbWZCO9CaT9Rhf2fZyvz1El8o3ev9aT6L8uBYoXR+EsU2IrhRCdY/beMvV/Shk
7m1WoyaOWCGLBkNHeN5m31y1Nufe8qCfnx7ZyGH6Xt1Zz8bQJFHc+XB7N0cVE3IamGIRJkPkDuzL
PbJNPo2UXnYfAI1KF//Z8wd0El3OXLqJPaCxIafebI5DbSutwvthdFHFvLULEqjVVj9Yy0DtTJ+K
e8fwJNJ2SSwhldo+2xrs1X9TQX16RxJdE6aKNMmKHRebMg1guQ+F0VITsjOfY9NQKZKkQLMRbuLS
0L7qxBYeqSIC0YuXhP6Zfb3ocs5pJ+G8o+53khv2j0TpZ/anNQ5xQo3D2WU5ILi/MR76TWmuXdQg
tBfyionvkmejfhhLaALPl6Ct+vjsofke9j7rKowG6yUonHjzqf0GZk/GhnXG58W8/nZaw4Dm62m1
di/91DMlcaGmFDE0tWwZeyZjarvvrmI++0j+yBwxvG89Bl0Br6n6EU5HLJliSfHChZUPAqt+Yep7
Z+13c9w2GG5jx5Dvd8oLdvwIrwHqOHJcjj2vc4BwYaA5sGfuJDmvFG3rl+QqYO7TGR3nPLbUcb6d
uCkTcsalrjyVhgZlA/om+FA3NeWIEArz8YMcAJ5KsgekfOVIVPjaLfXvbxNRgqhoyKw9eUXgugks
sC0VBOaeXDRdJP86t3eZcDyZ5+UDbOL6M6w5onkUyPOpjP/3t3bqslnY3ch/yTh4usWiE26hNtcp
c3P76aUGtug/4tAiSd6IJWwt8NK19BHF4NKaHzofpRCPPQKNLGgBzgleNzF3RGio9lwe03oYB56O
0Udek5Ipen1Xyc4YFhAIrCgj+W048QDTsq2U5mVzW+EBAV1rt37E9bnXAdpzgmEdQQK7j3NjhBoe
565Vguq6GFAbGKDJKWwKBnLPzQCbuD1Oh9r1ZG/BMgu91Ud6aIPQKWWpn0wL4prjoqNdFGWm3DeI
CfKJeFo8c55gxTcDc7USP8ArBQNbR8MFWkgF2uB3QIz6quZdRZiuwBL0/dAPStxT7hZbdwYmMuLh
5Zyiyuk66tS6/TQVaicOkbLGWd2w7w+Yp1BwA9dpaapaaIETewWluCFFMU38k95ZGzikZG4K6jMw
cLdxiheIuf7iODwskZEijWRhZp5VZKCGl1btz3SWL7njk6KgMqck2ZFIwy6zlpcRFxCyf78CtXpL
pw/NfW+64JX9MeoBhX1wsaQadFm9iEf1Tv+1U7RpdPq/dFLiHXfD4UWMGw8zcxFiaQ12RQp3Y6Cb
AvlM9Y1Ad2A7acGzPW4bQf6KiMml1avZw2iz5GSpKBHyzr8j+kaeiym4BxVlX1fK5IWFTQqYc0rd
/jw0epDOv4hQt7wJaJ0BukntvD1Fp9wKF50VFsbkbyAx2skSlJCGBKXPcm1RP25B0DvZz0+bQ2TX
jhhcoy/gQQwdnpvop9Zro7aXNg1IoQqr4HjQgN8GvOiealPTVspBFRqCuYhS0kJ9uU/lxVxfLCiM
3g6dTS1LgE0d7S9uzEMe1tXN4qVigGn2Mi0MIsInNOque1HA8KcfJG+ShKNebPT8GtVHUHOCDYiH
hWQEC/LSi6dliCx18OT7ShBo54q0hoII0FanHsizxvPsgfMgxEl7v+Ps5i4hmfysaNpdcc+OYIVX
7XT0evItsYQ0J5kP5l8Aqa4tabO30vmZP80+nZ/PMFHrEys1rhnyRnvSjfTQ0z1gGTga5JvSnDuR
RDsENU3KC8AJvxU0nOnwQ5pOaybp2NXNlGYAnv7A3DG2xl7284sA+TyA+RL1/bDcez+Gjx2+YPQ3
kPVIZj1EPLYrwxj8Ey8zxkatJKM1wNUYyezUZ3wO2BUGfkQjihjcT7a9cBGYPgi0ElbEoUuJCGaN
QWqjVJRBO1bykasCyq4Zg6PhHjjWuIU0RqLrpue+VFYpUNunZcDvFfSix5JXbynfsEuvqD8n6cc0
BS6bbr7miag7rR6YMrmaorwk9ykUR3Z5zLwHPrhzsdg2yQzag3vAxqrcD3a1kuvJ5RwVe72soMUz
K03KkwPDZLSy9TxY3bn4tyDBZH86J2c+0fbZNJeCiTkU1aPalzH155ft0q/hFMv8Xnk+JTcHSH4P
dnQcThL/TjvlRRwi1A+hG3mLGyxwBXrJuFvoAN7jyUXfoDMzc7nnliwcMmMNbnntO20J6i3PNegx
iF9odULoMPnT3Ktc74fxEkhQQBpW+4R0twhpXfmbb/ErMT1iMRzoVJUiKKEZT68FndffjwhxIeGy
WdyyNyKDuFbALfPGD3W5tQPm7a5cHBy4yc6OuOuns9odHErrVzQA9cV/r7T/5k0LSTbSjJZQ0qsc
8S4iAYnueRQHuJpYJVB8+a/jdGgETvGg4SVf+tK1yLb3YthPdFHDnpbM7kv4KnwyBEeKC1elwt8/
K4/++QNgL81kimYmFIpR3HCf2EZUJEjVpOMDW59yO69sPYa5zixW6ho7Cuk3MnDiFdpzqBGVS7Mh
Q/sgGOaDfa7koigaQm2/dTTuT1MPTk2kH7PdyaN6o3/VhPt5PGuK+PlieO1mDIwoNMYyqhosNd71
tvcsAW4Ffc6tnxJZNZOvVI7IJXebK8ym/JATaH/2Dhaa/MY1LKF+pF9mV1iysrOJSPECE5zMgtcv
pcrLG2mHyxGkGcLeqFBIudcKCiG49jMkD72QQT6hbl8s45isLE5OXEBKviZ5v7d2ok5dnIBZQbHf
3+ziAblshPaBbl9bf1/fAb2+Fef0h8zCQV9REXcIPx21B9ayeBBk7dfeBttQm0vsma7+23cjOuPw
B79J0rkmxUBnO9jnaOaWiimHu4L1U/0Wkzhr7IcI/AaYPRmfHS9KuFOldXdlt0l8wVOs4MhJl8nG
WUwovDpXp0zozNHQnXnEK9uz3FWc2jpXYvTwtQJ4R8iPeQTu7iJePxVY0XNTvtRbae8V5z0hQmnm
X8rHuR8eqA7l1OV1c0gFGQ8kxbs7ed6+Is2yjX/wm88si9TCNKXglOnVg9P+kwD2X82WUTeAZYur
/AWciPDCeMjB9j3ZwtOuX7MzITKKpuo2kmVdpRh1OCnRjEaZfp5iEZ4Lt8I9yUh3gkWieKhwKd2Z
PHn+Ex8rOiWbVqykUmyFLRlcRagOwhz+OBiYEmF5uEBpcATYd6DZPHw6dmdByko9qNPXj/cf2R1Q
fVSooHAp/sRcGAQdJBbqFg5S8aJjagJE1wMSkbbRiIiWyQtzUjsqEV6I/UusWnAE+bzUsNqAH4J9
m/+3UTi63k3zaOas15DYFFOOL8sJF8p6i5dX2IWfVEO5tHlTV7sqScrHOf5kRFg3AhrH6Kv0QSwb
2+Vw21i5y+9cKTRoF0WS8Awgm5H4ILXHpncKkoMw5oVqL9rQzcGMQFbpf/IkybyCND9xpiS9yq4H
Rhn+o2yn8QLSXi135l7GRgOdinUoZR/xh7cPYD7T78Z4zlsl3fssRi2tuvlB+6Z90nGgoYcbl6Uw
j5+XOn7c08V42MaN1fhIZLml+pqQA757D+hDd6YKZZP0TCAc/E22Z/fEmMY+194Y5NL048R/3ziH
JtVS1olcZynjUJz5s5/TDIX+iY/e1KMtRic3Lp/cvJjf0DM6IvKhDeu2t0yVDZnvzQk4MLO6JnQP
bWwaJ4m4ciZGmN6lnPk1nO9JH+eDF9/5R7hmKZPc2OaVXPYalDgBJLyNlIAeJe75woxBo6vO4Y8l
ueJXLQ0Fu/khBrB1s77V7RuIh2aNWaeQE5fc3jnxZa8WDH9zrJjQiLi+KkSj1R7og90wmU0kmIbC
jj0PuxRYvXCJdsCBvAZTetFYaF7hLif0aUPpgZbMuq2eoZTow6XfLNCMdZxqbMaY1hKAJLXW4NQW
RVrbnjhcx6OcZZ0UXX2yrh0bApsU8QVDYTGBRwFd6CLuRPHRE81PRNJKCmLt6kDNLYVOF/zVdMs9
Q0ESEXuCTLn3R1U1KxjhUEeUAvjWDcLS3pYt8eyFaMBylxeFDP3vG0P1CQXeMtHrmrdsh6CVD/bc
fX1wcDWk4FXAkx+ba2D3MuJWThgZioBUpIvqQIOzWB9mZ3I+JOFcfCeR1ZyjseGwa5vxiWSdOTLy
asAhcqjDO3rsRtCcR8nQn0HedOdU8/wgZdIREYyR2fhUNPN7WFL/94PiydwF/B97k3/SVW1yzyIN
KQ9yMyWPeDNOCM/DIiXCYqSPK2mwKfIEcDo827efB0NkPBFiG7r4/qUWzXJxV1FeSlSzByCQwUIH
htOHCigF3NrM8+mukmFXFZBVN6693+O07Bmtep5pyDYkiAWgbrocg9k/sA5p1sCZVE4KZKi69vD5
4/qghnxHtOO9KBNTP3osrYExQNmJ0cK67pC/WHQlnFb9/FMWOJjQHwLHWHlr+Ik6WRI478N15Neh
jl79voru5+5Dpfh8HRbhDXidu6m3sHB2nOEssvmYNpZUTaf571WQeDIN9T68yqG9tbqwGSZLfS69
O3TTNdwOEdne0VjoGTCSPtQL49IhySrwo+k//bozgxHzHnTsoOrCoOaETkHVljbdcD91GzOKIGoX
dcstTWtUe1NbBnXcAh5pkCWsSGUFUQhxnGWywPG862BQgzu+kiZE7Lg4iltfQx4n8qhWIyN1mjf/
gIfbYBlGRZaUN+S2E02cjP4f+ICqbl+lMCQ9Fo8zuBYniFg4WThK4jMNH7swI9hPD3qhyuAThN5F
wmwAcrlSKBuvJjR1GzXZREwHy7PCFQKpdgjDxvzx6DHXWglQx+sPZo0e80gTsDDBhUFJYSc3Se+d
pmWsRKtxLcsEF/a8u7SVhF+sLUrRZypm7ueYg1jgG8dOWQBRMh95pm/BGvCRc4+2r/1KM7MX8jjj
4/U81PjdguSbkAPHsXZsgykgJKDndsOy8DbscLMWpHvSI7khTxtzS/9YDIdJ6tBlKGciQILRtIZ5
thpdbamorWEm8zs59jmwiiVfHSR6ZkT6Asswm9Gafll9M0Rxcu0KN6sKrCXft8PYwGOX9P86EIKl
hi4jWSKJl1WYELdPKWiIEuKLHmPMBjvd2Nlg1GeTni8O7i7dEWD9LoVBHTiOK6oSXAqBxExRdIvc
yD60H26nvy5/7l0rePQQnBZ2Z10zk72KP9TyFl474xDQhtjT0GK9CPKcmdUuaWJXKCWJcMt62GNl
coINvnPWm2fai08yCQJRlcCzNMUZT8dkH3k8JYbLA/IcEtuWjdG8eMV0lLj15OnkXJTw7mXkVEW7
T0QyBwA37hUrLe2k2SjL2A7Ct15soIXpjFb3h4N10qpkB9DIHA+JkH1aohBbFzKE53wZHpRQ3Uar
uXD2TemDFJU7L2yVdgeiGAwtEHbPmZBkPI6o/+dtnNvLn4Y9tHRHFEyPHATaY8EZCyINb63fNfhd
SIUh3I0MP8yjcxF1P40GVsMsdpgyro8B0bfiSFF7BMBQidpilUju1HIlS4KAuEZkqrm5Rwlb+fXh
SIeIWBUgNcleoZENfLtoJeDnn0xIM8NNPYZ1+EB+cEfw+9z+h9n4v7sA21l0DQDpbbD5pZfwCwbF
USUawcNTL+D58hYPPJx3+yapUpkGbsNOz5psvwDceB2Lq5q6AEdj8t/hi8KOLyMdVLCCg+tbiTjb
In89nMEhAJZ0HhyyPwF69AORRFYRHbjMpJ5fo4yEQKbAFaW0rhmJQiHnxkepKspnZz3v25KsdDzq
Co7OxDnaq20/Iy8I3OV+dzbZNvp845lh7Po5WfM/y72OlAWtnAQF/rorfXBUu9S/IwkYau04thMn
bUdnM6/NexMeMK8wdMAXOayhIXZL2SMkD4UjFk3JHu61pysUnP55wC2FgRXCKy4/REMm4+6Zu8ws
QoopKFc88eJLfOC8oiH6HtsjXhsAInrkqYzkFlDPirQqCqbebA2LCzToIDTx2n6TEbL/QqpJzSFL
LGfabz/8kNroAw7+ndc82nHILMhagvYW8bysWwO1xDvmtf/NU4RKSWEd1haB9aNS7JKwIfptDb3A
SaGhvtwrGEDLRe3vT/1enrfUlH6EZ4Ws/MyS8qqTyC8kx4AG+c8sr59rSrgxocXOdB0aeCAHiByc
EmsDpTtWxs7dVaiut/iSAce9wjENjsa6tw/YZqwYUUAiGbI+qKmJ2WjzooyOq4AqFEL9zF4Pm/xe
iRyVVhhM/vH/6AA6KgCZ8fHusUrDK9+3dkJ/hPFUHAyNqYyK8lYCY5VgYJqfk3QD7LatdBEDEUPF
h2eUiUO5mfr3qyT24uWCItCsNEJBXEj3EVxB9NVYT0UrPkqiaQreEbIbcB/1h0VcVE9q6TSXEEBA
OJ4eY9kErLns5XOJbryqPwIRr2vkS9+n0kI64LGkJtRi529NIMoGLVLNsafjjS/ZGMuKpmOpVYVk
/c6KM9Ud7VtMAUqzZg2/i6XO+2TiryLl5KitilU0O8S6zNFwM4L0q8N4+lZahdQ3ViaJietWg2uk
TNdL+YSeZ6VZ1jPulC9sBMAXyutMMmx2I/qjOvteaSSX4TBnevFuJt/GA9MNZQbpO8fNP0Eg43Cx
H8rXYzj4RTeRBTufiwEptzD1Dn5Qi6n4dZQZBzvV2W5F/G4e6WLR03xwLtaCKxMOr9sp6NahZS/x
Wvyu4SyjZ2vKYvyCLcYJU4yTituxzilLSAs+wQLOi/T/ZZ5U+xjKkRdzmT+u8C9qXx5ih42YFlTW
6kBIqR/6RTn3Chd/Wod8wttyO2P5V6CSlTZhaJ2SiqbuEOPT0Kks6J0W6RjBbmE6BjUODdULLxGT
ODW1X6x3Bl0JAOJeA1Xo10TVoYnRL/0dW+6uS9s6Qx60VbOngwZ22CK99fPZw9qUAdO20I+w/bN+
LsCDmjyJfC2vuiojFxpXj0fIGdQvCbyt0jLSFYGeNDKI+f8LeqQeQC8W548jE7+IwA/CMmUMKJRv
iOTqaSOMcTX9NL8ZQZIRFdTnQnk8RerergX4jB657vBSysoi/eTKx5Q89Vo8pU00+JCbf/FvWPYJ
VTFcZ0xObVv9LMEMC2LpOQyRZlbkYMcP9fm4uOn1RPeAXUFgvgFvZSlqRrBc806Ta2ivyAsK1yEE
Z8pWyp/YNn73wmkIC/jw6ecxl1MBPccfI6p7g6ovFG/lS8T+Wi8TmS99L2ezJv2sHZR3emnNXH1R
uLPxlIQ59XuhAEF7v22QBU2dLT57nKwgmhzPiPvQXPAQoW7httH9Y0cfhQ2nJMZ7aaTfPWKiRMDf
y0x5wBBEnSbbAfzAZSFtJ5Mzi+UwBpC5PYrb/9ypBVFXuAfH0vugOamtWjn4ubZRRXRXmbM/4F1T
41zxM0ruVczZul+agS2yjz6ElMmqZiqGYsD5UR7PdSq22wE0VCgXb1ueUrTHzl8EDvJL3RFacTWH
Wnt/mdFpNEbxQsQr75lYCickG+WPleM6wMvM5C3Ne1g90gRP7S1QZ8c4lWzhRtSljMcQOtxUg01e
d9whU+oD2DctPL+pxCQD9Fk6SWX1p7LJG3k6zKFP3lSjxqi1CJ55OKTiYPedhE0Co2uw9WAKONE+
VpWVrsv8S1fuR9/t069RCjsmc9gyl+ztpppMmlK/Q1gSQ4NM7euusBCv8gQF+/dlMcHzwljxg3rr
gjQwxI0e/o599izsHgmFnxKWNq78wMNYAnOV5qge7Y1gfFVd9OMkf6aAauOnu3d6ipfW175Qx29l
MCsBCHbMushBSQQCJhwrbrU9y1jZY+qESYrG5bSXYuZWb9kEylrcdKXKG3aZjjXnjQS025SfY9Rr
HtMYazEoKkfupHKWGdB+gP5zAr6UAFCs7sfb7Zv/LrMCYk+R5cBwwzTiYNJUn+cgwUolmww3fIXF
B/vBuWVC4jOwUeMwaYRTLIHx8PtSXG+Yz/jWyW/fjTUp5bYZVaedizQ8tRsUoQUq3FHOR64iY3zU
3s45+GakjhsvMGTsmGXCZennzjtcPxXl7J1X0ZSdKw1njwv6RUpPQqbzjPl2Mvfk4TZaiZL2KtlS
kDkoOmyj8zfhHb/2cwM3kOfzaxo1dVicBkxnbW5pb/pMMSYmSRrPhTtt4byMc1lg+TTUTu/ZTyDU
JO53GZ/cXlc+hC7zjcF0k61tqbvwVqagf9Vpr6gynG+fm8jjPSQKR+9cmURm3l6OlTVrrrG+8T/r
UVMRPP36MVQYHLqTNZWQplstdSxCUgy/zHyExUryubj7jp2A+8T4KeJ/x6rajzDltYw3pMfUy6GA
CFkZ42QUTsLrMmVovat1j3ffUbiKrhmYzFOFZKqklXx+UmwGcgqLEafHBBBNl05OOZGxj/cdMnVp
V2lIIv2QME/+r27jqp1piZLck39G77glETU102771zwEyO5z8ZZgZRPhbjK48sNkt6YkoYhp7ita
6M8WzKb9xmsoLZPodrXWS9rbV34wUwPCOuo7IIKx8nBxcxx19XMt3ET2tbCWI1irdYB+t3s7nab5
R9qW34bJVC+/90x0wDcU9E5koG7uTXDDko8F/CttXVUIhMcUu6g1RMIceuuMK88PwVIV7lfPDdb6
+Eh3P6cOhTv8iREgWz1cDvbZcPASWqIjZoM49d0UjhPaKLy+FctlA88jyn5v4O+KL8dueaQCX5cY
UxLnWEUMvK6x92f3FZxsThSvZInzeOXx+WS4NmzgPqb2UUp7PyfdNlRSGFbKZNAUEl4sHxY9bo4I
7hKqVH0wCc4GcUBLQH/CLCoiZzNVCjBsZJVbeA6W/iuvi5C5H5zQaGq9tl7vlYeuFgHW7VRIvc1Y
PT6gT5qL1JrRmsgxncUp2LzKcTOBQD3YdtT9ivA5x6PcUV0I/CVB8bZY+dFlXisjUBD1A0oh2Pq1
04F8WxfqAX1fgvoUy6FjSCHMfaMcP+P/G46qb38MadiI3e4iExi2H6MBVQWr67qLdFX4w+2gfjK+
rbP7uKAf1csMudpBhCLPzmEdnwkROiXeNMOTkW+foTeoSe6XhuPWsqdDSb2d+lWMOpx6g8XkkMvv
FM2E9128m4qr8C5ATdwIxUGgnnvVLqUWNKvDc4s4yPRXCiyatsEEIg1YCGewrJ23TryuKIqOjMGy
/bLu07kwG6YfWQP7VzKNZ1ElpcHtOdOTOj1rL/Cd6dzlRJVSepZRUgj8lBnbSO2SKJAanko1SEqP
PFTxun47t/CBq6rrB/W+UhstxFq3PBgVVQc/1V0XbzKGCBzG8reSXzXuxnl/yOoBibgH66ICOesr
sEF6cSTHiBUrhfLIZuelxbDvXrBFnYgJdmYruFrOTW72gNJtdXa6DXP1LMj3jlBu/8TlJy4+qJon
PoMHyT4LAbZOQbNbHNcghkqEandRY07yH97pyRUuo24jG3bgNdANm/kJM2MQeIl02RHxp6Y6hsXa
DNjCmsvBoEHG+8LK5H8SyTbjCuqZhZRRHZQmvBFJpf6i+VANQ4F0ilKxL7JPK4Dnef7bcbZEs1GV
ALHBtP06RlGN3n63umbEtjW4wAHJZITuhaDyAeYp0DAbywSjVf+0Wx50BMUev9W4K2ubCbmb5IUC
FQmxjbgYr56obuVDxxGWpdBAyhRx53LqdjAOCGjsLEezrmbf9K9JE8SB0qTn+vYbTYwCOKDaiK2i
40d3YaBay4Dz0Pycjadp224OriQ1sBKOnwnQgf1egmlSvRopdUs+uJDAzOuDALdcoPy7+iK+xO7d
oeTIZWCt5h4Q3YoE8S3sbOlq5TCouYh127Ym88T3URGfdD0ni6VfhOdBFA/Fj/jiJ1BgfclCo41v
M92DkKxxH+EZaBaK3+jBmIQ4ylcPf3HsexUFm2uehoymI104L5UwsD3e2BZYUarcUEnIeVMXlklY
4yQtl/yXl4/FFhGjg0zeyKtyovucnamszakXJxOsmeKkFAMAKs82bUi0FfwXeUd50ZOSdXSDzhjV
SF0A0CluWr5GJfcFKxUXFEzNgL+06iUBkPoNUhVe2mPcC102iwg+LIy13ujJ6xrESpvcRtsH5Xor
grrVni+WiX6P2+As4Ue5B37kkvcSO1mbr1lnrpZQWFAFBsLlU5kqk9ho/wylfUPob7G8pIUUEBGW
wJXoc9Ne77/3K8qtRszzBFqm6T9bPzkc7fTMJhmaluglmiHXvJ1h722EEtFnhkvc9XgYeMFtIRPd
N/0Ad3fVfbHuJt6R6GFDlrLonDA3KKj+eqNTifvP9Zq8vCPQMtgHF+jklDIDtEZV9Zzn4o/JWfRK
Axu0kzUDkH4xc3WWu7Z2nWENhGsA9caaVjS/RZ6KoF9jCauCd63+0dyoieVYQ6ByLuT5N0HhB0k7
UUpeJj/J7rr6AUWpDg9J54RB8sLnWbXnDDfRmUlh+kcmIFx5s2Qs88nwZ82eEcX3YHuej2aysoX3
G7CXPhqWYVgGmxb0ivHLOUvtYxPHz77MCdP/SJat57gOE+Kn6d+/Zwo0N2uyWlgvSeT8ku0ESebN
lrhw2t+ypyOwka7S59SsM4yjouPcTOvcfW9BYzOB/qYkdUdiC6Y1yKZVDKq2wmSkqh+M1E/QNR4o
Haxk5zc5YVTEBd8KvGQAQ87UGCnHJq71G1+pactK96nSif1dsKkwdYiH6hyglo8N11DGvbHFEGW2
dmCmIe6/Q+1DuvNRhWavQo/USVS7IrBd6tnSo/ZTHhSrD7KrL69EK2Lx5WGzqrInDHOrtFjMVsWT
wzxHYRU27JfChzhN+As+EncVdBQR/zs0TG2yv2vjUXXxhfXd1N+UJ6wmwkC4uduEe3Rf+8+n7FhK
Rn9SkKfvSjcHifKiybaOwgex2LddTM3oxKbUVsjghzO8bBmot8+qtVT2OJLdAIZ5cCjmbPeVynHt
rQbCiIBOL6i4q7bAXVzwPd/6B5UVlWGPP7az+1waZHujPMM+ia/bJlGCn7kbYzGEeFV68KKlWtVa
FQeFmt1sklBs6E0aXAOYNfjsAoDh+WvGbfcSO2uNLww9HZKD9Li0nQGVx9TQJJFFbbGbGgCzuroC
jOJO5DL5zUhYufjEIK7ZynMk1ldq1LGvM4GmsoIgOHQF6W2EGrejDu8lyQi/Kbr5kfhNBy85EEBE
O0ZNiDl03KyW7UxIo5862GdvbHC23W7UyOklygASt0eKVWHba/0YPX8vDwUvbkQjQ9FW+pgA5ubb
hTq6ibcgYx8oeSlMkgfkt0gNubN7ygqdhuOc2koorBr3qRqP4+avyY4Apu+qJ15VtlsRuKFL8WWr
KYXexQtQq4MT/b//s6d4hIFd/9Q185iK1SZwJ9I7fF2gFSVlWESqBN1yCZHTp4MQZeNep3pBSZXZ
GXE4Z8ThNOXGFGVPerzuf6PYoHy1wj4ObnGWvVgkL60/d7Q2wJl/hdCN9IqyaxK9sPQU2CTyIJb+
idKEoKsSAqjtvWMcJMC8SjKBfEKR9tJC5VtHo4lUG7kzUHmhsZPRgUEk8TN3I+0rBuajyuxDLu9y
REKx/Gewl9/2WG8bxRkKb+M8y6lU4OP6EMp+luuVeqswqutWbSKjmv4ScgyPFhH+1Vm7mgdO+UcD
akHZPl0+ouokE4vGq16q1aliCE4hAk/oLrH3qQVsFqKstic+3RNouQOrQwtqJ2qFiskokzx2kdn+
+MItv9o80cfo6m6vpzfaxM8IvVTPDJ5vAopqtgVtXKaKm7AgvU7hGO/AVZp6j51H3XaQ2x4Ugysy
QSWDbYxe7xQeNiMidlB2BoOKeUo0K3jOeKo9gwJOog8kxiKlTtj+Hp2rZqV3fRidCLC2hDxxeu07
AjclBgLV+EjKRTJ/+60hmUBPm6fNkk8PEdjD+iXsXEopK6djhpyr3egwLMrfSZ6ysUYhKzFh9mHS
bAMp7dPaNxRfATFeCw52NoKsNtZdMM0jFpOR+gachriNkVFtudUwuk9XjdaH12nhd7bMS9HECgx7
myT0UGkvwWEMUiideAnatLub021p07cvuNB4w222vyOWUEn94N+IC5Ud0P4zNaf0zwvJWXTh9uqc
wt5iEpUYnekY1dA+wNQ5carAeHZYwBT9n2WkOUpzA90JvMVMopKKsJLd1JLway4e3K84gubGx9Vj
bxpuiowIXuR2qzhcYiZbYZZ3EemUqINT2D8sw274idLh5aJb0p8qWfaER3xUycatQND2Hx1UUe4V
EggO+UH0Ga3CpSA/uP8twZzpJOXqW4KkEDJyMb2SwgQSU6BWuuwq21koUa9NyCrepFVDQQv/jkt/
TR5/q8HVEX2Md1funv1Uy94vOX4krPeh1Et+LO8B5ALrnHz02XzbMAQcb0Fn6vQUTLtPUyXoXM4t
mQYz08CwMwvzY+xezkWuG8DDGNi6ElY7i013IudWVWe7SsgTH9kk/uv1vfsK8+UHO251tOa2GkgI
Uo2hGHbWwO4q3aTuHg6e3QsnoUuFodRXxCkeqO5zGkgaoh1bDbExsRXiIp04TY2vcIyVtOJ+6ocE
+zNYKtonelDuWJW2K5MQb2mMlPO3b05J+Xhqf1NZ+/urM03jzbEuvTG6g9s/XfXdiXuObEByOPrM
nyyTELNDKkAMJRRswCMBnVzyA2vZEgtdsFz3SJyHuzHobiZ9SWV+Z4NrTXAPws9nu8V0+Ysobp59
ijJWSjXOl/AnUYxOmFKQLjrqRtedWsj3WbNTBx3aWgdn+zZWy3qvgVNPLZsmy640+zAdOXPes1Ib
PbUHpBwzaBJfA8c2DkqpVTqnsF/+Ts+0ITqVmx6ny9YYHlHKwk3P6gcs4/wzYubdrQGeTVyCC8l1
fA3VEao0JUqICDt92XRFf1bdaJJ79TqLoIknB98X+mgdCPzO0uefrQ7K57LV4h7Y2KIPdzvsuSxc
X6xtD3bLwzcfGSj+j92cxRml1Ldnp4PDGIN5cqiEas4zkAraaMNsc4GAM4dQpl2RyNPONyYdgIs6
VfSobFKvT/Uh+FAe3s/t8aKhytqQmU1LqLMhITHF//krgwNFhplinyFaUaMqDfqNO+Fm9iXS3Iy5
lzjNUFdgfETr3Zg1VH9BTxSYUoLoZtaXKV7BAZpHy3hXvxP8vh6HIS/DWEEh+rbNtIR4kZBKOfLW
NlDtNTRb8i9csHLu5gSfj2zMJvAF5SiAOX1JizUoUqtwynxMCGEQWSxOUX6LJKDrLReIWXpFksM/
tiLxaRrD7s7+iLnvFs+jywxIh+xfqhJjFrgVrR44SSg70dgm9JuDncQq9fC/jOHCzOXNfosjfaD2
IvAnCuzyjBBJmHmERX5yfSDGz18qwd+FWt/3tBJq5M85x+cFZ1rBDIT9qHDdl2z34WP3YMLZTL0e
mcgTy9Ef3ZcvEAjikQ0/FU7eGSdshwnDGqCia/KdWKAzDfHfUW57XkUuueEERwOlydERU+a5tDBa
Qo0glSTWXRzM8kqa7CG9fWkEztryJg/jHztoh7oBpIPwnj6UJWxosby0m52szP0JOV9XYqTAxTEu
ajnk4BXLJaa0hyy95+v1xC02XU3haD7FvYyxXS1NJFFzGOIuOt5HY17DcrMzRJ0oacv8/PD8fgpa
/BPnhlDJTaiCqQj960B9IqWL6SiIrFkL8kof/nJPL5r1xAo46Hpz1JYGpfSd6r+61mIj/WFiETUw
/2/r3MHPVp45dzy+inn1mrdkAmk1uRtqdrfgA9FPWg+KhKMAHj0q78hNT6vKQ1MOD1qF+CA0Pmh8
1jLNkSCD296u+LayDiv+BtzgHdNarLn/8cTupZqP1ULSsO207IanGCX2zspv9DmuLP9r6K16buTR
RwnZIBx717dzNjttNM3jXyZD62iW+al2bMWyrXNmM0Q1lCsB3F2E4UlSXT4O4ysLWc5WJJkm9Eb1
kuiY0iH8fZgCXKmcRCnQxYqAvkySOE4k1LGV9KukuEDYXWRX0T7QShn5BYbjoH2EGMhU4ufF0sQD
KZIQoYX950Uj5aYsJn8YsHAxBj9E/mNrg1Gofrjio5lU/73cJpNTj1aTHluIAJiaVjDgmSQKfwSo
jYs8iE1y7/qEXqTTQOH7Slpavcp+ssexO8x6paxXxhs2H8t7Ht5jbQT+OSn8BBfFLO+YFkov2Swl
ewz0wCch6fBCrFT9re+RHLKNJgp5RgNbBfBlbwOuv93W/2qhGiGAMzVvWtqj5eH9qKVXBLksDaeN
hH7QX7uHKI9nY5ZLqMAqZ89M9lYa6TtEfIxpQZUONTXnq/ZF2CGOp8Iwr4bqXOXaqGI7aE3ZCNEw
XWOLQuQqJjMoCyIC7Tm0Gwz6rS+Mi+ZFhKU5seCpiHVsd9+MkwYdE66xP8/TnRQ4VdZQvTtvatGr
G4/XJjzXqHD8tHqQpjekNfLE3Y8ar0c+UhlnZTCjW5VrJegHlVNKM/+6txeF8Y79vVbMPW45s4W4
oyfW7/PiharLlntMuLDWtYG4AFQhmw+MLfGK7JlHFvRpDFZbHzVE5Cuj8ZK6FI/CRud+Jz7ygLG0
nHMFGGOEF5JeRYPwoAny+nmEXZv4xADFxzTd6MDU8Udwoct5xeLNzDYaDpGDemoNArFKz3/X3nxX
tYgbcgYHZNqF8lZKqmiXsTU9Qm8kFlzO1RUYOedmLvmFKTA8xh3o0YmGHGXxNUhb4nKuXR9lF6DE
KE/Cs0QYYYqk+/Oub69siN74ReMRSjzg2ZYqdAfXN1ukZBtEiWksr4UagWzFo4i7Fd/kB0nQyBDD
hBuEkX8NUfeYp6NciVKgaeo47R8iRMMXXVvLOim8GdI5g3LK0gPygI8Q3UkG6qMPihR07ijZx301
9Hlmt4p3kxnC/87V7tkRuecwCrlDQOXNeBNJ5b1TjVO6+UW0QeKzMVAqqzzOOVF4tO9OFdA6NCYu
kcGgmfX1R3itvbHnVMkkAf5l5nfSdAOzp4qLguz5oGd9bDlewf484igSx2Y7TpyXF8N+8q01REI9
1Rlgbry8I2J44ZLkSz9/wa2VAqlZ1NcdevmL71VECj+MHyjYHau2DjHyglKNQvDVJtNlvsihiFG3
PYidtBr1dsFjWL9d3+Upjr5xw6ixuJ11glljbbH3IpE71nWKM3GTbVcebZcQJyOXpg0tWQgn+mrB
p4/jWAH0p502eIEkqHBqbUgk+7HFiZmbivHcJmvKWGIdKJ2+WmFGAV11mcfIiWVBhWvRDiCjWjtu
C3BswVQ9+xnEDKB1cg8UdXSGT1cZ3Hqc9KkyHiTmzZgR2pfdF6xlbMCOx/cVk94TumnvouIqKWmw
18VhZrm1DpReC5Ws6WNqcK/d9Po2CqOK0+KmCQ3iYHr/k2OmcRttK/3OPwLrbfiMdK5FCieK81yy
70sbDEMNPlc7SUGDyUv+W62+eO6Jz00Hef99aiGKuraNXEdKg5H+amtf1ft4BLyXlYrEuWiWh4xI
ECSSI6UY0CGlTa9CicgwQg17CztzSuL1pCyVw5E3OVwKCA2cw9bGT+HIC5n34YlMmucjqyrXUqEF
ncjHF9rL2uT7F0PXZWWdcgjY7bCBf9dob+XXbqdCfT23v0SYM4YmPcOzexOexxwFUiH40wTlErnh
9eoRWmtQWcjBQHaPXKUNyVGJ+0foQeQJ5pymQspAejyUrjG1jGtxuwRBUSoggmac3LiTmIwqiMjM
qiSrb16zDDFSgyfrpf5DwEmowmPpkLakB90w2agMWQz7M5dGSr5pmwPzbyjZZFEUSrKNQTlFlKlT
YSevtBKK7T4vDBo1bNocJdXCZv2LoDcNnWRJLtuKSf8k2g1zRr/HG64TipNaM0RgE3TvrUtm7bc8
gPmqPIDImInyh18Kdu37xfnEU33O4/DQV0BsINw4NDISo7mY4Lmh/YxEMAQRLgzKsqynQxdalw3Q
c0CDTn7Exz4bd8UDRgZ/DW9AsdDUKDu4OmwFMD7iTC/4nCirZaw2ODOxJZ5bH5MtfDJFTrXFMFbn
JeMpuT4uc4HYVXu8YbFWW7jwNbwIouilR6ktUWjUMxthgCDPrkOdzAHe748Yw/QPTG/nb4Wh6PL8
AmZELZxuHtDW0ChP59kKx+OhliTk/CndYYkq/AbNijJ+4/y2vzRqcFSLDKuPMDGPO80aLCt103Qp
vIA98VpL7e95Ywu26znbLQowYUMRaSSWDDSVCBG0YU8zA/ic/JNTpW9Uam3FDFFyADp2gPOBeSVB
q7yOoPr9Om/yvtqlW6QwEPxBvVzY/Ge8DkB2GSAJnHQSuOajRvVZnScldEorAHnefplF/9WF+386
z/1MuV+r/ltT8OgteN3+Edvi/mVAZ3F0v7Q18EgtBXFirz+rwMIh9Afpir7o/9gZB57GGrJfMFyl
28v9cWutGFcciFU8yinDViTTx2eY1CTzVpOXtcmRT7ExVZV2wAWe/gsbfkUW/ojhLyw3IRNMydpf
NdNLtwLDUVYVOQgH/gVjVYJqGuNXtJPubnW4yWPEviJjvOv8LMlgeQYcYH6OCaKVH0DdNMhQyDmc
qPyV/9lZcPhRGsbWNqhVzeb3vZAJ64CQH67r5fO+SKOi540VGhR3wCxTzm47Oia68InsFAl1Xw9r
kmofXR+CY7bEWaoo1iL5c9BGjrKYb4Fct2LGez7JNoEy4jm0zj4Sjf/8vzHNL2tqR44X3ghENrhE
h8sj90jUY/qGFt2ioQfyx269yqNdq5P59WZMHhVcnCPEaRDRLwr1oRwF6AJH2iVuZi81HI/7g55k
SFl9mN1GTgWDl11w8AbeI9is7Cup9iOZlGyize7DqPAUwKEGr+9YRA3lP/hKdgG96FYCm7y38LBB
fwZkK+stGcc25meiFL90cBTfJXGsT/S+NIM9AoL6LFYvxaJ8EtasO7kN8VeDXqrgI1ydmuQSJxoG
iWv59vxyqc3lAOaZp8YVxELidC9Ha1uBUsKb9GEv4jQmAPgB3gByZ0UeMDeeIZzDjFMxUM/a+MHg
YgH/DzUXdQzyH70OP6Bs7BI5HWMdLDaM6cIpZpbiNPZtnHPNpKmTnhz1WNjkFohgeTgvO05xTjGM
T58EkXqksoziRrharNK+prvXclIHhWOg3E9Z4STwqsCFKhaIbTqB5EmeownCIW8y6UFt4MprXgJE
nNGUsLTiGVnObDBRUrMc7OWNWgxwjJRbh9Pcg4hrrJE3OSy/qNRtrlgsbgWQ2ulJA3bI7mxrItZt
bQo+jucdsX6mek/P4I1dSWilsHCUotTTSi2R5P0gTcQwxDhI1SKYX07eG12kL4PQD1envxtwjvce
Dk+w0g8NgFIEuOFS9QF6HSa3TKiOVTnFdyIuGK4S/uYC9QJz3S+DXKryaL0KqY0+/OhVgxbGH+6b
jMWwja+LaY4Z3QffPAPjwpQDqxCEpqerK6AU4vVMBNCKCQzQmU3EjrSrOpg1zftk6KY5AbsOix8V
jyx9Bqf2xcOEiCIfCym8DWQKUXfV5XHP2S2LFoeLdQ7bdVWLHsm7b41F2lhpt6+OqTgyNiEMgXPa
Dzoe+KNK9zStm7HpPr8g2eD7zgHnoMGa21vceUFICJmTOZJOg5/nV63O8rPL9NoQFKCNpZAJa5/i
qsJZRF6QbLWLwcqcu8yeRCJcKf63kl7LWAePdYJjzpoYg6QxtU0hNq3u1sC2MdnbhWkcownBrqgI
h+iXvwuJAPpC2vA0Ssx2BR724BcIRw7FOHDJeqoGBFRD0BmrpNlQ032H6RQlH4qNsUpJ/NBUxdaz
mn2tbnayBCKenICtBVXxW1qdXhyEHE1LngSheTwEK/Mi9IHfCW/+sgd/nG8n17abEWnjqHgecp5o
SjhFuliDn/UbMpxhXUt78CJlMii1Iye/9q3xjtbWoPZfYd1UeKm8Os1UKr/vsPURW2mKbT179iwK
X7d3gpGPt2MMNza6iDuJPCQMRMSjFeHddCl1Nuq24KK7RFLVq3oWj1jVTomO/U4vteat/1QNfaWC
7MJnoPHv0AuZb99dzim9ilJS33a4V1VGIb6iiXqV6Je2X/rnJGUsPVJ3DJlZxkpFVk1l2rIgrGVO
kV1Z5QOJwszUyKhYNSC1bVyCZy1TnZp9kANo+Fov70lwPZ4z9b1vdPvdnGfSCR5U1BwmVLNFSwyO
q54KgPe8erLR4JfMDR7lsONb02FqfqxO472MNYpQrZJEfBFWVRlA0jEUlto0XZ0ys8yRTcnSkJ/F
0vP5459Xg3QBG1NKIbOs5279BprkdX8FwcnjEQJDT0SYnzmSiiLh7snifE99/avIcHXfcmwH58TE
dyuU6QWtKTyndz7MEVxd0YhpmeChE5A96DyZGRjJ2l91M4Q63bKYXDb1FxruqkqIjR4+ezUVLDtY
tljddS11FWW114FWy+S81ImqpraWotI7SPtAKo6gSJG0t0WGm+oGbIserp1kSxYkw/qC9DYulnTm
JrIVbgmr1wiXMv8AYplvmbfr+AkreCSSATki28RFb4BjKBDu5VG0PEb8+yZKmOCxA//WX9YguDv2
IwNnLeRavffA0yEYfMMhaJnb8moig25F1FkS+wqSU+N3KQEA6SIYllDE9yfJNgfmDiEUe5qyi/YM
IzIy2wLKRjTw9wP2tBJv3DTFfjLOrC2vuG/MmQCX350f3n+GLR1bhk5Qw7GTe6ZAZNaiUqjwVEln
sKJzokTTTgsT4fuatLtEy+4KHwImeEm4QW3JbruS+G71GGKFgvklGTSfTCPpdDMEks1Ij8ivOl1p
9+MjkbUsPz2Btjw6XrbENG0fPytOVl7Aq5iLL2rCVJL94KUv9SgxzuFzZx9cPLflMiuNvzqvRXiK
XodUhRa3kvZxtXusgYLG+fbOggCx2L7K36N67xPsXV2fZWSFxXXy5OlUke4/N6lfPJGq9hBNI9Ym
V9A4x9tTSF1273RVXLnTRbpFzkaKNBsyIe1lQqpei4ikeWZVHW2qBXbeenIciMp9fsUnfnlL2rox
LDJa1lydrtf/99gIDsetdnAcciACVIVVqpkf/I6JuWfcHZUWkrGsa5kL8KLZaOYw40Tkg6mws67J
XUM9Lvpp6AMkXbv9SLynAHgS6wjw3190nUmJd8lTAg+eCD4ddfUxny0pN5Ly/X0F/zMRuY3HFH5m
xRwFzJJfYKzkJ2SQoMVWldghGSXkbI8ZUm/hA8BHwgdx3VhecbRtvFtEP6tEDWmrgeSNctp3Jiys
ZkFYB/pZHh3zDqktmI5uLay9iKQ9t2WvB2Duf263swK/wJcx48fvKuef/LfhDRtNjF9uV5Lm+uFE
036Aks1aNcXvYlNcxCBn7ySYeUNT2u8xplj4O7l/TDi9879VJI7Ea+ACNEl0A7k7ET5J04Wk4rYc
ONpBEkRlNJiwm2A4oigSJ4usoTdw3RVlstLE5SNIYZkJwK77+eKeBT+Fg996IWx/72Yl+TqoieHA
ChoglVaSxg5TBA/lj2DSsCxxqCJnDUaX01xN6dFmPfD7VTpxk7qwhtkkPLSITNN+1KLm5Bjvs+Im
AJ3Tjig/5WgAloKOw4/+HtVLtfT9ZXz3Z+gKmgm6r8OsvslS5Sajkhtjz/AiTeRRwCCknM/4B0Pi
lm15+DMVGufrDDAEp9Dq2owONWsq8D8u3hSvBngQ9SHRUdYSVlDBbgES0TKFeBTqlwx0teyQ6ik9
dTIDaFLgReKzwtzH850TpoeCyVnHzWnRkTge4WoT0A8P6KWwRgbHgbBZzrw5Bq0c4Xr1Fi74iWAG
bRm42Ax+DyQp5fK0lvqmRpewDIk4zc7XB26KmlmDp2k19jNc8wM/Bil2wGD8GVf5froFZHpbRxNS
hS33z9aAKKlGTiusuO2DPi+x9x/QPAw3XShLZLysJsXnuuUodmB6UfcaQXQp/KCDI7Ym4lMiOhy5
1m08Acp2Xj304awvP9miYnOMyFrXzoqcS/33ZBho8dWQ7zUtJU+/R8S4nQzxVWwQ3e2u2gLUn6Jq
VDQsPo3+jvu8IitAVeT40wwnY1uuMgYcQmjY6qv3a9UGQWt05s7MGIdhSXUbl+7zxVW36fn2I6Ti
P0M1/qVQgUEVESTo2V/c21YYgOC9AZZ8dqzYQHGp7OesBYvkqsswk5vdw3wOc1Vzli6togGqyFO1
0OKjjhJuodq7pL393UHmPjzOJZmeiI4RSNciAm3Wm8T/7emDZw128owsejHZWEbBieKMNkKLrRyj
gVbpBPcLuqgpbndQV/QYQlLtrmZExe8bwEmGTNlAzbTTYQvF7U1lOugTyp8ti1T+eST2hpgdtUF8
azFtNHlFQWegv8aZhBZ3QzhZ7ctlCFgrVCDXULu21TnLN/YA4p0qCY4wh6DhZ27IWy15OjMDqphV
vDnk8Y6L1LXuT5Js+pvG5gEIpHXX55xiV15cM3ntKiuRIH+CUaUzYD5IEENi6WvzlKrpw7sM7aQd
jhb5v1NGAh/8/qF8zDA6vMtLW/p7ydL+RlYPJjnyOQCFRfikjz1APImQp3xX5ad2KjDF1bVwdq+a
VflVyHlK83SJlHY9Hj/ko63OsZlR613gG8Tr5QR5MTMMavcSfv7249osmKJuOqBPzM6p7Ie8wK0W
RDc3MfFBNOffYQkRT5Wp9IfobV6oOpqf7cP8TkpCQQ2hXBPU+OjG2ckUgrsxcpjlzRF7mkWGBwac
HNNjyxVtsIIYOQWmeS36kiIeA7slCXgsTwnBfQq7eEhFip9+dc/RADzXAL0+mKwKf9wTIDob/Dy8
Bq/WtuIqFJgb0aMKewIrI9jtysDhkHqgWfnitHJX/T4bytVl8XVjhwVw6x8xkd1sOVvu5FJ3Kame
Aunc5ReyVgKjb43F2zgf7OaT3riH38i9Zcoygdn5U0dGFMQNNDyp1jjG4zKwDi7qFkS/MjzPjdGo
gExB8f9QHic1pnqJXHiHcsyDIYG82KjNdXjYJtdrSNBhZE09ESu455Bzm+zrHtON5I/EG5KtdLR2
BNORk6ap/xRWykoddxoXzN9u9MKAupdm3EgEe6I7EXpLS8W1uF4n0XYFucL0IibWhapIHm7Xcdzg
y9sAmO+KcIRk1IGqfla3tUrCuiBmUYneRsxy6llzaz4JPd85wG/31QY4PmGhfIL6PUcf27S/pyIW
VAV5pLZtRFnQcZCfeKoKuIylWqhtOCeI8OXjzUhJm3dJs6ybptG4BA0alI6kkNmD8Dggy4zfELQV
FTimVO+k7+p+SznuB471SsdNp1D1E+YTwStsurvH4fp1xoGgkDjPWeSbu7XrdX3p3TUZM9VYkjr2
OODEbJVP6a+nwQrL1lIlgWx4XAtETTWoYwW9RtLQT1pJ8C/KYN0RCb5e4GPvRXLe+VPViIBlZiZo
imIBIwZRguYr3R+McSKSD4dtBknatIdKn0GgqPGMrxd17qR0lviTJphDX4HtC0bkWoWH2AlWW8dR
8ETcF4uAgcb6hM4t5mHaWPXvhvdoZ1j6m83sCvInECqvFaYam8e7b0+ga+0B5HIcI/A4bkYUCGeP
AXms6wZik2SwaOWlsiOgosql2qTongnlr9fT2EnIfoVHAOpY8B9PsnYjjSbnJ14/viTY/3ug6kLZ
NprvIvDAdZBgCqoQs2LX/1CEDjEYkKFIFwlaUDtuH67qPggMhgy2qdazjgEAQu+dZirRD+ioAB2z
LLC2sOrObgfBeS6Gc5ILUIV4qgnrqk18qTtRJheVkHb4Fdpfa4jOaA4l+aiLh7htRcI7sTUYJ8Iw
eDOC3eIVjAJj1r4y+QkWaAg+Ku4cb4m6tcsb4M1PSEM6aRl/R81KaE8b+0vmwCGFH1K97ZJqs3lG
j7kLCp0+VwYQ27gFKop/vf86b/nvEiQtquyTQctqBDs5LI1FD40NxruMwGrXChoUrBx+8+jHACbE
PfncBo92Q/3b637o1RyZeL6a9D7X92FV3w19UutesR//fMGyYnVCGHYr3NGVYiPLoPMjn+QBSOMb
xhudR6f4oNcLtM2WT0T+GRl/H4qzVouWrRFkTUHEdTTe1cAiYc7FeKeeFCnKQRNvEec3Q8Q96b9d
J7mP6U4cPX0X2UruaYY/Z3hE202kIzH6BSCdlWhMraVoqMpCsWrNHdeAbF2ltFjXI89JBiYujo79
bsBEiy+TGEg6wESOyUftzXFgMeZe7aNPUq9pcijskSE5EdwLfqQjaawaolp5bL8yXBxTYNViMVmz
jPT8q/GS0utVV8xwUMZaNC6b/AYIwLBWR43X4sDFLBEzMvW8w6/3mPnU2oDPTuuNATkQicxRhxLp
NxyZmuF1kT6YBVq1wF/0ihfgJicQll9CWHVmQzKNOn15+mCTsUt3KSbaDqrzmlRzO0OXzz8oqII1
guA2HzouIxp67tewBXKQo2R68hUBBXIHgpcQ/uCDPehRzj2h/3nU8lqEwZSRfm6PKSVcLairHPCl
lCtrJ53yCC1kRujWy43ks419Bes5YBXKd1aDSOx8HIS06sYqkBByTgqvCA/R/hDaS+trMYMz7LUj
S0qsTQxDam1D3PZhE88TZ+MGwuSbb5H2JAWdBxFWq6RJTIZuEybx8VhiYLCHZSz4UqHR/PS9l9U6
336TWiIUk4nhENE/h4X92wEPH80tyVg1mwBa7fQZzkAbHCNikQhQB9dk0P07DSa54M46XVMujQzP
QWIpV5VThh6aznZTRQemXSzHHMnd2Y2hrLGhQItxBF5ExymysygSLGJJgRtBdGhxcAkSGPvC896o
1v+KUQp2ZZ1FAkRwAbvGDI58obamF3FM7L1IcxMiWILfI+jZkZneDFYmOiL5C0+v9Mmo7b9W/ZHQ
wJrWjvAdDRpZm0WK9HPso3fcXp4kgmjGfdnltVmMonqHNbLjIlHRbgKMq+LWcOBx/9p7z/VzH+ho
UW9F/lEDdpNNSm5vUh3XtnwvtyRQLFoPQlxar3/0vcOCix564bNsBV1cr8Ulq8+fJkTY1EdZzrxx
MFjXi7Xr5B7Qj/T3gL8516ixrI2leT+snDTJ6UpJaUvmzbz6XKP5F9ys3aUtkaZbO2C5tZUHbQcS
iG8dVGNec69707UoqGbQgXRRLf3sXniw7HT2qPuRkIXg9d8+shDNhasBPyw17LuOYdRocE/ha2Yc
rn02SibiFNmr10NBJvWA6IfcMk9ZipBvMIbScleagHtq+Bf0JeTKV4T19/UDLWalapSdq/ZSyAbz
PLmz2fLdHQ11Zr2wuhYIL/8OYlSewDt32HGii95BHOfOIN5d4aVl5oMThfgUw/sEt5wAO4Nn9X+0
AD8mhXVCTqycwmTJZU46WFgVkpobMxpRhH0n4IpZ32DMDIGecLyL4jk/yFP+34U4gH5g73BX6W/D
X5rPzLzYXJ374mW+o028unb2ql2IQfRL7FX7AVClHzH0/qR3XuwlF4pMWLMv/UyBX0MrH5xRtujh
2wvjS8fXIeTqPeOyb/BlDfnxuYX88Fv7q3AWQdzFm5dweFM/Eo/WAWAKd1W8TYj8xOGaQcqoIHRN
al+CC77+k6TlAAdYCJGDc6am0fbyh84VfIzzeLTgqkIxVwxJrGik5+ISWCWDyBwny1TaBpaaMk9T
oWwboNgdEbbzl/Ho/jlJxRlWLzaZ+v0ts1KD34m5o3WKdqVgsdj20FQEVbJNwtqfbAHF/EnYWW7r
PJVwqstouu2Vfe8pzeqQxVDXvK6ciER2bIVLJ14i+Va+JvxkzNYOFN47bc9DCxySbp/2ufnlqx8N
qqcE+fV8fVaAZD569D0b0FvIGF2TyL9fSCef+EtWmDM0OJOJlH/JYkWBM7Q7zW7bJZgMNDUK5Yrl
u304AzrLvlE0jujz4LGK/GUQxZIDf+cMMnbJ78WsVgAJHU7slvR20jexYcow7NiBR4nF4cgMt/dA
qPBzl0jmAKcUWldw6DGV9EByuV3xW0Y9oNmCKzIS2n4s1poYByB86UXn0lRafYD44Qhmv6z6I9ys
kadscZyNLdqJfwHQ4mmsK763TcX51LOZ8Iog8QEMvOyoDW3qTzp5h4JVyFNu6oMo2r+Ns4uTjtXU
xwZWgEVNo8NMYYl6rKeVY2gMCGAVemdKhDTv25VzLVNjDwoZTf0kkALgPz/WJnMOGOFP2Mkd1XrQ
n6+E1ytR3XtW8K1tCNc5Sw0OOE29YwfIPP2hVGl3uXx3uDEgqsbqLKcsF9VaBeVUY0c3Na5qx+t7
HXsnlxm7dythjYU6ZlZ1MOkKJ3cmx8m7sSSmYgEpkV0uzsUN95c3j/XBfpqqK6S6M1At6LxWGfKV
I/lkMBMXeERGiyc0KX7wx0mcES8A5rn6snXe9Ilz+jasQpgUyhf2URu5Grjpb4nUVbgBBb6fJA1Y
GdN0uW1/BlwNKAahQgG1Hrtg5VYmByC/d8xOgY2NP98rppYvK/y9KjnbYSHTLy+Qaphn3sT6bqCu
ISQypNzC4BqAOP8nw6EM58Iegfp0vTtLc3tMYQ56dQ8VwgLu4Tsh77R1xIuCp1vpxXDeGMd9dIWY
ya9Ao6opFqpxNfYhw2FgcZzVIjzHcY2TBN6pJcLahgf+m077DK7uAQ9DE2Gcn6UT27EYpQamII0M
4N70rZzu210ZVMCDfaRFNRRMu2tg/DsliqpSYKDB9ceG/IU18/1g5gVl8kt0mXISyYyCug7kDZqw
9GRlUUY+Y0T0aRikq83jSMf5dqBg15x7QeAQ9TjNywrdNVz3vwqdlYMKZPmGkBBLp9lwCgACvhPZ
K7E2JFvQ5OkGkPxu7O+sbL3m4cXnPsHKSsSxUHJSjsjbl2tfGHU5Y2Q/d8d3moIRhK8sz6aZV53x
S8R+eH0k9bH4MFuPNMXIMsZ6ribFu2e2GrIF2SGfZEKEiNImCLwgMQ6/1VnF0FQ5ro+cQkuejy6u
zMgq0kEjSGyj/NvMGWf6rQtV+fwDiXFlwQ2YYAv0+RBp00mTc9ocE0Yo5b7wXYTTWVfbuVeS1H7H
V4JZNLV8+YRmb82wQAjvoSwYsJyoxdVHkEIk8WIi0KCCU2fxSX4Q9C+99kEdGD3htiSlzceuVm4U
/SI8wA/FknTKqnziNwHNey3hFRErpH2Sd40YmrEAx5wpc/r8TkVwS00KaCGO4U0MgRRfWOytdaCc
8DXYNklrIiyUF7d1EYzabSrC1XST1H5eznXNxkS8wISNRdHAJEX17ZeuP4ZbTh5Z6rabr/0ysi2v
1GqTGPvnCiPfpbohVSTVmeUI/xEjr6oK3pzYtil9pwq2/p7mxtxNcCxYXw23TsmRcsszPHzipOAu
VCqAsPKH3d3qKITYcix6PSQpuDcM0RhzbUOe0aQpxrHNuerIMDerDdp2pCQ1GDzUWVdU9tV8AI64
I5c5YeWfyuetygI0tGUCXcyRUbfsjH22GYGsdvHmB4jSZT6I6Slz939zpPUSc1X0cDuLoD0khQXV
J2GJ+rzglK5oUqg7SdInP0nRp3EcUO5/gFmOkKPWw36qvRt5s4sKq96nJiWWDf6LAaHrzrjPTCqn
Tdm8wYgOp42pwXvHlbLCzOSts/h9DR1FKQ9HKBcW6EDQ8f5krkTdCdbbPc1kJM7xnCZQiI2X4Nns
TbSEap6mAnanq2qqfvhGUtLfhu430mwzEUgOYX13f+gML6e1YbMjH2/cZNMmsDbLNy5reGzZaiPB
hQx+MnbVRjWCZPsbp39gwMhHbqpPwxZhNMS71hDsHHSHedFym8xi3u5zURl+EcsAwZEJ347NuKnL
JfXjfQvJWiQi1YLlbM7C4dbVpKZcyE0//Exun8u+9I7JiTXeQGTV4ko8zAFkK6klkEjjntCG33IZ
kIbvhOuO4CEQwdr/DuhQO8aFnF/SUVuwGZTFEhJzfyZYKphf/9vHb5Jx0rGxjtDK19NgsAmSKSQJ
HtOj4A41+mlGf2stAWan8qJr+s9atumXIXFlT2E9bwhSQDCat1i8VgSzJWdwGcRx6mTHUFFceBUR
JYTr9XXAzx2Ee6NJL1wqo5xbW2BS5fpBMZefLlDycnk0FJK8KIJIY0xMCY/EvtMA9bXlYRkw83zE
30vIz+SfX9BzBWudzWNWfPFUY1ApN2Y4BypXje5s6fgM+Q7ARmb3prUxn9FQRBRKcmbJF0Ax4F+5
N2TMyWapxUkByaGnFnLg8n4xkUHI+9zVVt9jR+X/Xb4vKdkKyjbGx9XEenHf4AT6Esif1beetnxF
tOczjWNPL0SKDDEzyXC/aWAuz9geH6WXtDSuuZPMg1bOXg37YEVQCTWL5yeWu5j6dhSTpisS4jAx
BaDVF4CpoVAvi/VirQLNLYbPCOqia60O1yoH0eMaFbcCAmkTFW2PDvtZS9vYc9HxhNG2u275BoUM
zkthJSglcbiUCFCqwWh67sZj+xZpyn66AhOiq9l6/r//yvb77/Wxj/YCAzfa562xBPRfgBYxQCVe
+ZA9vY2im/cfsG4xnhFtJlrm61FkD2ztDpPPgx9U9m9/LiX/QDdHuJopCtmGNirfUFvRkIpcFXWr
y4AapJ6LBpqAlYV9DIob4Sj9VVAXycqZmKRkFGAX4zw2i4bdwtIy71tgSrbC2ikjXKefewfiTlin
Ma4q5gdySE5+9p7mfsADFaUhMYJUeFMIe1WwGY9JqZmAd5cSOrd7Gp+16qQgGLxoZtE+gL1OE4HH
Mr5SHZRJtXGd54tHIGsccYBtcf90aDhwrAKp3RwzhfciFFzzvP8b81xqNJ6JGwcu5+I/5pU7IF21
vsnlycYhEhX2+wFDqhj9oujmhIwBpBA2rAUgvSDJ2A1edfGzMcAZSnn9KxEFQSbwHoFo12nU317+
pjVaxoE1F3FRhgqb0LS+URtW3jnbYXcjinRHoZ3I2B8oVuRQRgBn0ZxVLR3EYxY2k6hKlKh+RVoF
AKv70xh0OShTw7LxZko89hnDmXRhEAEnKaUaMyEuBiOJw/3vpwTfeErhxetXGtcCGFtC1HEhszpc
x45pugaxUp2g2UDHBQ0YCAIP/XUJ2lAH4+CVJY4mYpM3sJL86Gp+5Oer+CeE0ZiiX30MUctro/z5
vYWgheN+LuAssmtk/+GdzeSak5LJ+vuav2FOhgjQ43bec4GX2pHmrQMsCr0QrMD04E9DsPYXRufu
XMUy9PzRUvheqQYgRK0dxJbdbde6wFoOCOBu1vNNxPJOjvN6pvoXdozP8bvgDMJvMANnczxPU8VO
6LGxL+OqL2pxR2VD3WQP8oSluFky/6wCRrt4B/dcGTvTMmWFMe+UgChBuuSEQ08zbPREOgfgUn9K
Rnz3ONFL7wVBO38TPQahm52Ade/E2hKcWh8g8VG3W9C2eMJbkEi+6tUpgx6mKAkLoLAG6Y8Fh8Cg
liYjYCyUeKGqKRNOcY/Dbo08mQ97+oyUHQXmfGB9jxea9ERT1EcLd+hEjv5mWtDJXezCcZC7w/Hm
TuvLCVGFxFbZ/sRLAsqrFLCo+elEeNCGmNFGKnHE0Fqw5o/MIYBfIRB+lzqTKEVkrstLx1AGXPq3
NlqPSAZAZ0zvf9zWk+FoPvhBw+l2lKEaRy8uFXnRHeFIAuubPIfLZzBV2/ItxdAFPNEb7Qst96mS
BgNuweOGrb5LUs2h1z7d338zu5KSN701CV4mLAvF3ur0wVKTJIcYtyqZeN1j7/ou3V025IalAIJ8
FXktt0C4trq6oZlnc/EpkwAHFjx8UKbOVRPr/7G3ILlmMA/en13UKRr6OP4AIrNMkd9L+o2Jgmkw
QQhOOyF+CCsg+D/7eDcUOHZVaMuXBYwm/lhlhWrki+kgxHvpXys3U3kBy7j48UiBoYZFm7YGmEq2
0lq0gLB9EJkqxmar1IRddQ/oDtzg+U68Yk9I6l5IXoCvS2uvn3IzgYlg8ahihe0hqpTIpXr25B/u
wjK1cFQEGo0j+qfRuNeQq7sOuZV0EoPmk7qNTQbSMwl2N0tDVvcBn6W5Sl3Mj6MTOPXa1D+nXvgu
5n9fmnKkGtMtbBvods68KDCHwsTguXz6B8YMPgHVmsEvvlz5JJ0KlH4VlvtmLjiOHSLIy7r0X7Y8
nyP9OCkSagsloIeSZrdmS+D699BghbwSLVqhv9Y1qP2EdocYxGMqcDU4cK9mGj4iXN15oZysvUdD
KNDIiTIvEKtzYVHok0KA9/OwOI0q89l0ABABPQ1WCTrRkdCJFGMnz7PjJawE8umorh8+EA6p/s4J
gk48G8nXychTlBwgtdpcv6h9HN6ND4avHfFM8osY4ZHmZVZWsn8tkwKuuUAm29RYWftPLYMnyKCt
ThL+xiyn7dpjC4M5ioarmxILo03kdhdy3Fg1DmzTK18MmgRLE6fCUafw6j0ZBivePg4bJA45abMB
fANJ2S+tackmFHYQ9geLpj4GvIuWpFyZ5Gk/2D5pdqRzv/p7l35Ad5Ta9uVwLogWnHemupubQ+NC
Eqaje2LgYdmC8csNirgxth6rh9Q1FswLQ4gxhJJQr4gcRvWUeBRN1kAXxXkxh/WbxTdoeTCU3xQS
lUD3eX4BrluX7GERAaezmtpQAUzGRoOsUn9KhjaXn8iJTuOWQlsvmzaAIZYCjsFV5qEUQ+C+eSqz
bOJtaEbmm182tPiwISpTZVKbt18hkSNUkPkl4QzUhG6G+BSi1n8aADfOPpVuTyKhGysNVmX60UkU
BgDRSwrKk5DY6FeaIdETlDkS91FtJQ6yJ9NKZu2ouZ+bcBGtOVQ5LYG5f+P5oWVrxbN9DCIhh/Pi
Ivxw4X3gkaJa9d80/yWoaFsUjsd6pGgPgcwz/bVfIKNQohuUAmNofFEOwTI18mOo1GgvR2BBBhsK
66ePi17+dfw8oTYYtazETZHQD4cMjDb23FW5MXfW3JzX++xc6+wD7HS/5YMIZUmKRyAcbGC1JxjN
MRvbbf7VB/9Ed4toXQrOU8wLiG7pVECKEzxtsFkVt2krT22AFkclbIPOlm/0hS27D+kwSakIF3Hd
31W+bLTFi8CMlBGrN9IgTXesRztRiufw1uXeIMpWUwj9zKXuc62gD1NnShTr2gxgGSy5hq9a4tTe
YmDvnX5yqZ8W5dmAxOR5FIbM0f8n7/qNP3/xi2YJDvbZC9jSUWn7B1KN5f/DkNc0XSAAUYG87CIn
9wOxsV6pQ00AI9JDAxEU8V4K5QgTrRkItOEQdy4zPDezbgKLPOZUKkPFcME5PBCCMhGDD6vy56zU
/8ODxK7S2Yo16qtoxnMUPN/Kd/lgkLZ3wjMBmhUbq7HG3HVhbJ717dvYD2FjNTLHAtGImWJRb2nX
GUnmghkGatvELVPAcGnm3L3p9hhqSMvTIiLykILVJWXyszcD6xNhEVbbpUonwMAC44vS5oDSz/CM
VLdUZKWQvr6u4dVOlQTDh2+h8NmbWFzZdeA1wlbyEvUQSsfQSQEdDkJGarTbj4J/iGK/49OYsok4
uID60hOeNQdSKJWhgpI8ZhNm+5KfMEYYkfHU+v9GAU+cvHA/PNqLVXCQMmjsddb0WSDlT6FjLGAf
pvWFlz9dFueiuqSZZLePNwRIib28SY6Tpw0m45b8BRQEpsP8fazFH/VOu64cG8NIWsjcMEvTdHwb
f/NFztLJApCZkvmPCMydl+pvdKNOOZv9kggHpCmRwyxghjd8eJR2X2yDOqaFISCQ0Y6+Ks9BLKtp
CL0QLCPWl9+XeqHCv5OoBnnhZG8jYdoh1xLxlHx3gKAnuth2gG7hPZP05HiccvFyHXroqp2F+qNN
HBQVo1xEzuGiVX6dAYoIAjIQcVFJ2TsStz4XUO4PAT8dNzydfcBUSEAC6yrAisWLYcjfQwo/DtCH
nubshjOpVroUjcOPI5vo6G0OHonz95rz6boVYfX+Ytxm7qkIFxadqZM59Hxhgja0WuBojNn0OcJX
zDCWv71MZAku9rTl/bEFw97Z/rszrCWZZPmBU7Ud39tDu27yr+UHmr3GklaFVl3bHwiWsAhxlRdI
y10Rn9Q4XCcrS/s1yzx0O4cSQJ12O2DAVuEFOfOzt9aqFobyUfT4ZMqzliW6+ftD7O3uSyZu1J13
L4bMxbl7EoiPoteskW5Z8UecYBQjOJ6fTD+SZjovcgeGcH6ur8bjdgO/IDBkAl9W+9BEfBskeuts
iMAajRdOp79HyTJeKBKPreqHASSctNmmErdwYEV4O5jWrGaLLpccHwtNfjSOhhC5PH3Z6H15EamF
wscY/uk2XD9rTg75QxuGrPGdZHT96YGKUKBOhK0buCItvoo7xXwSVH+HlGwUgjapFj8yOzxrgAe9
cHfrrrjhN3rLAaO7wkShScvz2R13Uk7cSC12kg2XuEI1CqhzPd6je8MoUM5b08AgsiSNK2ZLDhCj
N4Cfm8FQEe9cXJQ1Ea5egTEv4dGba7dAJ5b0LOxjoJuhmtM4kleaVh03ycbd6/AT7RQxBBbvdv+s
Iz8DZa5ViC6yVvcAt9NdZ/jnQKErf3+uF0RutBxb/+ryVB6nyRq8q2pbFrZ9pTh7AND3zPRJwH8U
hS4UBIJPQBKM/IoKVZLHVig6Bv90h2SWW7au1Fnx2/y16SKtCdoFh4WBw5lGSPA2T47WEJIy/I22
cADt+nqS4JUyh5w9oLvQ6AKIFS5jew6UaM/7WAKl0+PD9rtYAwKeuoWPSOUGxtg2fnC8SIqSl71P
o5PTOKEDqWoond01Vcb7cgT2jkuRKprecQ6tzgTZb9qtHuRi0jZPeJAyotWSrCnhDucvKarnrSn8
IPg5vP8CZ3e3HmAW2YeVsaowELEwVVNOp0ZGXvPJW4IEzMXWEVSNO0Pvmvm8tzVUOjv91vZteLB+
S/Bki30Omz/FEwD5Zoad9ei4duof0jb9BXFfbkmnhNpI7bFU7Y8Z9qQZ2Ir8RzF61xq9rYuc5Tf2
UNW8AuEwhHMzncZAEQT/DGol5BEbp/rcoM78tOpBiCnGGQBmozdXuSVIXKGC1LARctWYVb0M3Gvn
XDa4aG31tcKiKBabkKdvF8YtPQxF7wzxNFgYdiiQVIqQxAD2TwON6kDuOotuP9Hs2ZJQUy1FAF5G
9p/fneAF1OiIlQg8tXBNgkHshWo8v77y37Q/MhnXesRm4oMLXe+EhLl5mfJ2b3YsAlyY46RcER2N
qfXk9JkSzKojLwfUfBQShr4zD1hzsSfzv9Co6brlC9mfcC9sbyZ3+R0xh9e26cyfu3anDfv3zbkz
+eJ0hO84MjQByiKXFEs2KOR6+BoULSVei17vcIwsxZxsX0BThjotNV7bGdgAcrMCOtxCOnzKkIjt
z0vJAvjmwbYEA8G+4P++ISOTlhUXEzkTq1aY3mZxCVmOkfZEU6MzYINU4mFijX9vrCGdz14GyU+L
IDgK54C255+6XW7qEObpTT4dXFVuE0YyqwkmM6BjrfSQRwbyiJAHJVcI+U7Ru2XRf2ny4hUVuEq3
K/sAQscH6tAq1dUaWXV6MXDi3S95sdaIkT6wChd28bF6OBd7OliAFEdqmv4dE+OugLAv7M/IP6Kj
K5O+UFg45OeU0U8bs0QK/qPKZlcMfiw8/qEHxA7WViarURlvZtFTe5OBryOSn9z7aIyvX+guQLFS
FmbxyMAMJBDjFoDQe3lxqmWAqZLTWAVIuk29nSEJPF4fA0hCls00xdGcx7m0OnWr3ks+QjJH+5Bq
bmW9ZcksAgZAyGfKF5cW3ajcf9nJAnJrYsbX+vcd7Ufsdk7ie7QZKLNadJsB3icRrOjDZQve5iC6
0CnDLS4BCocvJAGOVznAAJEL/qwS6lD9FyD3kb3kEGUJTNvksE22tYHh6GdC9j6P3R5yPmxg3Wzi
SWDNwFFsbZ0taEhwuvXyTPP8yUJypn14Veod/1aZXsyl6kQN4FseqLOLA9yu9kmpe9nnCnzpA2Us
m8g/pfOcptmUTrnyKwzTrJ9u0Nl8A0uJRmWfL1zIh8ufaX+czzvmSJrqZdMuUdrxc8TttEtankjq
guL3LQpzz/FghCLBRS0aZ7YuyF3xPZQuwNsJCBO332uMhqIcsuYLbZ7kzH5Bv8qtWmjvsc3XEaLI
0RQzFjOgtTNNJyAF30iG1a5a46ROS7oN7+vTYJ9E8O6/fFKcv8g8iELXUKGwUKoUP4mz2tcMFSsh
1c99N6Tl/AUHJNmSLQKhmjYTIimT6xwON+zyROBo/TzvoLEb9tvrj49/HnL6LA63QfpmkhBWThYF
Ys5QznpOfJRbsyvCuaSzPCJhydr4lGvYAsBWx6EoxUvJjoItxu/scBMKkqW8VL3hbMewAcZOSJz5
YfJvOy4u54yZhej6kbHUNKBu1ekkZIWLYOcGazIXpi/TGROl/VXHqUAv933Or/DqMTABMh8/mqf+
hmmX0Cazb0mMGAoype/Jp/uBw6931gNIR+QYj2KwNf6kQwaSV0vSulVdK0cS63V+LCqGQR2UqyTI
1WEzeUfT6a4VpYx/KUlKf7LUHp+NJ6fZWfGg4nukcbJk+aN60MVzjk77x6O5vPYb9pcj7dt3bMFB
rcsuohpeLSJgML/YCqwb0y8UFahgQ/aDVN9TQminY7qrEj6rhrz+d7mtQ4H8/xdLezJM+HcZMieU
M19SDfNV9V2DQ3oMzc/5pr99PTaRLeY+/BNzgT3dPsRFYcmN+RA6uJUyV+zxUkMS5zEkdQv9lRhV
cv1N+HRLB6ba6PhyMvO5dkwFNbjChM9wyGNDbFMreqaOaKVT8/vrLh2trMrTQ5TEpOqQyvgWgM4M
X2U6nW1H1FWJPF7OULNWmqIxTx0szL55RCPNl0jwWYYKXM6Yf42VdFmS+YuJL6VaDd85ycAs7LK4
pu7ouGSHqw4brKtinmxkOcwBBBLYzAU5K2SNOoD1U5+0RtoSsBYFFnicQKLqa0DGqWLUztzBm5X7
nFZU4HjdtZiflN9Lltv0v7VaRo4+VoLFlfyNNY6pcCt6lS7qSuUhDLbDFaJ/+VO20H4EfdLLfI1x
VwZdxxPM4rQG15BbRty1lZeqapAHeYAyPZ9xFRwZO3SiuGj9aSPpXXTnovJZ3sYJ6eYbbsBMoq7y
pgLsXyVs6q3w1dZ/o7N6aQSQu6BVE/v5FiQFzoimwN/SOgQdVFRsKZwCHh+90uWjkzFptHG/2W2p
QuWZ0R8WJ6aGu+sRc6qzQCT++AsqIRR0qt8U0UekOZeeMfZ6FHENahEhYpQeK85uEBmKOT+dDxWK
yWuGqTyajfHg2OW5j64Qu4mq+7ROXLWX4uaHOTCnQ0xO/tMGnTc67gC0ShGBlp8igX8a5c5zXk0d
wjcqV2iNhGZYZ7AMFH/XHnhpCr6NqrcTnK3SDF0nVdci4KFm47PV6cPuD02m4VZxJc9HZgnbh7Ma
fx7wIfbm+TRBLSP9n40O9eADyF2ekAvm2u6zdEaY03+YWOxbbLH6UoQCyGw2YvgjHkyPVffZ+35E
LDmDpZApWN1oQOn3Bu0tbkJ7pAm45GR9lIJ7np1xgLslb1ydFuPa5CWQ1x3qyHjAYJt9KzpsB9M0
N5qwapyNGyq8i4l8S/TTGDWU2nIw3Dkm33EMnUWjFCvbBcVl7hnH1IvHYVMXL3TOSUcOgNx7hysh
C6bLa0YwhY0wETPj3LDIgW5WMGm0Vahi5n0fVepJqjWn9LWSf85Frvc7Ixa2mIJLv6GfEQmsnpLC
cNCzv8fsmm4++7mpakGmtsrnGPgBPR5L99ES5rRpFfyikr94NxpzXU6zvMlzSpS7vALtHxd71H0W
libcjSHQIe2r8c07MPB+pnjUwbcbOsIDbkJ81fL+srt1GpoqpUaPekwo0kHzrT3WTsyHjkWa4nTS
zyxZWMNc6tKUDQHHOjcZ7v/J4nAuhopqyV9smhm5gd3wZVtpTiAO0FtPKPWfbd7+ZCsnNSWZs87i
Islt3+KOTC8rXQaddKw1yhrcPm0x4ibwrtpvNiEJE+IDa+CIkqVb6YwmP4FzHsV3v6Fmdt6gxAs9
mLG+reVRbeq7VlwpiU+Xz/vv8UzQrFxjKNAZ/yAVI11YqMutzXcUEouhCghuG8oQX2irmxH0+prJ
iEcSS2J+yTvXkAyYKHR1B87rpT++UtRGzWsjAO28pDGOtlxur+5uYjBMKyLsrLSHZRtpStLfAaPW
uc2HEEDs37uLdHOIoAoiDMNFBeb8FuhK45S/H6U+E4PtPZZ8wtXB/nb9U9hi0NReZbtOAS1Qg4mO
EBWUaYGD+GnqzkgGRziLL1U+aeq3i6NyPifXorFRjcd5MMtejeRBM9PjsvCC0Ie6eWmkBuCaWO7Y
IXGEDSXyO6U6OiyT5GQCaiR0KCOY5wmpjrpmb+ZEmJcoMP/eShdYAczpo/1ej7zB7ep26ndcGQ1X
P8KsUpJ6KQkTbgTfX1YHa2baLg/W19c4bC8vVex9ypQUlfJyW5L6CHCqZXpUZg67QjDXeb+bLM58
ncuTeTWmN7bBIDmpREbo7h53qxIAY11cWa62ams3SekolR7xbrMKp9GvHNesNkyAGTqaq05hVIPc
0G8Wz/tC00bmTvEpvClKsSx43FM4aS9Z+9g6bTdgAkj0VYrKqZ5skrLh2v1Wkyu9zBwYH+22tLaj
LLTWXGxLaz4gA6W1VOdf4eHVQ/vbxXOXwlEvpAxoD1zMgBJQkCV7seV9Pt7sIhbES3R/RYCOG9F+
SC19xTZZjUQ8GIMX0wFQWFOypjWkucKu6EVpF5QHaaX8b1sww9LNGR2AgQP/GGS5HCUL8eO1znQk
TYcghIgZMn9xswoerHGvRjI9Z3i7rbMxBs6BitvB5wvjTT4GcRQOXFOdLHklVlrfHtF4gYiKPhFm
uk6xjmdH98MXdhalROZ5YP7/Kp7EzDMvL9WB/FKkjXNhwhqW7VZbyMZLKHczv5fHxzwLt43bUPr2
uMrkNgPMh+4BSdiY5CRtP9RFBFbYmzE8rvqq5VyfrEowZyELeeIK7QhiMKEO4NvmSJg0xlXb9h4A
xQMk2UkxREqNyFlcMi2MwJgWq97L3YZHuqMHgtqOoBnWKYNXGgTGzLCmolZxvTrxMFeyZ9K+1TwA
WXE40UqcRl+wYfqeR6yGh+ODlMDEdUGjzKJ45+wWYwdEWobXH3uBobjlRoO9qhSEDDMggwhHgEHn
AajH6O7RItOE1Gzx7ppvu/zk5bMOGeqtq/8fhZlIMpyjYy2t9JTn1dXPxn4/Mfh6RrWd+z2qwrD+
ZxOHs5gMs879ad8f7ipGlx4h6B8eRUFBm30HK7VlxrdWBlaJNq1oesxjs2VwKkhQiB9V2MeH+zIS
fEj0rnndR/kjZChNP5TKZtNRRrLLrkcZufaKjEtHy+Uy8CphXez7YZDCNChC9TMwy7RauMa72Ib6
R7qOqQH86lkDzmP7sApxNpcrw40hdRevuSoILx8hIMgVwwOWvECwmDMpSIwmYqeO3cO6w5X9jG+G
7vQYvDym3/U4xcAdmbwKJNrUSD73O0Ss3OQ1b42cT+79NW5r8RJj/35gbe13fOwdMij4QEXqI8Yv
tOoA+oGmQRPzURPTwrSwbUThdX4eXJ1q+DCTePd7mLpYLVklahiLkGyy+qNQTHFFlzVKJuZN6mT0
qpfoUxBJhyDce7MPTQfoy9K57YyN4N26wk/a3mCZ1EZrS/nFW/awbl+CkPnNrzHZ+xPlzg6Vq8XY
WJKA/TOTMhm4kusrJHLpVFgs9J31h84gmybvZA33LzDbxgx4McGKHputmK2EL3QgGWjTN5kvSzO5
pB4m7QoCckv2URaQW+/b4kH6SO6WsIkMgeanmg4frGQrrJkxC+jCsT+Aryd+jakD6Eh4QqDpVil2
44l+qYLtafGJV99cHEN1TNqOntFMHTgYoeEZK0WykTkn/aGxUKiUUR853dpp7ncVX7R4TxuTH+Sy
7a7Twwg6V7YUKyPy6El/l6IhwiHHihbsD/7OZFr18Od1HtTUrBTy1Kt+Xq+JQgvIu7G52aZfGje7
N8uyT7OeweO1y5X+GLnaBAnTc5JoK/LacR2NmGPPihqpLjgtjaw7zoTBf8occyC27ctbLUeYZepj
zCzwX2tSG/lhq/UcI064OILs0YBMkQyk36LpSELJ6RS7U/vcgJriHWD+A/E5Vdz4MOsZ+l562JyY
ieg+F6XAjYgzoGGWSKxUEj14BfD0QUD2aVEA7fT+Ax5mSJ+hDyaQcO3FA4kpcOQ7108Pl77n7X/E
GsmbURWjt/kfG1XiP9VPPYFCCwPsJ1t9FXXb/tCLacdDgT3x7gLwUWWIvw3eHgWCAAkKL/2QIp1w
2zSv/23fshkOZ3Li0Ie24JBRec7eNRNxeEwf4pO0KMqwX41rx0bzqFXhbKVH4zEXYovtuWbkZQ/K
o1TFhbI+fy2SzdMM0Fhl2IjNQo1wjrwcVtVN//eZ8TJn91WG7+5Vj3DWJSFsqERW6cp7mqEbvBE2
TZpOBXNqZYaMRG5ie+GLGnu/SSKryf9uBDK78XPYQ/uyaLolTxlfcNAAZ+pLZOvMbDwgyZglyRG3
5WoAOuaNDUIn+fYvfGSbnhIkw5w8ets4L9VBbt/d2viY5Kzb1TRcZ0ZzSTHBB8J6k7fuPmSlq0X+
FQ5cswlRhBOr8b2WSHoVZzR6UysD4kAtQA24nfY25QJlgeDNU4aGZMt+zvS+uGVqRHvhJb+XljXu
gtGC3FB1TPeyiz35vP1fbyttVA9MdoQeOX62iNMzgDbEeoLqtVwTvW+kWekTf7efO9/zXn64TkSz
y3Po2QsxtHw3s05t/k4Lvr04I8gkFpW/FXrwNxWbnmXT4QoWF3VM2jcN8Hfn8s2zdHG7Za6XKZDU
wzqvmp/xKcGewCm0OqnwkzGbOejeTVYqt8lxpg6CyOY/f6IFlq0QCj7++3DydP6k9NvWjqtATPMZ
TNQqyxVRdMCydCp3LQ08SMsz+r64iy7wVDWChPVNOmE+TgW197ZqW6Ye99JWE46y2c6mpA3IA4lo
/5QiwynfYW2ejeb0AhkFfrBFkDfzUdmdlZlbj9hfLKA/ZDVg5wzUFzCOVGoec8Ye/gf5hzz6jVFg
xGBau3EpFe5Ie04ZdQLjxdWxgdj8NE5Zkbinx2csFRdN8BNseaSpZu3Oi2rwecSPaiUr6DuvLDm0
AxK41Cdim35NkKmI7p0mQZQX06aoF689NESlAGqPS+MSPYbooq0JGxnAqKXLbk97ZWxRRgry42zt
+02YL+ItGrFBkioN1wr0IK+g0EBiOt7lNh/1RQPAKKzD1gFu4GPtJJLIGq+JX2kh4lq7me+kkG6C
QeuQ4su4LQVETXCfNSYqz4LA304Hsx/YfLPTZb61pVZVyS8foYHtzf74HiBCW5zQvCLzxsHXq4zt
p7Im4+GuhXB9t6nFtHD06C57F/hWnkPmoB2W1JdT93BDuUKLau1mdpcR81e5Ay56yAF+DxKoH9Ck
gRP28ZGjuS+rt4ILu7w62370I062/5C7cUeW+ipAlABXU3wOiFz/FQQ7PW92N7Ud3HHR/Qz/Zxn8
5/H+pX1b8Ryrdhf61Yn6bjFW3giSPgimBecq4N6nxm79FqE//BAb3VJ2JNMiaZcq/u0aSS6YgtNf
g2LOLGYmBvlptAEqzFcWVgv4IAUy22WQK4Ak1+t79p/e+zgp13GWLBGCbueuyKpxxgjNH+Wi9vhL
ETpHMoeJoX/VyLLI4EFR2qubgHIJQIbzM3TwLz+WHfY7jWul6fkyA/jv371GcS6LVgoxUpS3dDLP
1AYMjVEEDYTrR6VPV062s6TJse96ZIprcDkcdLkMtWRAwILxfpzszV94uahSEXs0gRFfCMwxP3zT
QLjlVzHkPRe1euhxpGSqPA/9kWci5T8Y3x4N12im+MTrAuHoIrV7ENoEUW0aKkQhmE1u9TyIg7W3
sGBU+0or5Nc2IHOJ51vmGkQiRo0u4xUdGQPgIK9tyEYFOVM+H5bf2baI1YMpwZsp0mmJtWGiirfJ
WYi1Vpuomys579RTa8JC+ymLWwvr9jeGZ20DxFrVOanqmo65FcWsVVfty7qlZROvk3O0ur/CC8sc
PoGRVTVifZq7DmZk5oVffjxFEkwaccOY8v74UXJ6fFSVRksRmlDvLcOykC+qDBHpDLQ4IqnSF+jy
rZavv+FBiBsYZv079dFdmdLDij8XJHM/yjPUh1yoEN6DpORzDQR8G4PIRAeBF0BvR6Ed6Iy4aV3Q
v0obZt4fxa/zb50D5ceivhbVHnC01waGNa9hmZhkClX99EE5vxJ50FzAwa4PQ6GDGwV/oHMH/rBE
o9GfZ1+O8D3kcpYQ4fhQ2/Xzj55JxezayyKeLsTw18kPTE6wnr2+QPIVaCZy/fz6+HamA0fLpVH7
M3i1HVmH48t/SUV/qQAC/gDsy6QCL5omkVzAXX00Dj1mcKwdFRAMPFqvgIPsDD3tb1fJUFLjBgyz
9MClJY2i+OAVGHnPJIWy+UUc9FOrJpo4zG/RMQ1wZzToUIFRfg2U4pVoyhBevbx5qXF3akP8vfsP
LFAWmYCnmo4WNjaMRr3cOUGFpC40kIWaxPBfg/G90TLuOsg81qdOVWC8Gprhx/98K/nrcswQNwTw
kh4Cs45OXUN1lksBMbKzpbF+zhT4fwDwAR1197VueV7PtnJupveNQz/0ZvVd/ENfseje8am2HqbU
7OYo+Dbh9y3m9/DH+MvCVaQgbLYI3SzDVtM+0ZRaafUidVHn8h9jNRgtDH5W3hOTEwDoD8Ghbm21
Ycbr2bXTZ4PbZTkteU0yrCBNmKdppAGheSQG4+0cymtrnkspcIY0vIxJ4HKEWVyqGaoSInVEMfnn
pcfU8RE6hixJFK69aRpOJoDuGnxiEGAF/v1iIgyLFpnfgYITqDTgCuJihEabCIAje6a+u2Gw0/hL
qqG85VvwDXbQZKLGniSf2Sc033scLUI+h/7i6MfJj5tFKPbnOyRzSqRS49wGs9/TPmjFez6AlLKB
vtUXCXIP0tA4r7v9mvw4urTP1tCu/lsYCusmv4TVEzZvnkYkXB1MsaGVX6veH6BI8ts+QEGWtrWl
kt9kCasi35pQPsdxh6c4eBqZOONzBuT79dHtuyoZ+52Xf4f5gWMO8gXqKLp2R8USYhVcP7Yzq5GH
JZ00/TPPLjZvtJM7Dajra7C9I+yIgYNDdsDu8UIRcKmAawVb1U3kNAdQm7di81qevLblAWtoyJ6e
QWaoBcoEVwsBd3jXy3UnVNzPMPek/WuINGueZjgyX12Onc/ZSfuu9HrVb0b+SDY5mLvtafuxK1yr
phiNVPiqpt0+pIe1ZttIyKqEQe+9xElex/lZfQIQb29G54KmjTiBIu7MfyEE1WNvg6MjffGMnwm7
B8NZiK6nYE8KRM6e6gl7TaadyfVA7Fqugm+FwTuKl6sY7QGEEAQkRtukP6a+WJyfo2Q5V5wa8XM2
yE9Y0BAU1TSPZFVvk5s5GUPpGAf7BgMnQ9BKx0oIXxDVe7P6o+hVC95Y9ZhkuRl+sIr6D/A7Kzio
iJb05FGntiDcT2UVQb8CK1988cAlDui5sYQ61YUoCLM+op0+7/A+c0H9foR2a4uK4cjQApRWnWmC
vBLchHia7hDdRMh41Mnrj4tgpkSgUcAbeYzvgLSwqJPEu6h4RreQE4KK6XrK06rz5DQiMYuJ75NA
JBTDhMmOLGigkiM8cXefEsAQhTr+JXtkH1ayrHY0YJIgNghUrRQ7iBoqHrKnyqXNO/Icx5KAk2lE
xMLvujqNxdlHCeat4YvQcmRxGWnm0DPb2DlGKVneVhzDStOyGhJEWAn2z7+n4mGC0Lr8jmn/VdRY
HXn7X/RKGqukHPCMKnUx8FLa3Q/lrW3BH64TejTZk1W0dilwoV2xzQ99sxr0N4//F7n9fxG/MKP5
xLZ9Q5lcbEExJjRbPl2fHrczwGfgr7Ud3iRsBzSrqDeg0R3SK7Y2jCaEKjTy+5M1rhSP4PzvxveO
XealQgjF5W46UrN4YHp64+SCjAfiWj/Fm52X//K7fduBLfNmjL1pl5889kNPwuDliLX+ZwVQRgy5
tM3VKfqTATP/U5toFfh7f+PlqL3p5gW5PzOLJ+CAyJv4ap+t43Bx2S5grwYDPmhpvtsw7CIuc9MY
0WuboSaKWTh63ePbLFaEjdVovd8lsUMCjdEb53248ae1YEKkhkUevUrwyQ1Gx8VClSWW8gORTZsm
Ldn0s7MaK1+Rl4MHPp+L/yEs4/XtWbRaWK56wbD6JHDcyCjllE88kK44lyVpwLVvscgB2aLUGnRC
B7/VAzSli0XcDrJvb7lm0PQ50MEn+4HKxvKn8Gn9Cc50dhTDbcH0cFtVHL8AQo1EGh/oIcUYDObF
pe+Cul6xoTsTpU64sZyEXNQkJ7tuzcCkp7kAmLBEVnQOhKxFx8LTP66r0OCHTdVbSxBtv8erbLKa
nT1nQSa5fYi4Dj1i6lNhNq/6EdkwEehIJaiIrOJTAWSfNEYBl5Eb/Kdh8ueC5OZMBN2iY6EyTLQb
4Uhm+eNEjkPacOxj+kkVl+n6PWJKaN93wQNP9u0zP8FNlPd+KpapD4XvE2FUMzELjwLIIw2EWfUB
4ItbY8T7VYc99HsMF47k5QN8YCNySMN1a7wFfGKnaf0BX38kW4GRe/TQkJE3QQa4ekrdRGvXdWTy
DIjLMBd+JUfBTeyCnLgpV+yVhhloI7T2epzJlgbWuo3yZd28jDwaeIQ7tj2ayDwnU3RsSC+XJHM4
LLgt1C80Qbz8FoAVsN8sjoQSdt0EsdWL4F29FALj98zwmDwYo3+s21ojN/+uhDohh8pddsZ5w2aE
xnlN0UhU0xp8E7/uqfkx++Md0xlFLrhxHZ4DWtYMZbL5ewzuqOWvZWp7yXZQo8XQqGIyH72X1gfz
sJrznD4A1Fsm7oCgZqbxeF6PDsWYpryTnXa+/qPKNoKaCLR2ZlGjDBpZQy+LsAYQo17sGZVGZ3+1
1xV/1cdZ7wsRF5WqPO8RsfbZQivapLPT0rDfC+qOus1WvcPusk0FTiJcbCF/FDAVmX6yex/1EQoF
+sWv3fRioySetVC5syR3jsqEVHB5Vf0T7kOuHL6yQa9kQBgisS8IGevtpF2ABiMvh8ZruIOZ2jX6
QQ0kW+YBudjPezO4RRtQjPm6xEpv3dGsCCihX4qojePtGGw7G6/u1xNfFXm+tvRcNeHNx+ec25B+
mg32fI2Ld72tqf7Pls/k8gFU7wJ+msIceF8N2MOlOdbhE4PDljRlGsGkyt1/9jbkc4hc+Fm9+LI0
3Hba5GYeg7IhuQR12qykYV/tIOXISwixxG03aECZlCkyxbZH00CZGEquiwJ3IguthTSH6bp47sUD
uCGbQqbQoL/TR8iOJ+tmcZg1xAdQXabo/aQWZQsqWbZWsPcdGo9MxtNC+3ggGnHKHZSbwouWCrF3
2FmlG2KWlGMUoiSfBES4fmHu0nmxq9+YqdZTG/ovpAtTtElWpFT+zqEavPSn+o+Lasn48enVS7oJ
8yxqSVBZm1Cdrpww+BMNY87rl+lo9TSvt/4t8ZoJzNVNMwDaAUy9SgSsNzGe9QDxNgSGXNQTDivT
7FIz1bsTKE5c5x1Ht9FficM04MtLh53I694g6aw/18ellWi5Aj5VbYLOFCDzlgjQn8mROBnF0Orj
Frpc4G3ov6ACFTTBkebIQwBGz+IATEl96XyjUEmhOdtvNjMWQ/3r1TrtXWb1tgOaepF2B53iqiNf
2ix5BbzW8sob0SDxFJQxjlgE7PZcpI3LtwEWR9azgnLEIgVRXYZkOaqikNMeiCBFGsh7Kyl21BZ6
lj5zIag1kdZ399tXln7CnRPHP2EgAh0dOp7K5wiaTDhd8jBb/nl30eHGqcI/4aTjfyLENgVonxAo
XK78DjL7xDbKFn7e25/57BvUBAOwHH4qWiaqK9PiwrzkYXLA3+0wl7ddDtQYudvIXphyQXFEDFI2
hbsMe5dg3S68bV9mI4FopfdRxPSafKzxln+7YCZwWY1oRnBMe++nUI+MYr6j0Q2Tb8z+ZJFmKJXG
HOYHTSeKT37Oh0qx9vBlclVUrifjQRXeFHgW09ZLOjSfU7Qzgq4+/FmRuSAHyNPD3j0943nebwBQ
4J1GUKnqIIwv4vUaYW8Gu73s3Wr1weIyVvuVD42+2SvKt+78vmDo586mj5vACRgEatTo/ohxJyWQ
Vd+4D9d/WERuNVKVrBNHeD/rV5S2EF7dXwOAzxKrtZRqSIYWTbv58dMYC4jxUIP5xoH6UsEj2RXx
TO3dasJSTfLoO0PyHOW7atcT6NT9n3MOUTSHUo5dvjtXXSQLw3fiiU9R0jTrigtg2GXOyxr0tuMg
fRVLeximA+XK2gu5ACtVynzMClcogPMurJIODEEOc5ADK/9LYsER9r9q4F8rnfy2MqYl8fRXvgP+
AioyX3wKULK6uFK0h+6foFZT3zLdvbMPmvOUvXfS11bRNaB81JMBiGnHWlJrcV5bwRHFYduBbyBs
QUj9gCJOdbwhLjbUzrIJPGhO+gq+vrXZ1f2Ttvte/IzBqu0xN0hLwZ1N499egAwdsyFM0Yv00cjv
J0IG9alyfWlTw0zSSN61u9dnd8G4G6lQ4zRLQxzN9+jhy3FZzJTCSX568Yg/KSIk4K34mOtL/ZMU
xeW7m72j5HmDVWFg+1umr0aa+XLo9+cgMpji1HWAMiMSBIjkmbATKDl5t1LisPkbaKwCUTlb4s0y
6fPrLBLlBIWkQPI2+ZH++lq+oCP7W6s9Gtpn0wd6NuQHyx0NQ5Lf4QKyJ9AlG1j7fR0qwumCsDbE
copvy4rgc+yrAFfrxRKmFTXMoHyLbE1diFqr+8og2IXDtzvnoSKR3HgYaSS+yDtn45n4U2U+Qumi
+/Sl61WKPMglU28jX0FrslLr20p39pHM1vtRoQDB3Vbcv9w+Jj7FcUpyRDmYyYn0XTUGqZBNXqKH
IoT0/s4vmxwGRXbyii/EAp4stNnHR5cyyfLSQigEr6GSLMRY8ElE4eHaAhc5Nd1iYOwgNhAFPOEF
ZFcYI8CL9zPMrcgXzh9pp/0irUvIeK8jEZmhqSJj3NVSkzILjL4zo1Ur5vZLBtn3xC9jVzn4oiwR
hTR1VYMCm/hRasbLJvRxZOdAwU6E2ea3mxWigNMW2PQtCCyTaWerrdey4Gd/R/oDJnHHHoPcMOtN
XUusHQxG2Yu7f4fnqgsOrE4OmUz9T8jAq7YDb/KQDKP7JucfErrITlDI7+9PSqKj1PWPlcsyfHTN
6vPzIZJztSdO5utTpoyQv+3Ce/zMa/7dIeuK+4nlUkMxC82LZskSwDgyPr35Co0kBkaBuKw0MDbS
mV2Z9rfyKsYrdCBe36cuZcvAY5ydSo0TEB99i81a79Xb2ifJIkN05fL/JQUoI7s8URWbEFIpzNwl
Pvc+eXsKcc3LtqfQrJd/qnmJUT0DUtZ+nPSIFTYP1HGLzag9OtW8uunoU9IW1H77PC/kpVr06NLN
HN4nKEXbF9ohD4kct5ixIHWU6uynEA3Sz5C+WLGdI6q6XgGRs9FVf0Es/FNzbNbv60EGbK5g2SDS
SPlfUccWhvtIeC8taWLVQggjyT78Qu56JxHhqIZ8M+77Cp8VJqNID0dGy6djcF8Yp6jqJHaWPQ5C
bTS74lcKMx2HC6mCWQ5UUW58Ji/TJNQojUKpUIjWcIIlaZq5m0cWQUrEjLz4jKXpbHGoyjhq3/B8
+zgD65Vkzw3Xrg+FXH6g3QBV0ktsOYCR+FEHPTksVahWFh4zUWxMaBSeLd0aByuiOUW/SRcyIQAD
aIdw+h1r+ZSkb3Tg7CWPHYS1VaaiLIGinRoF9Bi+8HMDRF32aZFD3HDeoQxlFV/g+nRNFd1uZ3FF
jKKmp3r/adXVdIro1JDv7HJBN+SC1iIEZ+6lmMC3itrqzuHsdW664qc3JnpyDQt1c6j2Q8Evm6oV
ZOlXWU8kr7TYrDRdVgmaJSWqb2v0tfJcW/Kexbz7JIzpvP9w382DnMtm6FHPHMApa042uuniVgQ+
01Rujktm2wzevuT90iHizpiNiJSFgaXgDGpg0tku8VpYHWJJlTHfCla9D9JWcZu0C9dx9S5Q46xB
CTKgiSwPDniDKGDPAP0i9g/upB8AKdFf/ofxgmh/NmPGmRokp5yQJ+nBpX0tQQ83QdkMnxSJPhtR
XPD5I/KtyP0GUJS3j1MLItAqzoEWzieriVizFZQpv/nErA6RX36kmN7DC/n0Iife7jmKqBeKrzj5
PAG60jL93hAPfMjHw7N1GqHf4iC2GD0+MKZyzaYpuOnUjJ8oy6N94gANQNze4Sc1TDy2gMZLrIri
+FN+NBHPH+0dgYyngn08DxEPGKjvz7oqnMcRQPp6CUkQRxaR85pOhkJHUPTSAqNsEXNHGEKeOe+S
kv2HeMsQLjI1YRxCXXU6/abZETXGOVtPESGo0Il+JeU4Cv9BYEDsZA+bhsG+l9Iu17esMvEZnxdL
3spILWZqv37evq0FrFxuCxp6JzwVuMHCUlsuHuOfMKUlMeoEskSOenuvuFfV/rGuFlCFvKgxJRql
xl4rpB0OXQi15o4BYwOMbjM2Ag7ZnsM/vrYxrqIfa+Byn1qhDqsII7hVWA0Y+yuGsFerl6NeFSX6
8kNSWOwEWZ531YDgGleVjzM5ve8yVK0E9CST29QyMYaK6mTnGb7657ymLW0foZSJCgRI4TwBQ/eb
xZsQaNEdCCLFGz67e1LfC+Ug0wyBlqLVPrgXqup1paEm0wgcoe9PPrCyc2ExaOcrWd9Fz8gSlLeX
qakTH6Eo4/kXQAW0E69F+/mhX0SZ2GAtdduZIbRGTazqp1Sk3nWDODMzqc1fJYM07FxlvClMCMZb
1hQ3O/kl9bY869FiyJTzrcgBy8hz/U6n3upO3M4tZnW6wRdU1sPQKVcCsiNn2b+IKZ5Q6kUp83h1
rabZbP6u4mBe0HHDy6G8USwVtCkmehPAQmh96WNV1SSB1fPbJ+JpAIaa8UbhlvimBTLgfJBwsJf5
Onm/24FE5e9AWWlPYJaqV84rt3e1QCbDnFrnVHWKQ4/HreEn6noWlcjJN+gZEMKCMIt1PkSONFQu
GaaFe3QyAiGY+cOD5fe0ZL6ZMY1lgREwa+omQu+O8ScgTCx1/Km8MICq87S+EXUZZw7qdAvLHhIj
8QnYfV5boSMCMOrPnJrDBK3ehPWSKNuxTF2RU3kcMslg8oGynLtP5gY/5TzSMjg+ZficZAVsGg5r
n65gYKNqTwL4HCQOmKZRCfnJ3rFywjKcb2Fu69/A1U1f+NVojW7g5VNYv+hOkNBSgKq8cYkP0wd7
7rNO7J42dBBBEYk59Gx7A04/gZiyb15De4DH9G5ToFPgU4PeeOPAEvfn0/hyQ7jkZ0qhEG36qV2t
nZmz1HfVpb9M43htHLaGwcdvAtjkL+V3u/EI1oO/Lg6Gn6fYDuan6pBcQpfZCX9DUDXcecEV2LAG
ASpYJ+JM/t0S626WQT8f3PdgSHYjcD2XGUvEUoEGrZ3Q5IQrgeYMmE2NsxZiOrjNWMCPplSBwuqM
+yXukrmmPegCENYv9Ta/R/Ig9qeYE9B83lxh6Rx7tz17Ap6btG4DlckU8+W3jD8GCH9j2sx41LNG
OFgw7nOJobqzPJnD0Iorce9UlFCjuIZlbST4Ec8OLcuGI543Y++/4wvdC0F03mFpdLxlxfCIPcIT
7j05dkQCEUlDWAEPaCZManllLNOArFAA7pRvLPyxAtirJ/RtcTeiTwOVgrl2Sc9yZZk42xJeD0Rj
OFV3/ibrxV0KzNohloLK/Ld/hI01CyZlnQ8TEDu2/whkeNg5vfT8rHvYlMAB4yr41D8YSgOGoAkN
1+A988HoOiUrwkKrw1lolNxev5HDKzNe9OiZpNGLlx2k0wgewl7udpMMCVdn6NQ/frRzK2tkJ5xX
CAVJv+KU5fYr9L0sWy67F+C15V+EP2/P3XAcLAskwHvJzQC4ovjjt1B1ZS61/9pjWylJavB5PAxd
xzX8YEvIa6Vo6AAFkdedCgI8taTh4uHmMIByJ1It6ByOF6CAmwm97UCzEk0Tq0slshsFxlE9QZ5r
Izf3pc1W4iFjfxoU7hGg78pJ0yWwhsPpfZE1WnhS88sBAZS5nO/7kIROh/O4HI2cZr8AXMLTXJ3I
aUsUb1dmORQn5R+FLDMVW84KWs7ERybk+9yKslewxw3C+MfR1wG2PFV1NRyeDcjKrI2kDeppOomQ
9bAnxVDLlSiEdbwiXmpcvynpHZ4KMKbLsRPz1TOtQAJvmCCGgx8y8IF3CSr1Xbf5FnT+u2s8mZIB
7u6LsAFokS6KUbeMqlATcQEpEZ0uwvXS4DgnraZxxwFZkl9pknctmvSxeQdz0j5Mi5KWYgSdfMzS
sjLnGqEnZ2u+UvILU5kxZ2QYIjcimL4ZZQo4o7i2anDeKXkzAtjfeudGWqJG6QImWAmysNg4ddkR
30epn/ovgOXGHChp7l00DoQkp/vqIH6xVCbc3adelxvJCX2Okri3cV0XK9jgF6dcOy+w+Q6q1ZE6
Md9XBgn3FwMmuNiOGmWbarb/AOXSnbZO70lJWyGQ80U2vo/TkiIjNipJY4vbn/R4FeXvFZFMv23e
akLrqS3dxovU2ZnPY61HLXWTdfyHBaBYPmDN1/5gf9H5wbtIjhKIQB3p7hCyjBb6ZmNtuGuFJhkP
6CJAdFAOYL2nIfjDteeglGRAPkaSG3Gh18rkEdcJ0FXsaT4pm6Kc3/+uJymoAR5yzLaL6dSpDQ1r
/RA8JYtwYxCM7yTQMyAHp6X6cgaYjJVi/08RqUH0yMxm/dfC7qac1zsT1Wjcuv37F1A0ewsMgd2V
5v7DzL5v9b/iSTdYWgY3i5j95LzHjwSIJA0L2LNKXr8HqTQeC+ZZ1+OsKooxkv2l5LbJI2ElSgQu
crT/N/5DvMrV1bNdoUYbPcIWZqPX3cTj010wq+afQgdh2kuKVYDFHz+89LaJd+08InPjQ3JSZ7oN
E5r8YnnniUZKZ0XNm6XHGwYXY6eEALiMzQTSRup444nvDA19Bu2UECQ2MWoEkhHk7rPt+OOdwBvF
pjSmV6jNOyuE+oBKJWZAsVZBsvituBpBvMiP/NONWOkV6QbUgIqRMUuQInyDp4138qrqKUKlXcOk
P2cfytyPxSns5bU2+q3NNebE6c995KEP429VRq8cTCuRfNoxv00XFvqX3M9PMWxRTLb9uSUAb1xb
CVsnRdsDCDTn891etzVyqZO8cS1KLwPdzK3Tn0UBIhmKg+V4EM/C/T13ITk17TOnqqV7SxvJfBzX
ke7a1qJtCNLMcLDtx6IJYFa14oBWOGkamuEDIxIoSGcJKtsk+5kmJ9J0IYXei8KLOzuio1s8p8EG
9ClD5EQKrfO0b6cr7E7o2RSjjPHzWN10g/w8dTzHvetqnXtbHFHRvbL7qSNxqiHBNPQP8CkxJATy
79UWqv5hNIJQgHpHOw2FDlUsrBhCQZXHruamyvVKN9WmiH0ZPi2qYJIXwU+S+pjZ6FGLerKLF1W3
9ASJeRO/tZ6KInAn7Xn4O+VCEb4DgNWhmLiRKstBn0PNMH/hK+PBIML75ZjDth964ooSYmZIC8Rv
ZINcMF+oiuU1qFh9tW8bueNEg6qDH/gBUcTWKvtHg6WXfOycgysY8Nmp2QWEanGdPLFg4PTk9dQI
P+lc2jIRJjFJTvuPlUIns7/NWsVT5sb6RJf8NlV6JmlWsaxHZit/xu9BkM4Q4AW4lueOSEwJmh5n
BOct3KvEIFrVJ142Fpm4L8dstuZXXtPCHyBSoQjOkifXMTyngSHQTuyN4J3jjpf/BNi1qFdr2TWq
c27oiwy4phZZ42xUCuvYJCiKsTefG+VC9cC6ELnL/oomHxEewE1Uih2LmeNv0nRo0elDJGj3DHOz
ltOxBSzTJ/D0XXTYBYZi7lqyMoxj9hyEQ6wg0wJsPX/hsTqy/I1NA20dtQBR1qijBkCXDI/LjgRa
f2U8K5BvJpUzCYAqVGvypt9HdhUD/hBR6dbmHq06WLnkKS8cdBLVrgsDI9qA2Naxc1G4CQCypeHd
Xx/rHMTiQoA2cFUkalXiBba4olbg1/Y7Ztm3bsVEcL6Z3CT+8yhPxMhV3MBLDHg7/QEpFr5CnKSY
XUY7gaxkucO9d2qV2MapTbqu0vtdxmqb8Emb0POI+NQ7qE0f+/vA9j5IeKRQG0E+irA3y7/QBknl
w9DAGS+DS0b9WvlWqsfRAvZ+Unh4/cu7S4vlL05GOh4Tq5SJ31b342V80PNZvSUGFwxuGYJK7Q8Z
xnCnY3jsoWunX2rARZZiXuhyxekQuKQG5r2DIcSFIXnx/LQHZN+KbIkYtvsqtaSC2JZKOPSC8eef
Sle51K4MVnTOgDbv7GejgH9MLAGVSsQLWJsvl86tLrWPONZoPS7KE9m/czvIh7FgCuht78nE9Q4k
Z97IJZ20tg6cKpqJAhmgesmDB4i7URbFq1e+GUOMkhX4ZlM063V9zN5Z9ZjOUbPxwknkYci1Ys9R
R/mEiifKBspLB6zG1JZspkASQGDgcnBbp7WYHPSFCHuGEPyxdvLwLZBbKwpE1QQ7s746PjgeGFOQ
Q8cWRQnI6Zyih4ZVmfdppCOHfJi5AvBhLi44ddpTo2sl9hnI3/KG+cehg1I5iTzACMSxrNK9II7B
Tm7xiIEssBnvqViQUCdiqSsxjp71NNzJHI/Qi/8c2R9doo9FMfYm3cm2XcOSPZVTelaq8Fx2uOZO
lxa+aD14pzIs6tLHfB5nNSOTpBXP7mCoqngxsiQAegxnH0nBcORvkHNiMnhTYR1YSkNNd6c+dqci
Fm3Pq94tNdxaEtREaOB4KE0uri8c56iEFdDMzJQKca5+r5WL+bgvKcS9bxp2faUB0u3cNi/XOBYG
tBmFYg2VYFdotSeh8Y+K9pJG2oaK6iN+4WnDVu43KxZTTcFhZFreYHtDqWPfe6huHlHDr02juR+8
Va/SecEtPo1EOxh2zYvRKSUqndffnlmNk/elJiMrv1p+Y3UfwPMTPNeo+R/v9CJ4OoJff9B1+cMw
hdIulnEgS2d9lek2n8Kk+kB4K6f4zDU6qpW/8IxHit5dZpHZnOeJ1xhJbKgG2v+ad5nlLwU3dqlq
7mzALCeEa2EUn0ker4RWT5x6TyuBpo4PvudKfyCGcyLZrJqXNzsIQEWL5Zkj2yGRQOzLvfkhbzIT
D3gF7ssUmw1/L3Z2XxZ7M5CYdLVZgo577EWTrJ3mJNK72AsroLVqopUttroYkr0p4gtdF3J7Nm1o
/KfaQyu6xBOYWKaScfueTj/ak9YsnZBgXO/Wp+KqbJV2Cwwt2YsTywykJ8EopGcBr5qnRXdkLB4Q
qLvSmmr08zMq0eFKNHFQyMI/VQOl2oT+hgylAbCCHiRWKnI0ekal/iY7+sDosY+LVYQRw7smyHbE
CnP6APIKT48QdvGBtn53v6qoW3rOc5Et9zmqAWu2nJ2SCyEKuAqe4wOEcOuqQyvtZoWt9QiFzKbH
CCNni2b5igSG8I1JPvl1QG8Q+rYRUdd/27nziaP/FMzsI1Gro8DzYQT0ZDLpjIhMElHk6fvY/a8E
Z3fG8YHNVZxs1hVlkn0/3X9pCOyhAeIfr4jBtFxLyZ79R5qBQ7fORp8WS1/HO3dNJ+VlbD9QhFwC
SmH71zbsCnp3yJtFE1WCg64xGSXB2FU/MZb8EYVOHMbNmjiHiIeFlNIyCCaqzq9Pt/rzkeveDLpI
NZ2mm8B/JTL5KY++eAy7ZQgDIcBj3RtFPAT18br0c20U1axExljpMUJ6xNkiKgbCPxDj3Yi8Kzso
ECixIU/YbLH1k9qnbkJF+fZ22xkRhJKsnq1/gZ0JgGS9/cuEnbLAcuRbuyMUk4TUQY5YLfz91PL9
N/A3S3Ux972vHVSOHstC6VDeEcTZY8Uao7nGT3+Osilfc7svhYEHJDbw3voiqS39j4+w4GyLWVgs
be6/ywXinBBARSINbJQEDM6Ji+OOhFSEQu8cG2nxtCBdH7UNegVpL6DTrD849BVEIv1SPnRUztHf
s0VgUbRa9Z5g7EVatO5aYQq2ZGsy2t5YMk8knQKdg5NA+pHUgCGiHOiS4VrYw8U+w/FkuWPY1s/A
sIcrxQywVj7llEg4hTwwdcxSJ5kpTDDQUjjJ9Gia2u8TGup21iuTECC92QTCgA/fhi2FTslJ6MAd
2sLnhKNjsR6EQ5JXVUiWici7xvaFBuguD/cJKxPVrXIBCis/dgq6yBhtH31ziITozxGKDYMqCATU
WeDxiawHQa2NCCh8zPl/COYJ8z851CkjTl2HjD0T8GvQbslgi2ABzmTZnr6xZrnFyZvrH5OhW2D3
WBQM+efZBQuPT79Sa1V8sHuCe8HqVZWK4qGnnNLABhvhpR1qWyyAyadkTSC6Wo7lWagKl7qT9ceS
Y2LIjBO1fPgJ57RYzJxAdXl0f+tve/oi241kBbHAnncrKzJUjD9UjFhrfEVVHZCzICzSg/QAfb7H
Jf3HQEIK3FrPM8TzCp2nQ5yk/Sf+CIB8EnFHTizOsOVoLDbv9aKzq4ZSNbZG6HBdBOWWf4QJAmTC
OQXO3NbMtVH3RN4vpkpziEGjK2JcJmODuc10GHp8z1G3Y8sge8Ch/pYExpx9a5mA8tJ0b+n9Hfnq
NWvVPYBzoGmuc/4IpQ53SBM4Ew0SIB7AjxMws8SUl4EALh8D4XpOGDdXxlfyoKSP0g2iGuUI0ylt
YMsK1iw333YW68cW2fQlQaqEBtODr402k8Yls5mIQVATB43LGjbBF0RLBC+h/9UVhqY8kz/yLzLA
cbyZCY0ncb0NPI3YDZ8RsGqPQ4yXXjMzK6/FFWtXAY0MuX+T96mrbCje7CgeHfS+TLadOrfnBsY9
wITNEbl+PsUi8hsK5mzu49MAbQiWkq9OPse/ejOWhpGAjUfRbayihfNARRRdTGAE1OIp8LgOPkUT
+Gd878Vk8vCFKkdrBvKjsnJMps9u/lX26zZBt8+wL8Yuul9WK9Dn62a+kqfKcGXCwrUIVTdT8hIe
1/l+ULMaVLL5CBgmpmSwpn1bnPKa2HQ1w2B6vJ26WaB6xplVjcFLgG0usnad7NwOGXmFm2F9hWRm
S/22zSL8ZsF7CzMvXqXO7vkdqBib8nVl51u2Ddk+qoJVojqUy0Ikt2qcS6wGeOPCeYIDyEkFcMC1
Oknvz27AOIDOOiLXstighyLHnYcMpt/QdYkWfYykrgxia48JFhGZySXuqiiOESTibYVzkCkUkeT4
nhXnYnQlgnGpsSfQkENLktIlgaXQaucFmx9aen1cRkPAcsZ6s334NW+icpus923Rk0m++H9uMQR8
vp1+25ZeKrlM6fikRjM1J1z7qS9krElIk3YNzSFkY1yheyaAXfqsITBy60Rh0JhIVsrpMWSgWYVG
j5c7Y0eMqdQodii3z5p0ibUcavRGHsB4KKgLIIzEuZRQvWpeVtawtO+VpOrboxtqeJGEXlTL6HEk
FIU91dOI/Z0z8XlDNQS17Cjdjjxm+u4jzgRSf3I/Cis3zgncCy3pAGZqvQW97JzWtAqLZx645NjH
4yMNek5Yv7c6U+nFZxkRPewNuwtjr8e01rGBo+TO1POFieKnWtqcIJUQbFaOBf//kKKetxlImSQn
AwANKx45FG5kqTzefH7+78c3ibENTEnmQY5JQrPMNM9tJFKGzdFw+/jn0d8RH2VrEWOMD5gBNmed
j/Q8kQAiy1ShrFGQ4MfKGqJZw3PBsAKY43juDTrCDZC7RdJXiO7JyYp0cxSttGrx63EazyStuThc
3eJTeT0Yq32DhBURC5VlJh9T65IHwsc7IO19v+kyUeZJUtxK6DuwcckkHXfjmeEzBlXxr10/8Dm4
nZTj16FKQlG7hKs3csqe/TElq4qGcQwL8jhUVStc8L2v7FufRXjv3djq5eaAUKM6bG63AQK0S3Yj
Sx0v7OiT7/LijKlWJ8TGdRhfOp2sb/ofPgthm5VXMkYWEIyuRJF2sSPnSDPS+rCjSXg6stAqlghN
ULgHpQWRxFtwyg0zK9BhAV5SA1p2Dnahnub17+1dK4ftUkMQnl0t1cGKkKgcrdkt6tRjN+KG3ahQ
ur+AbGyRKAALSMchhb2S9iFh5JSHZz06FRogWASNNALVOWeWrhrRC5D6FiswRwXTGW4A5iBeE3IV
in1vnK81zg2Oj35qjWDb7jO9Jd7LiF+Ubf6rrBqJhC2rPpFuL/UdQ2K/ahqE3UexYvFklFzt51eh
h/5fjoRYsLq7trkc8NwcXlwcortnrnM5QOvW/al/FZbJe9WgK9SknFJJKpcK6QtS9fQOH27bNZTW
oPZZl0jM4xVuuN9El00cjS09oJjjCJstNBNPU32tCgPSO229yLKbgCMIjjtaDg5r4NXTf43/y7hK
aetOGOa9TI02VeqVsFaq9KrtHJNhCTOWUNqru6sJ6n24gn/SG9oo2ixK8NfNBPWeg88+BxcM2DUI
fM4fyrcsEoETarqyNRwpNGKtAMwINpPNmQT0CNBvzfUoyqD0xkD1ayGEnGNOk7f+lKvSrvJMroZJ
OBWEwkO6NQEJ4OS61QZldUd/Guj3rfAXBgK53xoNspXdmKQxiasfTdx6nsI1VkW4uMVfATzOuwFC
58bjnwQpvaNH/n0AGWvDsofX7+6QJYlkSYWBLxja3vrDGMV/KMZv9TivnV5bHqcz1p+T5c6PatwU
Mu9WnjBSYpO8OQUYoE1jsMyyq53it0TFL/fnmPUyzhtYqCLFIM/Q05g5Rmazdzn0l+mZ9BQENGiI
GAri2r97Yx/m6yoUQouZ9qcvefM/AAKy6SnSuRZWDCSCtVO3e/yI0554sOPyRbMEZiOT0coo9erv
qzR7T2DcaYQ5PKWPgr+1QXGXYiIcCyKP3zRWcP4ZYbZKJrYwopaChZwYtXEJjmTG4/0A07QkpHyQ
P1cBgP9eHNXAn4p4e9d54WaG0htSq2BQPVbWTCipf4nmN72kP1Unm8mjdx3SKT7050fu9b5xq4qP
kVCbhdGmN4RlkUtcFsKzzhBg1mLXv75wVSqoylg9wSNaxFfD4wuTqQHTp7rts9ldHUCHRIQuhxhI
oWZYELvXXqV6t6vpIyB/CxkN7bvzcIwji4yBsZQyT6KkKgZJstOcxg8BePonryWbGx5tF5fAiWjr
i8Hbmo+p694Tj5SJ9pXyDE5L3iasohx/8KufLAEjB6ECEUvulUd+ouL7k88Y4nNAo+4hoPAk91Zh
a9ZC5qGegvoz/VO/wq2Xy7mx9i+U8/RaCwT8UMXcNvDcz/1u3OEA6FxpjvmCZv0h7CCNicl6N2Ye
kGW9xEi2fmSB/t9QTaLF/D9knBufDYBlrlMMtt8FuIxPVC5i1GHAUP3X62lGITy+uIoDKL0TVwrL
DVvPA0Z2IgRST16vqrm7Ehz03J0hniHvHIK48iCt6uYm70rjMVq5nq8bnfQQBsz6M54lg2tbMddE
oXgQp5XNDyN+XC3+JVS2RCgEUSRTtkPatj6d/VSILDNCN2WruIAMmHSTPQL3yEY0EjTc0T+ONSiI
UcLExfR5atdDtt6jHDgUUPICCOXF1ahMBtsPFj4BQRqNA0UFNZ/1kzawUg7eZ4PC0HmVeXlQaUD6
ad3OtTLVzETh2wGef27vG6DVd8CocyckjV8EL03aSTakRq3lZeXPdZ0/c0S0PyCx53+gAQTOttf7
7lSqAEVUGc8cIhj5/K1ghaQbWCn4FEBJgHaEoCNNs7+WGfKb1iG22iSw7Rm2Ufp5JUKCYTyg0NaE
RyZdo0LTJ+7gTxWTSNwHffySfv3DHEtqg0z4Pz7LOLeWk0CiLvUVQQp4lJS7LrQndfseFu0XiPTQ
lfpUV+fxi6w6G6jSGWcBvZvkG29bWYyuwuLmtfoxypckpGdPEOo2VQdQfh5NSgUrTdpLieOoYCBM
4+MWHOmgUaEiPuRTW2kY/2BBoaUGMUFMmEphAnFE53tsr/5p4GbuPudvBxSqa0+7ywVnNqhT9VSs
2oaHJTESwCq/zYN5eHbTK1/pZzWGeaW2xXviUHBDrCV9wK0r4r4dZK1xgaZo20huUuau5R6qiPhh
d8tIoaOa5cU+7KqpqsKdFZQUcLiREQ8+tDLr6E2gzv8CDLVyJpaaMi6P0pDKnbxXEU6tE8t7v1XG
R/6Amu5RfdyJ4Cu8EiNF69uDL7IQGOhMYpRxE08V+VrplhRLgjyhqL0Y75d59V4mSEHfyIQESakM
kGVh4rwANPrTb9phEcqAXOFfmLkqheCR6pJW9yz8sdAS9Qbckd8gRH3ld6KYk2hp2WrP2EEqg6Hs
bdxyzWFqMpZE68ArpQtB4vAUjLup4Eccu7pCb9bmd5pEeC5Enkhmt0dM1IzAe0XhOOITYCm0R0rI
irl/AasecSK0QU8YhNOCFNfwKSq9kAgoFGOzvgQXJLU87p86CQlUMNFVdqibV1e72fyyM8/aTG6W
GF77HvCFd/JcbqCt8+7l+ScCmZjtlkcn79MZs+3boC4Rrpww+igcHtCYDblrfPZ/RB9AbaA0/FHU
AydCZUgJ183R8V3hYAtPDzIQztWKoskOBVsw60O9Nfn/6F/rre2tzzkeXD5ayuwWZEKCv2uGqK7y
2bNIQ4SM4wTK8sm08/aVHnXqmFxcPaEg5FOfXbl+lrLB4LmmfZ6khlu/ilKl63PEPVd6JYYaVhQ3
/QGuGXjWqsLVRkzZsYX28LASLuq9x1nmItlL6OFb4SO9AoSz5kCmgcN5pb3nR3/ex+WX5GqvWeYR
h5hoCt3pL9DJG9hdYbK7QtLk9X98W02zpATU2i2LFqQTAjHO1BkgqqkaQGwr2sWnhwRRIjRa/LDl
Ve5jFWey3u/zx8d+P8GPewkW5ldTzRhk1pgdpw6qNlPIPVo5t75BdVQrFqB2Cx+Ixb1yWF3Uf+Oj
RSqyEWVttorQr4215d72pcEXSB616+bqbCJqmhbMawrPRCmxzKtmidna6Yvz8HNx3pAq9gRhz//5
rp8/rlQmJ9CR9tlfgOVD7zAXLQFrQ5JSPXQau45IBCJ6sJ5cVEZiDaB3SrsQ4yOaIWl/33Du+LsT
wkVhYz6nyEMljDVGZj9hDLTH+ejagMmh2bE1bF2M+hs79t+nDN2Dg8RxYPyYc8fokqJ6GzdY4ujn
EslXen3kvVGgymXWNNTZuarxSGkFL4xsQRvkXAH4IkqgROO6+/XNsDcj/fKQzb9s+O98nLYwLd6t
94nTzHNB0odDX39+9E+CjcTxLBMr5cWDZRscVAEzGWLXtU660wH2tZzM2QXZkk2+EVQd3Tl9s0/Z
nbKqM/U21fEB/pt0fGyLLZaQFg736/DlutxXWkDzm80MZiiCLFDV1UU/TLcjLz80shQlX9cpeFE6
IfYNKFIp7TydwqMSHZAbpZoN17lqFBX8paDJgN1dzJJjfKqPKjuRlstLeKWeAo1ec6Jz1YAyY/Db
PVZkH46pTprRqj7eDYoSxQ/LfjuAZAYeq9AKM59sLOdn0iPSO+goass+Vp5dUaPkpObbF9+ynK0k
ykDzIXQmk7QqEXafmsMh7RbwV5qg6CTHD+VvUyplRVdKgP4muEdfLgZB53UzIsXiaXN77Rw8v80l
n1DGF1gLSVnj7r34X7mHL3+4yuKh+2EElr6bJbSVUP+OJ85OnBlR1A0kymQIUEDYqOgBkaCftoK6
ZY44MA5kSHuY6EH7L2OT5L6iTdBJgAPKaiOb9uNNJ3k+5Ru+shNRrDpK3CapKVJ/Y2N1fdJEHGJ1
IUUbr8W2oIg1N4cmj80P0kUd2HpQV6wLbBUEg+QbMl8+57+fe66xMjf1oPg5Dhu9UuzGXvM8ldrf
VNK55uLp+jOvJWTOO1PQ20mfcxDUDrykj72UDxTB/Pdw32KWwMTgWgm4svyqbjjYGKR8cfG0oB+a
i08aMELoG5tKwElRAk68YGtpXJKcGbUNINfv82JwWNsEjXI5x403cKuByGZpzSW5tK1d3ABvBSe5
oudn6KsB8y+8KNkobeapGIuOzl3/EUt/hslUm8ymluymsqE4nwSVgAIy1bvIzEFUknrtdRBKiQEh
Tp+m1h3/rmxrH08V5nYgxG7G5AOQyu7PFTuxpjC6bm/LiKDQYCI+OM/dSw5zIAMq869II+sRnmix
8kp5T8v2T6uz9cMstMpUYB4ENGj0FxZQF+XWQ9wVCRQzIlAJeQ8Bbq3loBsTdzcT+5nRSdP8BPmj
ldq0D2wgaz9ePoebZ8uR0th0giCwlKp592ihly2XMgOPvsaKfwWX+xWan/C9pxLLil7nNgw3yo/M
JRx4jwGky8lHKUv4xBbZjzJHrSGuctKGnNnxWHQXxg0ynNyZTsXbbQ0yxom1bniWOQKiQwv8Zlw5
eQjbSB2QEMNYB6P1yE+H4bGTHYbo1I37lFzuvg/lQrETU94slJVhywmAsAXbSlJqCDS4iaQlGkLm
Z50hPgMyUDfRbwz3mgH4x8OC6dxVeY0HzIoa0KVSChZM7GH8/R4qWEhXqbk5NP2coplV5dID7TE3
lMcweTE4mR7oJV+5FBijS5flVQBAtFcmUA5ncSvYUbiqtZl9nkcWXh09eqZhbx1fZ8qqInsNXNis
J4i6g1DHIR9u7hGYnrF5qzQ0ptFky947wB22NpoR8D0CJIQ/AxfFd0lKAZxNa1meOWBzPLqMOPQU
MUKjXxSUrbBkq1g9I4BEXcB9yMHQ0KHTurY8FCEqhjRdq3ntBKcxsZ8A7AYVcw9RTfVXo08a8L01
19FAbGDQqU0TbEZ5uKCo28tbM8vhpoi+xL3OvuQyjerUKJwA8NgntelnbHF/lKS+Tw9h8WdLDH3a
hcGwakLVYGKzzCV0A3PlN5/7Y9pbBvLYNOsI2i9S8MKHZaeLDNSGRZzQ8QlvVV3RZDs9QuwpeTBj
IoLHQ3P3yoFJkSjPKJ9WDHYpk3KSFg1HTpJV4ZbchreMCX5Eu5h5WJKbQUjLvCm5SNfon9aPcya2
+Cv+ZmKSwNFyNxGxRWjItLSsAAEXm1m1cghGMtRlHuiilcwpxnuaX1yc+enXm5ZGAlQz9xXm/5dh
fhn3UYMR7e8RO9zTGGiQu6oWL0WMt1HXVgxFLx5bbEtRqTxMb5mhQoLiDl6A26rmssNc4qoBdaQN
vJuODg/93QSXLOd3UOYv3X12kj65UyQwCoGqPlXiD7OkAU4F37zFGcg7qEyzPsZmVTmAiOqGNYeW
/YaJBpEm8s7PBaFwbsMhiVPClhDcamQ7lfYx9ofdMkW0FlaZVpMkaEAaXqTyQDfVXkWvnIB5Sp9w
6uPkA/YNjF9PI6ZFFPLDbWU6cLE/3gSxJxu59dvS4dxBNJSpqllvLjxvZagHK7Zu/iHwtr4FK9Ds
UEJhp1NyX5yu24eAKEXxsR3XHxEbt/rLF2Isi9MWtlg6mpma6d9hrp5qrNBlCJp4NDAPtNu4KZbc
k0UYpTp7cRfGUm7Kn3CDZZj52GG7hQ1a5v5HfNX47h+7292d5jz8SQ3lhI4q9rTK7jtaE0MFPmiv
KnNgxEnBSiIUq1Ji7Tk0reQILDTCOryb1lSW1jnoISQmxeVm6WdyV0RDYYoXl9MM/kXV9W8blFUC
eGa2fVYPOHn/G+tukXxVPvmaqUctuyETxfgfbPNofNQQ1lC0j8Ni0u3Wn4hTUR9IrKv663mdmNl+
idynfvrShhC7XV6VFwibL/3JY7XoSuv8o7n5/NemZmCDgC9QnuBOwjYaqyj4QlythfOJ1gLWHE+3
MkpOxXfO9jKNlNPKGL8ZkdmZkXBzNH48by8+ExFcluHwhKYeF5yzReXsWR3e/Y7vODm3SjKxEK39
IPgKKds7hKgOg71dfYTx8wCRxm1nO0zpLFs2kQVgqKh00xQociEP+A0TcSVJrfDTiX2ULeUADBJQ
BQXV/keW9NqTppLAg8F0kHncz3N7RLJBTi/PNnn4wTApUsTwEv/XWq/o5LfV+iAbgSPjsUL0moqy
fnpwk3sLR7wgTCHb7SSYgLrCZNpmsDrv8rJhw4T8KDm0XDu39CXAWP8ya6G1FPfuqqw1sl8Z6+x9
uk/KuKiw7CJKdf7qQHNXcRKW72SfYQcpJnbLOMCseGqtVQ0N2q3E12Cv7ObXNLULsED4V2M1XhUV
Q0kooGMA0XpGRUDLU8Qh2fv+wvNonHPKcQCXj6j9FRAHQEJkeybT510HATsKEtwQIVbssgcxQRLi
rn5kRL5UFRNrUbhUrvGiv8VG+yIMpoeSg6yHpbDEM6zsHac+nWOvYasbho4MZgeVSNtEvZOAW3l3
5/Y9tdFJNP6jL/FxdF+IgzYzIYBhiYvtnkNXdJcXLIsdnrhrsWAN2mWpzFHusSA5pyn92Eo19hjV
YJUnWxLMjrg9nrxCPQxGQrkwo3XtK18c/l6LMzFeYst9Gbu8QZajaJ+Xp6JFbjwZHtI2a0HjgGM8
ey5pBmwpgIUFrCfGYrmUsFSr6xfRbicds2aLQwDUbLxLZMliVgkrQZeFhtf6hQs/3El176J0syKy
vAjrW5cqUSlGL7SRtG7xbdBcpQwdnV4K0jVMjlJndmO/0KZ/saGjMa0K4D+t7iwQjXVR8mmtcRiG
oeOgPAwqYAR0OVQbDDh+4lVrK0H5eSERDu+Xy8Nv/Dr+2yMnG7pWUOGMD5SZjepD+i8noBPrWc81
rItf05ZvYj8/I8CiXwz7olq2JdD2NyBsFavlvj6GxVdpYfDzQfdN0BEJctU0GPbpM2lD6Orsr2qi
kkfdXSRkNzcYs2o5xdLFcYeNwGCknmBzA4vZ8cZ5PO2n2o3FdlvKew0riQ1rDGHhrj8HdmMkpohr
c30WDsu+OQ95ubJF9PM2nhJV/nYboCWu5PyMt9UEChtgKuQNSRAX7kJ30e8z9ahhl0L8PzUFaTgD
5OA85+2PlPaeMSAa+VkiTX7eu3/45+beL7AX6lJcQYYJckS8zeQKyyzEVa5Wp8jBTBZVcL5Ooymb
F+5JfCKd/f8S3Qc+sEu929oOnio29sIyTyGVJUu72rzJ7A3IoWaVeQteIzIi1+U+GaWj9542Pc6R
m56eRASIOCoKyXV8kJH/Fquls07EWfv+3onhf5PaDgHwbk401jW1nBkHUZdisAAcFjReYI7BOSI8
Sqh6mqndy3hjtiY+9S+yY0Rg+4IZvsyNRpTIRZuS4lBQvhdDCSujlTXvcTCmeJbNmjdXGvaSrRYT
GwYn1mplaFj+AqsqAmVjgX4a2lpnNsu5HjrFFH2UYRnewJm1chahyLJCR8CdLNnhou6ZpglXjq2S
cDC+HVFIsBcN/TZx3sHSy7Dq9sjbIPEx9oc4Ym+n4goL8ZQ1zHEZuT6v7xRFWC9C8E6F/dBOQjE1
9FyZfUtluYtcqGEFM1w5FtY5rypnyJtxQiM2e2ba9J4pJ0MuoKZJOpNTlR2EX1lzmtb+urL+bjur
jJPJCFeDeUKG8oDvU3MEg4cuSjruZZJF1G5sRZm7GvzCpmFjQUqFyrtPeZ7i/tYOpzOkdiEmPdcP
roqwZ3m3AkA4jYLJtEhHrdokZjUS9nq9exVV+MNZgr53v9vO9SMh2vWKJQk8zcIlbPBQFuSVyPV6
tk4/yNEOFqnx2+81mKmKWHEfmZKkHVOX0kW/Jkvh4h0yIbV39iQMD4C69tqdMy1ybjAM4D+k2qRL
0Z4jSr+UwFiJcORdsQcaF42X/J0fCKnXk404SPk+NUQAGQFl5ayix1Z47bMuk/yirjCfkpUCpgjF
pOZ1IQ91KLxx8y+KOra1CeQZdaFfk4P3vqb/PTCLBPxNfkORIbuth7mFyPJ8MIccFp39Y/xU97Hc
sMzJlKWH5nGzasWWT6kbvMXQpKhLmZRKkpduq4GZV7LPoTgY74U3c932FJ3iXBY+xSlccnFlHubz
fT4N+WzV/1Rg+QuSUuw0wjeaMqYTcMj1g0I75NhCmoD26Jkt4A85yIctZ0G+QdQStxS3OD7kmATP
ZUbdiVAaAs64DZ0D4ZjsE2mIp/2U8y2d6qi9z4q6yt4sNVJ64gxZgTvJmv7cwrN/tJazDbAvwAak
hK2yJHoH52V0l7MDOnVyA83dW6cvy8hmXcz4nz1A/LgcLrnUVxHIcLcbtmhHFoRNGzIv8l+BTyYX
bnMWmdpQXinOlFz9GLppUOeJKk4WeGW6YyzPFXvq8KPPH4QcagfTJwEKCnn75NYJoudNNvj7RmUq
pbU5G8TN+URS7f3n3Hmpdfvhkx7Upg322Hsc0kb7RMla5kkqhcBERvDoNnpu2Xzjjl5di927Yrv8
FRrhQdb+6Dt9zXzb+7W6co6F+kr71BfrJYaNOapWaNK41IgvmhxsEMfRnK9YzYdYa+g+MWTcNiIH
ogq8bGZ57qP8zVyjw9OzKWDAX52ZMgZwCusEohMGhMpjffpPYzt9h54WpOjtjJk38TvE5lyXBAXO
icaK12SLWXX87NC+KqK1f6UcYP8VJILww0MpAS+teyf9EguS8bFtZzk9XB42GpL8YbRQ1Gc1XYjb
1Cr4oMdpp3pL6rEOleUvm5eOmPIax8vaxxYnJdInqr+LCNlNjrUQoy/GEzyJxewCHzKo6z9P74Zb
F8n2WDk+rRGLjiepnAQkyaxLnRBZhGU9GAKQXOVHRL49PwKHCJx/p9aH/EYZt1vogf5e4AORdcgC
GgQY1RrY6wzu1qG4M6VaN00GsRZFTYKxAriL6Ruif7iZynXelGrKqL8+TM4MyvcTgQpbHSPAO4wH
JMi8Bs2gVNfsjR9cRrJhfLjj4BMcuxQWCiw/E/w233bQWM5/deAtbJZ1W+bpjASFtxhLsXuxLbzx
gqwc5jH9y81e112N0RB/bH4wP12GLMhRacl979NWKKCWo9U1pJf7LRA4TEW59rWXEy+w6l3oycew
/25XH7gI5qNVqlejplCscJNLe6a7Ha7Bm89O72TCgqxe60qCHN6Bo3h5k/XL//2KNgbkyn/bbjqa
m3zWbVV1EqgjaCTUtPHqvsSni4eP6gFRH6XrwNoBoStM+dx0jUZiPzYl3bs2AGf0z42hMkAAGyxg
3gQObCLhE575ECvqZbG+RyzcZoDdxcpvDcP5Vz/KiHf2CSsRsEjosFhTN7yiWYHAusWKx9usX3Vc
RtSy8I3AJBRae08qBcAW9YY0yGd13D4iD5yJwfD/m2hfXfuyCBbJkdnIgM8o10eOxco/zK7uUw5W
pYPODTTOMudfNcDDf/1utnO5x6RRVfZTl5jF3meC0OTob7Fqg24z96swocUL2FykJDs9lR6dl43Q
uMy1PNB7OVsUOvnLtsgeTItiMivyR+qJJ+qM/0B9pXJd1EnLg/8IalcuZr1lZNL398IMaRoBv40a
U155y9jnbxnSk7q/FkytNCr9s+xIZRY6iclq7+IxPTbIL+pkvp+wAM1PhNhAcpxvcXd0prnVlcx2
OBF+8TDLzCN24eO8P+SCZI7Ag09RxS/mP3uIT1mIe1r7co+ZGmeSLgnyP/FlhvbAv18LO6pRLzoL
7GER1DLnhKQadbHqQZCbV1JdxNe9xP9MUaz5hmLhSIqZ7b2oWOLgFeUZme5aGejtneABBkt4veGG
5mdMS9igOxj96GerA+h1utk6N5PTM/JaNKDNc8Usxeep3t6l2+cFOileD2ZsYWU2L1qljwJ6CuVr
Rq7YZEVrdiE/xNdG4CQijBEzoZCnWDz8MdBxOxKFPVUUdf7amut3lJEhHAcyQVHP/7NBxnSmU5+4
sFO6wgVToleohZHJjOTAgIDZ0BmiDRrp6tmjd2XNSzej/pJyempmH6uzspC1b2s2PBaL7FhMX6VW
Qxyg/s0sYqJ5+EZlUePFZ4gxOXxu5hU7iNPxG2ziAzNQUraQYm+OV9H763tumkqtcmYlNZEGxqvZ
gPOiV7/dFbyYVey1zBrquQMAk6NAwkDGlM4UTCaNCaZLs1qz8EFd2iArDTkxFRmT8yhxCaSy+kOl
9ZxTicAhE4HNNKefLz8fw7EEi5RHXzGLMAEh/9nrm/WUpgtS2p7zYnEcuGrAlaJhgMMchmH6PZM8
qf9zCxUcZZHICMZF1l/b0m9ciWHO2wi25q1E7r6zZVmw7qhCxZKIiuyclEFrIrlSPkQRwmg5LRJc
Wi74dESRYFFKuOksh9EDOZ6zkLl/Hob/cT4NVdxQVfQxEhfoO2TVKElT2QsRnC0i7Hbpn8ffTl4+
z7lYuot+PyxYP63+aYF7X9NdTQsOHAHsDq32HIU5we7MlYk+JgI/Fw1pqKkCGOD/FuejvlXJXP+C
rsi5ksGr75zqExvrvtIpnIuNUFhNqq8DK4oRESG1bHPp62EwwA1G0vFMDKqI5nNAiQMFmwlClaTO
rXGJL8zRFd0gTWNzW72jP0WlQaDu9K/242PPoif7abWuL6lfOCrX+sXVFe3nWzcjAa3dRtjjIPG+
5ooUEG36wuFbJuCsu3+6iQAScEN6r37j0+Dl2TkL0vpKdJM5erFc2dT9RM8PXq1/xRHtvvwf5BnQ
R4gsqiYU4E3aNfGpjUzAHXIfTnUKivmpkZNL3cMlYVkWjQfq3za+cDp6LtT0+ptwC1AocfFPLMSj
avAWkwsIqhib9UspWTNrf7FYRvNw9Rg+qr0kHLaXqj9z01+ewNl71J3i4eNqgpzy7fbe+guwYdJ8
ie2i1AeBQtnacSlppP/VA/tvK54u/iMaT+jHIX3Vbn/VCJVMq3JMupKrmJbst6FziyF4PBwD8p7Y
k8GRhDgYkPrKDYO3IF20HJAk0ZOE4EXUNRUc8Lash+w+dTC6JgORkBPK7Gny1in+2rkOnSNkekeG
wzuClLQjtAoX2WbgpvUHeJalFfsSP41m9SgoC/xi0+iDbLo25cHYPgGcCbgfbZXuBJzJV8LMhqPa
quZRE3KsDs57C0w/2zXsETAnyaWSNsBy5eiVynHSAdmg9O4AxuS+f/syMBZkgfh8zKMYlKO/hAP1
yuOg7t/NsrbPAIk3Tp8ZA/GjRVNKJQxdPdmPZYIJ/W8jq2Dw9gqjYyBm3cd/S0NQ5WM53PKBinq4
O4HVQT7onBR8I1AADXExyLKY8bcODRuT/A4KWfpqn+0w9oHQ2+INiLiBt1uCqJ/c7Ev3ZZDo2B17
dnh2NiQzDyYZMpIR3OHwhc2H3pfeN0PeCGpLnXIBm5tg53Yat6ruVHNJ0hu71DzKaO1DOoEqGmyw
wxnqUg2zxMV04WGuni1i/oF5JazJra3ONHlrfRkPE+GeSwwuMciHrMbA/prOstXETZv60y+QM9Ho
m+kBDIeO61t9s3t8HRAcHWCCd49ZBUOo66hgJ805JeIQFAREfXkmJKCM74K5uv3imE5pGz2TjY6e
LU0rPsLi8DGGy66gkjrtwLoB0buwB2cSrwZfSyXoP01TRNM9jMxBIMAXq9FnBLUMaCrN+0fcbpbZ
y3JNJJCZrQq3/BXZd3Vu8d0bcLJYz9J9wh2cmEsQDwKH0Vb7y9hZzNnYhw1Py4SOuTAEFkhOYJoe
Eu12wJHWhW3smrYPpqZRkgeLR3Ai5j9cErI17DjF9ynW6G9w49QS/+ceA7NOvC/remwZcVk54taF
3O/mqZU4DwI1j0+8K6/D27StEHbbBYUGXKlqn6NC8ItUg7Es0bljzQFfLBo21iVCbQvE495ONwiB
2kAq3GowGntqR0FAhULGBUOMklQwyLKcN0+nEGUqh+dD1jR4KwFdzw3NVm8TA51gR6LbPD9PFGFv
YldXPhyBnry0jstWyFWG8NPsql+jmrVNkr50fuEy6zVWpateGBfKTR5KQRhOWRpUMMZmnQM7+sSC
VQAQalORiP6Z0/JSvpQQ85bAs+5ynefRas8g+I+Lj1AjHJoS5gafYR9ShHYqqFeTo6rX0vha6Ex7
OeK7rdXOHlFA1l9+rUywhqN6ssHWVldTvNhoRs1PNgUI5a6KrIk5CSMcppyl7PUaE7cwsWveepyo
j64ma/QguMrZziPqiy79puP+9kd7DVfqA21UrlP8D/gVbHuqUlXv8Vv6Ee/snD9uU0BmGVOd2w+1
5ftbkF6mTYSUGIOKmUOduQQiQP70NA69cGHQGT0z5viBTYdxQxU2oYHlKflljCViDwMX0ek2d0Gi
ZDkZa18qQeA8yNjm6JNt7XJeh6J+uaSBS4Oz1l5Mi5Q6N29AXCYz7nFHvvhN9nykDyH4q4k9l388
om0dwjl2RkcVvITlHdyr3lzO/ZUj0/sMqaaihR4pto+yWiOHUC/nYKdjhJOJjhZqztAXWPWVpyLx
cwzm+1l9tuHutWzB2VLf4R6DnESFSDF3eNr8DVngufBAu3WzDWN8Pp+kclwoW81TvSJqIelqOoX9
98T9DrRPINNfc+/KqPWQiMr3UfQt0e3WNplV63uJPVbZJl7mX8eDei2qLoHhveUr8kVzMSBNZaPH
m2BQA4jy0lyRDMd6MkI8/bqQNiW/KbzbO7lDGJAVQMYmor12zWrrHerPJKvAie77mUFi3TOGFg3H
Edr4uo/E2zAOYoAlKTssek0fPebK1os6iQgorqolYz7qz6n4efYF8wqu1IPDYRsw3llOLhKrnGSb
DkksKOo9/TtXSpV8OXGcYXBBQcF/CrNxOf47b5M7qrH3LTk4P0QGuBFgDfwhPprpL/NNU/dB8llb
6TKWGrMFtC1ZEpgXeyLDCNsRTGRtBWZRGPSPwJKCSjHJerGQsXYgfu/LpGR97YTudvV/hcq3Aeqm
/azhLcEJVQp38RLjd/Tqs++IjIa9yGzzvcZLZykmm79MjVIXqbA9uqh16o6vIAPSPtMa0Ty6NxXm
1rpY1nbWCj9/7lj0+eINFy/JjBFjSL7NGE4LfuljRkbEkoJnx3oQE8+VRz0NyC5O7sNmYdlZzfui
2+VpLNzjJElf3CHPLWoj/xdVDm96Nk8i4pvWdiVW3NiN2kGC6YecJg6h/n/CqkQCIe5lgZFUri44
gsGFVrckaKbHe4GsAHKTfnQvAQ0VhfhD8egciklNB3yrVxZDLR9SF4jlAgQR7vbCmiFLYsNZJZll
BWuoKG5kgnGUT0oM8S9I+5ezeaS/Lz0jHnycFDaT7zC7dUDMukNzcV3IOVtaZc7WPMATaxrS7niS
9FIuC8undEJ+IXlZmcG3FuNfo6itQSoBJIoKLGuBZyBl5rFiCBdBYZhKiP5GM1jvTUj5C+D6Ey8z
yTyHtycJCcW53YWUCLgVHZtbJj3YkINekn7ESOEQmFtbIkxpI/ycIMndDMbRNCV+FRPyM0aceNrJ
uWX06XvyFj8iqc4wNzKxetz+gMYQOMa5DkBG0PTD1B5N9gNQbz2FMX4gGr7Kw6PEoPfUToqr81OR
VXOa3Q8Up4ZS9K6qHYnbK/WndI8V2YalrKFP+JMtRBYEbXN1Xi2MocXRFhGCmM+JRTmVN3/nRg5z
N8Sx5mrItwJEKeMnUkfbVJmoaaKSXhc5fOJ7sWGzP5KdcRs+VJyuwaxAlMh8CY6d17r1Bp7XEzYF
hm2hIR2ZzLIGj/skrVNQUiQVKej2tQxSFQpE9rF50aCu+xngMKeny7MVAm0j58TlbkHEXdsxAC89
ihr6vny68Uddc2FQmNWUJF1n+HC9Q6xQ7S8+MYyQOw7jY8N6a4ZkPLR/cW+HMhIP+gGDS+8iJKxE
eku9wqgsE7Xt6oIkofelqF9MWpqj0/BdqNcYFvmw0gp7F7c480ZAvcr+VdiBCjh3+Eh9ZyUUpSzt
hsykWduYjprEifhxEL5ne/kBByBsj/WwdeR8i/PZq3c0uyYy+KVGCVoygPsPKWP8jqXPkOBluIQv
UJ2LtNW68gqKiK0schio8cOtA1oFn13PRDODE9+UudGI1RlaPjhCCkKh8bCCkHBnjX+07MJp25gQ
XNvz+Mi8+A7OX06fRuwySVhRSu0A6afQ9WtNtKH0ypRPiAQI66qN/970MZnX//tOZDM4dA6JM+J1
zMZE6tcxvD+GCA8mPoJf/xv9acQ0Ksz1nXG+guNgLnCAXUlp4KKrKhi3garqkfF7vkzrt8zoy1OL
n0w01z3J3QTZSz5E4metPq2FfI2YvEOKXwWhsQYH2ofKVF/fUfAmifPYlN9aPMX4SKm/Q5kt35Yb
sYbwV6qXw05Dm5kJ6q1WbhhFR5iyz6gkiegja6Wo79+hS+jIAW4CcJOTmM75HwxpE9sXgGy22uij
N4p+nCnOdFQDBm84vRiB4rKdqxCzQFvGpGaZM9bDDEoYLfnh9oo2U5QQ3n0BptBGU98HJ7LyTM6A
euzAvtQs9ZfJngF5tbn+uNQzHSQhfpmmXux93x6ZQ80DNSIl5ruEfaj4cqffon1RB7UCEND6csDd
lJyA55rfWRCCw88qWlTSH6m6jN99nxYXn4sYyvxTwXl2DySCYpP/UodhIzPrGSF2676MeabJAT/B
yFT7YoGlkoIBVL/LBgyXTztbjaQcmF22r+BM+/219b7fNznhz7/Ru8noSxyBaHisnmfa8YLfRwe2
nlYHkGsDfNE8xP1Ryw29PTSiUV80sy1DgmimzSFisq0yGtR8F9l1VhHoG7eQNTFSsn0PKcPuEbmU
Ck66ahKEq6lglk7qco/JcMM5ry58vJTeNzomqWdYZP5jyyemkJRGTmi9JGkvHynIv0a9ELXB/egv
UO/xwJiArxRE1/oMLLXz0GW+qMFc4c0HLMVVEEjWpIkpARr5ikNmlkTqcEFu5Fk3/oOlToijr0+0
qfgQG32oBhjiDnglQ8SBEiAW84ccPAlgDAziIFOqWZA3KQDioEMOLpEd3Xq0Mxfe4Uy5TkWHoAH8
LDOZkGyK2KFpqoTLbzwNwQWzWM+ulwJFOnaX1b9azoiIja/6nzdBhZyK5RnNqF+sZTnlaWkU6/bN
M5sPBHXUryF0HnGym4E6yNycCojJRVr9HY+gNkkR/rahC0u3bUXm0ttuU8PkZOLB5ir106no5dUH
6EZkh3K2a5uvL718lu3bMqPakQxK8TaA3q+RRagK4RPP8rfGXzug+B4STfq4tAJ75S09x2fi6XLM
q+oFaTEEtaN4yxMNUa4BKuUJxsOzK2M2RAx3si4AYZE+SZ4mVDiqxhsW6NAabaeMpnRL2Epw7/YO
hNjNciNZtdl+KqX5vvHH6x3E2z9buC0fx/jb+PDYAkA7IaKZfllO7jhJcmHKYCoY7zsi++IRClTf
GIwxhD2X6XS2lC2+Hwt0iMnD84yrvYHrhj/qqBJVQ1tIzmDE3CGPPh/cv64UWF5oE4J6K3UkTO2g
/G1LHgIlprzbrA0GIaWLfIQZRD7riSkgeCeRuLIB0VHLAwJeHyxXtx5O+wIAnqRtdVHdm1swb1dN
qCR7h01qM9dZpz7wix6uC6gpbk3kb7wfXpVU+Z8gPwwgIa02cEAJxqAKnhJkhtTlJrKRtqOvS2rZ
fkURaqX8VYhIkuMvNNM2jcovvxMRFDuLikNe3Anz//9CTnX5H3xrUPISs7IX7VAY1B4+y9SC0kxw
mbd1ZF2ZJ5oA2AeSIMvzSbX40rFIylc2yNUwq2xE1iuDWH9ap4ZL0Ar7hAUMyubpYkw4iJZJ3UIk
hLRA/XOVMRtfyS9PY+Ckfxh3RA3v36P1CQ2Zo38+PiF40eqUwlApPKvIO7tNdyCUx90dBtOKg2W8
Iam+A8PVM6vcMSyVaeAM/TtL6xkvgzxajEk4RXl+fBpKFIqQ1PFqqVIwSSt+OH85tSFH1xwY9IaE
74uLdYSlVGm1F5KjQtCZVU78pO3nrXqrjAW+HcoCo2VEV3/bip3WDn9BOK8xIUT2aRhJV7asY1li
9iSB+bjpALpm6N5Mc+o7DsbgEspqVZ4k2qwY/CKMZ3aYgK+iJjC0mCBv8XAVBtyiyr3US/U68um4
DWzq9j46xRgJbWrT0f3wpwIUjge0YnT1zRS0mrzdhYMfz/zQQPGFo2VCiyVG9nfJBa1kwEHTibIn
+6DQh4Yjzoy3ryGT6kszQbXmUvzgw6H6RK2uYjFrZNL51syvKIVxwRODs3M7o1nx3vWLPxBPg9vr
VYnpAXcgvorCmoUB/MC+v5TOfVPc42JpuXJXCRMqVt7YxM1jJBDyID8YkPTOpN4CBR1KSkMXKI1C
DjLv9W2mYJtap1qX/r67jl5kVDiZvOTBWaoZ52OqmhqytBGJLNHnug20r02biWUGXwLJW4Fxkll1
NyLCURaWtobf9d0eRp0iKN3SQ385D0vEf7/vI9D7Ufs7eN0AMe0X4YKqysAo0jbMwJrynGglH4vz
Sf9NCWm7INqTBcqIjGi7rt8gnaEaT4o+4Sw0M1K5hbQe3f1mHrU6bT03g3Ing4pCbaWCdRDSHnUw
+I8K0bmnp+G1nr2LnbrVogzFTAu8nsnKfgj/Hh+01S7qdtpUCxzUI78g/Hg+skWB9rel01uJFbhA
LYhtq5exzRB5CZ54vxZnJusjTRVIdt4u+/SRV7xZuBX/5MTzbBuHCzofZ6wjlLGzGf1JVloA20P1
c2L6lCtBts9XYik+/frps5lotPZnLuqNDJEwQ+thu9SM/ylcSssrRInB92Mh19ENh0eM+BGSD/rX
SLRY5gcm9Ifv/VXYObjuGWE+HOMob8xpQLiXoug1OJQcB2HrEjIWJUP0oHrBDXN/1hrXWuLhGcdB
ecQwyfr0Z8dMiPYmYfotVZOI8RtvHSr4zfiU30dqN4h1YM6ueUc/KUZyg3CWTsuIlQZPOkp5aRds
bhQ5cujthp7n2XkjNo0zLN20fVUxRYnM82iPccsxZrevhXkHG7hODTpjY9m0Tv3WBdUDzykVWdlR
/KVvzAwcYt+KDKFZ/6BxBxxSsgBqTQ2bmlQM+X1dbyo+fRFuWgbFEpQGYmGVojT7lIO1SG/ed+BP
iwn+vMVo1LMAjf2VP7prSLeNN3k0fbhUmCEZF87V3Q28XuvNb+9fCqr7l47eJ8qirp1C5tQf7u68
hTm01xwSppVdwYihWqYSTVhh1PDJZhZyeutmmzYy9ABswUMOeV4H2xki07EQtHPlYvm2VceeX/+q
Kimis/B8HAWiAkJyn3aOfMl+Eka0eSc8icjX4E4gWGIXEe0luEyr5ztxqB/XCqS3q4kP6Aj0GQZh
NXTaO4Kp3y4zIvCSyezVGVYN42adZlcpNIPVWBf/HiX/jGzMTmKWMtuwh0N8DPa1mooKDolKGpUI
g5rx3308H7lJGYIYD2ynsJt5qaNBAjenB6M5E9gp65Ukxejy/fFvG+IKvqF04DX0vDmeLijOEI4+
tuEbagqzfCsgUPgASiUL18zjEXZ6/ygWeqA3oevASLnNydlTEVkzS30HpoeFq7E9DJYkJIrb+E+b
S+Uve6Ybchu8bYCKa51F4rZ13xYsNfXTFtZ4EYtbd2jWieXQiu9Myg9FOGEGXcgfkJ5kVGCDV1nR
NGgvEq9YKc8ItjvFBbjSKZigOjS57XynXrHnpslrlS0TQSAO2hTKfWn1jugmCQx5MIaw19mjfmA2
H9BZZMtePzNrVEXsqY5VicXikUhO0MeM1HxWuUMh/DyNQQTIxUdyBWfDQwYC/JOGTtToRpC5XOlV
6hHeenPyaWhHuja0JEKhkWYCmIAUqaQJQCDtaE+VH+P4q83NK6qpitYvKiZmA4CtgMLLhMa7Pz6j
OPwUm82+1IYm6FoURrylJ85XaiCKHQ4XtC5YC3WAKxIf7N6d13Ms7/7hUcLIMYKeidRJuuq3k3sc
MB2puHGOgrxUaFrYX3auY+J3PElGwgbdi/eb5/jSwLZhiHckqWIR1KD8LBrXSnNSodTvZXIqET1Z
UHICsxRMXEcPipvuyuTVKDqjQ8udwG4yMUqwYBpLdNWh+hU+uijZmUoBwtOyXYfC92kcO6/TCQF8
NjCbdts4RjB8QyT0ZckJ7XgOtyAYSU4crxX7vqBEufIV2Dce/9wl4gBZJoCWClxTlI0OUbhl+R2+
dcsutwNbS7Jk8tbt1aKlymZwDtq7vQUrfJZmDzH4vUBqNqNfEowyVfHILbPORLSHXobBbYhg++yt
4NtT5HuH2w3t6EZbhs5Pgu6S6dyi7r3XPtDFH2QGd0Az8GLytTK3OOijxG9Qnkv5bw0YfeZV+I6R
0oCWeHz+/xjuCNiOqF5WM4E8wY9LX87UPXNYayf/5MM+vmOCwAbi+PTbwhIfQqkckGY+UDt4A1i6
DFA4zcQHVUWQQIDAXNsLCWNKLh8V+f39cYskxfvBFAEPY3uj1Z2xBKvVfdj24NZfPe4Q56UK8mHv
HcvJGXwflKdO9/sJgYZPe7Q8h8jK6hMXSzm4ar4gDGJAjHK99l3cBKo2VOfIUv31w6PXUljPzp9i
5siXJcMJZyb0QsHCXvz9QOnoBfoxAp5qEve91LDq3J98ea4UZe07q/Pa4109OEVZyuJFWY7Z+mSm
cUyrAgRc2JYObcvCkeUg0hOb/9kGbdGWjL3/9Y6poiolb98LItHWCed0AFpfAJ75QoIK+c+zipKK
izNTR/80IORm9VPEb3Yv7HFqpFhMG9IoKRx/N9lEskjs4iQNmqk8yK1Qtx/0Q2g/yCjXStrGzl9t
+ZufhbvR0z4nPfjN6d4OZj7YDWycYkQrE7YrEWlHPW1TvqLZcb9XQiz4SRiihoDfkMji3OyIEXLv
plAJLsnaIe8xeO88o8mvtQWTbZAKymhebXERARewOyQgI6V4u9EM4Is29wrjo+yWALUetUmxNoeU
USHyLeKNQyb8Cjc0AuloiaysloVWlt3XVcJTAnFiZnw1LxPrEB+F7AtkFEcep+ERF7qQz8iHJJXN
lOa1VhRA2c6M3EMnN72g6rmrdrywPxSMUJ+WFley5i9l9nWIYrTFACbGvA5e7iygyoIEK7tBbKyf
DSpglVfTgSAJ5AA0Dac/4GP8gNQDGCgsdGFhkf4V07PxqSPVGqYOj6kvv9gc3iJLecD2MujiU0tt
2ztNeGxcd/PLjLbqz3EDbBMfyz5oeyc70IQT/TSmZhy8Yhx8wBREcu2XI6bMHSh5mifkt6ovtCOs
QG7XtoTAyir0q38/1ANVQxZ5BQ2LmuLD7FbQzOjDQkEnuFDr7cL2mCfuNQW0W6Vf/v3EdvNSctrb
bUpTRHzLbJYbykTrt5nE9l2jzamRR2BZjGyAF6IG0XX9vU5lPbTW6dMaG2t5GRvu+koP7mNwvfvK
T6hAVKrsHaMANQQHZtms6pMd61jHOvazCmuKpzGXangnxi/KSRxTeL0e7M/dWoQrbcPIk56FLGjz
uz9KhOTHHyHrMBweOsKZ+UwDAMhnK9cmIt7A1cfOKS7AkQS+JILloi0ljqAm46LqO8tIiFwKsocJ
3UG+7+RAvUTclIAsrHfbTwik7DEhMM43T0Z5mjl/f/yhbCHOVc5T6oAGpIv9AfuzfAqUwwvi9Z/c
sd7szxAM/FoVXzUMdfADCCVSs0TD988Nge8eUy9Ddp84PokOLj94doZl1Cb1VvSPPO27m3Ozm+81
6qt0Qg59DljGSpfnrCy7psIHFb+ncJrstpQ2xMDLq9WXdvgmCvIAtuI7MsstSmV8GId/tEUIRI1g
BcyOGHSSl/k/QIc6BDoqvcCC+XREElDcXSVCbYFoNBQwS3rb7uSM9iMLhZ6PSmlA7RfusJelDTJL
Y+oIwogcRlIKo9e2HsGwfZcEpOkC9A+KQj7Hnq+v0Si6yh5TPezXC4vxJwQEgoFbXT9+mkvyUSDc
7mwG7QhLqS5KDoodWMlgIuW2rCSa111D6pwFZ01u9rcLgr+aC3Rn6fmsvtCI+Zmu3Fh3tifbXusb
s+zr2lA4nnoeR189F9CfjrPq9nkuafK3qgstu91yiEAocMNfbZDlSyC2xq21Wk/qV8ZxhF5rYaa9
xGrL0jo8cxtFvWO3Omh+1168Kjiw4bk2UTDNkIcbcLWfSFNikjX9CGA8mxOYrtJEYX4v58uua+iF
nvhFRB4VQABie4Pt7ynXKZ/S1ImciyKZhlJJ6g0F6KH+PuAyIHaS1X0ZaNwAorzA/yRL0/7aJp8C
3c7NZERVN9K0rsGX28S2+jKX74xMOWhg/hrACwgIIhxwmZPW9jnmP6GPLP+devo73XYYkvRfkrqL
LE+Yillgl6jUsr91Q3PwiwcYi0R0eNk8rO3ZTzFeROS9FbBflTlpDJ3PPh51Pp1AcnHDuAnnF/iy
dUMvSWzkIslENRZPzRElwhbR8ozKBvg4gHKR6LSiWnJi5MKh/SKYIvIPxnZYFqp1geNZqYFIgg1J
q/dymoFKjh3+UahJJcz84Wd/5icaRgn6ElRmY1UilS1g9jgZ1+ser2GQelbspW0TUKnuiwTtR1ZS
aSZBfNorZTTFayO6BnIAOJDhgX4MlpDYdXfjlqv7Z1TAKqAUOj/GexQ9YsY02LhGpcTIXpVy0QAs
AOWIjCaP3qwX2dndJckgXkTDXoWFhzodN9HE+1mKVh10xCriZW90oXwT6D0AqGqwm6hkTWYOFsvE
dv4JH+sb4d84Hno7zMxgJOKowa3/LLPjyFSZ9dUWsED9qImMbmoT5A5ntk+xzgNKK12gpqDXg1/4
JIwPdFTE7qM0Em4sgjQVfcdRTiLWreBwh/8Ew8T6L7G9NvtxFwliDkE1XnCZWMDzWbKyn3p+qvIx
IrNh0QJVdbgwE5sPrWcyTtbAMo+6j7b+WYDGbVN3Til5Pq2l3x7dVBbA/TZMmtMf7skHHECaW+I5
3gs9u/DJXe3swfC+6diLnrubUeik4qMnk+LJQPJfcHp48aKEiyfLlqz/ykrJ7VKphDnmRZl6KrfZ
Rexh00JWE/wtrr3674VcIQH2Q6D4svg9TshCT09xbBZ3bDkTn2mDc0CB6p5Uc1zxmviq01+hAG7s
chkBKSya+1TvOaIjZ6eTQTKn8GXpCXmNorKJPpqKc9461mVxxxyZjACbNBz0usrChYJouZ6YyOZx
ZhNpDtbyLsPYAzVeAHpotzuCSQzmpw8JMc2knJtSCAMLvrlRn17xOrxo2R0VDR+KJwCZc8zLu66o
tnyoaAn/GXQDxLHeQTJ7Ipuy71/KLk1zmvssRSEtmY3Kc6fskL3/xPNF1d2ehuavnVVirmEG1cxw
AwgsJwVOI4uw4gfVymHC7HDMPXq9HtM+Ky5HAQzcM41o6ZG9+PfcS21AywS68ybblgeS8t0NU2jY
lvnLaqEdkhQ10SPxyCXJcFt8AkMlGJMQL6sR4+nojDyJ/dCuVA7Fx4qxKORRuzOKaBIpKkwsaqtJ
uki45kxXnO6/nzc/QLKw8QBtEqwwvm5iUGHifmGr1ZwgCeGevA48lHyG8yyn5REAqeFTu0Lzu0YA
KNwh7Ieq1z07CC/44zNQqB3dPMrTuSbUN1w8QVnDzQuNQd/gOMmczx6cyuIA5ZqlhoVhvy+VM1kE
3vWMVFH/0tqNb65+WlyF7pROOPqL59zhEiWZzB0OMhOkVBsAZ7oPB0q7AVlrQ8okA645/qcOPX7i
8rgr1AhdOXADhAiKCkAYix5l4U1wzSgL2u+Pk3T8AnQ9akn99rqKt/8YVFYlCA6pVSGxxvKjafws
w+vQLD+7L97EqfjWXliKH2QzqIEhEjIqP2nmJiOSAUecOZJVuLhVb8OLA1LrX10JSDloCJdIOtT+
NhLnQo9H6vTV0hgHk+T/lECoiIc3086QRDgZAcgv2BZNgNo4AimHtmeqFUi8S4nBG9B0dLe2NfwO
o1dxLvDDVmE0WfhyrL5tbEGAmi9fnwNbhdFBP66pVFyE2wvZ93lNasbA6cyUY/VwLEWDvtSMGh3/
XpKe3LG0DUZmrx4acvf3kaJYg/ufrBXGtH5gANG3jPsAwvoNHLKSrMPxBPoi5wjUCPTVCDyZ+zXX
Eb6abxDAeJESHHO1vVt8hCMsyh3l8ED10W57Tx2l9G+FAHx6CgAoeSJEl3JCtpr/S0rhSEPJOW9d
s8H6neN4I8A29HZS7tfyE1DDpSs3eJsP5KtaDZBqSNFRL12DMMXg3gKr+M60R0zLlvJsSAI26jce
avYd9jTmTUvejTB0JxculEkKWG4q9ciivgdOxQ4MQYXDCak6a8Ta+KWhKL54SLBdymn9N7hs/5y2
qsy6SxL3uBGjQIVCF2LiS+fZ6aAgzoezr+0zO3aT0iOq+oGLixsAawUTOpQNKJUwLICFvBERSuvq
mWGaiTuYnOUUnZz/xt3glGpFGe8iuq96xg0zQ7r51xnvi3t3lSJ6xgSKoMdi84OUw0cNWn1VsMZj
A2EgFzaVfoViNfmyv2mF5Vticjnmy5VPGbTIx+mPtof8rGYAX6iPztTfuNoK3Cyd02dYV6u3/hhL
29l6ZQtLt28EyjGxefaO0oen4s9TJ6Sxm//Z1qOfroQtr4ZqG8gGzF+AWllbXZQMpGeiORTiZdAh
f//quqB52xAfl5PZpAAnWcTWXhuBZIuRwRfWGg3ZZnqOUKzbcdMZxlaKOqRLtK2wa9H9a6AHE36Z
ZG40XqIVWX2vN8vTGiPhhQujuKuJHHZG/RVZ0BXLm1IMpKQ1ebi3A9L5xnjQlpGM9Z+f2q9Ym13k
0sERUpec6MsYuUQfar9G8Eoqq7LZynp+qGFSm2FeoE9Uhv3B4B68G/lWgapMZ4oAU+Gv7XTw0opf
fbgiEEq3ANZtRlDVS0jXHPFpIS/ueThg6ix/54RzbbdJgyGOkgczcvyiDQmGTHuYUO6ONgmKZsDB
wz7RVdEMCAicJlCkuvOhi7g1hpXK9iXEIvccT6aOFJU5MrBcZmZ6jc53LK9C11NEjE7oS5yC6T6r
LASsFVEJzDM/tIRMxQoj3dxHoM7s93RRZKQrInGfEOKzI36JU61+v5LAVudbeCfogN3gXrab8Flz
KYvbQLa7KemdXLQzZEbmIApgtR9GtiCAhQcQdOZhHKIjEvgxw8kKjXptdw5ltrg5oeBYga6psojx
XiaGBGWokAQF/aABaC+RZ1gOdnjskoRCucT0tfAn+sJO8dKPcUcb1B62l7B24OkbKAV9sI1bfYpc
y7rfTBV+ZaMSEa6Oug/PPQ6AW8A4gJV5rLXcaVyP0jGwYVArRO1Cpsd82X+TbgOpN/pLTX9l50VY
FWEBJUKF8717qQvvpPDvGBZSyGhUsy/Etn19Tn7k4cOUYU80RQTk+QHcjsn4gsAVLjvnxc3DxkIY
Vr0x6JoRI7QSf9iK1ZORYJ6W3QPdhpSWC6+N89Wv4F1dso1gj/5FxDw9V1E6H1ii3LWBza4x/MD7
E3Ol+dAM/agHo95tzneC8rsn57205opw40wBoFOzpFIE5chkGzldAazeASYH0KuH1IinVZEecjL+
miHNWwVZtYgQ/0Ngj4Tp9y/qX8ISmQWRCgdxzeYHzhyRhMYwoyXdF7LMDnB87KOwrc1TfYfMEQul
N16zIGbu6q/Lm97F/UFdNOpnmTFdIYU93siDczD142Mc/h25kyKi5X3TyeE6kg6SKgRifvxOieuR
8U3hGHaaE9nY04sa5gzMUohn/6vFB6myf5iYOeutHu8TlZqzqEsi9AoadoeOTHrRGrnQC4I+33Ld
tYlakolGwyFXf04Go+f479JAVRJpR3i668dGCVGUBQ+Bk0NIswo1gRourr4B8K9CTgvB2T889WKQ
Ho1Nz7qbYYCWyuU/THw09AXT5rQf0CHZw+3+K/cEU9CVewe9a62PlR7Km8K/jiHDg15s358/YWSv
i/eOv0DmPqRhtXIkFXVh/gXJ2K5QAgdey0JK2IASUBrjmttRdajvX1xp52mVQOKV5gBhcQjPo3FR
p1tZOmvOamAeq0+1YNRT/dM+xgk/IKlGdOKimdZxQcAdv4U1fkME+aGU+KwiZq4kHflt8+N2BLj/
ud5yIbQRFr4AniUs8EXJC+wK3fCwSsYi1a8Ek8LFL/c4sLBBNKAEOuOlMsoQLwyVySVyqKy3JhF1
SOoBuhszoiLxxpctC57bRgY1tsZ8pcvFMtPTc8W7+sSlm6vSZC3rjS2vU9pQEDqnraDrROq1Vtq+
VdM07mdqgSvPLHFuHImEJEmQ4Cv5yDFQn8j5O2FIPiPf79AF8CTzAygeO2QbFXg+fXdCGMJOjij3
pWNsXrR5BX2u9foTTnZcCMYCfrBAP2oWcxYhqrdvG5oqddAmigbFL5SN9HXagW2XHu+JVtaLbza9
tJAy9ceiyIQ+8RNh/QJHHmVoqqt2jUcaPrjWnXurfYejqPMXG6qZ+K6S1UozXAJnRCYduazE+A9e
WOBO0dht2z+2Uydw+9AWIyHFIbKKHKIzP29yqxEVi/wUAUNAyvlLR0KZ8keDqrfM2uigW99EFfYf
cxhdjyuvV43qe84otKd1BmjYfqHT1VaI75phKW/Qc/Kc8UOY0QmXeAHh2z3rBOWX1vTPwJY7IaiD
tdeAKDLvLrlFPy2R4uP8l4PEAKuEpfsIh/OUeFO0bHZ3/KpEsymMqoqNObE5ybED31BL6vPcFh0+
i6JEUDc1jVgc948j6SUFOUGVbf5i4mOJlSkrppJ7RKoL89iTjInBJaGyV4jA0FKIM+g2NdLtOJ2P
1U8L6T0ejIyI8MZkgjplBai+++m54IUJrlwJA8fGro7I+JY5giaf5zH8u1WGbWS5l+crXfJUhdi1
E4ha7VywddWJE3a4YgLsycyuDGmcRXtYVLZiiNBzZKOaoR41pI/hJhU5dZAMgoykpGSkrYWAQMfR
nozJyiNsZ6GAmFMH3dTSkmpzUZPQgZahffqwXAxvo16U6nd583TTz23/oOnf7yh5LOIqu1BgaZrR
DZnGBnNqGsjosnc2+T8I7Hc5Osbg+O8dMsoQ7Dtx+YxzSW0oyLAzS+G9Z++PUfvBsRVS/tVX7tE6
i8ff1arJcX804x/ffcVdY/haUf5Dia4J9i6sDfTz9Vv40IvJdqoaObvjiiTa9nuyPTVniSmot4Dj
lNy/CR9+UYH/KmCf+BCO64G7fDwq3A9YU7lf3JZssBE485qXY5qdS3QaDaQZ9ijKvGPHqasuMXqq
ZnxbqmcOqNDTlZBo5FtFH1xfAfPGYxzq0XVWJo/uQPfy00L9GHwRGaCqH2af4lb+6WF8qvwSXV+f
Hc55l27ce6kyXbWDhnwaJLMg1VaRtAzZfb3okDQXfPjmrmZbd6IUhdVjc474RX9RnpVAJhVwLOE1
gwkcY+cfix3F9riTXpCI91jIcMYZDiog+3zYDS8Ut+pqb/MjDv+TP+9cg7S7Ystj35OVfXM2++FA
4j9iKgcD3JmLLwXaRBv9uPviXXUV3b+DBClzfnobw3R/w5l7jAFLYt+10YEwiB8bmE8jJDHXiv7L
jOQMnY3exTK/Djvftjsg1M2SwL44Qz2yJFUdNEg5xSvNht7bOKylDF6e93PL0FrelJxsn7z3SSxO
yW8BWsjfp3WLzzqMDQHfPV5j47nYulN2BgnG2zgDPVEcItXLWua5CieswPXbdnyNRSSUtBE+J2nk
T/nqKOQ6c2pFEEZ/lx5HKHW6Q8ulmwQJZAeduRvSER85XAK9zJKEnS4OH8mGBKKyIZ7FKy55ttn2
S4cBlQAvPYxNaLHLE4fEQiUxVBARajgzqoX+JS3mtE7zB1RRVK81eXWDuL8VNzCivinTCHAXX8mY
oxMQsWqPlZXJplYV9Us/svhcIRol52I3R6FTdlQjPZD4b1oFbzzGTtzeyG9P3KIXJ4PZGLxASkaj
eFm9sJyIgvDHLEgDhlFP6Zpg//UL4ecnUwUL5KZFt6TpoLdd7WGFe9yn0kGq2D26a156jBm66+Xi
CIsFop8A3X9jrB4vBIPjtyJ/mmxXnvnmZyLHLXffdTEX1MExWcPRCw0zDCZ5DJobrpPQw03RqOIJ
TXSHbHcr+fEjUISW2Sp7GJoqhhANidhYwwMWY5+rcwN04883hgzAhkWVEBgeRcL/tkYVZKS1igRG
sKp6yyyLywbGsoCRsJapu6dyReplQcd0q+Z1RIBzv9hL/Vv5BepnMQSvkxTq12EQALvfpjsK6MsJ
chnvxY3VhsqobSW5v1F8oEhdlP1/7nr2fhj88GbLr+DZjiZz9n7Zxm920sz1b23uyj1eK1msveMJ
wbEdfKEEyseX3NCBV/PkJW3KJyF6373e8G09ormryGHTYuXtypOXWO4MuIMAaLIyavxcEhugJxj8
z15BW5sBhaDVdREBXa8zRdZ7WY99cJttDP7E8ziEY6Ms5f3yCFkSsjLzw/wl/uO5RZo3mj/H8UX8
9lx9SsqiAS1nfFYM0hlwpf+10jCvf3i80g5FKbbTAJLuHoqG9FDOVTSJ5IjgXXYVMuUfR4wu+f/8
dIe1WW6dkF4djJCKuuIQQuHH+A0caTQGPl9NYiByBwSRU99Sktei3DqB0RTNedj1rpoPhpO/urRd
rjKue8nE2ekHV6SXc7MOjs9WDg7mRJA+5DXLZv8GR1xKlymHd9RUnBY2jIEU+o5HSUioroNXebsj
u1jY1yQ94wXkaJa63cw87irDXCoicu5QakAdBDs8B2tbm6ZFVhJGkcItYsIhtZ7voxKPh6q9PGuL
8Vl2tr6TLgruCVplG2ExSaxGAnclnBJy27HglFbqIkfjtAzWopOh0tIeJ7yTk9bAkWOErIc7mR4C
PwcAUELycmzv6RuhuujbP9KXBPswBcz1aB47ixNLKtHDBL0t6EezYz7lOfi2L8u9XSrpgDoxVSaW
s9MkB7IT9vBjZEnD61sAtOUmaNdvtouBSsRhonf77TK5IfqWslCPoazrUwucA0qUKELFWnrEj6w4
HVKotR4non7hKPDTQTC5aweN+7uOcosU/I4MkAANM5cjlX0FAbmzrlBYlQX1wtzDIsbGOYz+DWB2
JH5+wmgSb50fLyTW6ofWd2+Ubs0/VWbrUvD6HqMRMLoVqjj7d9pui7ivv1om7qWDNcSF1d+P3qoH
8f17N1e4OrXt5KIdBwakrTfo5qDi2U8bjcwNW8z/7LVKJB6wbQFnN6qcfeSbh4qe0MTqsEFIDjbV
zgdizbC94Lvi5n4NUKyOr/Pxsw66g3U66P2NMOPCPNzhZYJjmyxNNXtAHnpjoacZAzix+EcP9exp
Dq9gOIgloc6nOyb5aLnCQOGj4t0sg5XiwkWurzct6xTmQ3BlzWUxS1bSBUeK6YcUcrwZ/zNRfqne
CvTQ2UnPQ5Y/yiSRf8bebI/zlJ4/FrlUURv2sCYjco81joHzmjcZ9hMp288IhOPN0WYlnL03zQRq
a7/7fCXI1EnibWpliE/O+sFa+ksVhE7P6+dX5Brw4ziK6MsV/pXYZxW9m/5JC0RN3l1HKbN5V7jT
R3UnVRGlQe0lmTn/zqQWROEgLZ6aqZnjtTLgBgZVyGAfSazvUH277huichDbGI0Bh5yFPXXYQQ3S
7tE5pRZnVUDd8ZAGtRCjNrINn6XV4ObYTs/4Bmagfl5wUBv/61GSeFlIUjkr8OHhokv9vvxtlTwQ
Wh9Kih38jrkd9/2KEMt4+e8IcLNmETiabhkp433l4yVXeC0HgeoBj/S7gZOTw4rqWghDxCcCgrs2
MEX8/fEL5Te4XqARztSxk8Z3pjH0g+Eez+OyI6aq0EUiHGzZhWX7Iq0u+z+A2J9ZejlQWjs3oG37
MrSY4kRvJld+gRpENEJmdypdx7JBE68F8K78XUd9bKZ40K5actGpx8xAiUV70A/2+XwOBdZtL53F
dvdeSWF/rRoqP8CcrVPWw/zvD/DaLkdTSDoYd3lHWbR+9DZKrLpKj8Udzt4Pdvnna5qObF7aMzdI
gN9SczXEz48Rlj6DXTjC7XmKngf/G0Yy2A3EYNe5iQxCqrgG8+dslAfWTpq552OgkofJTOr/9YHL
hJQM9z7wDU8HcukW4Ad0tkfuHZGkOQUgDh0Km5gDUR5kR7FKWKUZ0ZwYbbkcMU8STIyjKL0Oh2R7
zXqXgts55wyVIEVC7IsTsE8RTfF1f7evdCwIiN/Y8GTYGl2zG2LWCAzrIY4zKlKB7WGyQzEjlKc2
V6mARMrnwUSJ6zqihHlDZMGbPvrJQ6eZSmQyDoxEQmYWmRR+Gsq1WArTfPWWFSfKjK2iSj3iWyJn
mmC7vaiySbhY+1yu4gL98QaWPKV35m7yynTxhItqDhd+AYxZk0wZZSXGPNZg//uALDetbRCW21sT
CKWhXWbkTzB7bbMCAyrCvuGolHMjgGlc1gQkBAfEsC94nPXLhQ1pFZNj59BM1k18cX/M2gF5Spl/
TVQX8oAR19XEBIqxYKFAsixcLlabIGm83WXlAMDhnaieNGjaSKe65FA5eKhoDtDRABeBbXhZdXNa
iv2/jjbGNKtrT2ZdD0p3QwSj0ONOte3RjtvatmSU4b9Fdt8pwVWvdaJahqkMFaO6ZvMwV5eSCbab
PGqLH/HX7PdRpiwpMG44DpmpvAbaYLPaQyNugT/iIRYSPEh7yYcCbMAjg7kUa/403/BMBdbZ54gQ
3kOqfDxUaDFZreq6q3xcMf9F6E/wyK642OTJSA09AQXVZEUQaWJnm8sp4hGHmbh8g8XpxCz69yFF
zAUT5ozr6BlZ2NP1uSbsKhb2Ot6Ws0RgZ7/UxMTlG5HtKFoGook0HyUkvykN8usCRjvj8RWs26Eg
BbN+NJKPupLkmcV7x7x2oCuuaXXvZc3dfMyaqDGDO2tXERa6HpUP+8gwDNjgsUq3SnxggtiyvpE2
cMZECsZUr0JdxqFnyKLNdLJbRq7Ycy2uxmTKZCeMp/ZPBe98S/qjOEi1loq0lqh6IB5wNTsEqEWQ
HmYkyBEoVHyTZErtpUDIRyIyQbUgwQHVRPO9DTTspE6W6o99R9iy4ZsDzDGDEj4A2BjcFgvzhLUE
/I4Cql8C1kOA4ZgaIC8vsffokYB8GBZ5bTg2A5vjvnPGfejNr90FtG2u2O7bejhxzS/45AYh5B6B
13/I1nxCrPCUPNSy4n3Kim4eY0r7pEdbD3/L4CGbsDTKbR3DkVrjzy+lqYKjMgAVZDd7tZPLVgsK
nZdKYp4GZfOCDy1+wr8Q/FjC+q53Sf2auaiKyHwxv0MnzTppCPD7lJXS80gBr+S6a6q52hCCqygJ
7ydQ+T1qDLoSV3jxaTFIgEiGrnhf/OkxgUcpMTZ21XcCrLTTU6XSm9NtcEYDQy9NMRjCCrQL835A
CNk7J7N7rvq2VooVne1OvRWLck6x8GLj3KCqe3HHWnVGgRfpz9crDUkuKj3Hl4W2DpCTjzYZ2zLs
2IogDHaaj58rbjXm7xbm7Z36lB1mqmdlTqr/X7rlQDHfCBCftXMA5HnebM4IfPChRE/UClnlanDR
8mnSSIyKMihyzSIeaO4rmx6YnEyzjXfGIeZie3Vvb6+SoSbNcFQ0n/wtf1cvPgwhzctNIMsYOnQu
H37WQIevZWlXbAl6GZE/PHHw3pLUZf8eO9jVQi/lqy3EapStRs0411cpIzfDslmJy84Kw2smBFf/
VzgAumfI9gQDGF4m1r8dnhzuWAh8z1df/VA9QMB5CrDqw5j2BZcMYOUCh40DPgVR9p9oE8gAgKsz
ORufawiJ3FysKMV1H5geu7TId/BlYPcE5V6pIXC+mWdDahs/XCw8uwfSh4EcwM0eQGDzV4okhA/z
EP3IgAKPc/8tij7DswHAEvxEfvLobXvUWHZFy69ylC3J5PKUdmR+KFrmELdWCoj2VaGb5sa9dF49
fcnfGbsreEETJC8huqGyytdsKLLE32CQz7ch5efF80HuZLt84cf3DnPDC3t1fb3jvd2DAvMUQLCn
lhQGi/4KkczHjc5tnMn2JltaRRL3e7l0+IOmN9BFTnx1Hs91kYasLjVkEr6k25Ewan0Nln5S9YE0
9fRjTVpm85X8pldS7zIPSeCIaIGzNTZHjXeB4p6RcOkvnYFE3cxmzAuRn2hTyJ54dkWRRdj0slUZ
fQVKhxTB2AF3kjwHB88dApGHVpyfkmXMyPQP8kpLTjj9//KFKLcbaH6tJM7DsMsShxThecPW3JWC
Gkg5NM6F6UgA8amK1s8FTsa8pS4UmThF/mskjPbAiofbKbg4lLyzqXnTDDtTKSiV8xVkU5/M1Yor
m1IJVLk1YC84hKQvQb1wAsrM+sBCC9tSt/8IakRwvFeuVrZUi+No4j6BIOctWEr4yguSWdkXdzIF
wABbJWHQZezBtnrrJiBJdUxc10Rz/KfTWoupRMGiRjrMQ3Y1y9SOp1o2NkfQ2icIzXgPs0MvFI3Y
9Uhls3egZ6riOiFudgGaPzDh9h7PWwMkSGXCNjSqW8+9hRhWcRB88MwSZsWLC+VXC1JbqUjWHJJq
VoK6LH4n5L08TSBv5jw+KbZt3llasxr2616Q1cA3qIsxyK9vEthqcNg6yDnfsDHbUdUuYluxqoIT
xgwpa5PVUS/uZDa4fCdbgRRHHpPA4EXYTaR9qymLGkcrKaOuBja0vgHApw2r3F5dljHWgZZ97GBn
2bzSi7pEZJ+tjzEavHQsW5ceMPQInbmeipPSwifp7d7hpPM1SGpnFfmzWAH58jq1vp5PUaKvMTos
4Ka6bj0UdAaf5USGQdWuni1gACg4w3LZpmh99kaxV7+l0ec88tV0iYVDQf19MoNT5dE4wWFAeV9V
uUm4EuLVuIionHs+uNJXlU4DDHtuXBtiSTWZGGhtt4e/ZtQFAo3Q6n/DurHWsi9xb5KK8+Igj7bH
wdnYtDPY43bv9SPHTzalpYf3QVgICTD4Set25wiNMcQRUdVcouUp8pXcYJGgsBuVj+DSotP0KVdv
VKEp1M6r/uXH/3BQRQLtMGZFrejxLU7IPlPNhjmBHMcxLLMCZJlfPOAoGDss0hHx1qvAbIpam1km
BGKiTc2pXkSjarXJEPWdzR3E484qnk+mFgsiXu5LFJ8SGvwuEzkm1Wm69LLyfXk1B/jBlwkiURKJ
sz+ha6lrrzKxUOSoUQ+0MQJoTgIQb988dzG7hct2xCYJYedGhHJfWDou/A6odp7S2H1KDgOUsRPL
x6giHYKcXVuuDUnk1jk18aWTuKWwLmmfFVVyMcCDQDQpL/Yoc3a3jsyyBGcWyJ5Sfbst6pwmGo/C
Z0L/f+vgAUOmtxKxSY+NXVTMEX0VfxKcf3odEM5e0abzrRJsYbx1sklcx8Dr4uwoTQbJCMAqmn/f
pDMQj/dqOoy9ywcZ600+fh1cIWDli5cEu/mD/cNwNFUEXi2cF/Deoxx3quwIJDRXf7o0lwIzVs5F
eSF90+W/YJb6bd37mlr1V/EJ1LTMtCTbaKEe+RQlT5rjpYW4VLO2paP256lKAO+BE59y0eY9q7Fi
Z6hTfA3IFBWaWviC1/n76fVrmiDGW2X6O5/pc9AIJ5XTPMeI4Wu1k607ZHKAPIWEMAqKFn8mN31I
I1dtnSB5xHnaCd3l4fX5OTqd36sTCzj1v7wicWF6UKl0U17eaIg0N7pUe6DhN/taXuPwHocIGpJy
9VkQCqoLvZF4Pyy9WojBNhcQuEbF/XEYR2Rnqu1SOUWOw03CT/1Vvmgw9S423Y7e+xAxyLosZIip
EZ4oeAYMDaAjtk/fQDMOIE6bVVmTwnAwIYos1qFwbhUwSWXXFq7qdjD3POF5m8ALXdETkc96bd6n
KlyasR6K/ymSY80PdAzq0UxD4RXGormpVMcbi2+9m3s2F9S44fV0ucLruNRoUf5SA0zAn6z46kyd
02p/fj4TpyAsaSfdI5WPsOyqhr45yGhkJwbnnZWwii4AM/4zEbDaRihKKKU2STKvZIsL1/0fTvW2
el5uONVzL9m47R2y4DylcK/BjSx+B0VyDfOK+fqaEX7ZX5D3cVAIsTaWUiziU2mJUsAn2Giz4uXh
wMs4Z1n5dCmjMwHbyrFK0I4zdeWG1w+Gg4rmp9wHZjJ0DDDtKntM/W1C6L+4eMAn4/POrxJWOHko
SJho/8gMYvRi8MMuQi2IU6YvZ9wmSpNhCC+y4EYUK+W6YN746X159z7VCWm1sqz37aVGoTq1lkNQ
H/Cm3wiubxCEF3ypcLe9dn9dhjOXOMI7A3QIPIuzeb3GBg8EE7ESqAFY8XfiNVxfosY6+hGaLUjX
8E4yZe4lXsHorbPys4C0yCSVakUdl9qy8s6uOtfVVOm94AOrBwlz9+8Pe2IP77N3QYkv+AUKdRWy
iDC6oOWxK0pDPAfGl6NGh5gj7YcN+x9ayAzqMztD74w3ugOD9FFHWhOOoaAgSy9FKYfd0nVAHKOO
yb0HWeaL30vYDALjqhcDqy8/PMjGAThQRq86xpI25lM1hGGgTHxkMosij7/lT5KnSvyAjSfJaPpo
O0htHLV+x8sGbRv5u6yizga5nZXGIwKCfy1vwebyKN/TfoTNBQs2YK0QSevlGyf4AMOda8fYjAlY
X3OHjosrccmFEdU7nCzJmARpZFoVOp1e7TtY+EGY7lPlQzFLaaHFZif7ktofmsJp9gC3KgkUV43s
OUoBEDdKMxG1a2IgrQ6xvWftF1OSxrAcSvYZyBtn8oWjnYx6p6DUD9Iiwn16ie32WZcxalaMYsi8
Vn+5QFAzzzqIyoScLNi1KpU3TW7396LKtcDooHavS6Lk1hacA9XGhSllMpzGwHuJna/RJmtBIlJt
ntKhpEkCnbjuX8m2jr5hh3XKpwxmTcQgiJNPDwqsf7agdrD8UpvlmYigFCOvwHVf6AEwbOddk7dt
mBOJsG/oVOPfyObESKD/0gC+xkCZ8+PPRqApIl3LNETh49jShp0DC2YB78qUnFqXIr5kWxl2vlAf
tc9aFSEl+aFDt0aNKcXEY1icapwMG35eLXNcCNA/BuLh9nj5sgVGAIswwYJM0eR20QJ7HUPdxYDN
ssgzQutgOXrLhqHUaA2PxJAeBXd92R8iSwvsr/hktpTx8oKNBdbrXnuiIkYBafiIOjHl2Lb73qso
mJO68zmntEfbD4yvv/Isd4miY1HfyS8aZc/Qw3U/pIXqjFRdGOseW9ahCZIPvWrN0cZ1/bLia/UC
mE+y158IHLeIWdF4kklCuwYRGhi0wXh13n6/YfXcdounSmhb95Bpvc8z3O/is5+hT4/isfKP+nGa
I4a4QtO5EW/arBz4ioMgVSDAUiD48W8OdPHNiMGzMz0pr3JO1XGk2PTdkIDLqVBxCgJB9oFLtTeh
6x+ldTvOHMTRPH0mAFsyuq1h0j+MIpjs7Txq0YnlJY8FyXLMS87kjM/oe9ptwl94XpRA9vsWEutj
Xz7DdqSdb9dWExLiTAXE/EUx27niowrt1dsPwR6Oa80mxG88Z8AKzmbmHe4FAxoSNzVWfkH5fug8
gQnyLRI8m/KtPEbgB3YoDyU/2LBWo/BSfNMo8OrSker+GPQhgJNWfWO9UaTSJHHaNkthH7hVx/vN
ZsVI7r387eujen9FXI0RgVwKlk1GOlOp3nJpxoC8ocLr3R1QeYzEOon29FasL7abr4K0BT2Fqjen
hWhukH7Vq5Rz8MprYCWJnaTC/JvbW3seifIdJvTwJCx8ojpxo1IhebuUbnKG3hPPBB6Wl0Nn16qf
fVFVQrTQgYV5rc5jtmtNLckvL0QlYXr9VUq0Zg3gNbLi9Rqr6ZugjRa51PcetYjtEPxkPdxLaObe
ABPkuOsJg4nrY48bXe45uepl2nOGBsSsa1GsLUjQMmXwg0PevCt6bB2+fYehRe8dhq4CGI7o9Q0n
eRr99HTZmEmfzLPGL/0ARM8JYI8V0MsLTbwPq91XeMHh86nEbZ7LxH4YhtNZEXTVvib5lPS2klXe
YxBWcIMLW6fl2Kg3AHhIwL8HzDq7PeVd2XRmj/p8qRVEnuT4ENBVZoI6zlYQHh66g7NZNqKhFV2O
LwWRCPAcwtMRx/DUnzoqIfjI6rFPontlKFWoJ7eFwwolrFG6gulv5FF16gHzapLzzIbmNEbwTs0n
AZnEKQM+BIMOEqeaTJ5uYoLzqhqlHnDURttPDQun4+iiRQDax09qjxSIfVXkvLL4s9QcgZObyO1N
1QE85nbKQ6X+hEDivNIaYToapsRqgK8+4gZ7ZFcI7HFalUNB+ibjy6bHGziI4FRoreMMuD9qvvSj
Mp5RzaMhZhJdzDKt9s/h2J1ZhkT5480FSf0qeMKKtq5y4Vhf4fpCmH3y6JIqKKpz7ZEMAKHNAHIJ
bv15NCenYebPYcTAUG6/rv7ZBkjIOGxTkJWaGMH3f/l4QwEqh9jeqLcepc91P5wIhfCqvzIbeAl/
LZScbNT/x4mqsE45RF0qDEnHHuwMpaj5Q2Gc3kJCHDCg2CxmlkHTpON8MhWN5nTmIfzWfMR/okGd
P9gHteskruRKkL02yXTw6+BP2ba8fX3ctaAWWNl2Kx136Ub3X5RrfVIJbV2LdEVkDv43urbtsCeF
kl0d+Tbw/uEtZCf8Tu2YXnFp3ltziNgIKFW24FAAiR8fiX+P1HNjAGPk6JvI9YleA2iS+t3CLclv
bOFs1nxOvqwgLFL1+vYAJhyXtqkNofFVgmQ65RyERtxs/sOSCqgMJBm++SCVaCF7QimBv0R92tt2
LuDDKLgALt8Uvpmcrpp/OxzLuB5o4/6/O+G8wUQ0UAs1VaYkKQ4F0dloCx3fyBTuHjMcoQzXzBBo
XR7OKemhfVNYENJgcCTg4ldCdbpaWxv7nNisrZ3VTaM7o/CtlvsPRQFO/lPuamVEpjB5RpibatB+
rCVmLugXi+am9ubeGUxDs+VCYPflG8wGgRygtODjsqv03ZzOEE8mWhw/1jceQQqRx/YENVA0pzON
Vm5fxv6iJlnzX2N1eH2bVU2suasYfIGoMHyR7Y/FkczOb+NjbMZtOj6DXb/2ZT006M/mVKJ5htue
pSWLqaothT1NLgCoDMgC6m9rxd+FMYaycBKztmrW2Xc+MSP3vnvaSO5Gj6L18y0bEU/ywG5StHTZ
e2XWte1/xOusW6AdGNGdD2gbBMKsj4sG3wNpWdIGjQAW+oM6LJliQ35hXjQe/lzxyDa/Us+SgFfY
TGMv8uHVeleEQG0+uJ8Jp/6y3AwqKEEhOEgp9EYsE6V2+gxkP+Hq2GsNbv5qm3dKMZX8DRAaQ+MO
5zMyOKNLxfU9vb0CkZCymdL5veb9XGtSZJzb22+K4UZy0PLPKzM6Itnb73L/L7IK2TFf6mmBdMRN
2fc9ftYrF9aC21Q678XtPHuQF7zI5xCJLMNVyXPF+aRSexpFj5mIt+sCK/zDoQgFmfAZlUnu0404
yFgPrbFrqUe2HePbUCN2WZ6VjdZfBh68sg8La0xqkTycHq31klR5UO+i1mommRx9xMzf/0idcvSu
8744Ilf7CtzSameDZZQG+DaWkwNzsB5zGHjhldCUZR8h6OLKoyh5vVyvYeDzJPgfa4pt5lHAKOGU
I7oJBPU+dtdW8y1HGySLUt7RfrsoofVr3WuqoZKQSzl1KriYnX9d9piOyKPAATr2l/kj4hQqmEZz
FFl0bV4Ut7c5x3y0tAK/yAC4MWu2ewTwHVED7DhDs7aPu9oLs9mdciqjHZZ8bZJTlJa+VydH2Ld1
NIJH2WehtGf7e01x5levtmOX3f+kJmDJYPKt9IdbxKsJtUCSwuIKnFpfzZBQf/xf8bSuyvnvmLs2
1AkrC597XMMryLEekwyqEswOl2ldTsAN1fIr63lItv2Vic4O1aWEiPfj6jSvVrHjsMmyi9mQJT6u
6tA16y8shY96e80JOO5Kx0T0TiNHBoiXapr2AXZtM+PSIZ4J6J068SFI9AMImrcE1BXpduQTuo3S
4/ZSISMxZ6ppI7WwFZwZyaeBXqzNsFIotZJVQ9+2MfFIMnK4sGmu6txYumMxYAiJ7bcS+obyPO+Y
NRX/9xC35a5H4yZXpD6JPts4n7r6NbkF5dhINSiTuO770B99aqlOCI1L3aD0zYetC4ml99yRcDGE
Nyoo/KlZvX8VtvK9X860sKi6rYmIsFiKwXYErK7UyRXScmxWAR37BB7rA3CcHMmvz10ntqNK3pOJ
rtdm9NNggxV2J0Qj4+dxb76/Kad5sdxYzPW9G2DXframcZKEV/1wTS+DA+9wtMT241ZtvDpTIMm9
miitCXVm/REHPCggY4EEhNcYe6aAB1bLEbRfHtDthkUgtVJKCKjbmDHbxc9SiWA98E6lRy/b8r66
oAZPOGeYd0V19kqBoc7Z1uI/78pqU9DASJjOqmsQZKnDoIfyD8FYPX7gsVDYTYMTrvBpUDgkxLcM
Uia+dCTHDxa76gHcpQEa2GPM806QoivBppF0fcFihkNMRX0WgGyVcYf28xDcgOqiOcxwC2Llzclq
f57OIR4D6aa/s6Vl9n3lfSOQ1KHkfiwdkhKJYQkJ/nyz3y83O0yPqNoRsl+uWsvfyduqiLC56AI4
qhFV+0jWMiI6Jwvf02SYNK4jf3cdj9PgmVxnAVGfkMYFJn7t2loCYwrHzA1te3LFJ5H4zLGHZ7Ox
1JKi8neBdD5led2qd/sn/qbVmXRMEp2ZiyvYek8E8STcm8GWD+Zo8zB6fYOvXusBOnRHKtr9LWep
EzUqXZxVoBG7jzte7RPMDwjOz3AHnv/u6oaB5mUXFPLPEXh9sH0N3j+zU6VTPmPghtbub/8PLueU
BDqiFMDaRRbp2JTJ2lAKXR1Tascz/JoimoRXOnsPtWFtxMTvLSjL4af07khEHo+7QMSfEx3JV7/C
hriA0Lv3h007Xa9/NSNXP3RbbpwXBxKhvMvhghhncKEnO8ZiqkDyzCenHH72yv6FLrYNViiRfhP0
Hhjrxf6SDtLB6/euG8FxoGzHRgEFj05g2Ib+Zdkvqk4a+5U31T8KnpnfaSJhOG94k95JEmkC1b9j
MVcX8c6HLOhnOdVXg4pOry0SUR4QnLeWXzTzmucC8F10KXBG3OhA3nCW4pQA1G3HBg2zgQLjYkwE
lv/6iYxGH9H+1efbOkySykas/s0lTs6/xYrE8MsCgHtAYNhdM2PvTjdn70ywsG0BK9p82KyeIVfW
D8BhNikF8dxH/9ihhTEeJRidqmqjQtoFJzx5PRden7IrxJxvil5Mc9uUv7/VzvnJtUU6Veje5+uy
NHEqmmXZ3tlAH9IHmUhWit0blQzac6jYDW6IBpVW4ukSiKvnfR4/brLEG9JJ1MUY2Sr47rWm5lsx
bYDBC2dyORWSYbjhrsO8wtiK3Bre3XwO5nMSEg8P8rUeTmSpBzylBWxigBUdoSHsWA6OiP7F35VI
QAAqAZRDb1Ucc786Wj29RGYxBnvG9TrjbV23/hYn9AnEH9seInkyF7HH++eol5jksNNYX+z4EFPZ
iDB0uiT6Zt3oJXX7n+iP+EdgR13U+D+ZlRBphEM8VSWblwvIYrmuZkuskf4wezsGILYzOHXB+2vr
taUAzIdZ+RPutXYDEgo+YygMhdaG3fKb6vyWvcH3SMGvUOJbcdlHTxC/jmaUKXNHiHUfrXOwjyhH
3dkII9uEwC0DryhrvDs/BQpNtA7dIItw1787IJUBtNMo3XkOy15GTepkP71I/qyHfo7pIWCOq/4D
wHsjplZZbU5MFea9a0CltWF6uKBVbBuJ4EksnKJXW85zHa7Z3+Lhl2wrJzIHqw9hbaf22Ei4ahDp
3zjpg2MDRc0ivVV7fpQB9F7rowsuRz+DlP7a0VZyI7QokAxvw1WBmWFcWRlbVLBhil9TRwNApSeL
WzLDqj+lh5xe6y7G2HCsV4us3lvIwS1Czj9ZyJZMXBSHUCNFW3MFNmgGEphZMnFrObdi+2BNZe/Z
C33Vri5S5E3mpoWGNAS3p5kDpRVzUTfWDL4Jvtrzbb8LM1db1kmPGVxTUaU5Tmfz31jkjVElRCy1
hxXR0K5F7P9L6VKQL6tpHHpXnYOnX4jrXPeFb9QEDFx3x3nIUvgviWDhwlIZ2/WCWpVnqEMsXV+4
cC+Pk2xSi51VfPlFXoPJRg0dhZNmDyVI9ndySb6usY+ppjoedBcqDtxAcCVnN3OiS9HiIqJ/S7+0
zxVnw/VuhJ0hmoXwlC3kwTBS1636PXShAx9SZTstvLoDhkkDWiSeZDWWsxePbPiGFGiIcBwEK1Lg
2n9bqgZIlJ1JgC70bs0AQPfyL4RTlwp8aA6M22t+BIy3DpiHEZ6omwSzstkLDmzajtAwyUtY7zSm
whnuquQMciKEqR4bwRM6/rfsh3zxRGsluQCOImyl7ZsdTelK4Y3icDNIZTsDNwgrIi75ibrG7a9+
8SJDTjSLmpRB3hXaQSiZIEuT33gqeyvN85E5QMd8aVWnHAtVZdgRITaOd0UWYAZeb/zXSKparp0I
HfHTuWHsluRQijAdUsIQYQxLwiwt0VLlAEiKHEUuEBUL4qC/xaZ06M1knAsmpwfGFXAbrJoabFBN
SLMVOcy3OXL7RVgh9OVfmowCHFsf5AH8j7o1OjbAqT9XDu8n7355jrTocxjMACp5Pqmp3jjw0WE+
V1JOwrxUGpxox+5AysRvx3k81SEzVLtieqB/0AoLVR6s9Dm1CykQ57MdyBgn9i5HvkEWwRqm3xll
gn4XUnaj4MrHa8Rqiym4EjFYtEKY03DHaGhlry/RLouWrCDH/YcZT6bgFPRNXMF2gpWKGsCavpDJ
9fpvohOTkShIVJdPHtpwJdptAbJZbhRf9B4+XfnrYVnj5pDh0mFEriyLckcMvhGoHmpi1fXZi+XL
PYx7nyc+1YFkvxEOfuE3ZSnACftGvesEW/3VrfPQWozzyMPijRBn33/uaLiq7TrZsD51I0rQGPKn
n9CpJqqg+VSvdJb4CBHWzeTPhveORL9rTR0U6OFQBHj/rrKuSXMBnqbCjuA8v9ebhKLgr5dslapE
9Mjiulyw+blXUgO0mGVAA+A9WxNoNjA22WxhlQb9qL7Hz/d2EtEE8xz2i4ReCLtoPjTtZRNx2YTg
4k8qHS/9W9nKVmeHD8BtiA5wU0fDA+5X8ni+iuydCoFRZWpl1vTBantYcM+HzN7YKrWD/XfERrLy
u7Bo67dPT/PVRcTk6fO90CA2cMeZUwIbQWmZXS4LBZuAW4+gsGqxpNfJBKOMDeW15xrJrTPmX4nK
KgYtcMhFDLHgQwwBgG+/sgXcPkFWExhh6GTaZ/6QHpO0Dt9YyVoiPajoujSis+sn4/9vO+QbITnV
ph82AHy35JxXrCsQARK9gdB/rP7UmhNcXJawZGzlU5BwaoqhIVUKXJvnGy5CV0kVc/i7d4SD5IGX
opip9Qe0UpKlC+OGL9bb7T79/gKvYCCHjV0+J4tp9vCV4uJMtNUkUU12aD5/jyXDJWnlOkaAd3bJ
CilXunvt5VOy9KUPoZLimffTR4SHY9svnUhZoXo/CFu8lWuLlqnCu4Ja6ci/fKjCAiuKDe+E1/vR
GNiqkKFggd9wpzprl3A8TO3yL1GUfZe0syf3RsXQDIrRVddYLtPOo0ARRjjW9vLI5cphJoIML+ku
ZAfBWkXdN6Jf4dBvr0s7tFqzo6O94Xd8jYzI70Wdzz9vCpybC1fdgGGydj2V3fMYckQSnC3GMbXh
BsY/iVLFXpEYfhG+3lPULJizAQ/B0RDfY3RBpjcbSfD54jdEAzQexC8qP7jkShWF2hw+p1HRiNuq
3bgEuOVenflw3vaLp6gl5hJz9PEuoDV6oRVAuDcfG1LR/QbYjUPtJH6If0htuwkFXlh/w9tEFrEJ
y74OYn8CuLkNNNNjJ+O6CnbGJw4sdGdNZiZ03b0gIaJMPTiXuMMMiDg+BTU+poAzr12TsYj1ZcPk
eNw4gZ1o4e3L/6hsF3ZfH6SyblcoCL5v8agCviueQX2oxSBmSDGMbpyxYNfFJL3Jq9ejV5I+gJcg
/nnw+IYEsDvmsmVjIp1yk+o4cOUWhplJs6S+BuBoorFNZzF8z3K21PkGoNQjwOBVZ6cU0buVk6tm
mkuQMGj1nOn6TsY9LrIucAyNL2bRS66u0xqcl3+YN3ITNcYGznrZpSPoX0ShcFoG8kZqge2kjDuy
5N1cPyoJrH3LRecUmpwV2Li3E2NGB9TmMhvfenmcAbQ9C87EKHbM9bewKfXJ2xUkQGPxTAc5IP33
J2ppW8S9TUNLSipFrnlPaAUOI0YnuKr82VHLC3uXZZHxVw22SZJ357V2AMFzFW+VDcV5aUp06sC7
34e/OCNkx0veD54+JCEmBO8lbAYHNV8Qga5lYDVI0wNw5E/UyVEFq9sHMn7n1FCN6liFRqFNtnQI
lYkx5JovP+jYjQz77tg6sEjsW0uedfRPGdDCN5lCNAksEtRen5DGJy6cHjOEyp24mtpl87AZmCbi
0vzk8YtV9mfdFPH2OKTSR5oWxATa6xSYfrjwLuhjADo2NZdr9KzzmbFa87F/zXrl5kNo5Sh4AgUO
MZFAzdvOGy/6RNVr+y5v//akxxjr9Umg98BaZG4il4jsD6x+JsIXi/J7fln0M2RrD+dXyPOJWb/4
u2ePyASjFEg4uCcPZLECXs6qtPQElATn483zPHmkzWCiekt+bjDGm1bSne9sAtEqPbaIlwPRbQJ/
8h6hQN7xiJ18tL+NpaWY4ocxREbZ3nDQCiefXT6s3QQojcX7ZKct6tENHGKfPc3NkF88IwSDTaz7
84N22Wa04ivZxGGTsKq2XUqSl0CFq5yAVDX1y7kAeV7jjVGQ98EkdjumjHh3AjJkcGoFIoWaPCZb
NYDykrPoraVouVop5s0CWn5dEuPHG8FEv5s98mpC/XcLAen0RVvzcc/3C9VdYnpN5RkNeAQpSOGb
gMzG8IEGWbsriCUMAq+lLrc7l3j/o36bEPzSCbf4ai/6UvkxldaOR5zJEy0O05wqWv9ZVN4zlTP1
maBqE3U5O0lByVLkzOlVXm2ko5z9zROqeWpJ/E5xk/wVFfRPCS4XdxC8hhjKk8AN5Zqy6ICkdFVL
0xK8IJtOrw2qLj6p56NWwPj4b+IWFe5d9UwTXNqpgrixWSNQukXZyHvMYa3kBiJs7vVB3mBvHNTI
I7jancy3fOGRu9NiShH2NquntQsk3LkSuB2HkzWvf6CKXlZ13ysyEzb9GPDJqU/YRGdv6JedhwjS
b24bYpBLk0R0yQ5qhq/b4jK3qGx8V1drEFtIce3DORQ+P1Jz7HBXT1zqWJW8ghwKnY/LnG1wU+Xj
QMjF+obqoml7KFsfm6cLssV0hZ4zI4emdq1fYS774OZugocC7Yd+ynCZbqBttl5nIfD4kH9s25p5
QF/RwMckevt5E6MPMSUepPLaLZ5CpD5HbOPc4nyO9EnCrBc0YgrKhtY+OMr/3T4FgOtSGfXefMf8
ImWnSoEvRguy0xUSaS/LKZWg8a59sq1SOB8LyEsF5FGnl5K/hjvriKRRx72mi39t1ZQoUG0/nrmv
3EliSjJ4/hvt68U2p7vTuMZQAU0dyADtDhuLtyrjBIKdYLfFm3Imms1wEdqf8oKMDz6l25hEk+ir
PwoVt/lyAGdoA27EJhKFkNlO3gRcZM2OfoFtppErMWqqXpOh6ZAhO4sn4h5BD/xYCEDi5hXgWuQv
gs3L1Bqu7QhwTgD5OHJ1Y75OGXXRD1MTDquMqRvMpIqV3+A07ZsabWgLPTEKg62S6dYIlTuuhbgz
mo6HerB3/68DxHEjtaAwPHnjqcGQaHQA0U5PX4Of4vE65JT6t9fymO7ThLFXUI6GZrcXwZdnz+km
W6FXkJHgYyoow1yhkv1TXJ1cfSHUKKVYXg0uAJX3ElihevcOuQvWxWaO8a9LFciZR8I4lSDEaOiI
oyoU4nQ6EU8Xq/wo9ivkLTtUmopLGRpKshOyBkq8YMiuim/oe6n2Vi/O4v85qsCEII04Pm6bei1b
rtQJcPjRnRGBt/GGerakjWjxoYFROMKR+4cgFQFgqEaRA9uQQLfnyjGdYc1sxibrHRmHi9HcpQig
ag46fGzLU2238NPEeF8bhd712GzzXDS17wcDV3Rp7rvVMocrVvXfC0lYcF6MZNO+RTv+2qamGcCS
MYqqDyhTyvxvv0NGOTEPj6gf2YtnYRENMqhN6l8IE7cS2i4wEv0lTFAn2ratnVaA/J6s1dFH0oUj
HmrkCwGY6eIcgiQoqGC/sdzVcEUMCovL24WmNawDJ4pEYvjpOguHhgN4InArRqXvXxLiR/XCvIQv
RZ6sAmegLiLwrxYU1RqhVMVjX4zQZblXfa4VtmYhfDbQY2TyQvELgj/6eqeSbh7OWL+kaWkwoqbR
VLaW7awjKlijI68Eovcu0RcnqzMKzH2DD+iyQQleaEmnRt7FNpz5tPZMvDYHOveQI6VXkifFRrT5
feIR3xyO9RG5E9GphYLo1yeIdsn4JevdvDJThWgFXNcYhGuYLNRgttqpLfW1fNCf+gDF6ap64T9O
86+PGaXrfOcnkEyULIAEt1bjju4/PPguNnoWMwAalxwfpfSMr71KqIupm9fI2iEZXYHqX8hM0+52
XYICEqlPuzWy3+Y+Ezoao9WAXPmprWqsC/RefpYpm/bgivkeAtTK6a4QwrzLLcPiOvM0v4FSFDuR
VUwy4rewhixuJK8tTSiTi1ROFT72d2hLlB77fgmgn/OxI/Ev5umxoS7TrTk4l36mszSrflOjmvRs
O+v+wON64xQS708hvJzg3hShGqBjbcFEg0ok/MB+iZTOhbDplUJeoP5MGAOF2pWNEolZxneoX7cl
go9ab3CZmWD/2j4Rp4YpHlTH3yPDLpqu81QW+1k2hUstixbgE5LMB9WgLWbyqUlFunpmFIf2LXO8
Ejz8bQdohyxe45IL+LSiWW2PDmp2hPHyzTWENnVNp5aEdChdR+FrXlIycCWXVlcLyXNTs5n7P8EI
GAm962LrreLBTP/t09RtUbYmXRyvXmNr8a6/RbYhvS9S6rGupaZ2nWViSo75wFsBYlFVwrijZ8qC
G8PdVKJpKEf7uQpVtUXU2ULsn1MaSd0FWvkraAuGa4ztlTIQSbsBoOyBlatnNy0KhAM/8i5lKtnJ
E1n8p9XYk3L2ewISSSKx5eTkdp3LO85P8hfftL6mP5gH1RhQ3ypjSbliz9BOrkDpvfYmqc/lanVc
BBhJ82CXXhnxXhJqqtTKgxchMKuJzXAnYS9YevICGQtGKWFxZlfkdLqRve8p+HXNTnifF/UNCx+A
URBVGMEFQFD11X+XrrW7sEcGpOltlHJbIn7DbY68uuNOUFaB7O3vinkre5j/Laj/KVRO5VXxXm65
nZCqA+pCCEM6OM2rF/RinDcge3R34C6Ws13LCBpnZ+4vNd8TobB+kCmEgNPa1YQ2z/vfvcBpvM8g
3+m4UYvmbaYHu7VqDiTs8xKU96St2zIKuKX2Zn3wMDTBPZy9T0g6axtfzfmkKYL/dXCEdbX2zTOn
veF/5VpFALniZ5FlOee+KroKo/MKF0JrImMK8tuPgaiTkVHusWMk/uxz/VvLRKD9i6Omvq0KQF6v
rKYQSKanYlfzkjxh3ityvByYj4fCVOCQfCKHjDmJlAEkTo41r4JHAW3wle7Asw6dA9jSB73QRdlD
eLbQBs2hEu5oHquNOSkHcEWzvGKODmCnogZmoBersdRho5kaZ0e9qQOUsHacHX0yMuL7JyWrvA8A
XXt+3ywsfwgC1Bl3Y+oSfmrdYJ8yR38te2t/zkmswNxrX0F6HqpXb1xyf2GE8ZvnTwalI3OzW0hS
SkfcB5XZslu7NCNIzJ4DhakGvqMtTGzIx8dU83O7eYGLCNlLyUSWFKK/lbL1CUFli5n0ILFhQK+l
PWLwiQQe9ITSYbbL4F2qK05q0IbOJVc8T3eIRAJ5sZnSmCWBQn3RvxtxEtpV5EgdCq5LIPVuLIr5
vOBUznUaBJz85zJHjc5bnr+l03ixP2enrAdLK7b53j/0zBpSmcEfOZni/GyVcY4WrJDECWUAVtX1
zoFiSB++lbvMx/yVtfdDMrzid1VjML3/vw4FN1Rq75QjzgCWnlCl+jSKrNbwNK+RclrCx2VYwS04
G/suTC4QvG/WOHpwEGWm8zCQeHBE7SDWkOy2pAT/w7JJjTia6OyDkLLC1+rQYO1xSA6Gc/ZR6tvG
x8LzRN8dNCz64fGrXDVgl5L1bPrU4zLubCA2wo63XusPLEMHdzL1hwiCGyftfITEkrGPPPzZH4VX
enmJd70xTydKyrI3JlC86pKzjCUkmyTvT9XVKWfdbbyU6hRh9mhHP5jrbMaVPBlSnszjptR9Z9CB
CCAs+4PZs8Wz1OCvQmQ5xRWFCCdF7O6pAuVoHJxoFUDhSH3fasSUcHVR2dECDfJxkyM3073JYwzd
xggYMg4qyiVr7OYomAANqSTNvvfGkzt2u3HV3sc+0HsYVq3HzlQydL4ITcCiC67lnWsSAixiDBWJ
eqN0QA1EqErcrqCalHlqfIJCrSKsd5TDswquObqrK1f1XMRJ4/P7UbXJ4mZf9AptBBsDlzDB8KFo
+CF3pwB7l2KHqEtxUCXaI+XZOsOSprhLkLEkxYnRRcnwP0a7jKsMoa06g+NjEMv618xTmsj6uSY2
kUSUbh3YJmo52D0S0w0ISGXumYcBxZdylQGdfKEHZXOMWegmFM5hPNKRJ+mSWbmBysAzi0Zbt/F5
BghR9stYr5x1MgtMXxNyUJ+vjqASzJq9vYJjV7cQ8Q273sCdK5ueEB9eBA1yrkumx1oCfyW8RF8l
S5y7Bab361xcU4Dk17pnDYHWNH1vCXISV9jOWTigSom9bgOsDTqkdAdpOM02VSXRTojW6brA2hf5
LOX5K1jq1w9oHZYz1jsORGT1bl9ZrjkL1VfhCxcOrnWbjg3VdGx+RTFFvLOIv82UyP+or0dgH48R
qJD4ccozCNNenZp8bpWsdT6/BfKgPK9ZqjhMyahwsybiAMBNNBIi+5jc/6R0vuR59ju51u+aEliQ
Xgb0YKMO3T8nVtDqQbTTe/bg+piYWXzrVKNxIIp/HhTFpYarEUy7A56eRyUWSYvYrYlc+BmsFaSm
TAD8F3UiqOX6snQ4n536bA/9UfetzSnmcbzJMw0fapMqNV+Xk5Kgv9L2rgWdNbPnp0gRCPEl8Meo
xrZaJCVojN8JBdPcMREJbt75ffVvlnQXrRsZVlzNw+zjh0q7/z7hloPYfloN7FY55sl7J7r+dOVm
b9OyZLJO9X0QCEus1gTYV29IxlQ0k2sYdrFG214mIRUqS0kA1rUn2kQ1C5TmPooIXHF4njH3KgcO
QPArBKFegppUSyLXZhCklT2fE27ieDOeV5Be9ZS5qjj3kmGIzbysKZkGOcD80Dv0gnxnloiLfu6x
DQ8vgIxlKu2/JaXptjl9z5LmYc1qIvulao42D9+rM8lJTdjysb8rhgqMeLsYDUonThejVO00baPp
XQbgtSItivGCM7y2LZgWJ6SJQIebnYr+cXW02mB5pYZeOOLAilVg01ws1XQvkf5+R/HLgk673GC/
nqBfX6BNRcDBO38mIjJ63CffnM2OMxWkvrL3AlWtv6LfVzSCZzfhpuNTzeLDXWYK8lpF1w3aQf1B
Q07xhIq19vjsVY9O2vcQY2btVwt/a4pyZ44/kW23k+IC4iPmCQyF5jM+Vyvt2sxVcE4UiEvZPkVO
s7gUw4+UP+3Ucy9XeTexLcAEx7pTv0H/MHgH+HPQ6dsV9qFOr0pD03rf1p7r/TO1XnryK9hefD39
RQTHubxryZnJm4Se2MV/9PTwl2A0JUH/XDoX0zukB5lzhtGI59krAW6f32RTuvMbRogKnCqspozQ
yI/D4F2UgG2dZmJv2M1pjDFMLBz+cakicQz/J4NK6wdaLgOOxobWJQeuYilT0Y01OD4kHxlgZQWi
BVASop1+U/7rrwtHOIeY1wut7ZyT/VMdbSCelXFf6Iaw9Y5nurQqivHQ93bLvOkitKuw11vI3SE8
R5CUoytFl0CVbMpOjNmwlx9OE+pHWH3hMcrOlhmgKa8krKWzYd44WOUtTPBMVQXcKYDdFSlkGds9
AQU5FtkzOD906dg0pkZ91FpHpwbfycKYZT8O2NbMnCmsM8eaUtYkKwtIf6mWBp5oOobNVoeyUpOh
1DLf9Zy3p+Bb++BV8MyEEZj/vpHlBOw6R085YzAFOnCFS3fZSG2bjZ1h2kP4Ty4DeQXzEgS9AQAu
NVlVrG235IP8pXse0IbwEKGRj7ls/+FoCJBTWdPjxL1RC7KqG318FVmJxt8gE1Jze4WAvz/QiHee
y0JTvpqrlf07VbFmDBtvslekNxdNlZWMexZQc1c3V2GJKNtzz/WkddpHzeChDi2PL+qreuibumbA
KZqJALqe4SWrjC/05KJOy86EZbvOxoxNwV904y3o+1GwrQid6Tr2tkCJItU4ocv27dDqM63nB5UT
qqf3RfyMb+u9NMKnmt9nJmHMR7rs90tVhlvqWomkpp8SsmETA9xbqYM6sEf2G01QYJtgeePzcLSi
MDv/NBGMCGbBC9Cir8U+OT3pYheSqRuX4HYh5sCRB9x6VEh1A4eLIW0G66/2Dk1DK+2Oo3dHj5Pn
kj/9/en58HahekYQYefrjNYkYbKFM0h+JVScKHvTtLXERAz1suhu5BIwibGDRSg6LI4tMsfaOyi+
uQhSGVbE9lvLHKTzNG6D1ChtYcJPRtVuARXARLyKUpwuvt6bmvOGoF7qAMV4G2qxEyr43uGQbKTj
yEpkTSWicSV2/V8S/3pnK+4ZJJFGZq6sm86IyMzq6NwVvvoSwdKxI26/qgP/zmmlNvTVWxa5CmWX
I9d3MP4Tfe1cwtxyZs4UlfeJJllmAifBll7XxjU/9jQv1FgsL0zcMLDkSR7u6iahJAGRZTH4trUY
6BThU1pj20zO4hwUHWlSTzGsNyqi0FzLCK7Xl3tEMAbLf4JN0BevlAO3cmszY1oYuymxpgC7rmrc
3hkyMzUJ2j+0ty/M/EysavVCxEixp17xDsfdifFVduAFn5WtxufzTsjwTuWhxgAfzhlUGrF8PBc4
mNrxrKIT1V9cOZWHsPBZQnsPjYe93FZwulcEAnKHhmtch1AunzkF2WNwTXnOr015gbnc82aRcgVG
kwWA6vS5JgF4pJfugeLXCJFWlK7FhhjqgS9KEWRzahgHMNIpuwT1uIFTXGSlqzBHOu5NhUtaIcPt
CzqAgQwglZFIfX6hH90ChdsYsM/C4L6PvV0PKn9aNyC+mQOd1sY/lfV7MKHRJEX/SdYvq3s07P+n
ks9ZhY+oKti4oY6asZYGTEdszzcxHN8zLtCC50LtzbBKyJauWBroZE+oqm11dAzjFj5W34Zdzs2n
D1zeo8sNV9c8lJDlNVg8688FUlW3/soUbrtldypa0tcHFvOirgUWrf0wSmt1S4ns0qrFCh+hbHsr
4TewKET9JNHCAJUyJJtkaBjJhftOWS42Tvxo7hj6ngpatb4oI6jobTMOTV5aIGkvM5V7ZOk2wlbT
fo1VXxrXf3R9hw3poMAgM5EpJKPkMwdGsujXZwHxcpgnBJR48f2qb2rNnAUucj3ue8ftiLNGkd9H
N169qUbpWzRMFvCdoaCegtoqw9cHUhilTx3TGYYEgSIxlugQi0jQmXH963/SxcBO3iJbhhFAPw49
y24k8klz7a+DQFXmrtjl3uWsNtCsUWu8artFTjYvX8E/aJNrlzu9Ztb5hlwS+wxp3UEThdizYDC6
Uu92u1aQ0CbSRWqItbxWVtmaajx0hpi4YcSbUF1E4j6D3MQIJtjxWy2KqrBYmYkH7mnU69VWcRbf
Aes08IDZpjgkvObce0uHv3ZLWxAWLTb5nGBTAmpbED5gW3XTxs1usA3P1nDkuAxUL92ILg8QnCXt
dX/KG13E3ZstI9I7F1Fr80+2n9n+snAgnY+3zvhnC3osCBWpX8smlZigOrVOAi1kRzytfZyreXKU
B3Sktkqm0VtjvBzgSO0Md+K/Cxb3PgldJUAsS4Vq+mUX4R6kivY+tlwM6zAP5zegk2xe/WQ1tJWV
lnPHXzfL33cnQvW0EOWlVSLnbWw3bDCl5UbWcdfg+/x2Ro3A1hNdAqM0qqaz6PeZxvpv2GwnMWSB
BP0dPK2bAbu2WowM59Otgx21SFDWe8XU7bIGcp8tsVh6i4zfyfXUxRWcJkhOjDUdF9Yzpa2xDX8C
o+oAE5Zk4ZBhjWaOHMdpU07WkYZB/WBkX6no9WBK9lVzuE994+1mwHc9vsHqFTnXPTLIWvjHlQ3/
F9XEPpoPRGe0dOeeMa37IG5gkkm1228ftW6YbzqYCSdAX7bhAMw0UfNoOqAFEm6hxQBrlZv+T3aX
UnGJsuO/5F4j8CDgw6C1XiFf1oQtKO2iYMcNnHrCZuKu2njKTE/EJEqL81cNHKnuBX1S7hi04R3y
BgD407xoeHzAND8G+Io1+gBrbSzY7xWmQn1Ye3tHYq7R2caLUDU+F0mGOidNycmLcq4zt8l7suGH
2lbqy0J79YSgFmySVtFdSAsV2DyR/X7wg7leXKYSFmPFRnp3P00Mib7wCjOrwjIsFDPq7MwdcKQf
b2SRZ/3t39owg7BygupZZZ10RtzIL3iRVOnUxL7rl4jJTSRxxYkVrK+MiBZhA2Hj5LjUDadPlMOy
DwKwPirpHMKi6zBLK0aeqbQMld1I4hYiIcy4NUu/TfpoA0D5vWvdaWkf9/xxKX/ggO9MYhvDSLXl
dYDpC4q79qVjTxWJPVt2qXMNSIxSSn1jbo5wv6dQKOkapAt8DD5QQchnBcNDiyMmnp1M4kyUkPmB
75muB9HdRBAavZ83qep5PKFYkBiAc0ceeuLJ6Rss7z2eUl1lmxRT3Sw54F0WEbTXCAN5scMCENuc
oZeypNvbgmxaRuZz5remCnYYi0etnVf0aZ+XhQ7BjRpw9CPI/IqHa0vSjTx40wfwYL1XTNJV1jjk
iCCKtk5knmIBNweNf8Rcnh3v4MOy1p/oytH99ELlSQJT080/QLEad7eo2UKB0c4U/H3HlkMCN6je
ILP7uGxJSXUFjGcrvSM5DYFrhTqIUTNh4kH8cukcLGfCrVwXbkgvxQpq1Q46WDzIl0DPrEOLYxAm
6znWeTm9JejSuj09wKK1k+DHu2HK9f9hbk5J3R0XzFnJafK4DVzIJZBsTCL8vu8867UebSy1W/aw
RMcCkmb05W2pQiHS4Uv8jbDdusnWZOxKzb4jMODY8PD17DND3IQt/uem6lRSJJ9Saer+SCrghrUX
GQxmwzGnhMokOy6sQtySRQse5IdPnnqY1lRK6dEiyThmwVh5wnJGPSUuq8PLXVnr0TUulCIFW/KC
+e6SoXjCRdexOC+fg+5hQdR+0AsWMdOxqfdQnPS25V3vGHfrH5YeH7lp/54rj31bcP2aiPpbQSxJ
lFAGhObjnHczze8o8mBbDplg+HKbMP5P2Bo/MsiojedZumx9wRBo4bvHCPRt2Is0EIMDggI5uGFW
pDObQ8ICkzMcx0J9Qjs5LGZ63T94HBPWX7pmzvyl0MzSiCCBlnAN1lVWZoLgDorhsD8DtQjHHWs+
i2QHlx+OA8qxqefHeNjKPjBSWapg6T1bhyu7z8y+9sQHjk8LGwuTe4u6idTKsejseQ+f+ADkkuvL
HcN7wvTPRVexLLkl3TIQRidJbVVdo4r5xc83E7omMaZhejFW9AKRElpANsC4JF6KQkm53Qanlp79
jRyPD+MZT4PahpKTCkmrRkQxvfXvBW8l3x0RxWijokVtYhuCR3PE4ZnCRO89pWuufY3GtKQuktjm
gTEoOdkRF+QtY8WBO356t/+u+sPws7I5cJC5VuovjcwZs2WX/4xKfLr4zTqWEufHlWXi5tBeclry
fjAPKekza8R0WJnlx+YnLnxT8uHVNJ0qPJuHMkctqJ+sV3SnvMk+cxoJIJy5/zC7hXZAuw+QnpNH
kQRYRBS14MtqAAVAxhi1eFxzAYSKvpRxwIah2O/jv/FIpKLCScj7DerOo6pfpW9wH1prlC9KbaoV
bk7D3DBczWQMsZY8aApEnRrc4Ec1HqBKHIf57dRK8h3c/4i/oXSYUIEtW715A14zSg5yKfXHrC04
vN/a6jl6lJrc+9B27PBIbkylof3/MwRvh1+VdJVpUUbR5+DaxAiRWr7XO51y16itSlVGqczIbV9B
x/jiMu4BH9rYonz2ISva6wnbcp9GCRi5hq391+R0z/F3jH7NJCxW1oMoc7DEnV928X4Hky4Jv5Bc
F8NDOBskc9thYazgNzMNdhxMQxPFxnOUjEgSZUqJVeWNyJchfZH0YcE/LnxnL453+NRcVjx2k95s
kR7tUGJFj6SXKf+zatkD9ZW5HfXT39pxTJOfr7V3c/1KfEuCihB8Eqs66SO3MBMjsOlXniw6lfPP
GflScNLxlZ7lJG3Qo5g/CyW/zYp8WrqR2quDO+rK/PPcmpdeEzDz4zguiyyyn2aoFCUHQ7+StQZD
4PeW4L9TkitUv+OqKjIQ/fj8KOOXBo1jqUoyqmhxc/y+9DHFPO5nOwyKOuQuSJ8kVEeq5cA9RA6b
l1fASy6wgUl1dM9UhEv6Y4wgbAmkxbGMvFmu8MTMgnv+swU4jXYkCo8578RQkCosfLcsGbGFDwa3
1nnrlfadYYBu24UULI/dAtz5ufxsnJMyu2uPlFFpeVO8LraLHFU42nq8QO6S9Sk8z7Fn/YLgEfmb
zaxBCOaosgcGxavviIdNVC/4yYs2bpbNu5nC5YVA8/d1y/qjklzkF47nqz5D3PwHhuWOqhG6c0SK
ZSDez0zpaseQhB2+llL0kporxth521CAiTlVy8y/S/TK3BWaexuE9oQ5VS7a9HuwLpW0eJl0LdsY
vRCyXOZ9IzusHAKUAU4Vhmw3A67thO4GHXYJwoLbrq1VHrPrAJ8HKEibKleRGYjccELVe85vvIEH
rg5ajWKUcB1WD6R28m7CfMqiq/ymRVQ4/cO4ZfRizjC3Dye+hE/sk6kRAROkRokpqP3kptEbKuBV
JFi0mwSSxbN0PBmsUXZd2CGNrxcHkctt3TnlUo2tYzOEQnGhYwbAuU1OxJEu6bbvsSs1D8XJj5ag
m+u80I35av21xuOB3CzSpPfWTjxfh9G1AGnnBh9nADUwoi/dPOlnxxXYtmNoVsL66usrb9Q8LfQO
cJ+uIzE4XMg8xPPN7PQxaOXa0bJ5I4RoeDd7ZI17cQmb7m/ncatUv6wysRHnWCDIWMrIEacgh1wv
gSU0lAKAns+Z1dLB4lFCCkFQdB5Yi0lmFADESaiRIDt/yayMQOqlspDOaAVMqf/bvX2o2a1rm2YD
b3D+zS9rkmWPVw3jEpTHXwaZSApl37GZnpJk2HM409TWu0TM/h67kLn21NQA4ATgJ9fDVBsU5gJ7
T8WqBZHbXE8pCa1zqeHhqLHC3u31Pi5xPQbmnkWakZqBufDuvb/VUDlNztYALGz0rkbVSyFrPXUK
UOu4OVg6trsW4LkHBEgFjUjRpU9VKoXp5sXZs5aBbWoid/cd+hnw3/zStbAL0E3hHFkJXxGg3JW5
Ym6FQxUUAOf6L1KvCOcJKkRzRLkleYzX1/enMdV/qyQIXvaNNCJWdI0oPGS8FLfPEFSPSJyzrLRM
KO85lfvgEWPYsfYDzVgGW851PIRqk35CP3aPQygZr8JFxk+Bx6BZZOLwSYy29neEYaZLJtDPIVyt
ONKl/eBOm2l6sxDpccHD6oXnmPktf1vaEhC7knVIUlKQ1NrDWkUXqrlQWsN/1OewDScOAWH56sqs
dO7kIStJioDRIM2GyQpvG7PV2NQId96PgOJFs/tJOJcfhnjtXZ/CG5Kj0lwFhvX0/K6dXvoeKsdb
lS4BESaj3DDE/bjhroARNGkqfi3H7ottAJyCt7Z6Z5j+4E8506oyHMyG56ioa5lNOqdNnXlhkQNs
dmjD7f2YL7tJwdJ/FUX2XbF6OBwz72lr080tapksHMiOozlCVw+ZQ2AUXqmvSiRMOa1giTW7mjzD
3MuEqXDt/KFRe1M22dI6f6/gy6NA9of1hBhgaH9nl15PQ9qzwM8JoEMmzsVzVisfRBHT2C3neBg9
2N7uQVD/uJoZ29RJ/bZ4ObW+eb+z+FKvEFqtscwSjkeuajpRLNjy9jy3GuAZi+X//caN1DQinGld
rnYTkkqY7TAW6Bg7uGiRn09x0cPXyhpzVtQKf5BoL7QoaDEMQD6mYRt7oGLIT9wGXoWN0zocOmDM
Bvj8dhfEIUTzv27l6IGrqrXXRC5UuI+umbSW4q6nFthlhoeim2eXtv2uZVfltgi/zeGaCJGqkFbW
i+V660BKGgfWbsRgn4wIEdDuQKHJwSz8OODLxdvl2/TvJlnCmnYTeQ+kXDPHl5vE4mfqFzQ8OZD8
64yvcRUU7AR3UvHyID6I+BCg9/H7JvZqOTVbvHss8ZMFWKNWmWqfbR2ej45k0rVjLAhFWAlfOe8b
oxZDaRPW1eXIMhT3R6nVesc6UyaVRa3mft+F6MOBubyvVqu2pvGO7Izvz+GL0p6XmBv/OkClazTN
LJLjh/mBezGPcQV5pcNv+719pWhoQGUAJ8xIA2GH+Tp9Iidsq9jO0WWiifO62E2Ma4ppw/jUcY1B
gLmz2DXYab//ADZyMfJF6R+hVsgCHQ2qv9EOODGb2V8gJuJBD/XGiJBM1jwvWXEWjur9qq9Wv8Dr
huvTkeK0x86AmFjFeKQr/rnA8A8xo3kMlCWPsKVJA10yr+M+hxo+D0pexhaHQ/07ynzVVwKKtP7D
r+vjuGTWsntXnhZOQmFXnRDZkH6fBGZq2Vk4F50YO+69O/xmmKF+71Ewsu/qS9Z9OlgILZ+9s/DS
s3MV2+Af8cFRgY9YMsHAupTUa1Pj8JgcKA4J38y0KfEtU0qQdxNJahTkWLYukurygNmueqkOSacm
yHVfFNNlH/2esbaGGHiFupMNdaaLXJUhxtAgfY64U/sy/dWRFZOhgiAI24f6BrD0du8WinAcA44c
41lnXPQ3y/yrJEVCruR0weXQzLM9vr3pfAP85kJ6J2v7E/XZK3TQwnjcN0Why932imDFOGaNcCmI
RS9GOvpNnpDfXd9Of84tKePhc6jJa2AMAm/pjTCSHdQs1DwEbvBkq2u8gNZ8gwmzjq1pAT78O+xr
ivMCHrnhloOog74F6wPQS9uHpRIlt5GA1ZandLlNrvARULaP8OTGz1dQF8In/k0Hi8hp9zRmBFce
NCSADIjPvQHwhZAj6EDwE0GT4hqUOrkwt5w8sqHqjb9qmwS1njEnosntdou/vMBtP6z/TT0PXnQp
h45EraSrT+9TNj0FYsBvLseHA83yAGdkJPI6ofcql0xeIamK8Uhdm331tcT6aA9bwSP0OVT81kzn
XNHgQhzo9ZqNDyub/pma52Te4W4AAG1wNP92LkYFodfE+zRiPOTD3a21AtautMY0oid5dLtElIUh
HtX4BE4dO4cf4Hr34hhtxOwZlkTGjXK12e+aIIFoSi0FLDwxIQna4w4fmqb3aQezfbyJAmAyEnRa
DPu1Ugxw2MJVy2L0r0K5neSLGzeVnx90N12wcOy061O/P/Ou1H2S1GwC3hr+TaVmVp9/toO2oXgI
+/+JPP6b5iuhSSM4O4U2vPzJTPrgvW7Ejt1Rt0RSouKv343lKiifaYIUv5XkWnIQB5HtzpD2OkPd
/U69qqfrFoTUFUx4jyE7ikyJt3t8ya2Y6Y3Nx6HGSU1kbWgZUilJXdABOR7aWLNq7+KyB+LypSI3
cF21V8Ns2oO8Wfr7+wbUMo1+N3y/Yc9ivIpZTdU11XiMaclppTzM/YtbxCNtl34Ooz/1PMYXDMaM
Kor5ESi3bOd1LeKJffjAueZxp4ISQU/+2JhadJ9koE7M/JrjzY6kA+GLmADO3s1OKSyTj0fUTwRQ
BAhpMHnk6HlmkAzMz6Fv7kDiqpa2uIc/vePrekLkDJ6R1C6bsZ28N5ra3C7FmjJZpPEKxja+/BS4
5vS2lif1L9l8UDWj1ioWMZJjNkAM0aXoVJFRI64N87bfCcr5FRimy4LAUGVjaPZ8DBuGZeXGj+CB
Z/92rfXTY1Y1eWp6QRzT9WMhR8lwRGVzRESBabzQatWKGNj7m2e2FXhObI1lU8m98RKEtOTsS7Ao
h8HO4wMeQtNlAtixY3HBhNQrauY5BfDylzDIP5L0+qXvPLUS7uBL2S7ky75ttmBrUgkHzoaLiMA7
Dsp6WVbXea6gfRvCT0FbMoz6CDhrd30dZT4ZrZqL7KtbhpUYzdMlzXoDwea4Xcuo3LH1ToCi0Sg4
7NUozj8ZK1aY+uhX827pc/tcvtn0DhB9GjK/UhXAIj4N7+KLMVay34IkWH4XckGCBdpBplkQmQbt
kFu1oFEcNuNTjTUP6fR5VAkd3+PEqoYDkPIuWwyGFCSh/TbWBBRQqnYzJPuuILH5ScLzK4lT3UxX
k0zut6uTjU/XHe5YVY2kQzggCmtzRje6TG86SVdpSlWPfhI56Y/pPdK+MytihdIol2xHizlGJSH/
BB0hwKK9ZOiVuQfseBxIZvsgfpWom1oW4vmHk9ft2t0mdHSU70MI8aiw2s/Vkzfxw72lnwXNN+jN
c701BmGtkYVgXzHeidUcQIw+YKvIk/+i1Aq6/qdk/CzfLIslyd/LlUbPSIC0ULSclKL8IF2FXTV8
46JoFV4Ue5hHQ3iIWA8QYh0wvmRjykxpgaTkb5XB7RaflKUmj3mSFEYs7Gy9YBPfG8iFuQpNfCZn
0NLUVUVsnzV7yS6aw4CiokYZz69CZJed60qf5JaYxRU9bgduwKgnWwf20R1QKLhS3/trSWCrRzs/
H6GeToaRUFim9xrlhqNqsmvDbRpbemurqWvz/FpSVSRZcQ9FcGIVnZ5+PFwL6XV07SuKY/Yxl4Fe
WUdaN1pO5OMqWPNjG1pPjM9LIzwGJy7jYj0x273O8V4UuGrQFz12aYk1iRlNSl3ZZ9r4OY6EDoyT
jAJIGTNzSOvn6AaEJAWs9uIILDCav23opwzCebFIwCpsTUchJ2NrduOeKhAY6tV6or3SnfGfmwik
N4dxt0hz1tgsfgwsyoJlCNruDzImJhiqjl7fS3q11aHxc/bK8dzelEnkyWrlagcD5zJ03g0ZO0vk
qJJ8s/FjWFLRjLgU8Z5xQqRZ88A7z1GYUyV3WxveSNtLXBahGBcV7YzjClpStTI/JVl2qAempFg/
5IxrZUfi0lnJ/HFIqxUjm5MbchI86/K9+Ta2r4JoZZbSXVqQ/GFmX67h/irMi7ttMsuYTcHjitwh
KWmaxZv1prSp/OU4Jt/3QikOAmDxauYsJmI820PWTRe1y4Bps5viwedU3TNUQwlJ8SZvRbo4BQ9Y
gZ3oOoVtWjPMksAB2qapdhnNLvEWLcZV+CKNu52MwM3wjBIryuOioDOHFNuRI2cCr88VaT2cB7+w
BunVz9ZPfjovFV9jzCSJhFpPKpaNdfBm1t89psgfjNtPp51tSsfVJQFlAKOD/VkH2X3la2Fut/80
OyVlrjP0hCVh+JKcF4tdKFarq3PceXDVHQuW+5A2Di8HIyKMkwEGrxUvtO8QCPbZo/yt/jG/vTe7
3fqr01EBPIpkbxSUEA7UOWjT60HXBSvuMTjQzTVG5w0tIwQNr72R7OL7roXecIFOVHBztNau3TT6
DvMX6c7e6q5k3zuA7X1S+UXkI8cmC5ZtnKcXL+TlnfInybiTg49lqJoke2b47E4CHXD8gxmX80R8
MarufOKcOLrQGbAJbhuGPCtJh7vqS8SyrJCqddLBLv6mwm/awlmQoHAwOtDmhT/H/FLhbtDbbKBS
u7zwR031+AtAsBCrJX0hPRoy1xRpIawbr9janmReequ5Kdck0BmSEVM8w3SjbplyLHhwglUYUwAL
+TzEIQh7aSTiPENEDFK+/5Z8U3o/Q6Zt7x4jB83FhX9R18EFPEMi6kpAUlUodK+DlDYFW03viyVo
nWjsi93Qrj0Ow0WJGGDLU9myXGJChGJ3AkOSYbp1Wgw3UMzDT8jqe+99QDsE0MIp4PqRcl90vVjF
n87oODnbsdX1dxzV72qtmQn5+mG9/Ti7OLD031x6NROV+UUmxdviDFQ8sO9xbnV1P2J9aoGIDvT5
a5dtO8wjp4Fpf5MSY80y6NCVypsD3/TVxbuUAQoRsc+KN7D9dgpPdsvwBKYfbghBDoR1lnUlciPS
mDpkb32B/nFpW9oRyJEh5XstRWcmlbXRCaOH4vyu6gJbAYB+h4J1SRs/B5PHPPgMCIImz/PI39OX
o9RYrUFzm1ueKIfajypCxrgJ53W6Du4PDdxsr+nreg+T9xP2icXvFGY9+oFVWxYsekwcd7O0h8N6
2MX/UFynFQsygjlN+7qx0mJfI0IxPk7lGqTEL0bT3a5+hxOrtO7vHMrwoKonkKLW9fKPlWposWB3
TUxTD/5q5z7jT8RJeRz6lT+h+Q+AsvzSyaD2zyxD5QC3bMiFofAa1Ccj6P6fcLc5U0mQOZvkRRQG
XS7a2HfunTBfr5RrjR+2HNw6n4xSSNpPwpvlh1sYLxW493EgT8BMQNnhcNoEpHRTzyc00qrEs5zd
UtuCuut6smV6ncXRybV72aXAIaQGK5fQk5fGnI60mZun0sgqxrLr7xtzg4lZcfWZPeNELBKbqmwk
ehQkiXGpnxtnmxAx2SByfHLqlu5Mj0WMfceTM0kYP81D43UJD+dOumcORVhuMgx7HMqlK1N0z41I
bp3b7xjFBztZ9I9Q975DIUrVhtLnL6ux0AEjCDEG9M07975klOIz+1+ZWSEInXPFek0GcbJe+kyH
hhHMGSuum0kN2IOhrdMvvA4AX/gxm/XC55DALve3xvwcZDFE8PDchm7d7jGROa0fCanvR0MuvGEm
xj+jnWyWi1pc/a2lUcOpULv9iPIgtk0osbjFV4ZvcN+BdEo3jstisS3pBNzMT3Kh4ShxY6ZioRVq
aLuOwiy4kcLlvIXXhkDYUbxka9EzOztCkiT0lgogpcX0ScytcXgt6rTbRo0kwluInBzapUhu9Aew
1GNce1VZNZwwXs9t/ulMmo9frOKNekWvTk2760APhZmMPJMOSInnO0gs39zyLLtNdMTDSB6mtMHP
hHp6PmtuiybweK0cgMX4/lgCZK4xAw8C4eyiQOIuKeBe7Ozy6m7X868JlLlYvK6K4aCQiypB4t8q
BYCxEoSpTKDoA5L53bhtDFDNgzNu92CfofaHkouHYuu8Z69V9RH/15qex6E3M7uNg/2ST0iFWQcd
i6OsWLtHG7D+azXpW8PEhRnVhLg0GvI36cv985Zc1otSJwj+JftS4f/Gh05o6EjvS76ddC9f4eST
5r3B34vJoXtQc4IajViHG2ypNWALvXPDcgF0T7ZvSg50IhMxR8RsYRgiWjJ3mebfCjf1QUbimqln
CcPIRBRIJVvS4TzeU/ZfNXcEeWGSxK2dKf+gBOHaLKp6pYwyD/v7AVY/zr7EEz/liTvIuy2pR0Jg
CpKZUdRf28HLgq5rKEaEr5NeUKJ6Ka7eVs9GsNNawYrfteEwQBUjuAsybXSkU6vsYN9yEyFFSqtL
DcoNhrkPAAGDN2zc/eme3z3hovUxk6NMIHoLKWZJyvL0mkj20NMEOsGd3SMqJpaHxIjU5+97rCvH
heUUheV6ybfGzYr2Ww1ebkGTrXYtQ4RAULluS1yHq5F9v0AMh3iNGwgsdnQ+hdpR+KZXTwzAEpXO
2Lk2JYRNGVElvXXYeTZ8QwFdR23NaaP1/aUreM3INjxA8oPB+JtNW1EecI4i6ax5g+UZBbv/uah4
rnd0lYs8r+lNC5dozv1mYIM9zxQ2fhWJjp1Rnf2ughpBWbdw4K5+7DLHhspEh09ode+C8tz5B3eD
Mn+islvNS/kseWkfch4ICAqhF9lqR7XquIAtsNohpxSgeNNb3/MLqJD9/PWbcjApErqi+XgGmMRS
hzlz67L4UKVZ0RSam1ztY80U/XUg95BG5dJRZ3XrncdagDPFN9oF75+upk5ClrLVZo96BfTrsmaR
6bgTYULbQkkThwAcxZcFk5IrMuT7EqrmyMZ9H8F2ecLJQbM+1hF9X/e9d97yli3CNqIaK+6LKXnj
DfNy5lsmQV733Sf3igqj17HybM1fnM/zOiKmuiHyueA6act+N4cGeoi41SRABx/HZxcrHzw6Qc94
ekmJxlb/t1fUaNztY5G1+++y63+OFqjUit1cKJHB3jIRw+0fxWDMwgo1Ubm25+a0iXXMu5hXWYHu
zcXVIJEG8Uvu0+TKPjM2JSikSNI/wNWh/BoJo3Fz+HqMmewWO/LXmq7lp8mwxIQIH+fqijCrNeKi
VcwFVV+3wyFqG0b1CDRY3WKMRTt2e7Nd1ZHyu8LmoyfSXBHuPx3nTnO6mMMSj+vtHV9F5zEtUvaI
/RCB9ZBK2bGAkJKE0dnTw1qlW3tR6KpoJtA5fCktoAcabgrUGGq2oDVQgY0Gd/QapwaiTuSxThOs
o7E4Tzqv//E8JKjRAmaEOPPSb4dt2H278CbQcgxKVe0Fb9qvGlCYR2MzQpyHo4eNotw6f5649xkO
5BGtYZuIcxehTNGUdFVQ7eXDMYUPQG/GgoQ5/ZiozqpUyIi823Hzxa4GDfQVeZiCa+P9VoyGotYz
NYtw8J5CG8FfIXwe1OvDYFOuABtE0z0lbcvAxaHWTF02iMnZoSzZlei0l34ebYXcIGIyeX+Cise4
RIiHwgs47jnkpl88w1kwKHeqyQ/Nk5NsCl/OWaIq7bnRFfkSnzQwiCZM1tmP/AQbbMjtB/7W1kVQ
hxwEAztb2XXMOuqOzd/KkTbTI50/c1UYOhXT4xLuP0LZQyKpZyLrFxlifnT9GbFOaq6QO3+580fM
6wdHoX78fDlyRVQFfkfGaLloeRe7crxeyHB3OjYe8LHrryOM3Cm72d5k+DQX4Tp2ytjAMjbdPK0I
huuqQ2d4iATDNWE/8rPiAQ5/8wz8feDFXaET6BkEITAO+NWdHegPu/ZCuwy9Qpe/1Tp+M16RMIeM
K3WqokooXhiIcel8iaNwibXzdN4osmnwL+3UC5rgob9DDy9mYfiDgKMjSGTNE4BtgeOXAKJAJSpX
p4VyFk8B10vvnh0VOPLeN6SzfNgumQeEsmzw7hA9y3efCutUIO8LcJJzK8GV8hc12LxNpVZnDJ5k
A6z78cs60VoGWoT6kw1bVwz/eirSnGHIhaIpmwQwk3Mw5WRj1kEJaa6oY9Cxx82Lh5IYRi/G4DZJ
pPWjeA9rNcqwknnQRoDcSVSXx5040hh/dVVPpw0Y34VZcl+h7+DZHofOpQCpRgHJOl1wlHjXOHHY
DXC3jamiqTYP8DF/q3KEld9+Xx5kJ37ctBf0oPhCznP+Y2ZMkKDaRwXn9UdBc5JZRbog9WmUDBTF
efXyo4CmQ3YW6wE8K47PdFX/T7n2+Zj0+W7IgNY8its42yGyjfDPtwM6t5VmMI/4rnZfcGWIhZTT
BSbNa9y7Pch9fjSgB9pou1M6pk9XN2C2vkDCGyv6VSzle5lYlxfw0m0iA6h7VRb8gNC4Ra39nggf
HyripurV3wHQMRbHr8ZB2fjYPouKvUroIobD8fxwR0VZmdj6vwOlNgha1uGDwv9ky7Dr2OodsgcY
mmY9IFbGoeRwnklppuP6mh2E5H+r8mza5PRWDl0U6L2JNQfb9Ael13vmGu3ePr8LYQmkyGGZQIRZ
LgYkJAHt9cG9iDzr909VF/BkAboukEVWJbpP20TItdN0nFre79AxojxzL1e9nKQ7NlMPnUzaS1Un
bZALdPBbp3JS9BjCm2TPl5XqQSF9Y1jF/AUZojS/O1asaw8Z5DJ67oZ/k6T0ko3hKsgrnSneOVLm
xD9niWL2foToqHnIpAUaX7SO+fnkxTpEVobOhagb3fMaxg/IlVKJtNT3RkK2/aCVjEJTxDovABEp
GLcCccJa94i8Mp2GqP41SWofQq8KZObXJW/mKjVPb+Z9IX7xHsey+324n94JyCK2FcYcg9pysiuG
K881EnCLKpbAo5Nl9uRFQb6i/Pi9J/TwTcpGYa3ZD/pf05HRklbi0dwePtSpwolajH874uOrqNJV
GsH/LJX3tp3KN37rg9bjNLAUkQe66FipVD7bLCnDcwSk+Xkv5EF/LJQ4oBR9MKq8svjCW6QEUoWz
ytIwrSH8DonZelS3uXwHweX4nCua78KiEuKD+c68YhzAGEtaiEXjOFUhpU9JAvQ8jtL+kqd71LSk
seztDDnmrlNDFicrJWGJ8isMsVVfaoxiWu14olBE7N3ZtmrkmNL+2ltpLqBEgBJba3TFLbK0F6w7
v22O+mx2AnMgUNmxC+/nSlGioKeX21cVZTuU1T6bBBXOuMQ5HF3UeURRUIxv6TtuKE+FRlNNkeRD
Zog2J2e9NdIolcG/UzsH5NZ9UNKeCYguLlu3CLsTqpM5aGTVvD8FDwewJc/63PBTlZltvPxx2Cll
Yb8ax7jxZUKL1Ivj9/R/QEffJgLGACnuiSbA+vXuKFbNgtGc3rECDEdsPlYCzwcX9Xr5jEcVXnhQ
WzpcOiD8Fgm39rjG2B0u+C1UvbescbYN665YN07qZZih/69f563TqHepxfM5JbFWB+ojhCMTYive
roDDrX7pNZuDRT8PylCsLFNpgb8Mr32zgzLg72W6ZUf8r/Ba9ywEuG13Rdx23z2zJ3ANmUd8xGxc
vh5AmXP//qASS5Z0NndfeHhMEjlpnv9dQmIFKMllLjT0/VA5dd5v+Egf4j2T9TdGRj2rnPMf3R2M
b+J2REycXEu3dxbb7T6l6gKEGRInh5XgQxhTFvZwsFjDZhMb0ERqsxxqZDlwkm75WjnZJXYoV7Jv
DXYniIkfPSiWCLshmToUTYqraXR+HTuVBRruT34+0wWAKZLFzKA4oWO5eXjfgwc0zig782xLslyw
iDR597ICbP4ryWAGbmiB2GQ9WQkuLZD0EJc707/zahfVrXPGP0quky9BYbbPQ4o047UyWfG+WVMz
VCUCdgmhbWN7LSrTE7hEo+EsGIq1scmKbgWjQ92u1jg8zaDV4VnrYe0akUCr8//aC03gyB9STStL
LvrXBapXBf94kyUBAB5IAtIJhm749FRASQmUvN94iFiDhx+S0zOuHZ3StddarKFK9YAr/LGu89PO
eHfO2XS+tzjW26eeU+bM/w9hZc/ta8/VF9jAiBv0a+CHfNPMPDUPWWvljX3Xsm/I40ze9j/mfyVl
Scy/SxzUOZIP/u8Y7r8h71O3HRxBNR7jJvu9RotPQXhkTAoCwvMzBN/eNSxxyUc8lCkvXNq3fOoo
m+J7yOCI9q/Ty72yaaU6tZA6zcbPWjdxgNtSA7W1u84T032/tuda+4QyZOmQnhbhFHxQOd+DUEBB
O9t4x1IsWVZ5P+YQpAiDC5nBcJrvgvoRwh5LhyF3nnT7br575QxoI9azIlmGq1nhMCyulBsyLRIT
+QK+6/Li5skFGRmoSrYSDnI2OzNtobFNjG90xZnRjzc6fAegnX1lUIVZ73uWZ/sxG35vx5WHJZpB
jDfH70arMEn1Ccm8KRk6OVa4LiotKA4Pu+7afPgKS6VDnxSEvxZRG3WBLxwGY6lsf1XAG6bh2PM6
m/1xYjdu0CV0Fxw1mnj12HSvc6OgyIBk3GC1M0SUaKh1P/SeeufgRXQg1CzrYYy+Jhcx7bTrvFC1
QUJVYkEfxJueDgVXIxgo4vzptXkovnWUoInf7id3JJSBG8d81nDmg0qb2LL1Ppmtf+dAgfOpaOSR
e8u7biaYaNGuI4i9RNTaYfJOBA40WwV1QmFy3MhKZ0fKoQPcDl3WaVhWmhE3Wzs5CXFhchciAEJE
SsxeVQ/QAqHlw87q9yZDLpwCdsXVrspkgCvKqP+NxKPqctSA0d46taFBRbhNEP7xhy4KQrCQ4Ae6
reLrrbQvn85QDXBVJmLRdKDJticqZJVDjkla3RLds+1x7HyNvmHAUc1fW9nkB1tUE+BYtnV9RQok
NTWMCwVA+1a2D0PcR39E0H1BGTDp6kWrIL2ewhbB9jT+EuJ+Tz9JoD3TRyQMSFqtyZuRgm9ACv7o
yLFW+gqo8n0ffB9xvqBOSjLs4xZXUjGuhbMGjNvNiVfhcaQtEz++jCaNQSH0v6dAJ3UFJcm6iyMi
t9g2dpH80OB9DkrADkvCMf4CPdWcMiDGxvxcI8JbxFoAgsRmo7/UDwgWdqflQN988JzalOwhCb20
iv7HCf6fZF4qcndkc5NOwDFCCJx8XszYZ5disb7tBUTxXGAeA5zt38x+bODED37LcrPvlO+JalXK
H+1cCD+ZPR5XBcLbtrKheAEORAix7fKklSfFGxo8k5jmX/7X+NqxCo14wO6HwJswE5jCqlQwsqz0
p0HXb8O2bi7Yv0VHwMcx6K8RlYhjVnZB5MmIexnNLq5puO/VWHhVWbGm+FNYV2MTY0zcI6P5fgVK
V8GaIo6WZBhbm4arPJNqHDzhp8JcO2kpywyqH5Ss2XXLKHHjhuhcsXuAxtY7smeK2uXYrdXuao0S
fhDDnFjOvTMiQ1AAmThjcuB8K5stWhOnxvqsRVZBjyPLH9bGZ9R2C2RKIhjYrNgQD6PO6P0qwW4k
qqR/9JBxm1PwEVkdoWqF4phqsV5Oar3jjcJ9xHVSIS2XYlTu8l8BXjGbr7GrEdXB8/7avb7SWetV
WNI3CxTZUeXsvzAT0umg4sPPBMwT2Up+Yb7DRGmC4X63aOvQCraXbO0XWKyCAtto/CwBJpoptjh8
Jyzql0EkbsnHS/eeHi3ffZTdwm4SHKjaTW9sEtHcuLQHNjzAXV7OIg5/DJmegzgZSZHBOIxRcERq
hu55IowNnjmvGPoUUPIn6g4PHTGQx0FaRAiyQVETveMrOK7erCkcXZBvyaHTXl3K9reGb8gyp837
88AfWJSYvCE6mtfY+TlhXPAiX6GZwTCvojnDo2797iDiLadntlpccA3XIG7G5eZrpCiX/NeG+7oe
idw+MhfR8wqugw0QXmJfUz3IQM6rEKIxj+RUrsbKuRmUBfLWdsiUUjWCtQAJTagBh1AjBsTI98l+
3tXE0tbR8hBsoIdzFq+BCLSdZnmSkDE2OqzXIOzz20iXAQ2wXKtPVNyMiSzcZIuQEZ0LtMo1rnmH
nlzYMaoj8nEQrQakYK60GyEImTWuVoylQGO5ogKy9HWux7T7TzXDjsg+PIUuAFV/uYPtE2YxhD+y
rV4PpKzxU5s1hml6/2knKZm9YnavJB+OEcJysDoQyoAx750z792P3RePPnzXMpA4Q+N61b0NW37S
xnqk+ITGl95Q8jyrSDo4yItlC+SyaPU2o5ZvPxbmLXQ7oMdcPWHFXdUcv/reFNJygCdaZsXWsPoJ
Y+Vsm1vTOMO8JAqukcLjqgyo+dHTjjDdXJMwGHgVf5FwTm48THfRtI/1zqPkZmuJH/66ig58t2md
/QEzNG5sEDAaFsIs5Vz8umbUw2Loj7iC34fnq0geROOyqCFIUsyN+2hE6JIxUi6D8LAmHRUtkZj7
zxPxXvRT009TaLWHy60lzXh64s9n2zmvVP5HZ89AcqTpsPZ0YB2iB+LJMGBSocT6U1FypGnTUWQt
j+oE3AiuUPR5+wZslWP3fPgg7pxkUAHWyWiUvXByueytTNQdA+zi1l07D1fE4PMdjSmbm+SWJOFN
wnRSKOES4nKgiv+8xZmr0ma3X1fKgPpiXHy18mru9drT1KaxyjxZYBuIlj1YS960lew8HFY0FhtJ
enDSTh2kEU+FSmXzyuJH6t4Wpr9Q2/BAbjhWaGsIfDplcUmWfswOkIQYXp2rd/M+lFBlZjVwGvEj
ijUWUJKXLuef3nVsyRk+Zp5wiI1mtaoa25QNr9mmTVZs0fjBCsgQdemnx7RAbwB1x0ND4qvh5hUj
BcrinufQCdmB26Rllx3jqCZiA2MfthvwllaZuWzeaGfaYdYJoOiZPrZIVO4s/iRZDWUHYHz71SaK
LFljGh7OHgzxHJmWoU6OmJ8XPNwSa4hPgs3FNb1HBP1VSq2jHiRYsbxh5UHkk3uUb1ShK5NXq0F8
y+b5dwefHzSL+wMyEoT/TfareMckvN9RauvYdyif1svBQyEYenVDrpJ3FANx//B+3xE8XL8L0dL1
xy1FNVJgM/tq/fEqZvdCGL5VuNAosTSL8sPLxdAoPGV3ULnDmrgKNLi3TDUhj12yunga8f/odtts
3s0tWJ3tSCaNAXPXeIoRlhV/mqD8u21tTZuSGbi05Sth3nfJ7kqNfuq24pMBfWvevQmDc/MJVJp8
Oqp1zfyNVNUM5s+fGXXbO9XqnWrSc0SbiDnepBUcwYiDbjA1PNcrzilXfXgjq1D2KdjEOUnflV6J
kesj2oMnahRxQfdCRzMjotAhWN5JQSswv3yz6lHqMSVepBb0UpadF1dcX1ijOhez6q5hj4jZVE+6
RjAsw6Pu/JuI5mS6GXM6neNBlS4ipcgz+w2fH6O/GD9GZ34UUT6SDC8+LKGyXbKDA4DrIo0Zk5mn
nxAyxWFrZBKlGIH+DJzeQqvWEPOc2MRBU7aYgH3Ne6MAfD4896iu03HrWLrha/IptsGzkN4rPHb9
vEiBiw+04bqp6gdrwX0MCvD23Ph/MHypNhgIwLdodugyykKFE1kPV1zyeyRYDi8QmckjQTdAncVF
25ZnG8uRljPqr96Q9De6Ab0fAwJJRhkUQ3MvgoEDWU5FLW16FjR3erHYYCySZ7Xs4CfkqmmTbvC1
FhpLYIp5n/4DdhijjW7D4D6ePLsxLoWCYtw88VrMzBZ8jNKpQgE5Xspq6HnCS8bd49EOUlJynDaV
HIeV4H1OFs2frNEYKDP2tUy+0n07fvV9iRv2HrjGmFOnN7S2dDevlCARE5sjIL6d2ErpMYPEF4o4
BCFea1deLal34Vv/baaNuI6okMXF4hnmzqQ76wEzn0lgBrHxf4Li+UEXZl7C80aHuHhPozjeSBe6
U87EoEnFOnYsFeLtKogAnAziAHXTOGn5AUUrOhtDWR1h9nERllQVLU45B7A3282Ow4Z9rlT3be6s
6RcHfB/PlJ5QjJ+g18pERxr/vvj/J29eW8CE+i4YSZeQO/PEwx2iZpAHuAFW3MuwRaRAwIpo0MVG
XFErZS4Ja9QIFGDRLdvUfZnX2ZUfcInw/O6uU9LAEvF3Ru4wgNo9UtoA6ha2A1ZkHHvhPgbIVAfP
3ofXeFCVVafBq+RaFdDpm1zQOm7cE0s34YPeKOO3i5Ys+0qk/A7DZIMRwcqBgjYfkIPBFQfcan6X
Kt6usK60Gv7V4wQ+j2Ff91fLIhPmXmpAjDzgnNsmyv5gTI9QafWb/0Rg9RaAVi+o3BjnOhRvb7c/
rMf6iZi3hAcncV0Zl749lt5yyuLf9Ft256+WqY+0K/k4qvOsSQ4cPpqFPSsKM27BiqnNeoFL1XVd
HAEE94LSm7JQK4u6+hvi2Zv3sRlyCi/1VSMIv5UqTmVse60WxJh0fU2A3AAjEkNQ1MoUGAoMTE5c
PlBoz2Bej+1K8E1YVIBTZyna/aEox7Owd9BrW9cvLSSS3MSceU4+5TNI6rtMcYlDz9EQBe8a6YIt
2rSYiIgWAkTezH7P5adj+bvuDTs7g3CIxTULnhBy817e3AHlrsB2w9j7ph5pOk8E7ciJkT6Wp4Ov
C0DE9w13fFLpb8EqiDKvx2U6EicXTNA5KSzpgFi2cuOeinxz+Zbn9XRyRKLWSlNdzfkHGSzme9h6
dYGaXCMoVBWtCHPyTACW4fHwaIgtmFddRuo8zuEW50xrdN7KhRoMi74gbjCgl8YuDseb05llqMgh
v44jyqyVObk/R9aS+elQky9ItUiq3oBFZ5OIkq/Uh5fWXuz8bC22VfieSML2rUEATu8qwgxqeBnw
Pq8DqZwcOYsy+jzx/a4zSWq4SaJSRCxyqtq0RKbx3LxTDYWgwoIgpZge0kWIW2cGuVZHNgJ9bpHn
cOs8/ZwtsaU6f4uN4HG7cr6eIQC7ga1dzVvAf7JWVM/c5dCEOncnybbOk7C4Mg3+5iKAM3vf52KS
WiMwyYsNXnsgMkh3f2va/1rdJf9UCJNE3BbwLQ4lp3Z7wiDsMUm6zCFzH//BEKq90mZjzYJtPOX1
BhCqz1AyqzU12jpBgB8eNAGXrmnAtMJbHb4Xd9VwQqYlVtfbqLU8cfCt7CiSr/IIh+kTBnl1to/b
wLzPloJR7MbRyXjyIL6kgCC4Y9LUVBr6p4q6TxxY1pOBjP0gYXvddtoWMIwvXeneatyJc1ojAPGr
9AtZfZKq+F8PtszszzMqEtzSbMWUJ+Blzu7lcsiasIsz/UoDFT717NONy0t1ZAagJbq6TJetHRAo
hVjlywomL/8Ij7QQeJiFwy/kZpH+ARGpMdSA7M99rc8mUwE/cg7ySzBMC8aYqJreGdGhRAboMLpy
+gKZAaG8+NXUt8jBRvcRq2FmKixH1nGe9hp4QD6wYL4uFemC7gG18RWR+ZJPUZPemNN64Ru1tj59
WhC4N9ocPVsR06yc5p6ol32573D0MYHRHVTYOCzvdUOvInuH0YxLQJyYQMWG+lLO1d/TVL2YTSNc
Hx/HL0ocgkAqs/+b2KpCuh1znrja8fVycD63omWErV7M6iPn77Lc8v2X/oyHsNkhvdlTd/iFzJdb
wJWc0gmidxQ8dvgxB0Pl9z1kP72B/lJOuWDP5ijpqH17dCE4iYxAJDqmQBnHanomP9pKOWT/738k
gX6FR63YqLSMvTuBlRwbcuXJQBPE4Ta93inxTPmzc+Zf3r7bBCMGwHlxqL/fNgQCDcoCpH2ls6WF
ifB32CH1OENEZnEtHBUGmFGcaQOKxADWFZYo4zmXIneVtl0scN45EA59aJnroJnr+MDgxJwh+3vr
VDWbwy9fJQXQd9+FWY66FcgDseBAOFBewiKaQVd5/Zuu8WIBpyDPKJiy3XZCKs9VSl7sOUtPwhms
D9clSTe88QcXB+la5/8fN+1+soZ6D5oUMaQTOyCIEI3FzwI7HN1rOPC30TYyWWm1aDwlAhjn3Ds0
elfEA87IuVoBx2EU7iP+SOkz1dsieY2oOj0xrH+yJDEkqj6xU6gmOqPsZR1upO9J+Xm5puOqJmar
HjRR4qWpO488UumldY2iPbsfaODBS0xRn1tVVdw2k535DWo3PMjm+6tytE4glVVYbThYXuqqC4+P
sFuNAWDOfJ7NYn/jkmleCNY5K6LyBu7OeH/Du34PYHRKVyu9qtLMnLCnzhRQrFM3WRrVa7iyYLKL
iwjfvkG7o8MuNyJRg3OYr8sTU/FuyAli6B2ds+39uyd2yNpPGQBmOApkfcHxo9T5hkciGGROxJCf
WjALuDVyYP9KQfUVSwATBLg97+Dke2yRmq24ySdAQDnDQ3Le4E5JfqYKnaLNTphEWoOuNtwtbHYM
YPbVyQMQ7ozCJv4BJp7rMvMTDNOIQlNuzC4o2MXNwNm4A1BSRdQYwhNmY/hsBeL+KFTpnmmURC7v
YLZK7Uri0+u47ybOQXoSvcU3FEl8kfA/7VSUY76BcUvTulm8MtuFDd4xfHlePFv3seFBlh1bginv
gc6FiAnczRseLIdrk8Pn4hiVD0hKt5UC87aUUs8+RwsMPR8ZwcHO1emCYFVbFZxrLOA9JdVI0F/0
Kh8UPy4U+o6USTJwCCAp72rYN9btnL6MIUpL5hP7NwtiOMjDNcQkevpwpiWLb7DnzdsaSKpuyOOF
mGEhyOlGsLAxAMdAIAsXhOyyt7R4xQnh20vF7aWayjm+7Ckuzo6+M09rhS/oOnG5l42RDrMPcsMm
AYH+GMU6QzBfKu6vCcA1l8Ua29wdbj6seQczWQxv93leKXkCq+dELY0iMeEemQOZCt0ypVvcxsoi
XHpQ+rBatgT5AHxRnT5spi4O+pN7pWiXDUfZdMzbiYZkcYtVSrpAiUjRWWh2nzepo88I3MEpqcWy
zic4XhEKn5Rv70/rZODj7gbL0xZx0S1Ck1sDj9Qpq4DGggtvK1gNZxR7ZNZqbisqy8AFjr6AIUpb
glc4HdLoqgtV/O9+EfHYG6HNGPWFGWdKsLr7xw6Vmnv1ChCQ/79I3XVMSut8fpRlSO/y6EvvWY1U
8y5UoJThEyy/d2NPwpZbDR0w/4u7dVzbQi7YVfYtlXklZ85tnCqqFDM9JMbr4oWYYQzBJO14WMRV
oG/vBoRLvjwOgqUwIzgW1kN1x96EPsaXPlWZYg2JZj0T4FAtbs93WlTvP0Qkipgw4WwBDeN3m2p5
n9/LK4NL2GJ1JAb8ZVahQaT9uXI45YRKbjOSLIF650gkv3aUWusjYrh6CDbtCZVmTWIjwWg5BkgW
P/0vx8jn1r+3XsuxPlJZ+rN5KBTG9/J1iUU32CXEuagFgUIQEUVt3+y5ctA0koHqk2haWJDgZ9tt
D3+bPbQ0FjJyKGpZkw1ZBWQHApXKmvcWcsSWVSx/JfaVIk3Mlmp7CwS03xJ/lEZHTSpT0MNRy+BE
euayo5wBcphHdZlR0CEmRev4vune1QRf1gxfS8DxCPExvjxcPeItMuXlDIQ7MkJ0XXFcdIhXnZ0o
5rIW50JMYaOkfO5QlKxRXFcuM/atNyfMdRZ0idwiysiviy1yjX6XP9QYlsr/NrbqGY6aqrY2+QYQ
awArrRCkFBMWa24Scd6/Bv4XMDrpbqcxgWIBYLSRKaCwCIJsV6rTsi9g2jnl1Icsj5+7SyCJsDTX
fyN/IpV0EMLmP/SUO1JV+4lioeYWjSByjoPsvLHlzMFqplUDu7d4QkPgHxaVCEpU0EEUvbXX34yj
rLV4z+za7ni48WNqlPoezDM382HLmT237T1LTC7/xQdoul5EwJVJ5dAkLSx3PJjYRpND4VqnxWeJ
QSsEX0zyyh4UyoyqjrTwYK+385cfNcVqs2g4+IuQiRtIKg1aLesmYIhqd3SY4LwgxpTG7wG6ARq6
uWCkvB+cIMArouxGf+JbeoKUuzjXRXT3SbUz57Dozn3fIW9kQ1ZnU4QwI2k8NwkmUiXR4AGCpOJz
3wacxP1n+D0kvDsrS/LaTgPhBCY/NTJgtuo3TF97SzYrikURfAlry23gfW3cVOOe12Q6tkbUv8v2
w/o4fLv666UszkThgB/ByWNAi2ip1Q/PKipI5o/PwWfyLz9mWFYhJw3/ibc3KHiS5C+aqy3cmZXA
t8F9nfzthRdm54szKdGZOLGQfSYt+qD+SviFfJEfv9D2oEyHAmD6hqFMQX2ZosYIQ18iTssLLmY8
ydln5hePq1FbVMyp+oKCQ/QyPTjYMKsm7izyjvPCcHFsYNlAieo3VEbUsBW/P/NTQrpdFv+YwS0N
Dafdh7Z0GY8+020SlaT/FNIFagLxlySwZ4EYsY81+F3Y3PVIKFjuV2kOu7rbKzbfGeC1grDeg9hd
0XPnDcMaCjsHWDCHeRs5e202b8Y/BH+lRpPQyKZ4Vt/YeN+hu8pazu6LWd4sUXt+XNm7LaFjt0hW
0Q8yXK03nrFa24sXxjkgOeC2qZiXMtM/LfB28pbkgZXMUWqaaNtH4cXFaDBeKfJueDv1KMNxU83g
H2UEaI1Y56AnfFCmu+VRAmd/y4N7Lp9RxgkiYBAgooysi76Kb4cY/DFvVcLvNhFjDIeLo6NwBSBE
EG8YfdCDBqRIFhzMAl1la+/UDmeKDUGo77DM1/5xEA+d0WHewpsEN3m5RNsrk0e5fLUsRBkEfbKN
JG3PGFb9UChDN4Xdqa3/LVNDTCoJnkjeu71w36QgpHYRL+1UgF9lvfj4P2QqXIEejJt6G2d6orsh
2B0BShxCFw0TWcVpjml9Y0lRH2fIboMgGbXjyB2ID6U7TdVvbQXnswfxDtYqFyNdBuuYY11sTRPY
bvVHMA9DdzM+AuffphHrbrotqtWEtD2713bkBoWVoOfnFefvAvEqItxgEHWPk7ruBDxANLhT2IeN
+icrg75U/ilMC8tQwL8tAYLRRCkJN8QLurAHuCaYQX+ouJpN/XEG8pCrYThk0QeMCUs0qlyQ1xAu
NDuzDGJx5js76tmFXskYmis6n9QxUe/kiu2qKMAQ4QsH7LXlz3kKXijbXrVZDSIa4vsy/XmmB8cZ
6ntBblqz7eC8X9gL1077ok/FnSK2D7E/rI8bI8EBX57LWaeNyvb8yh4TRlTuxvXBu7AujFAId9Ig
QkjixxJvG86mMNMN352+K5msg3Vy70+v9Mi+0aAO4eCiqnMn2xDwJBUfXtEPyxWuadk8IoWYVKf5
+iNN53Q+AF0yHCbf6gplDoUk0RoEWEgDS6cVowA2LwkBGj4ea/UfzRxXpEDVAHAl2NCRB4L4R7qr
HkpBp9eL30BHf32gUGWvS+JdlDE4ISFhV/muXRMKpsSjrBGa+U70vVhpy4HHGxh/YQJ4fZAB7Wtp
+jY03sQ9pX0CDZ0qBg4gbqc28QO+mPmSdz4Z1GV6aVHnwQ6fuNXlXr4FI4XetZz0r72xbPYZ06/S
tKCv2Tk08BkFY04E+6jZw4m66QKl3up1RHxLs58KfO6eSnLyFClt99uaj1H1S5Bb5+YZiuwPmNql
sLt6CfY1yTR+0CwUOUg4UeBEbXm5OMT+CMBxpP9ttgNFyy36YMCYyeonKpTj906X/TF8b1XWLJX5
+X/kZMaOxMu7GkmaInt9E34T2XZWWIdKnQw5DWH8e2u+iD8UJRngk/EAOdCNVuy8vpCTvUz1XOzW
NQln+ptD2a1YcPW0KswvfR+Rbm1KmQDG3EI9DuUVKg9FYyZMsE0RKKXekm9uUKcCLx27fWYGVUGP
0XvN/hOuYrHRR0zwQ93+ZHe6t6ThYJ3cFInARSQPgDRMDOraWlxkc0vTgS0DA8ukHp4fbh2OWMgp
mOsXl4/qlN15/2qWAmk8siZcUB1G1X51YbM+KZeArRxhY8IHuUjqylJwQp4bOgYsht4zruQWchAM
t8ZdgxJcgdNyi+EYJuMOE0Kb5gCSbmTATPlxVwckejZS5o9lUGNml3LVQPR96hHohvV8vCWPD5ie
qKPDVdpD6zjNUQV0lCfb5YdY3vpvttE42sabeJsAAhCEYjvqEBG77rwXhDLyb2kF/C1vNAu5u6xm
1YIvcZUwd6wSNd85BpQWm/VfIaepiIlCkhZzkuYiYwPTiRDyKcU0VMpSOxrcb/UzUu7vMLgIbuoN
uQHe2t7GJB/MItoZrdDpsuenAVLh4FQsqQwZdS1dTwSbjvxv1RnS4TuFZXIveUF43wnnRnFBoh1M
l//ay9/HM/uEYFv4W9AUq6SlMeS5Wu0XHPGejUvDJ48wKKAeTenfuJT5ueu16832IfFVgwA5d6Dq
Y/tfNIzZMWlL+TSYf6BQH7beQWyRH+tc7kH9OKCQdEH/uaaKa7z3NSM3uHUDlp7w0fXPvwjiWmZf
cw5CNdVWmjzSSgG+3PZ6PegbBWIhyuoQDc29VVIl46K2M/Owog6zVwKQhX7YLtjK+uDlYBDK/0yd
wqkiDS6mHuO9cwHmoQuiIAZGb7qsVaMv5AqprlfykjQSTHWp8liDl49EnHRkwaGRzMFBB8XvsT8m
Vd5PwCTA9C+B6u926woO+dG3EkPb8EpO/soDQ/80/YJnV4oHxLQ+MOlcDKmkCDnDKlDAQc4yi2xZ
GMBFikjAo0uAE1A8H38gejy3+dS0kuWGVApaP2dlXlvzEF9+LP6Cc7zvsw1WJLfc2waTgMK0S2o4
7Fl9bJwn45JV1Yco3x2b6VPdMIplF6Ht6pH3T2mT5zpmh4ZuhpfHmzw4OSh4ghQT1rfCQD9+cYB7
t8CsSNKjE0WMKZ6+p2EDQc41Jh3JrVHJ3aXClI93F2eXLNecGdYc2Rw8E5GVcmbKpG9axJvguAGO
UyYGDe/hyW3ORL7gGPuPGLVUoFn3+KtuS5Gm143/4/4WI9btXJyhthYIvqOPipjcN+QK1U8eWEKM
vmOOlXmZwG3DdNET6S8e1HARWidsSwJRj/rFSTGwW+MCOxVCG1crGAtVsiGhFo8GekcfxyM/0+zz
oWnXSlzGHBBjImXrQ8BoEOD9raMg21D4Gg9TqhrpXN9q+X8+GSuuzifbohomh7nPmBQlt/O3Yg0+
AYgC/MMLcUj017SWYOVV3XNnWrd4DEP9ZqnhinxR97vFFxWhCYVr+Nrk4mdFe37MpUhmHhtUokD0
wyoHlmTGU0k5KmyqXKUSv8WXFKR2VUPEZRadhE0YuYPmQ2p70E3j6ADAIgoPgM2Q46jKft5AgvtI
HMl1ZV7+G6/k4fTjOmWnSRHRIV+ezod/HwGVBtM423/F3QqjzDnGw0TOyJf5nWYQda2SZK5FTaAq
qwOers6oIWBGnwpSnv0Nyfy5SbcZkApd02i3vM2Vro8RObciptD9Fdr58c+P1TI+TTczpxpHmp3s
aQ3zyAXQgivEIaYlrZGN4kkq4jj1hPFBBGOojr9fdAh2d/AbYhPYN5O276z7eGjNJl9MygVIYDPs
iAOlQ/05b9XYbJCfbjru6Fu7xDOe5iytVY4Z4yUXM5WNdt7ASBkbEeODN1alANPHb7GNCDHdGufb
F/pLwB+cznoRJZDp9/Q0CHDnk0zBeBBDPMIxwsAONDoPMDWHAnUsgMKIL90YiqcbDa4fP/L9eCev
wRTbebo4J5qbzqIHEIx4kr7ta9za8KF4dLKaFHJitHP5JUva53v9j7IasM8rR11GYBF3JArXcTcH
9zu7TK5SNhnsvZV71JukdCw7D+2mf7bWtdbvnTE4LYvzPokzk7Kc4ZssGAi3053S2d1SEcTafeY8
Wpe1iZamF3ecoQ6dcoHmAuVPEVWnd8bRWhfs2OjG82lCOV3pp8Br/Xtenay1Vn6MWx96NGj4E4ao
JuGngpWUgKcOMejCSGJqPIgfeG58LgrSUEMREISWQ0XejLnor2XdGSpjTva4ErTsCIuukE4AOK1F
7bE7hkvdnoHf7hi7AGFlC/ClgbxDs4LNGJY/5nsr9M0QSdfHnxh9RZjGRu/0QFcHw69p2zLPluqQ
Mm8zmJHol8OrkZDZMmInbyPS9UnvGbKvAk0Y/d5SBfl8LgdJRUzP66knQw2vtuOT1ityD59rbv7s
FMuk+Jy7YQftXqZvuqUhtYzLRGSFjshOJ40cciQi9Ea0F5NbwdjYCCJ1XFWBRFpKpVHtxMi8nsWD
GG45vFaR7zLf6ObZ7SG3w68wh0GJWvCUC7tZAurboHSiM2bK/Zc2fAkEqX8KIgUrV6+aw/hIeJ5f
mfhm3QEQG7FPFkZTbEKDQxo9heshFdkliIwyYzmiI+vnkKNC75YVTtZkR5AE9Cwk8OBzT+ABAvnm
n1QfFONP9SK06l6jKVa/ZLYKXFOCop4TI2iGOVuvlYKS4kFE7uzRKuyfhbVbg3nZGpqpxZX7N1q2
9SPh44bq6QJTFXoyLtZ/O58d2VdwSMs0E47S1akfmOVS+VlKvSYMWbFtxCBw3rkkL/sXTZDQAaFL
GfcJPcw65vxSeuj3+ZgwiKq10aZy+xxWTACaI76ftnYiP5vWHiBH9zn8sliFZEwHfqfv+8UP7ELr
6GRXIh1HaL9QOC3EI62HWdWGV7GtUmmcy/FnzQQ7nNSwF90y9mhB1OU634pNzqLVkPOnayoVJ/jS
B5w9IXVZspiL9jrKQNllK1lqr6GcYL0IgjrjAB40jQ3gFsf0G8JaFGlIwvH37JJyeIwTA5yOd2ip
KV2kc2aIFSFyv/S5UfRbjGUyyH4cN+9jDxBkFEstSswiTv5sef8t0jMWyFqE5jHRrzRjy5ttN9en
cxT6xF4W5YqZv0J0AKvz6WXyM6Tho3wXY3RATenDYrHBw3d9sSKnfSPuwzy9JNNyvwyjC2ZhRCM0
pV9HJZTlkPHliyUWKedcqGU1KLAEreoblsVgCATnVvbpdsJ+AQ49zuukWe7frfwh0xOqDNPv+H0A
+3lHQ8DD3zWUywZWKtI53HkWsSwqzr/jMI9UPKwYZ10s0+1Nz8q2/mZHudsDBrjpdSznLCvUbX+K
joBiQRs7amHtXoUTfgFPedi0uIZIrOxqDluDoT8qYhEuKljGn/eZh1lANUzRIKzNaIICpd86JRGG
MMVd6qg7+TpZI+BYlGjv8+5Nr+1m+/0Yo5g7UPn19bh84twrLS7kTRn1vXJeZOiNYk8zI4ayXvEQ
kY/5n/nghfV4Z0d3KqsCM/aiCzbLp+i8sEABnnLSBSfPX0xC6KFURH8SiP11Rn6nm3I2GTMZKtlu
3Q8wRWiP5uRnIgdQG6jYrloWtHqUy3PDpBdBktML1gdhMBBPPkzkTaxZ+9Tw23J7ONAm8Y/Qnl/r
3D9DSna4dsO5d3pVVOUNfYyJp5BqLosYPpy1q0dmoCB0vyV2JmvDyGUbi9ey+Q3I06aJe0knUpUJ
1u7qymVib9g/rh4CdDq6eUZxTpiThs17R6QNS/v7Xa+F0ML3not1zQ0EDZAPaaq7i32ZvGLkoT6Q
HCI0vfoeB+z8+YzZL+/QuYEoC9tH5kWiCy2cy+etdn7dTd2Ma2HDD2Sd2a6lWwkCBcAWx/YVYiKs
mYUdqNW+BlUL3n8oraXAlLIb7OZiI1moAk3cut1Yot71RmTNt0MuJGPea2+o7jmSLkLKsemQNXzG
VAv8gQTP55NxQQW0z5KuJkEX0wUh02ZUMS19N6zgCfkQ4y1R0vGN0LrobUk5c1i5Uh1dg64QbW7M
bTxtXXYRBc1BsXvBUxfOrUXuKvvYzq+G0x+olqe6KNhrHpaicxUTce1MOcO+/z/MraYiaEBxHkER
KVAn8uFnfMdj/y9xQGrxg+a9FQVcSmGl+WQIN6Ve1KWjub+J2TQjALOt+VJV1UeOgx2tt/KbA9En
Ktj27V4xfRP79mHyKWHQmHNuqlyqVqo8sDhgnNlLWAPJEbOk4jSMPi8/hV1MuHTkZHW3oP8TuTA2
QtsIZ0Wio2Z20TB7R+psCKPlZeID8uzZGvxknggqsd4+Z/tolod/yKbememHLYYAjmnXaJbxSpq2
7omhwueHl8jyYhWM9o3IIlV+dEPv+LmkUpKYY4ApDZ1i2GMmOlo7fHdhRkOhbGPdhaxFfgUNRdWc
20k59/XXjea6zFbrHSgoidgADuqkNCleXxpQs0JCw3SpH0ncC0/Bfs6kfjiBeEgdBLKvcKQ1h4p+
3ErJ8PKuvCp5/G3o8SnJeYecQXX3FPyyFQ0JZqAnvbvPfs6iwBCjjVLWkPt0chErPCOCjSGLUdpT
3XGgEVJJK+xHKP8YNNyDdwkB1eT1xLRCuXjcsvTR3C3NX726vwLaAqz/sEmXiN0l9WfldzLrrIqj
wZAOGykreYO5g/H1L4aPWoeggTQvvJkxfeX6DgIXRs9WhUCJmOo/SE3coulXCR/DjEezK3Vgaq4B
1hcXlHDmmKPw6nhrGjeKamQTxgCjDOag7UdZjTfgYgH6Z95AICFWcvY6idKCaq2BrwG/fRdP1bzt
sW/ppTs7eZ7IHZXFVcJdZbJ0WAhZwJz7Z7dk5bD0u7lAlMxJKIwZHOvqcymFjwl9Sn8W/LxnRUCr
rU2ZVGaN84ZJ050vItlNaf5TFbSddhMvbMQ0eR2ovfMaX1Qv1mPK9SSkhXibVJD1nLJz1iiWz0Rx
HiEyGt6OSeUPjrrOqKtS7i/1h5951Zqxz2QWCJhlbZAw/Q9CROQ1lisduG88TUiU8Ylf2SVYaXQZ
NFz0qMqmT4KS2QELxjp7Ie2MZQBEJakoh1ATpBLNcaZ86zkmBnW7CdRKlHT40LpWr/I41yIQhloS
qIC7pXWMRC8mAkm7U/HLlwJskDRJMZuLwpGztjMa6bWZggS1/+yeI5sPXJ/+D8I8ehdkHDIjbrV3
hyVnDzb9uqsBqS5+CiI6V8Wp+2sh6rpghdSgO6swUdNm9qCET1heJjED62TSYXZcft8wCmdSlnqT
6ARS/1zWcfjWW83LcO/xy6hBqbc3eQ11KB2QAR0ILks2g5CQ5JyYE9KSPa13bM125PWzLggoeRrG
Dvnlp6d9U9zNK0NkF/ohT5vuz7iwmi35LMXbX8kjrKOHxDqEODCMcuDPGPzYLHJoyD8zFT2215lK
Md2LaZTzuoZmL8KAHY0HI9T5yGlCuUFhPcUYnL+reGU6gnIMAJuLE9GbbFuQXQZGehatYLR1VTCa
fu12vYpoLVBvFJzHpmMU0a3gZnE9UpvSXndSBG4kNeXBkv2ox5QOVQSilC8do63jR8rmkcjWAZEu
yslgDF1t/00sRjEkiiLxReb4vDTkDkQ7x1T0GhUWfDz1xMfMbDBSJrR3PbPvopKNmpv3otTNvT9G
KD9djVnpmey1M7RJhjNgqeVnJEWtBSJnXMm317wbhmTQBcxISTv7GgqDlaH6CVe2GlIrxiBmTwji
T65JNgr96HmK5S1mHqm8hmmkJehsxZBjWFmBgIL5zex9cKRxnXhUquUz9yhLCbhJ9mU87XQ5ajd9
jP4D8q/+NgbhvQGGXdHXl7wk++QF2+R3a/xWcR3svTcGbEWCQbRFA6zGOs+SKaYhhvH2wnmmlope
CqG9+h7psS4ovvn4bFF2h6skaaDQQilooUxwQNFRZ6b903seXUEAlbrgy4QRL0nRl2y44CCcsZyo
qtNstgMjUsUlr6cM5HMWkkPcm9VeQWKgkhNNemFGhZPxEmUsvxmYjBx57ii03/aRSqsy8cXqDoWv
VBHljDXY6xWMFBpTHWLfVKiHIWZ8jDiRt8KNsFNKZ5KHvt9w+2KOCu8aME56Ypp3oRARlKmwBdf1
r279oKnBHi2eugmvLUbOnJR7/vuxTqT/1B5V5+H2FKFlorhLjngnwQ9b3Yl+s2+8ZTXOjavcEQe4
AyPxx+og08we+lQlskqWEQDekjaWPNVDum02KczVD/65B1iToVZ1hNKd9ylP6w+7VTX4aBBveJkv
5P1F2LrQU/k6BqV6AmUJYlPYa0OqRX8G78fhJ9YOCiv0CIBG+qKeFQCQegodb5L4D8M7ex5aKqX/
CMNlbjS4I6NVYLhhX5NVr/DzBEFwiaUsQyBOgeNBlC3QcNRZ9xpWr+V/urry1KgihHCRHuUkS067
gjJj6KieiLnm2fd8gHqagsiUQ8olD5Hy59XN7VBK1+2FAOp1cFkia13C82+9UPYanTDKBm8hKUXo
i+yeGPOpw5Z6HCZ3jPJ+xB8KBc0Ai4+KlzWvU7XmmEMja1Eh9LlzUQ3YO7ypE8u62Kk+337Tg5sI
eRnecJMjFggi8stGAFEa2RGkfQxnufbAILbJArxmdwSUT/yxHmPXQPjjjK0ATaTQPr609mNB7s8r
abKtEv7VlT4wtR4hS0M/WLzyOwMaUz40AaRRh0+84Iph+3biGLTqRnJqaK6F9VBE3tS/MHqyO3uD
5Stp/+JjBa3q86pYXKiO6rJ9ubiT7Bv/zVCdAMBZb3jxBOr9UA8wj78oSv9P1ycBGLqheyf+J3cV
uSuBZUKXNqeejnbV0mlWazlGNTgfRvuNq5E7zxxspEZPV7Uw+khl9kckIXkvAUGCM5q2Xz9C+f69
mmpeEqmEDdk8myBIulsKYQKk373hp+GLSdd/YHM3NBdh6YNfeH7DzcSTervsjh/iMFR4S+NgDSPB
6Ed0ZO/7RWwbCp8PZxJfcMCTbBiA30gBd+F1CszVKtiMg8VCx+f5ZKuKYM8lvvmC8TN5hK0zluja
od5wWdty6gOWDRMm6JgIW9ZdkQeZbvk3SCyLze23IjJjEOiDTaR1+WMhnYCjz+sUA8TxIWjGDTTP
OHrWkbqzqN1E87ZFdBLaBIdBIqhu2x2B1zRVEvbjKlSeUcXgBmp8+Ca+x1Ms18RG2cL2OEbgM2um
2FX4Qc8FSzbupV+H5bCsTS+YNu/YxBQIs4TSXsDdGMBf6pqLb/l0QXFYS5+lWKuhJI4j7J0b3EfG
3BVIlPkC8meGHAqI8XkC4aZX30sqn5FTqo0qdQyoAFlQAuszRwMdY9UX/STja9fcN0xQquTK+tFU
pSYejichkqBQdACvpGk6Q3DzPfTp3/eFKNfnUjvwn1zqE3qD735raeeyZchPz1npp66EFTRZFpkN
/d4mJzTyu3SoLS0ptGOz40tXsblWQSJXtar2TP1fZCx9aeeoD5T/6PqMOmVQcP6vUAv6efoMmEi2
04pwdvazAWaSzvDA5MjCC5FC9IJ+8kaVgiciq1tquKDH2KTh0c/yvH2PSBBRTQg4OfpKgMYjv+ii
s7ksJTb+2g79nePnUp9Jh+qsna8UNHFpn88umbrq3+y+8T7uKaDOgt4sH1swM5u9mmS3xdL2Aipi
Y2CULS7Le5uTLKsFgVgcPlKU12AybhWZDwW5TJtuC/miAZw3lmWMwsZgnYlRP8atpBMLBkyWqU87
yIpakttqMyvaPC72+ajJIHsFZFHd5axVcTi+qpZhrxNtLflqum8/ULhRZ+StzLg/Ls4P4YBq8h6L
dkLpJ45St7mIqOm/zYp8ndwSpImBlrMr9M8cPt1SFnwP/djjaF00LUFMHGwJUP/1DrVQTAjYU2pb
D4ggn5yc0RplolnWc+7tlJ7+wT77QASCARBVz+6zUN6AJMhGJC9SZVanepx6ON8/1PZ5WJ7+Xw5F
zkG018cPlqsRz1Sx+mAIroGFsd/2hIMf0bZJ2AGcEr+06mFnKpLjHTv6xLR8nXFi7riz+H4Da/Xu
pgdNHF+w1/29Q2zzLMaOs9f3CxZ88x8OrcvuFkj+wz2e4vVmQr8HsITJbfNxJLA1v22XDqmdoRAy
NE6dah1yLTMy43R4IkrQLZI7Px2Wtv4i7Y9ryvmemgkZZsgXq5izoOk11n8OoRd2e1keoQxOIrkV
XE4q0FIQsndRSmrDP6Zu6pbhNB1njHSttmeJDex9wBXJEn9LXzEWTuA3L9L3Ofhy8NugvoQxw8Um
wAOgucpZ3yrYo9vWKCqYA/0jcimJo5t35UpkRHUtXsNMGPHfsNB0W1/hUm2RhdvOCrD8vnJPV88x
ddQrd7AzQEaasSrlFv5R3r8NQ1ysniCLhdKJGTHl0Nh3/qajbW/wZ21ejjvyf251SinjnE9fqAUz
LBaaSDCAENpFQKByeJsI+87xRNOgrMypng24C8OSMMZ6PXNmVVmP6D4lvMzJG9SgvoCntRxV4aUn
47PCg+bZPlE0c3paOCOiCH6sERpgouJer/SVxF9GYl5PAPmtAknfnEbMPa3Hjl0Z5Mn9G12iV6pF
SfurreNYneLJ2JLXlw/P0lzjv7YLi8qpZwZZjTwRZ4snNWRkIPJxqBbiSPz67TanO7soaBre48Tv
54FFU08yP3+uxa2rWzLZj12xnxx2GNKDF4Gvwc5nN8pa5ERUAYZWE3fEsMlrvw6JemJ4JgALZA4o
FH9VH2dYt6Bmj0iLtGj+w+G9sAW55jdZ4aebnl+dIrZJiYjrgzF7ckiUgfWr/6zMQDpdgJmBT4pC
L7qFDEhha+WukZeCsurSepFWnMn0ZcJyqBwLR/kpF9YaB7F7Vcd+T7mgz+pCDCr05GXLJ7JjhK1c
dRioiMx4x4ZMttL14CQQVD80DBtCqmZllb7VoykFeawNFxU9wYwKfpah73q5kRdXkZHRWmPQaVQ2
CUMbAjJBGZN3K7nhHCjxvGozI4d/UmD79buy2CZPWTSr1duLJVEDwdGXHBAFKsDdJsgFUL8gzULo
mwS9IOmk7mPxpAm3jcNPs/hHlY0sa5trny7SsrUmr/yaqN5mtge5JEurZPaev1AYWUfnt098xjrO
tvzp3tS73hx53cqeQ7cZO41kHor+CfDqvstBtfxoSOeQXjIhK3p/fcPlSyjypiibfS01y8YCJcmQ
8u9W73c970rcFJJtAHpfhgVGiRV1R7uBCdjc4eG5R0wCThPMpRlCYNFR6d+mfROLQSXbdgwy/Z31
gxYptWnr9HX2c56kXAUz2hwXCrA8RN3/mrkmwD9hgbu+aue2xSiixcTCp5IDgracd+NeNIJGWhom
jLC3E07FAc1/sVKvpv6GyWLdtsgk7mj8OzmCCGgQrP6ARm4bDlYBj2YKyUZC+BXGeSx5actHRkTQ
JF9w5K9COTc/yKQ78+py6+dD2uCa34YEm0Z40//vd0epyyepLuILntlV+NHxAOdlLWebGgAD7dCd
b0nn/w548kosIc11vY7kjhx2zCFquNQkk7iHbTpp1SJ5kuK4rz2JcqYUvnRgKA/JurgDCqIy9yfS
+9KJASBsrGdhDYii2XvUYShOavQ5yJMQ8ULcr/HIGxxgP+bHolMUlBJTo9EUV01/62NX9AvNf2YR
GTtDik41lkCM71nnnXWcupDVgwyX/64BKd4oHcMAeaI2kKXfua9MIZ7Gpq1e1BM4XMqExlmDUmbU
eOFzpiRN/byEpjJI5++X/4aeY2zsTaDIkaBD0N2yJVquop+X5rL5OCOEDfx+nP5BOC0W6MOZ/q/v
WJmeZ+JdeKCb3HpGOYH44H4/xLlzQGNCuOSJdMZtfQLjvDEpKN73FxNjbzv1jvIe+sJJtvWJbfi4
QRrFvf/4P29g7RkB4tu8X3Dq5veideIwE7wrllOcipB63o7sOy07hj1MQ2hf/YyqFk3c7u9BaqaG
zJDS+CUTVi2vG6swJNqL7xahARBuwGpU15GnMJhHFPot6yWE1S+/Kt0vtCyb7hNo+DxotVX+VzQZ
onx3n/6DJxsqaStr0Q4REN5eUtAe/R3SgyFqTlW9rN3riWfSNCPT/MVXMdPYqvgAmrRyI3IFSQDd
kdmHWpsGO+V/jUmacfBd5mOoPPWQqAc8sdV+tMZ3spCofanYKTDddwZwB3BQ64DffEis6rE6OqxC
6nV1ctmg42tJn63Spl9cEX2HmX9Y6FQYVWhzgUnz5UHmO2WPSDICqH6F/Ta9Pho89a7mDUzWBuwo
i+6qejbFtqreehMBzLxE6XftssWOdZ3tFiCEfn4l72kKf5VpTJTgr1Cq4jr1c8wB9Z0I0eIkoYFz
4w38qUDe35y/YwypXt7pqo//SadCuO+DKYuow3KzBXXH5LQ7Sf3HxRenwexL228xT6NI/Y97dUfV
kV+kTVmwrJaqWUkQ05l9nfluCVwZhb3P3D6QD3Ebn27hPfkk6w6usCg9YYC7B3EwzrJrLFIlVmFB
pNiYBwPogvQqgzSXjBxgo93pkazX8bAv55nJsrOHL/vu7yeVdpKPxLbZDM7cMNCgBRfwIjREiEtK
zs55i25xMEF+I0k1xEYX6sY5lz/sVyiHRbkmEh2cJ6nGcqXc9Cw7mSwSBeFK8+sXKuDn+xW5D1a9
5GbaWq/Q4+z2aB5Huj9oC3KqNW2J203Gdri5iFyFuSrt8oLihluv2gYOZxZP6yg4lHgNsMC6Glja
aOY6oOKhgSqtrbneq5dH5oOjwuvTnQ0N1UOqq9qjs5UePT6W+IqTa0Kd9IU2YfYgpzbY8k2z2Yu0
kn6UnNxdcvpUimxEQpSWuaogpqVqvq8nb+Wt7E85K2xEcCMvEYY3jKQROlWbdnHZIe244WMcM/bH
B6LQmvSAio2EQdKfXXDnZSKn6hB9jVQ7ZPLDPk4FZVRdD51B5jMRwAYfWUaioAwpdJjk4VpYaBLi
NszBmP0LeRV/n8pN/rmCQJ++JdgWwHFaft2JCdg+EMFyJ/nb/iPivaOHugVCl926NlPpReGfTGZF
bSZLFWnibkTZZyWAdUc7F3/XMCR6ayixOqVub8f1sMEIZ3wTTxQviXrRyc0T4nxAdpHwiRzGc9wx
yzqHUNOwO9nM9xUMpREy/xcMhHnk51Vi30OjwXu1uSXZfF7NaWywh5vpa/XQdl2b9/vMywuOwgt8
tvZsuQVVWKGbTlPOvBY8Np6ZqNP0pVpVuGeXkx1kh9ObAB3qVQJIBopqr9sLcOErQGqY4WWvy2aB
RDB32s3RVqAi4qMKbPBbPWBLmrgq3g3Wd2ZZJHHXdgx6qLOXN8O7KMKTkj/Zak1qqdgzi2i3WExi
nwaKbp/0NABBJatOvNnR1kDxZZ2WVBUa39U1JLRvyhYON9f4x2Wstl62JFKSkB+vDIC7yhuVBD4h
EoIKdEDkKFq3t69DluFxgNQ68JHzmQmIbQadIPeWfwa8WFD4+0aGZwIYJGMj513v20CS1VsPi4bj
JFfh52Pw5xcoT4Jt7QELbn4EJeIv7oPa6XN9EzSbzdcUpTKe1Em2ZJ4cxJApfvyrgiUNh6041+sY
h70Evl2auf8ORyMcHFsaQbQtbuTu7Mw5WcFfsfO2hX2TTEDFr/G/lQewZwjHHC3QYA3344IulbrM
wFyiHmaLOAmkeBJDKrumdhyrsy36bMrhkJWbZGGEyCjqfV7vQllkwJsknoz80izlGrmkdub72fxF
OmmhvSRNSVs87a8FWR8CHHh+TkUSpiuwRITrJAx3ah8FbeVttRu0fRHPt5rwiwu00iIRYlT9dCiU
z38NA5OtHoZmeX/L9bR9561AFbGpmWr28/y0krTEWBPPnRnZpHXez7+YFzzmG1KvRjjLwDmScHjV
Wc857O1ZGg3m+yFV5GE8pHyad5Ufc7JcKGC0DswU4tZW4PssSeTRvJfAwMYXk5u7p1YnxA0ele2r
k4PSvE/Poqde/hzreFJWBB6aLQd4X5pJ88IJvOoqexLeEy4fzFiqjXueICFfyrujqnSkaICTEUJ2
jsGsrzsdIJd/JFkfMRGVqrfHq6D5N1o9uw0unUm+TQQeW/+6ndmSf9KlCFibzfQ9EaI7oYC0UzNW
Uz+RsoU5NLG4ikJ0qpaMNLL//zFKKp5VKUVK2Tt+dIvcvS3h1l8T4+9/107iOC9LGkj2d5RJshDu
TTgjNIE2AS3zQHkI8SqF1lUJVU/waYr0ki5KqJeQLKKeHZuKlwTeWIx0wMltlVBz4jO2AQcGlW/P
V3wH3IaXCr3PNH0mnTEeKa4FyMERvcJ3DlR5eBkj3dGkxt450eI3lcVGVM0ifyO+RKP7HdMxTrNL
yE5MGUY9SAWcuUyKEzkemttOJQcrIDcsrMqIiTUFph56mVIJ89tt8iXmy2GdLkZuFR5oI4lERoLd
ntaesdV01s7mbdDwHxJQgOWUQ2TI3UducUSUOpAozvqEWL4uPKhd1L6faIjWqvQIER3nj2xwjumI
ZmYG2lpUgiqIr1eToW9tX3924ckdcJ09jSIN0PozFKbIL2tH9bmwxJ1orNIzqoah+s2qqDz2e35E
3+3fHOpmcTM/OCWjcwQBAWJxnl/FS/+PRcv8xvL51FrtU2vmwwc2b0F/lqeB6qZE1KGwGEPRr3Xf
6VuCeeSqHNFzxnjrBD+U3nMPPc5F0KkVK7y85qe5PQkARYSJtB7KV0UdkGqJ36/BOeX27QBcHEgH
VYQ5gDx+w65uv75vCDR89j9PLzw1KAB9IghUL2TDv4hyuS9M48A5U7kWhTpfOHrUOx3Tu4HhP6y/
9pcMJ+CkljooEPxSZgtkK78n2jGwbo2eBLdFeynlxaBSkRKt1IYxJYcaujKqTcdO98Zkpb0f5vxY
EEr5VY9SWqxHuHiSOdolOfqAtBYzW4uZq8fk6at+M2ZBb6T/LyBiGfagK4c2tCKWWAjBGHy8RDak
vu7MD6JaMtTebLsP9f9CHvFR3KUf1DZj6ttf1EarnCQVVOFuswgMUva1Df+J83wx93burEWG8stQ
ocNygUB9s8QQuM6VzF4Xm3gAtfOHBVx+9CVBHLsYNPv7XPrnss5FNWc5snhR7fIJftn6i0VfFB9K
rhO8etQY5I1sU4Y0FYHIfNk5pPfIQDzCL9r2KgIVFvrkvTHXMM02sAGCWYD5xsOJEvnrvylkqfea
6AX1+YGToQk5XyXHxZJwu9QZ8WXdlkOAV+zqLgpFDLk2abWhIhurkbfV3mSKtC7PKlpstG8eqXtw
MMyOkS6gXEr+guHtFUvUuVV8xMDzBQP6CLrvZ6AlaxzmzQRq2vzbzK/OoANPqoA9+4jJGTw/xExa
2quTKV0VHVWJa6h1IR2TaWmSKCyOpf2A6WK8Bo6Oi1rZ2QYz86UesusYF9W5gaR/NWW2iQehXoza
og2AGcnApsomESyYulBrEDMvNo7hVxo95vCGEoF7XFLNlQTMCpMp9FI398iFE4D+9FE6k47n/rW8
gkSGbkbUCpuQsNCccoGKQYb9rHP9Ra2/wHCT7Uw3ytE0UUy5Pi5YaLW9m7OF3S51WY/22Fo5rErL
ZtHt9AWjtxnPvPEUm6CRqaQhQmCljtzzuY3DR+05Wi79e596JqndmTuFSCX8ndce2XYyv0h5xbBc
aXQmJ+Ieyaa3mjtATXePSjA9HraEmIX2tiu1s74bw52CBXiU2428vwjRmjI4mPyO5EpGQs3oqdyq
cjwwkDhXjVXX4zgUJ4DNn1yVXBKtPdZbEbAnF6Z5xs8DQaGW+x/PyzvAV+NYNKUiP81XIzE6yOo6
a1Z61g7MOmeIewqUe6UiFMFE9IZ7RuJtgp/AbBxWif4wE6uVyiWvc74slPaZgvYp8fbrP7pY9yLQ
fZcvkhQ5OOqkHEc3sJ+RbRxNdN+5O5WtiWvjdXUORKJbhi9jdFZJ7ChdC7xYjwqtakot30oJuVjk
X0mA+K1jtehqqxGI2MaUoLO7wOVVpcPCmsrYu8rbkr/BWgffwZ7b+6XH3BrIia/vMi0n/154p6Sn
SGNl11v/2NjJQSg1QJyvADmCtqM5zaSCHblzl0PN6zsmzw7lvmX8xpR8mGYP9bKE1XPIH+E4H/4e
iXORUmMWpOHRrMecm5k/liHUJcHqGHa0HpE2+I82y54IIAaOd6RYVq32uXM+CDUfGwlBkS0DASrZ
QnTtWu6j2VRgDlQ55l5YHNMf8UrcXB/FPYW1rz1IU/DoVT6cKbqPpcCVLi9akEPW/CxyylBc/QWi
q6PYxeUJ0ndRTvY0+TdfgNQZo9vMO5JetYg4t0QIN3rTGnCCE/hon17OryBR/+IqfnuqQ5W/XfRx
JWvczR/+eUBCY8o9A9YIUaKygWRUFpVaLjzXFX1LVED2I2JTpGFR8lAW+2HEv1QxZvnTtKaSy7Ct
08TwlcmUCpZW5a0n5loNMod0KUmDJF0tINS5CtvTPF8TaQPhgsKauOXbHFFn8PMveucc8N0sET0r
lt0aqVeDG7kddn3letlw/tBdIMM/95D+rh6/M/tSY+/vtzeUYWbwZYoV5IlXtTLooyys/ra7zxpC
tWEiaJilaabrboXpItoHZZqhvm6bBO6cfEeLZl8N/aPs2jsq1HoQJEbwAdCQf1ux9je92c3Y/Xja
tzj6OML9B0MQo2AdUFlEp1Vp5+08KRCX9TYFpYdD9cmf1iUa1Z3pc4cqvE2Rw65U+LjpTw4FW4aH
NABFRyDlqhAnmy6S3Q3c55go7TRM0LMpoQmqQ8LPRk53SJ5+bFng5+WbvHOVHb1tFvtx8GLRnEBD
VpVoL0sFK63Kdlailaev0IbGTUsyDd9h0EaxUunJBKqiVr57BHG2jhwtcyDQ7twqOfMCwfUn7XGf
N2WcKEOkqzeIwHx9irhtp3yubIxhXDPIKEfGUEDehxAlmN/ZBu9bTCzpZCo83rGvsMvTroo1/R0O
+gC8Miuyr2J2PAzoY+DkOA+nRLYBLJazuXuZu0YTKln1bkiwOXB78lELUHGGu/RzhiuB5VUM99Lp
WeNmPXmvjm9SFBFfaUU4hE9VHiyBB5o31hQ7IVCcgFl1I4zkzgJNzIY4rPYr4nJ6Z2KtJbMuQotv
v5HKr0wSMp78GqqjDStHN39TDzne244IdNoeb48FxCj0dYzYNGft6h34kKKgmsaOdHNjhw1749TD
KD5Z9/IQ+djT9aH6j9w71/KnqaFMrJ9OswAI2rl4N5O/FP2kmjEF7SMemrwgzlVXNZljsl5Nhjt5
i0uWsxMcuD+lxJkov7KQ4eX5CK+50WTohjkHb849tdTUIO2slb1UgUhda16sgNSOed1FPFZLFkU1
GxpzRxAM1WXhyIyy9+nxTydYJfMByOAb4s8cD8im3IDgjI6llJUJuncVrsWIKu5nyn+rqBP8b7UA
2k0Uk+aH9iy6SE7qFhjo854veGCS+pwfG3+8Xk4BtGpk4hFh0/6Ij2DyIEURbR7LM8zYlzeP54Ag
LS7DKH3Uw5In2QH6UxWNGWPg8Yyj4GLM+wUNUB1Wi7hlv2kcO8tBFYPhHa6lBQOzsNg6MAA9I1sk
kmCBiTXfI8U/LUAUi3NvSuba6YGsLEZQWYxKgMu/KzI+bvmZX25xJzaavUJoUYnnsBjqxHqZDG9r
93jvgccUPc25jGkTPxmUQdzqiSZ+0j0BwMvXWxgRXWD8m4PTC8ZNPISTYfEwRO+5ZKXo/1EUySEI
vHtJwMLbk55QT+V5VKBa2LRcFALFX/4ma3lPm9O2ibaCFQBoMt8jGyygr6cD1mcO6Z0Rz1di9GcW
swT/TpFo2zrcbe4HIm1wNWFTnCzSEUojEspM4HUTBhM6Hm8twj3wVxbf+2B96qvPeYgGfXsS0y3Y
LxX2jk+UOuXg25o6PjLUueNNmG3IMVq9cfhFIXxlssgpjcMzl3r5mjeBNqWx8YkIwDF4BqBylEYp
NP3z7UTDcdE48vTGLPQyiCCzzlzbmvAL9Ie4WVYiIsSIEyQCkV3RoryBi50ISTW4igwtCLehUUgB
X+jbCvelEsxbAyY9Br7vvjpKVTjkhUgUd4NMlv8AXLEQNEr8zY61i7CHaGdM0LVoTEWYqwijfR92
7nt/DMxE/nrSMgMf0RAk5ldodot167/4orumiu7fYPo9KyopfSYf7d190q3rCxE+Qz2cY2F+z2Bf
yyhZwauP5UFfmINVM/uKXFpNXcRNnvEJ7PxsOyD1349lB2hbJxx2i8BYRu/zXypvMCsYQk/MjP6f
fqmannDopZiLnlQnqFG0boP+SqmEniDPXBzFmWG5EzHhTrBa1oYAXT1yDMK2E6pWW55bEHRSS0ST
jwIw3SLl2/EORZB1JjpGfObkFsZ3KJrzyS8qsG/6i8k+C3YWIlLulsm7Wm/KVu28vUSEfeluopc0
HbgTvL+mSIahIXfoetkx3y8XsHxNK/24TqaSiHXOBNGhjv1/4V2j2GhUTr3nfs6iEzgE3OCx8f/I
OBOF/vTSjsVIFywDkSt56j1sKDbZFPOw2TIFomDFypSKLrLcuyR5ENHsp1HDYPETtHL6gk0jPzCZ
jcOQ2smhNkcgo/l6nXHuxnJgNktxecMB9IwepO6/B06fzfL58vkEGsx/gJZyOmK7VZMIHxYFhof9
dg6T7/l7kZOs4JbGYN61zvQoe9lOZTDYsAWZbLY1rNJ5j9ypCYWW0DyZm/TpyuUT40K1tWFhYWun
kXxwanIqQSieZBpLGZEKMCHGnRwxAEqFVhctN9U4rO9k77ln3Sfk9/xK5X9Q2Noj11BEDmxgGg7X
ko5jPek9M3lFTquH5sNaxFUlU5fS/9P8wDgYMBLwgBaKsPXXRnB7P8kGr+2MFw7hcTqUCZfT8GVe
W9g6PS0mlP0nPOhtz5ArpY9GnFmf/MYG9a62bHf39dwA0Ubr2ngcLs3a55JNBJ8fEaM+DxZc7i6V
5wooQPVthLs4MLgjmqbPGiGXgtzpiAdP3Z6siZ2u3p90tDJu4nTVlqV1aR1q2oajwlsdjF8i/GBR
R9IpaLlij+dH+/ynA/7NGhdAdgtcQoAdpE4WOrC8xaiOYUDWEJIFXHg45+imEUdHU3WMvrzQznOc
tQJ7UWEXxCX4S39t2wJGYGdMZwej4c8BI9p8Sa6Yo1enLhHyhrGSPZm/zX7AK8TzbsaR5VObfA3a
z45ML/fvvWYFSticvks35YU6q36wqxYwPJqDdUDNtjLwpfP9WWB27CuRWbNav+nqVaZUxwC28OBb
khEAYX0McYsae6vzGkpVNJML265qW+WTNdrDctcWHA03d3Y1pSxP/BFk3+3oxZHC4fTDPElo2OuZ
CNp+nxKjc6Li+FxVTK+BFY7fMjVtd+K8m/HeQm5vjOLwCG6rBTR1QjnTT4nCI83zc+IbSb91pRIO
qsawTHeHSBIgRYinLqoVRo4oTC95lKAf86AxLiHpCZGLN8lZXqWCBUl/umoJdgXIcwjEEvccBAK5
P1imlYX7eXfA8Z8kAMCV+fBLxBW6sDJrmzHPrVBuL+sR37X1bxj3ow33FQmQer2956XI0CCH/IhP
ku2KgMKtUNAzTcB3rG2igcVOcGGEiLHX/CENcV4sqyWXkrc3GiVOUILjUUaV6tAqrEzC2Ozmsn/9
pbrXbM7eRwA3YYqnza305XtwW2+a/bc17PIWYB/9xwQ/WGQxBGXlF5NHCVWm1cSpL3UC3Z3ESP7u
V43xxK1NZh4K6z9ssKPf4WLUHca4FKyNyuVUSevPo+ASoHrL3bBReG/E1OkZa+RGkt4wz+PN9O1i
C4SWqVscva0Fz5HnQAFHlKLdmp8UwMtal1APDtAwyAMsZRpQs8x9YGPzgw/bM9fdh4Df6stMjybb
+H9+NFaZ8MufF2E2ye2eQlWVIA2FonbLgwpqLTNC4wESFrXSkzn01OsimJcqwRwBN3v4q7mzIwI6
qaGKaD1Uz4Wvq/i29geHHV+xcdODf6D7w/eAVDLC71ia3/eOvBKtV0+IehqUQWGmb4uM8XUN6/92
Rcx7axiyJEUxEINz+/OY5d6JeTKVnYjOucY+eWLgl+8QjAW9fmDZmivm8sf4p927Y0i/I2yjofnR
Om6YEYLS1IUHpeo+8T501Xz/phrPAjbJdDskT6piNdGmemvOsLR4OOwHw6skjuCpM8S/wW5N3Qd0
pijqGY1C0AyQVx6IfqHX634XpgZ0H/p45/KRlqQh/DdZmRrC6Oy7+pzB09tBPjgC0D/8+oX+ECmL
GY9B2J7HFcvd1/WICTR3x6bTPQ0uM8stLCJixQ3Q3opj6In+Z0FbbdAxkUksz79YEIuBjHdSCq/e
taDjwlA+naVIqQDQxnDptHmKOZHObbBFq5RyenXttgw6UtCDDKBjTuUOTrpvUbpfj55wFpEnenqb
wzPVgbxNiUAu0Muh6SzQLUXnfE+LqSDwrrcKdfBh/LsgH1sbEN/T7hENuQ1nvql1cURu/hLdq6yV
VztXivFg+NCTZ/F7/+KXCphJMIN44CGXN7HJg9wUtgwlxt/D0SuzLuQBrWZNGdhIB4TLOr+nAff8
GuECuykpsV2KDKH0PQfwVLGMRDhoQuIWbO3WV9+fdxEAboeksM3TZ7M0HVr62GfwscadgMYxAgbc
5Qa2TuvThz1ln8YBmVUGILSynztiWLW4yOXnruPZYKPcwHeeNPTXEr1NUaMTJJ6s1B7k5c7jQYU3
NzIXV6tzqC4nB4m9miVb5kjWwZ7QDnXmrJyFISYrgBhDOYqainrlFhc5YZ5qbAQ0RABDPR8Z4EvD
5Uma4YokuWpy4HvN2ngmBN8lEIzVK0N8pmAdF3SzESPIzuRSM+jNBmxQdnOv6MyAZMPMH8+xhojq
ynz19N55u4kMJZUF9+k65dhM4KK4AgKEepIqXswqkVIYo4caBw6fwA7RRU0prRv6ZnjdnnuIrgbZ
DGGY1SdtNpK6WmE9UJzUpiHZG09Dr7Jh2nJkqzZgcGZ+Gs9KWE9OJWu1aA6klpOGyv77GfaCGVDA
WFyQGJryyjlSvOtHtlKyfmYXmH4B8bjNmPiGQ5rFk6maTx8cBctzz51pyqRUsd9FFrbPxRMBzAEY
r+IEZvmZTW8HpD0Q1xldZRCT29wwdaOzD349sB2fRbgF+KK0H8f6Iw72xECPOrDbaYDC5IkD3Yml
eEaxCsf5LpDqZYU3sLynt/h5DlTx2AZ791/wDnJ3np4oo50BdHoPkpTQokUJD4KibLpCfcYz8IiJ
2CDGWt8gFyIX+m2V2QzoE/QbJJHMlJgP5QAKuEmlEXrA3W3q3fhT3t3zuTPVd7zP78pUfod7ieJ7
cmcFiG5pe62iytKz5kpdNV61snGP7FYg1fY43D6zhrgI/U2gqyb1IHpT+BzMbB4s5zNz7BnLqB5i
trkIuveX9tbQeh47C/jxF9SXvPGTJsOROEUh7HBhs2ZygBYmw+qp9rweT+rKECH7yTtKSBLidR4S
1eYabyngDmEL7GgCFBYlxL1UM8NfJIzMzg0kKn/M9ftZfF0O5tTTUbtl1m9NxQrQkKhLeseKhima
wAVij0Gicl6t1zgYD1LcZnGMCSwV4vD7NbYB2r3jg7GhMe2/LOeMt9RfZIDoH9pvgsjTnE5nijEw
ak+1Hq2vE5smwR5WS89vDmbCf7uiELf564hnjlAZqc3n3gpYUizRRDgjprOeXxECS9IZ1zVeNRBF
wunVJQaUwHknScwCKLoxUukOIGwM9tlwJ5lPBsRwY/dqiblSNtTYXSEKnNrJJI19WNthe5/LnVmA
ZiavM53ZqLmJHryOr+FATT/6NdvDwm422jj17aO6ZDE8c+ynIofsZsgUEYFyuAQVLDSgF/0ycoei
fuXRnLRoMNltkFNSq1BQXSL+lJGo4kB+reSu444lsN5Dgj3JiL59UjQKFqo9AhmTBgFgdkU+uIsD
8ObnBfj9KV58i+bPnkzw3/71/xQXzc8cjqeyfZW+w9AZfx3auBqSwhjZa/ENYky8dTq9sS9pL/DJ
gEeSvquiIeog1nor3EsxolKEObmoRaTK2vcgrX0NZ3IrfnQ3+ZRcGBr0L7PMbaObv5vnNdDj61MV
BImis1fYCp9bWysaZJklFdIIWDpO02eLoMMfliPmQBGuqDS7DerMGKmQKE5zzDNtsf/lnaAMkL03
cjDJ/pknhKgMtRGfAZV40LibjDZWUSc+0nUxW6zdBO+2zky4RLmzdt8nvxax4FZEpQjWmNh9vU+7
bcUisP2vyXmuYFPHcSqV9RolwjOSS/TOfkw11HuKWuolWxJ7x7tSr6pVUaC5eazH1+/4WeUqnM8x
Gqo7uQ2TMXdlmwyAz2BluOn9SECwZu56LiNyvHG0WWwpOaN6Kh/yEkX4ql0TtKYkdBBe8mdkQUN7
4METl/PTr+m8+s/s7rQ8wgHlt6goJUifr9WR7dqrjH/mYdhWsDvzueAoo4sdXRN95jGNKU64jEwB
Fg/b0BNnOQ8ZN+U/wJHDE+/Nbr8LoF6y1c+MeAus2CdeNVZwmpQNKXLxvKi0Xl5lPAsca7IvhDo6
2oYYCTYShU+3JSVROmvlLYIPDEkcpWSUhFeYVA3fjMx/yasPwVLSDN3zXMJkEUcvUDZNrAAP44nI
We+yxzemhyGtNDehoW7zAGzGOXvc9jhTpJwR/KPUYRuNrWBB6ftRh1O6klgy+YpurvtzRMuLBRd0
LckXmTN+Wc+5CNqWCGB8a1FZMnMz0aVsoHc/GYde9u35vcCbb4Z9bZ2atjvF4rW48JWPQvI0kg9+
UjSq+4KJELMrbXD8i9eEWgBIvPYLJSc2KpRWfYeuckEuh4LOdaD1BZFuvZjz9xlO4Ib/1zcD8o6R
4TkZbo0dq4nfYaHcD4UoLiPjXJlv7sBiQsKyyKcwulf+b206CER4a7WCq5wWPTjzb4xL26SQ6h0O
tvCHDNNum75/NALGRy788B9ttBKR7Bm9SqN1N+sFhfyxayc1Ey3jQPgpxlk53AK3Y+Ie31B0FDz1
Gg15IqMTYsV5V7rZ2xwrFNZUahldW8OTW1PXVaJ68bMXCl30hL7SIYCWjKqxrmGRh8cvLs9wibv3
Hfvz2j8Z1yyD6nMyHyIWCkpk102S4WumgzJfHHWpIfERNSfwiZeKkQHpW7TUiFETbC8KbSad++72
aQbruSIdwuChTaHxTtrtVPzBUhY83K8O+JbdPQkVU40Q5rF2TpaD5qz20KN8/LvOwQYtHlonOllA
YhnrsdUJSuMdOd7H72V4B+ns5GpK0KMCrhnbUkhTJ/sAlA6plSmtYnUAYped5zplNIUH2ySNZMXx
vBTSFk/18b9Jvpy5PsJhPqF+79zFUHgbnXriPUBWqIF6fRheobdQQYZNKcUE4seuxKCsLLjtrYL3
Uan+uU73F1NGvwLKNQSScPsQTrqKEPANw8mJM4XPBvOO1PchQoTXHFJpYl7Aqci84SLYR9LlDq33
G7LZ46ufH7XvrJBisHpjxuV5Rp5j3SULtG8hwApYiX0YUIOWhBxAXtuV8JLzkJX0mWTVeZrQHgWP
xUjMxz1+igrxWAAOlIzpq2nZxFRHWV1vtA6hqdnH8LhrKCy5wFXPrsfA46oAXmXVICcX7mHTxEC5
jpauj1BA0GmahnvgbvzmQ1xD2KHKFEbc9+hX7gmCBZUTpQbYqhRoIYsWnNknqFx9CBkWf2GT6icz
FXlhNJHd/P1GSbaMfWayvn2sMDYAdRtxg/4wxnGRvG2wesKgwiZ6VdA9FKh3FLJCDVrCLiXIB/jD
YleTkEye6HfIyct/u9J4KWu4DMP07otMQAdy75S1qeIRq77PJQxbZmWXkjqmew4NAaNt9PLvvXUP
+YQNxMtG8Y9PDuJQe3eXBT7EHLVOUeUnL+L5h04CQMhO9L4jz8s+bLQ26zvU/vlWNwpef1VwjCJw
7txfvUW9O1v0kakK4nsrDHKaLyXwaBlf0wClgj5q4i6Tg5H9SLIggGzz4zKwKZBx0aqZhkzP7bC4
bZzI7Us3wMR+aCYDujRpcExtuHjl0oYFZbf1XDCuzdnqh/v7HZs6E0S0v3E+kznZoS7yU/YVScuM
41MiuM108XxyM4Qn8zoLixcLW1AD24KwqQj/3L5C/N2Ff5J+zovfJD5PATQGdLIQHvnlPufMc9iV
Mybgk2EyTbm/aDXxMInUEhdh2CY3NBVjUY3eAI9BuF7bkO9qoydIdZ6erY/QfeB2iL4NG4XsqByE
hk4Z0Xj6yib2eAtLICUWkfHXo5zQZAbwBiAq8B3FwApnyqQ7x//cn+2bOtap6Mokan5AkXtAfMvc
Ycnagv+A30VjCuIxny45+TFwkcQbTg6gBgDjOUcR+3Ghvg+XA67bo/gH+C7y/QmJgRXi4iuUhAyD
i1QEtgT4M4YnuRWBYPSm9xqA3OGCHqmieLgu5V2J/TPAY8s8ctbUpzDF9i+M7286E0kpIjeRPcXM
JSnxSVFjlwypuU2kl/qcOr4GOwxRoA5Hzl90CdvW1PlAMLFJUAB1nZdeVS0JbXPV4YJ6aJoeGU/A
vGua29cJsop9q4KOU7Mgv8ruQ9N8zRffU8Zs55oVIALpDbjN7tV0QtzBRDIIBZhzLgY8fHc4zR4/
ZZ7XQ9gXM4XbVDTe2W8DY/Ps4lfgIw3Cnbz8Ge5DriBlQT5leL454q3o2nIkQJ495P67efLzRfPl
u8PtFS4jwALXc548E4m5OT5UNQrcAdm4jgCkrGGenILWV1DTSuwTJh88B6G58YiCQnxFL+Sv1tz2
JG1a8CsAgI68JRwVfHWx4KeEy+jTu3DP7HUIMp7EPqgdpEkHd7cZ10q5A9Jl8mSqdyC9WC1tLpg+
0hDIxF3JVXbGUz1RejzK0D8WKssOJO9y97f2NK/qr3T4gWgWy9XMpufbACntwS+dA+8TxWV1l146
OK9HqeVICPNOh7nSuiX93IxYu4MalqiqjECJL130VzhTqXoFxv6vOkk6Tqd5pRX/uJy6gHxVylnw
HImwOobAwjVcDZmMFuZY9HGDknxw84NNK79e4lt3N4KsqXBd3D7ee88QvK0gX8VU4juh1g0+tPhz
ifsvQUrj7hMGgpaFzMexocVnAstED8OHKstcTAJ6ug46DM6n55A5YlAi2o+3h7cg9eM5GC5RYZ73
J7pUnxvOeb6nr83MQVLnl54C36Mqb+ezN52VefUnCmyRgsMBSadCXppjJVnDmB1wBTavtpF3v1zI
0nbpz8uts7CvgxxJlW7+vjF/WZT02P8EIosD+137OWWOFosEb7vtwD0tV6nieURdmyk3ZnDyeu8F
oxPhfZAHVT8I9pqNgCSC+x1Lt0kpi635/ErdTA6FYtacSC5cSkCu2F5G2kGAzIt+zOyAgRd6VQ0p
Si5PQsHLLegXdKY87Q2/Gq1CthBbh8jTVAIT7o7ohYOSfX/xEa6U1o6bZTMW/DEAauVr69sQ72XV
w/b+GNVkhSjXwCuFjrd0kHPE/vz03EA7/Cv0jAb35wh8+UPvlo922jpHBcdPYI9xaRU90lbFFEjb
74eOa3RAancI/MdcjDRwO2u7bwOVULgn4ex1v3BixYQLLopoe68GE3+Sbz4i0TkncWu1XwhdaosY
Ve1jeelQxxE80I2KEJnLwJvjlpqIQZjVJP2+wZGgoPXyzMHCt8OaGwtRCc+NtXgiTP11vdP62Wq8
3hug6w95mQwY7mLVfpSbKMTqHXikaTPnNMBvC6l2atjp3onN915Co2tBPrdaA2ZkQsJqDyIGUQS+
BKZFaHZnl6eST9hFMG1HnHoQScL4vFWTIrifwMgXR//zo057zNa01fi0fplp9TB7KLV0EVFCFd5/
eBH+FWZ49ZA8L5JKTD7FKrDPOmDjWaN6vYq5poU2DqtpTdXk/+iGoKS6Hg2OKzn4yqTcBFQpTQGb
mxt/SxkhCAvLT19aauGuq7VAvTpi37B2CKKhRFaL4CTgbh5EscRqmWbMobippqQG99zuGl6jMI1b
suk3nBsAr9GhVZkOQIQ1/xWGdsbavpX7yXU09LDEZo3ExEv1deKJxM6KR6fkwfNmj/Sl3vGUbrdL
b/cR3+z9JL3EmAX7YydiFmKI5spOppmTWe/MvXCOENk2XZ7LVzOdju5vJ1c9nWicPkSGXF9RTZyT
YKNRnnVsptyN93qtemRFDBJ8GG+3VjQ04P4jasr4Y6qQnUl5/ENPotSBfjY8O4uh/q5yS9oW5WlB
fp0OtdiUUnGAu9uF8FRlwiPiy2R4IHZ4/4jkXbYWcK3NhOEY5Ac6w7lbbST8X3aBr93jQUCJtqLF
weoxsXNvx4nR3/GVXnmOekL1hdJfX2f1iXwCrskQhywnVpNjaWDzMpO+jTFj5Ohdq9n6wjYutEyx
2AbzoscOyiy7SgUGTlOX2g7XL909fZlLMfs8tS5IRBd1pAbMUgzAEzhxV1zOGTMC9qBvsyaCtg5N
JAKLudknwqcGJSvWbRb3Fsy/A1ERcjDSn2YwHtQZRD6Il4i7R3bKefito0/k0ulQcwG7uBYRBip3
QaIx57uetevqgLh4zX9oFfB/R9sqJlhLd5qOUHHqCpRAUJdo9EvvXIFilCkro12hgDH5BrbVCKIg
+H1FJE8nV+3YEpEPdXz1QZAEz1DwRr8zAeYTwkabZy8wlqcvu2VAD9+x1CtnU2j7idFyXTn3fu+E
RScsjZ2XpPYFGFArLkFfIttZMWawyPf0GSeKWigVYM+R30Vk/6zVHtY/9Dc+ni2RkQ/9L+gJ+DZk
f4IyvUSmR6vYMno9ohPM/Nt6svNrBlYJSivVNN8VJqUDRBRIGKNxFbAApKc7CXUx3M1ea9Th58ZJ
igMPtpFVTsoNOZDkMVImbKNrNkEicwZqkQa4010blVgZOsdCXa9ZO9SUbGl2KkgH1A0bUoK0ajw2
4crn48jAq1khgzK1gY3NKZk4WYOAuigu7IWrVh2/FXcsdH/fvyPB7iiUEUSkdukdZe9Silrl1dkv
5j9E1zofubwTTlIqixqm9C4qHfRvm7FSJX0JKbXqutJomfInwASnMFs0C/FVGpRyqHMNkCsfhqkV
dY/UgOjNrEG2mxPSyHRZ1BrG/z6R+p/V0ssfeSbubOG203Or+Y8nnx3GEekBpetY+EsHZdHWLNzz
81xp+HsIp6BqHfub/Puo6UkGlG38VhfSL/veLNdZHugecPZUpyOqRg6gkZuA5Du+RLLqZNC1Bc5C
osbMPit2sEVjhKwLSCB8mfnq8dIwFHOj2Z2Pnf7uteLvn+klsUs+Lv9v0/TQ1fmO1xzs4VPDNY9V
xNXSEs9aLy43uj4TzgW5VN5LDpDi6OyBMHJVQyQbxO2+TVYYRTYxPlaRDg0QigjEWDEoBUoYCZDC
Fb2DFnTj0Gh4/xOWcPJJ5a3LVtfLCR0HEwsZvFJrfKcWjNc1ViV8W3PKorPZMqUrPKY+v6JTe/dL
TlY8BKTphfFlA/V1CeQKZ6MzgbwsEWNdcIfoQobc7rDr8OnD3bho//A+gDHka8mR0oUVmpFsbM7H
o3bGg3JOBIt2j3c5ibPN2evRJcnD/uIUb7u0I1jkRFQy6UEp3kFUmBaQ5JDwzqmVKqraJO5BtkKQ
aDegSWf22fAHsI53UCWzK4+JYJUihSQ8TSR0G8YDC9oXJnmkZPYrvbO0bcqZ8eRF2GkKAQxttwDi
BSFbzwN0s1kEKQ43GZDLD9tOsV03KUP15WR9x9Qc4VM53E7HOvMLte3Ni+JTX5p+dRneI9u6zbyZ
vK9OpKPW5fnMTZyS9NXQv0yjPA4Fc5oZTYft4T75sj/BtuGysHeuVloCrRHyVti1e0mgdzOHS22z
yNK0M5GlsS0KL3LpEJzCLsXxBfd+Nc/KOW+W1Caqw3JWVyxdpTVscr2lkQArkDjzubpk4/5+q3lG
unJIi/3qUQC2eJHk8SKUbQVR8ah6AVfxdFaqRc9cztaGXVDaP9shozw6cZbNiqa1IOY/CeopEsjK
lWa1DtFZtgRDMoWH5Yc8wiOzDxO/jGsvPP4KdqT38JSVQ8Ra+xloC7v7JJL2H9iqYulYsUyfVWvl
Cev5XPXXiWl65iJIvH7Y9ikT1FpxHNIpCbcUepOOyBIcD/pzkFlHVreDnH1u/o9vevXVKeOQqay1
J1MzJzhrzn8gJODOb6r/DiYNAcp4mHGU2DBRXoz7IrsXlEm56gsA8U/wJvShCVwwbrK8Rag8TaKZ
4lA39IffQvlkJ2VStBwvonGYvmthxjOSPr7/5UAFOugIZ1XJGKGZEltjK+cO6aBmbS+3zwmbIZ8Q
hI/NytnrHrZAv+iYYaemADhcVx0pQMRWS13/bH9QkLGKcYcBBsS90n0dFaIB1wMq0xb7LAoNcRUq
Jq8Qq+vZkabDI/NrlDRRpSJyIGvCLkGsng8QEQl+QKG3x+0SIW+OAb576qAsagdDAptNVu8/7SKF
47NMsP6Of7n/b/Tny+GUHI9vcjCRly2o7Ej4klaULaDw4FpCe7IZRmHrt5FTokjgkjR3U3ofg35Q
9Xa8V+/kTCVKHuVW44IfE69K1/8QmLzgSxGWRm+5kls0gK6xAiRUk5Q/GzW4tgnzJebop43VQ1Aj
mQEu2HHs85XKDRO83S45w5SZNB2IlukS3njt81pB8mAJyUSqAwaKBVAfs+1JhWRECrp3mi44tBUi
kk8Pa9LhE6B5hXg3BQYsFVNKRI0fz9U6kc5NXURMFklNjqSYB53IBg2hMJ1Qy4QIhF+n0REhYpa7
2UtcK/Zr/6p1HSp51h6/34rhNamo8UIc/xsoVPPfdaSw5SPyrGIC07fgH9S8f5+lvEoyXdWkKYcj
xSqjLzZquOBrjYBE0TYRp6c++i+T1oC3Qzphoqg7yw9eLbexm855ac0n++MNpG1qt80vopzCHTWF
JNyWLfp7/Hz1FJKpA1Xc+u+PknnRtB7g7OKXBl978xvb9TyFa2fvLgsY/+lviOfEEI4tyVlWV1JX
6vAq8S3tYduXhk54YJ3jRlXE+JLAkuwvsDK2hAaFAOT7CvzzcjZcIbLgT18LYTgaVPAWhu5FX1Ec
NRQZuIvwEJEOabx1fzWsZ1dPZu2CDkfVA36RCdGKauGzTy38QrZLxG4CMdu12zQEPaNo45nrU7g0
PHvoYfjPCFT3XapFVoKk8iEMe8Tfb1DiTTP8kvmdAgLK4CS0ptnwFZ4Hl84o3yFw6Ws8AtUziHnA
+6t0U9bJgpQQtf3/5WcXmAmoZMAx5ZRCuiXHxdO8Hg1MER58/syhV1pSMBU393AFz4Mxa6XpOqqY
tH2133sfSs38k6kkd/5pvjZBVsxaFGqWgWT/awLhgrezv0WZL9hRUIZHz4w/e/kVDrzyJ6OGOUe9
SS2wLNSQPBu+2FBXVYjLKuNDw73w5+Kjk5wiOvIW8V+GTSUJ+FrKFhRjuOqiWMwA3MBxnDwYS160
/Jz2kiZwM5Y+kzpjwKdQkxo9ev9dFct5X42anwyaKiWzR0tcyJOdMnEoBy0B3p1Nrfo8cVmyfcbf
8jrTcCKemq54ntfIE8suF2nGtrxwxNL96PKKEiJT/JE+kj7gXYT96gPriau1RY0b5u+hJBCqndv2
BJXix/1JLpQblmgTxu5oVYuwJRAMqlV8+yft28nL1r6Pf0l8hJj6pP92fY1HDblktMC3IrImj5qV
54DJGvc/3kCJnukSKavz0sPu72u180R1neUZkZof1OiaP2vzn3UE8cmkARofIc+b7bvRzl/oJrVJ
exQUFelggTZsy0gSZai2pFnOijY57Av9RlcfGBxRbn9YBmuJHIfsl9wSZjdpW8FY6g7mQahoYytw
LGVBTpvzihHesVRzupCHdyem9On9fE2/Yd+dXxrvfewDY0YwQAzRaSY+tkTHNNeWtrGZ+w/Kc+4X
tx89zxOk+7NhfA3tHFvPwG9dS9ZCKKZDiyv1WP233S8iehnk8xyR/IyE5QVZnG9C8Q1L4cHqFdTz
Yo/HglBlLlHMx+uU2rZpTtyMwYEAae1PYrOasCX7U3o+WGqSn7oBxcxGbUtbMmpLtmkx+pSJU38I
aERLc/BevLmVQJkVFAqPvPkEmdeBqtVDlmM5LkQoatiD2P5274eq4RT6f25XCxKwcFYdqMncPm3U
2V8hfUBWha0ugE2W+KL1lWqq1JyabaQueZKCKYpAHCen4ATU4/ASXq8SRnqFle39GEOYa20TeAc8
paNtVORQtwZqAxDap5VMtUxD4KUpTOOaqxBZX6BfKTdSQUgKQAzaCjcfmaVkNagfBXSsC89wUHj+
RaL6m9P4BVJiNS7weQB0IEnITt4bT1CBmQWeL2l4Sb5VkG0Z5S1u0LDO5Aj8U2sy1MCdi0WsaOiL
s12XQ+yMBbZxhD6iv2A9WkzxcYyXg5kC1T6lFtKhzta8wu40yaFhWnNZsRsw1Ng3A6gVHWNPYSvu
SKd54jXWy7SwUMIOUdhpkcVOH42dVJK9KGPMwfdhD9m4TIxNRDzraGdckjf1Xa5w9s1vc/EDJmyC
UwWvr3CDPS7VRLz5+HEeeUpHZPYwUYSgdONGAHR6swNQ9wbzXqn/XAoAs79jZoCSMCALepQhkC3a
DfbNX5PcK9nFORGqT2HmlSNpmAQfsiX2S0priAhmET23woj/XF5bd4pRue4wPBVDCPwCeLs2c+IT
C/fulBsrQ338rt0z4vbRtvBJz/aT/nXFWzV2almJJqEWS52WEVeJmA2yTBgeZrRRJn++zFl+wQqh
vwvCwa0hD2UH1zSH42mNBvd6ayNeOjRSyEe6LDoZMzJT1oTvuCXYvO2QEKIhVuTQ33sm71sbmw9z
b1622Mjt62dqoDXVkFroq5r+9qrAa7HIhKQnebtTgGYN96Phs3sQW4Y2HFIYn3IQDJuXXDSbribx
cvLPuNlFAqdgyrDXYKMg4WIhsquXPb1k1H9t6Fdau4n66DyeC0QAZ/y+JU+0Lum4ie+HqNJYQCsC
n0Ik4L4s7C6brvvjNZasLlepuf8yqATThRw/ieRc3nwtM8dDiOqmO3XHQrrvwcf51WULWeERgmmg
AWxiirpMXWOppaZF0eqCohhNjRMEXIbNYk061uj8eVhqaG+jQ8b5KUsruSQrmcab5wRDAVJyG+Fa
Jnl89dCn7hcUXh6F+FLAC2hlhpXsJRrp4O+kwBK8gnPvisDhDJNIb1ztujBYkjoaj4yxC4MeHjvz
Ae+/sJ4WUBpLkXAe4W9347e6lr/AQ00296RVQ+Up6yhEwqqNF5t7GivOQnfgIEfbo4LrTWXpe3vo
amKaVDSaePAIpYuy0bJsz2CJjXoQHHBQc+YtScVVV0bjWPxG3kiXXa/WkuR0jB5CnKDj/Xh0R3NH
cTSgkreZyWW9Uzumej9eCyN7Smu9ZRupFNg5X6+H9D+Lo/PnH/u7o5RwdWP9e0kR5PPStTspWwRa
1tHeqQRjoX6qrc5K5DGSwuCWmSu2UkqU1lhVNL4C+xXdeyydGep4xC1ACL8O5OvMzMQT+nGURyCP
aiK2MrsWX8S/GvjwaW5KbaQRMSKR6O0nmAkb8oCvERdKY6TlqlbRtcNsMGuJTTt6b5PephmqO2i7
ZhIu5gBxn8wZVlQgJO7KKyKBz9TTO+mYGkGpc/r2QLlMhdIy1oDazlNaKLhg3ZZoXskADsRe3U7K
0T9O0OGWlBEyhCZaZSxjIrHtlPR4UAg2/yA7bCYQOKvbWjRkBv6Y8uyURL59ambkZnGYzhFu7tvr
/7X/Zz0XcYNz70UB4xd6DIqLidURFcsPZxfkocjzw/bFjGQrTsjptYhFQDBaJhMFMz5sKqY6c2oM
3j/FntAFMkqX2AlgAR9iZGLNcWKSYXiDGYehMzSjICqiRzihNGVBs/XDfJffd1y80KC5ibdrX14v
Fj/TihEJGss9OmvUBJ8z4lt2VL9kgI45GBOIIbr09rv3P0FJS+bLu8H4J1k2WUORHhVObs3dWZKO
Y8OLHTbm8qAbGpknLLsauO1pZZ3bJa0BoO0ew8wA/kGsJxSpKDGKHw8A8uCoVVIcFy0cbv38RvRS
VccVmFhgesOmpenxPc4F5FzhfZv5uigyi1ZEkluuVaQl207DW1ezlQv6klMFHipMVBA6iif9HAYD
o8HzwLn7nrQp+bIojbxjZsbgMLNiDzdohQpfWhDHGNJi81190BWmlkXq/KaXBXauuX/CnTxo5CD+
9Q4Jk3J/Y5IAbkCYeemNW0tc9m3jK62BjEEbeQmSxNpzogr4rw61Nkz99WBJ6ONEc3xoI8gd888Y
3AWqlN+qNhqoWzuYV9iVTkmjCwzPQNbpX9szL58tCDoyvD0etIvbp77ZM3V0Q9JNEjaibCWFDCvz
khY7AtceKiIPe4a8LHo5NXv1/79R0SruwgRYw2LlZ6cJ5oSuYtKIMxStfRZfekb2FpqCcgca6UE2
qxTVYN1Eds96vL2tonzcq2r+pqZBuPun9ISxdR5R49bwr4LRK6t5lpBfO4HhPQWO40euqBm01o2I
U5k72Q9dKtIVcJvdLOew0qCRONQzMAt5Es1ivmDOvoDQj0JZGH9RAsdr+9EtR9vMKAMFQOKheDfH
C1Q4B3FQplVOVXY/3OpvEuUBnJwKm/WMUN7pSaZIXtCqWiOqFLTr6tsDXM2Z2kraX5dFwm2yWow5
wiLemP1LHw/Z/olQuHPSC9AzS9Bw/ViFWJ9dYTVXRZCA+CBKEZuXy8OU7Dkzd0YbVvTpBZjxodot
PtO0L0206vusGnEaYdMGIxDtgDP5cLXpJp8t6A8HX+xLQ4dJw3T3yCEfsBS/86lBKf7ic6UxM8dA
LJQ8+V09lLJa3PT25CpwqGyWIIpYYpNB2nQjuOOqw6lyKw03w8iQMQQfvyCe4JWJGgxshy8wl+xu
tqYzlc8/YJYN18FwtV6Q2QTxYf03oziH7xpbnFriBDmW2ZAqK9gmQf2hEqD214moQfau9pYSZhMY
GXLu/iNC4Q/wp3+vNGjsNlBxq34UiX53Ve+2/offbcMxS98tJ2R1iM7+X7itNMShlJ0U8EGWMSJX
iXWVwAi0QBL0XN0XPa1i0lgnG8aIFo7P3OnL8QOxiBriuwyHSPxcW4hrihnLSqZCcLcfu7PEmKrW
jmZS8cXaVvbzWNY+1S2+AWqlA3fEFz6kxTFhw2El49qrccYur6Fqn/yYcqDpdJUtQI/VEKe7TUkn
+6ZP8dF7XI5g0WwfEjRMyTDZspasAbdeO3qH43Hj0j9vTO38OLfwtMqD9DaZOvupNqk2hhgeaXbs
TjyeP8pqgLUJgKlbI9tkM90wAVCDR5Sd7uJu3nnAG7MXsR8CCDwhmunw7ESN9OWNf3De6KTjNn/v
jcw2GXqHiTgChxTft4CR8NbD8vcRF5OKFxbblAqR9GsPHPdA1F+JGlAa0SjOtVILf21XXsmPYrBq
rwTQ5bLr2FV02erb3QoVCX0y7xf+xlWS4r8M0CFzubG+s+dJq9D49ltynHKFGmzZVvXe6N1ENS1t
OQoc2vidIels4amQ3dXSkSnVZNL5xeco5XeaEXdgl/DOOiO4E1KRoMqC4zDc5oGhwUcnLeOVsGM+
H9Hb42Zb8Di1z/YSt5n1gny2ykidRZ9hSq+FL2ZTPoKcYuUzwTCumBMIYOW7h6Ds7JGrbZowtAyJ
YCFQT0btWDE7I0KWCL0KXvqcZeyK/klc71I+vTTMfq4incAsjT9nK0rq5BtnCYyhaTZjzMAVCYMg
oKrDLcfxFB8Dx47rs39OLavh2ehsqPGbcgP5jJxFuAFA2zOXok7g0Aw4TIAtRiSFl3eOAlY1j8cT
XhU0sqKXbOwwl8MfJCewEEq8FSZjy9CZczsU6JJtvNRw3jS8azTY0qn/Rf6K9Ct5iz8rwLIF8JFq
/Y5UkxCrUrNsDfQqbtK7+4vxGEAaR2+oxdEz3Jgz5FQgiMbenBF7z9bCwdC75MhkYjNnab7FA74/
88kKnjcDv6XEOeE7R+O97oItb/3aVQc0EPa8tIysGCKG2AlXE4OgI/95IjzkLGhKHihQrFGatUtO
uNm1FuJrOt5OWz5S5UjYxImHYDQrmrPJO+9H7Gaz/JwfHp4TSsH04Mn60PkllpJNSE9iaTEir4lI
vjLte5Txp5R4PtyRCJ8L6P+Dnxqvjsr6HIL2jTZKLQ7/k3wkLIpfsDieaigyT3YyZSuGNfYpBsIN
XUCaMI3HmmfJrMzrE6PS6pBlnUdm1dnehyVicK+kBYxazrOCZxoEmNKsn/vnmlkInL5tC8QDqNxp
TwTkSlWjDgOn3Wy29tjwCYJ/XzzpO8CcM89tYbeT1gpe7NfQmcNnDpXgISP3RsIaXLLuyZdV1Q48
x6YC4MT2KpEnebV4DPARvvaym8h/PdASueLjEBvVDrPGTiO2WRdM3dkS8Cym6YUtF98JpNFh+IAh
DI4wvNmSIAEDAzkuoZBETCpCoPrt1Jr4GqC6u2DFT9BN0/Dpf0i1xmb3aeU7ALWAh6LYPjb17i63
MaU7YjrZlAwnL6VChVxpOsTxx5iPtowhY3+tH+AiVb7ruqCuuEPijxOLnkF0pV7TgszpQUTINP5T
KdEjY60J2WiWVGlCrXvvSOG1qT5TkhmeHTPu47ayPy/Oxw3j5sItwW5uHFLsTL79d9Ts4pEXaSzd
f4Pxxl7oJU0BFYwRs1gv5n/O3BnvMudxqPcV/mKDZvzGvA6RjUDIHvi7F8vpNMndxxVkwDyT43t9
+jVm3wnaxlterGAKdPlLon/G/tEyDAYH2epoc06oitvH0z77N2YI2BQ629q3UjbtBKiLLMWdxhad
0mnz9cRIcab+e3e3ipFeH7bY2hCzjdXj+6/erRCnkBIwVgz88H+re9+6tkDM8IDDb9SvrWG9G6+E
/BjSZacERXXDgvwYq8vDSTx+qrk+aLZou6XHOyR6n7d8qEdF2lBT8kI1AsgbU9h/VAajI307wtfr
kTJk48efMbSnNoHfbyAvozz+YBBPv80Yi8m6hPka6FRLmEPhDdi2/oRRWrVxC+CV2mDptg1etm+o
pUGjicES5wlYv3S2WLCQ2wEt7l/B5OdWYTojmpoTodXF6mj/6NyCaFtgbPRH12ec6rgg1dWWRMfN
2nKOkN7I79TGvmBB7Z+nO1znDc4jFlJH3cPMw1XQihOtbyGKnRnJAmO1jkaetyZyX1yj/cdV53yd
zREFV4/aSJp/JzNLX+CI+3UhC5mQRAHzyEuCZObyVb5SYd+rDfGIf26rjPgneMvUyVQjXvhtHuof
RvVdRYyTF5BLJACGGrFNf628UtvnF+Fo5keOLZmVk43WFMT5d/7CmhWCQc/Q7wT9mKfrDIlWSfN/
iXHnOqE9r4yPdabDg14TidZC6hh3G6KtalXiMf1zNv6cMV5IZM6A2tgis0GxcEGcF3BuUDRvEdUS
oHOax3KfKnJL8fR2hztIx6MsD62HSeE2pttKm0EoKOnLA4rb9yCsyNJq9j5dQiBZYT5XzUdHyugp
F5Fcn0Mmd5plzuC8e4B8mhgxXALXXMJXZZEDRQ0EUNCzcjy53fn+FejJeOhF2t/yNGyD1L6VKfYe
vqS5E+/vPz4/tvoB9G/GBtzpab4/NKegmKx3dG3Fnh/uoXN2ks7skol6YUWlhFvnDBOSlZM59nrM
46/4bNh0esyjUR8BDUc0fEzTwNVQktQy9kgeNsG19UME6qffxPzlGUO3FmDoWlKfahEKsbN11Me3
6vR1gzVZmIA7KqmNwR4+v8rw6y3uUr3nOhL/G2Cm8kJOf+9fgUdohc6AJJ1/HugNRVrj01otbk1J
3rV6Y2vJDilZCnvcUePbaHBOu1mr96D2967jdWUgpj+apGs+Lh4HNLG816tNElHPBbYGAYg8ooxn
nwIBhzSWjZUP3VisDD2OCI+LaOpAll+ycosxy7NLG2+UJEw52IonmQricPuLF4kLbr/1bOFHxqpe
0bkITXdv8TnwpyPnpmjrYoyaccgzr1MxiEL2gOOnJ8Gbz2W1o1jcQ4WM8kiGshfnLXk/Jugez6H9
/Lwd17Deq7e3hSFFgLPYUscP1sQR1LFCtceixLzHhBVLC3qNv+zYjc1Zd4SSouMRtnzXQRDH9zbM
RnRoqF2bFIoMuDEV/TwjUGwGJA7tXAxw8SfghmXoqM0zHlA4Yt7mr3PE5R2v/hz2M+E5QGsoP4s5
grl+XRwUTfSnxOICW+iIsGqhBhosuen/aN+7rDF82g5XqhZY2x+Po8L6iGdEZlFFFozh4KCyYXFT
EnVfWUB3f01IFAmlIrxpe2PgNNq6CJEk4YaAsFKq5aZeQrf6XA5hJRkueV/0OBOzfYYIRA75+zDx
yllWxIHkSA7A88RgXUVW94Fnc2UuIoXpLiAMTxB8XveT4kjVTRni+c4eZ+vxYTzaYBWc7Q2r/1yX
XeabTuBZrQepqJJz5r1Bu/CAOQGxltZzriG05rXq+NAGHHbHBWONLWLwvX60IxYUD5LYdhwReIYk
iJchxsTWgnH3i55eFuENQxgdkB+vJRrXK4yzUroWHaT0fE297iHU76cYsIKnXxNYKo6P8ygHn6E5
ris7MEHlvN44FP3z/Fcst1oQwOagSrIBCYU9jRcN6rhvxHMTt8N2Giav9m2nmm7IoKRfaj+dAq1I
nxBRMMMNZtZtsEUxiuZOxOt0SsNP3kRlUoG7JOC3vOhm3zQC28OoQZyfaLQf1L5O8Go2h9csfL9a
LQoU3jAbYa4+Dp0L14lDI4OLgtFCLkPX0FqrETZBTA7Hgl1UHkuQRwDEKHnSF/w+cGAhHVrgozLj
4dDHJH5gZ3NC6wcTDBU4//PtbsqQO9/xCMv1SHsTwka238tGxVI4wa375rVgn5pI6WWJ6QK1tt0v
PMOo80T6yQ9Rvv3tgpOFcT44MdwgpCIErQqmrPA7lWQ+LPRoOf9Okzg5izYMQ9a+yli5OHlD/BwV
4PSqEoUoW5wG02QlRHIQrHs9rm5ErNtRlgWp9DwFGmbpNP0QYaZ+4CrPEfC8TG4ah6bPOdDGg6nf
6AoRlFU+eH/mGtP6MdlswGA58fkNwlAMmr6tx2jkesEkkOJiBWmf07vN+GXJVnqGXmMWkk6Za/q0
iJuN6f/KVGYDPyHTXexeZEDHKalPMKonfVfGSM3/A6+/6zo/vBRCuFW5R+FezzVFCzDjfCh3qJJw
b2HHcz1ptXMc8ys9bPwAyTpgc6gvMYXTHT/AIh2RZq3SZf+VxEtyG0VawzXcKoRvl6895Tm18yZo
2t+BQC+Gk2HyKDB4ADsQKE2ioWBg2VhOHBgmGECXD89I502BGl3GWSHh0peTIM45l5LzFzTxd5jV
toQa833XqtHzZ8AbbHIo7T5rkhwTRdRUwNRXdJYOv9dmeycBgAxVjw87T6SIaos3J+RCUjk+UApc
+D0MN+foybOXELHKI+lbDXNioQmDOReSibMR7PrFbRdgnKKn+ql+ps7LJZXBXn419e9F+K6xS6JN
hvsT+xsMj3IHw2+pbfYkSgs4dGdM2AunEiHor0ys8/nt1qjSy71hlBYkzVO7fJjQfS0dGBoB1kw8
Y1fnZ4On2CDGI+36w54oTTOLa1oaALAYOZC6iVgmQmPw9fpgi8QdzmDmkXBTIkbERWrqU+cKgdmU
4VnI+bzLt1SFguxA4hhsSv8LTDLSXOaKch4Ajn1ppA0OW179v6AgkcEo3hrhhmZ1RFbKsUA1O9TP
EqG3lsbTD+6+pbqUlwgoz8JM/dEw/24wmi0C28WHIwozQGZ2Vf9OYokxRlAp/ShOXj2AGypdsbn1
5m+IkVQPUZHkzGibpot/fJIaN6xubD0AEXYVn+Ots3P/g/QSXBVANbz4Bztc8Tx3aYrsTW1gfUK4
p7Phnt0vr32Cy+zVPjqovjgKtEmUlXUZMEnwUgk67eQ7a8auUu3IHrTyD9TNRkhWddleVmWwlV7r
E2hr+dEoSdFlVdxWhC3YBi/0FgqWlyQuiqYIakhpduqi/dEUv70f9/O/eCKrb20ZxI6S9g5tPKc3
2Ujbm1pO/QiADua4n2s9aEgFklIK82lLcJir46j7z2CL1vJ3x+j9FLKqU3D7sv6l9GoEl9zODnKv
7CWqRlYiqwNHPMMEDwr3nWY8CnDjh5+gmDvkL2mTO4dCMFUmNZeYoPod+Ucya8iIF7yB/3Ufwk9B
y73pHB1eU2DVN9Ns0u6Hoo6vYG05b8vF1DYP4KYF4NB6O/KZ6SIr3fulDfhe1aiad3D0+dvmVBIy
iHNYsDW5mA7vRomCTl+CwKcn8Nt25Gtj5nx9Dy7dlbchMd7RpG9A9spBaSHtz3BCVARxmCdjJgzH
nDfQE0CH1SqdmTvsBB2EaNWO7DkgCXy4Q3cqElxZZmG9V+dVQsPjTjFRpYXZFN/6l1E5M1c1p6TB
kx4dd30UZjG+Un6S082ABgPbSXzK5aYGZ5+aIzOc79ukdDetGuhSQ4BiS7SK0ZVUySeisNcxgq9s
9QG82BTzIkKTrs5OO8xdKb96K7PkLBcFI0A9ui5RBlsMfJ8qTKZB7ORso0QFAoUppuGWdRIZjOp+
tOnvY5ho6m0/Nu1b9aMWkHCxgjOpKzj4DNJVv9R1fj5/EgtUqQj5gfRYFT2bkHHU8iR0z83TB2kD
UZya87DykEV66ObRK9FSyxsFpALCu1nLk4D/bvVY2gl3qeixafkNmL2y40Tn8npOSz1YpOCLywgD
JOgUgWbuGwyYjruaJUmoqR/ZfA3niLH3wQLoEtqvrctWUpdrJka1GYG2XQtllXP3xKHbsplVmWUH
WGhu14U9f1zIdg4G5zQnIRkhPASwMgA7dv1SR5qjad0BdTdsLsMZ+K4zHgI1RWjg7FCm52pVhGJZ
GU81c9cKsdBBTjNQY7TLi2/cZtc3AKU2MI8mU34N6PUt2i4nxvH7CXyQmL6rf/9TVSuEoeqk2BE/
9qbi8j/JXcdT+WZ02rVaDhglW1Wz0WNz7DlsmYcodEreR4JaUeyxafbEZphKJY4atNj6mqmxjnK1
JIaSbYVJVFHCE00y9zfXunNJXUs1mxxDoX7VjVKvQMrEZ6pGtEb92cI5JHgnzdOS3aaZaCSWYHD6
RgSQcWpXMxDlm3AvrGvZAFWkOXGrrxaKOHAEIRU17EDL2JgQ7ICXioLot/2e2EUrhsmg7bfh4qZP
8Q00zSvA+RDG+0ll1iTVvVLdjk+1D5wTPGl38wAxoV7/BeUe3aVZngwGMLGQyiq6yz5Lzxjs8lVj
1Y+nm4EZSAEurrfDbp/UvTfxoc1q5AYW2vqwQla83zoYbhLAH6dYwF6HZ8hi0DLOr2IpfZqQoPYw
mZufyn33QshRUfDaQnAXGTvVcc/bk0SBTumClVSl81bGTvTVVeETS6pStSHl3w4kvfp7z05tv8bP
wLcrYn9/XNu+KXInn+1hVKvNDBT8uCQJBZfb22zXngHm6Gskk/ajjRW+ndRAE5NOd8EQXRahJsuH
2pXWHysSP1eQEA6TGYMB03b9XaKtGKEOD1UpfLNF9vxYi75hwtsI5RBRoTCGi+y0zCUvKhPby0zO
La3UuwrCIxDNtt/r1tFB/VgeH5IaFuqGUS0xZZxddf9fGs7zl4mEdcTOah2dZQVbYEnKVlDRJD8y
t+JK6CSuKPuV7Y50ZNBh8rFvGsqwHd6ofDfAFZvfic03BbAW+Rb57LJozIVE7IVJ0pkgFiNRif5b
pAzFNTLJhBjDlnqhis7ApAVanP/s8leTOtfMAGBuDfg/jPK7PVtOg+YqJKbW0AJxJWq//tZ8lC/W
Xi0qIccj+XhMZmKNJbZbED+CoM5q+FA0rvAmBRxlHu6D/4xpgV9fgds55npKQ4hx4z40u3JWMEl9
UvbXkwh0XIaMrjX/vRXsh0wkVfYRwaQ7RSogEX+hYilm4MiKos1hnQLbFk7eh+kEazZM9ASblLsF
69ow+OsgjRb0uG/LOi7WI3hz162WYY9tjH7hoTonnQLeDON1JLzonHj6PMdw5T6JSQN9ZuAHa/q5
qoWH3LTtweQQZcfGp8ho5mTNc8A2rWQ/Put6iCYqXHIF8bmwm9/JdXr8hR3aDsKrFsEppbW0/eQJ
+LaQq6v62iHzPLhgWO4+o7e4Ema43JJQR0FI7peeCFbfDUD5CHiEM+2gxtwJ4uB8viyy4RSmp7HT
Hvp7hf8PYqaxwxoDLgc0SatnlRunWL5qmL00GkWD5T5u8Iv4bv7gTJHD7bM+WFJ37uFDIaI67vBe
7G65+2ujxHGxusWx8Yb4NWBP0zHS4Fzf3uZH78LspjHUYHuu489RVD/UmRHYDTOc53Sbi4nEzUeW
dFd9MOVc2PjRwvlP+btxvf7Jdzq6+97WsEGij7ypakxo3CpZPANPTlHk2chNU1Jec8BfjB2Dm0Jh
iABI56FJfBmbGe2ENSorYeGni1boylnYkh/it47zO79D2U+Ug8U8AVYRUjOOu92WUAfnlF0+MLhN
bGW5PZHXCrz57BrBI1YwGt68eKAwcyBqM8wd7Zj5P71/J5jGa/nAwxTZ7dB6uRXyAOZi6H9T5sL2
p6WQN0YRzNgZDBd0wKHlShkkMkUmBPjEPZ7bCDAu4yOnvE5f/p6IBxiBBU7f/fQ/dyX2TcH1de6e
kpTStbtvRPWvHnocFYqrvKoGDQvpLj2CK9UHcykdzfTqhyQkX4tgs87+/85o/fk2bV/ZbCA2kAG0
Xpx+wY/QBiRFYnSbEh0cW8JQ0oDA8pUWhpBqdnXhJDO4qhLR2HG0YKUL5XXvNAMMLGbyvQLK/X2d
cK8u78aOqq+XckobXeM+/RXMRXoJHuY6QZ1ynbnoPp8YcaU5/5F0hI/aOYjnOXatWsJ+E+SPObXg
kW9ZnFiHOdJLtFVdsqsQtL2CjFNf9gMUWlDkrsMfAjkM5uOFy4fm6RK7TIqmULSR1ock79fj0u/B
ODEKxdPpKm6ukIsKhNI233YuT7p9PJHzYkJUPT9+mADCVLw7kEfYrQP3iLhiDTqJFEyFV9T9Bk9k
7rVTO6Nl4HuwqWBEcyU05MemBkD/425DkRWayd+rPDf19w2byyICk8DhueoRf2adLc7TZRP8TMaN
lyuQ48qYOOl76cUYTDiLwoakxekBxqvXJdONIVJpcAi0sWHFz2HQIWDhxvp7U6N8o7aYEjL0j0BY
pYH8E8IbkoJAu57qhi5LI75TKEwDjAQ3FaRqkHYtk8F4ORnrsXS71wXzeZFJWhP21S8Pj4J6ga/K
DzXQZWpRdpt2Ln6r4rP9n0i20XUwsaM4G8xXiSJqSPvYzbwxOL+mEGG9iM56P63kDxw4dCNadF53
2cXr5YdwueGkqH/n/BT+arENrpdPNNCPyhT/ugTDfhji0THb6x47dm2tMVy97WrG4qx4JczUKcK0
Ceg8JKVBwtIlLzhImMPEjG28l671qEnylGiVkxVDA5iUaebAKGGOUgOuqrXfUPkgzI/lZhpul0yd
IumO670n5YNt0wJgCLrveEzn5QwiBXWNXWOXDygwbII9upyPasv4zXKl184PdXVF3YScARcL/l+v
CpOFYS0gcDFqlkp/DdCcJkQTgYy9vkMXr+79R2ZEVF36v6qGI/GakSA2tpfc7QFcQ05eNC/GPsiq
l+dKDjT4yRSBey++My44P+jNzPKViu0xBwg0EVEq152ElOL0E9W7wIfb+6zs6FtzdwYHqnGZnpiV
epWju4cD1FBpcx02ZMT69DRVUL3fctVrbzqUZ+IpsBc2bB4rjgxMZ8Bee+vQktBqAUrr7DqUKTD/
1pTZjtoimaIqV0805jhCDyymG5N/uFLr61WUrkREbpeWHnGGzTFCYJc+x9Svsl+P4yEpukdPH3jo
DsKitQJBAjOoXt6QloACRmiVF2GsetaD8CzVySoHG/qpSW+L1t9P/PuOHdPUukINXgUS7WrYwMeD
eEAVIXVNs9oZ7uIj/1juXLe9BQ0m77xhv00XdAH2ef10FdZHh3q6Iu98EVi7nP+BhK1RKsU38Ex0
gqBVsEe0sRn8Dd3oPyr+CDNOLbq5DG5TREl2Ts3qNYbBj938maz+sLjFimsbIZTe0YnuXxxmvqgY
2eYhTQZfLlBDbCdZYV5FeX6+RRH5sY3pMaVGuAAgp/FMNChhpN6lty/ckitnjmCK8XIqOZKed0uI
FqmbOVk6SUjfxO0tg2g1GwujrPWPq4UGGPt4Vhmb5fQficwlPSePemQXeeV/i75JHvXb6cE+47UR
fJtOA0M/0Bee0EpYG+jNb8vUTMtZ5r1EPwSDvMFR9GC/WV89Q8fcOXhEWS/LHXvbA8muAU0gqIKL
X1yTe1kkwLp6op0YNBFAeudiT+AxNbX9psz6buivz7uS21H8OGqFt6aQqviHTi/+1GFEzPVjoNjk
RxnpTFcCnpsfWXlZya842l7Nfhap0e5Rt5XH+fMkLZahClWl2AdnuOpQCK1mNhSrYyGbY/+szPHC
vuOj1SlyB/ZlP6HPygMCE1EUF9znSjeApI01vJHijIVsiZ8oT1om09zgioOSnVU0EGmShQQWS30K
Ce06UI63phOlwwBFori6Qy28l5rJxab660RYo+qf7FJ3Rn51pbVofu6anzOYVL4D9KnorY/PLPTN
vOI4mQOiRZuw9yNejbvYejfTREEuB+NaFjj5OAh9Xj4Ps3mGkQwSvt25BeN2BRaYnZeV9Xn6h75j
LC1iPzcdjLu9olZ2T4+RMpam+h9ZhjoBtDM0mUKu90D18B+hkyHFv5bmWT0sD+9ZP1P2ITk7Ye8l
pFZESIuASNbbyMtq4+lHy77KOpbprxjaV5s3Y8WbnnK4pN0theyrRxGKN1EZbXdgIxYYm7FUYBt5
4YbMciraI//qL4E8xjZnVH2nAez4guYIPM74YkivcuWClV6s18a4vFPGY8rV5mpaTxB2wAJSpxpV
4aIBR/yavQK0BPA6Zfm4VZSQO2ro7kECYczBwkFaqbOC9j5Pu9yZ83iLbskN5xPsHcp0VY4OTNRu
h/+ItLbkKZ0iM0uyJIHABI9IVaqBmo6oUZBiIv2WHargxP6lJfhaMHS9dxjBPyawo85fiZrb/iUK
9H9DenRDV2MebgQD9P9MykkhsRBXkNtWnnS/BC1zMmVMbAzEXYHECgmEqKAd5PRlkPfjZ45DFyVD
vdOv3ubejA4b+7+ks5Q2I5fj+1+XsBrOCJ3OQiUz/XvSoWBlPOJyH8eN26kRzUYO6GjWYbXWXiLf
F8NO02PCQAVwpJzRV0R60Hs+Sbd9e4NvdbakoPZhPv6Ra6IinE2tgM1ni9iJUz7/w58Zss/kITJN
ztQC8dg0zB2SxN7bUm6Ju0p42pi+32lKInmoi9dILZ+An9zM6ZKKN66u2e93dvyV6XbDx9GNwgTI
QFOQH3rwVXzggjpmgZDKfCWa3byU+xx9laiUCcVxoznRue8RASy2d5AUo2ExQ7SZiP45BwS+Q9Di
2Uu5EvyE6cJhxkEYK32YSnI1vrrqLEG1ThYl2uoHY5qS+3GAp5tfCcxInIB1pUL6L9e7OeS+uezp
pLs3cYUlBfZIurD7+JPW1lyYdnuJHJ3gqd8TQ/XqTJ6Z5HDuXzIG7QdFrTptIfO0I3+t5+E6+5KP
CzHsPptZE3Kt2IJ/7vNYUHOLK0RSPjC+FgSN0O7y9EJ2Q//hICzOKRGe94l5dALzVuRbQwGa4w3+
TOwNGnWaWK8X6OmeBsnsnemzWkDBgsdIczZVRpbUD4f94bIAwdn5BX9tyED2qFTYBuvoduioR6zQ
Xc62FxXbjZf3W5Q4pDVXRlBR+zVvnYvx1c8qrfqQ+3NJ4FPa3HDVkWWnBZmqFCTOn7Kmsbn1d66k
dB2JspNFUe2IDPvsht94ckbNEIvazB6rfw7qXh41QWjdH/zdF4x88UQAzVRpUFGEPLF0yAcO3RQQ
iOH8IW8sWCxPKvfpF5lsXYvUAQdYMInkEaWwanQ/jJgxO492rKRy/YdGOV6Abnh4aXhM5Rt9EwkJ
Qz8RBiLKLmL2m7WV1EzZFtkNcd0KOoeh/lT7lHF76e1WAvSCrElnW2Wn9vm9lqHhNdpAKn7GTzHf
Uk80obkLPVkYFDxPcJyCdczSEopTCZtFmNzPD6j8c0zkWmO5fk0hXQxYH4jGieMmIGJRAATaP5cx
D7N7dBnhF/i0PTEMrWrFnvjMOSEp8LS97tBVFljRpjHszXqGfzJ83E8SUb5yqx67p7v6kbF2aGSZ
0DscW2hdicdgPejO8jVyjyHFDNEejtfrvsGFEpu933U8znxjXVpRJmdAW5s9YZiEdayF32m86Dmj
TsQVa6HovvULYsfo3o7AxeAUpK0kfgx63Kmr5UIqABH+0fss3RZdK8Lbcgl01PN9A+bR1Hc9n5ue
amsbm5G++YtLvuWSfMpMghAlx+WgRYkgkQtb0qN7rlYpDNTmXLpIImlf4vdL4lASfJThYUiopqyC
Iycp/yK5O5eTwCmEpk664YIwwbc+mJ9e/XmUGyAaj9WCAdYDvhMwlhT/yDE58+Rn+CPnj4+4nY2w
pKei10xEaf+P52Pz1GFMjI1NVDHkLsw6SmFRUEXE3inXm0s0uZFWEwWzUPIiVmq6BzJQRyJEbnka
2ZJ8e6kLRY3bNgIrJQIX1Tx8ijkHsUK7Yq+C7+QViBs/2Zr25jtA7BjxF7sm9R+91zq4VF6OdxH+
kbRxanhUU7H1PhbZkDOzrolaKjmSoeqpEYvukGFrD8o9gkDvb0wRTSjJGnPSbQlc8uBuDOJW8Nc7
jWWTGyOmSex+YFybx2XXAXHH9c5suDCr1OcZvtihYlmCTq162sPImw+ikJC/xwl1jaCRknN29TCg
ERVdtCW8Egfp1jMHzAVE2hUtUKVXTCHSE9L3PO/aJxsi2R2eto+Uad8M4WzrIgKcTcv4C1g01fjf
hk3KxXIX+IEOHx1MHL8BPrNXFaao+NP2KvXF400B56FA6eG3A0HPAziaPgo5FeQB6GQkGnlcwFZW
QHWvGBpLRH+jjcI51256l04xixVHZoRiMra2VUULjZ3u0kBan1XyPQjoxsqKfrNE2QfCyXRm1DP+
hwp3WC+DdOGvOYKYjiBnkxBN1Z+Q3ZKYk2m6kf2jAdhTLW3T0jlLr+QDmgpPZl9qMyY6oZsw8GS6
16ZwuFMW1goluFBetTfXtLubocC3lJnhnm0W3iwDJuYN4jG//WtF3TSzhh2iRR8j7rPRDSKw4APc
zijM2gnhIHX0dopL3O6MZC7clPhsuHNJjk74y7EEBZT5jEKORH4OWYq0C5OwPtKh1KiPqqGGrMNq
w7mBLQnzWLc7qqudEn1JhBVxdumHuIKb4cGeT2lTUhc+8LTQ2mJB3/qQ+2XpI23EUdI3dAXqjLIw
TiY63cV4CLKEHD2fy5nZZisVMFIN5KqNwm9n8+PaI8C1LIGKrYLiwEZj5CINhTPA7Q7qKpqD9eNb
mAVK801OJA23tMg3E7H7HFKbiMT/GRkIHxlKLnz2qdnnvyFZNeSEC6BNIUF8H/dqnPsP5Xz4KniP
W5tLzdbyRiMwdH1klPmAXHNQpVKmfvE/XCOPe3MUcqgnCshl2z6ZjhcKa4CS0iMZ3Ss4zKUV//wH
0S7xW9QzR/A1SEWmVYjLt3DHfYtA1T4WJvVLk8pQzsDlGgZbjlNkez7XfMMO25zapYSMNSXL8wF0
i1Nilf/15RCcYc/gXGLPFpG1raI4fQ7IrqqGfW+c146XLvnUZA7zH088cCsdffswAa6isx1bO+Yn
VoNZL2KfKsSq2RhrN9yyBkKZwsfoiIRlV5KStJwcXkjeiBxheN9U6yCfDIK//g26rQb7a85KUw3c
ibJFoCpWmtnsjob1Xss6Aq+v4K6X914d/QagmHPb9Bx943+NKY95rLEKMolj9DSNJw2mpCIzn20m
WFpLE++dj/TlsyHMpL1/A+5VlmOpMHHynE3yeJRVcCjXBeVxEI7l3LOJZQ/0BPjYrVUt33tWOVCI
iH7GqDHKNzXPnuc/celAN9eOn5gVLlIcacfBRI7nwPGD1f70Dp14eo3o7intiKuiM+YPW5jRSlzN
l2PrD2eeYInyxlHwO5BzDPBR2T0dUIDUE/zy5XKuTIR52bmBLz9kL3LxPOd0NLsaVwgVn5xE8ASe
fIXJT13k/EKswGWLWK+k+PRn4m2zbX5NROECg57TUP1pHfGh7YJBJASLa8piCtV3kNVOFNX30NYV
cdIs+DYXIVQKXJ531txhaNaARoUu9mPpKG1SL421+Y0ABQq4+K4KpulZq/Vz/gtRixDhliUPsBz3
8pO1DwgnF69xv8gA6K+Gp+iVFy3CdMvB0fK18mUf5xlDk6dYDLgVvKGWR+fz6yFJPGpWmPM6nftI
sHsDz8cwdpR4mLNdftxmhNhMb9iwDyRxbdsc/3F2QF2VAQY89sP/9n0BhA9Xj5ALmFI4O7KuH76G
EpMykcZgivdAOTFJ/Mj4K8q0MLnaYbFkv7Zm9ZWQaAwHD7hEN0CwPyhcn5C1QTg7kC7OJnj5RrGk
5dAY7rmU3Z1t5PuahSegvtswx71wBWShOC5/H8UB9OlwBpLhcBMVM6AtKbjFkzsJjEuuWf4KRu9v
EjIS/gkkpFVzC77zukj73tKNttrnImr2fzIElQl9eiAWmFmJty3XXPe/5SjDv2IVjbo8Q8IGSVzj
wvCKn3m0QeX0jGvwItq+MeOBxSS8SPzt6okjPH5QZKWpsc4wlXXVunMrgI4JOBRjA13r73sALB2F
fLa3QMWJ360tOz1AjGHRNRFsN45G8+FkbRhbXUOy3zCrFqlVUD7SW78Q4siYlTLtBZUWJDTKwmrY
HhA5GB9yI9vfr9+KfTv2abf9MDjvhr6ET9EHYtl1VEdL8D7BSQR0gm8Rv2sEXe+9b9jyIQiGY+d3
nDfK9K9owkpCn1LHuA3l1lEGiUAd+j5QzvBTRSgzz86OAIPSZixQTOEbyM9GZCope6Vfl3Uk+twB
eb2T5TAucOzPNX03Jld7vqy4Dm0i8wio6tF5R4+MnrB7tNia12csVb3viNGBnb47hhnH++rlYy1/
tYPINmTBT+ZK9gztu1sT0AXIQHtqEums7UysEEBxy0eYBz1ZMkw/opBSglkdPlhjk76rxsNTc16x
ps1nK4s9QRoLfA4gJyQb5XxlscMikaWOYuQlIip3Nu8XnH/TdVtIv93yxO+FwJ1z5MHmwscN7xu6
SuLf7tGwp6wl2RJAJXoj5w0pJ5v0cgwVLvptrQMbTM8jxojQafyg95zGnvee1nW06ZCAlF09V37m
Z5RGiLBYzYwkn7UeDkDRWKyGiezyOeoGf/XQRuGUgzLJZ6kz5sh4GYP6C86NfCejaR2IS/x2wR81
Qj+jRjmrHrsMdEfI6WWC75PXo9U026O1hlrBO+8XpOt1JV2DEsYBq/hOhEDGblkSGt+BdbTc3Uzo
zvM9dG5NvmBEWOpXs6clGtC2o73YYCKjcOuFBd9K06swB+2cdZvcvj6euQAOnTw7wC2CKxwlvzlL
tz/vDS5LnqZCSufzvThHMmSE8jAeXlKylvVaFTF18vMbCUGLMHXG0YN/VWngi+IK8/rB39IKU9Cw
U7IPzvahC0JSK1Z2HT40/4pY58vV+GJarQCAf/ExU6Rd9Hag/A+m55VCp9mSplDW3s/636b3jf5U
80SxsO3TEuHmBDUStWEcjccGOweqhSb6/Sslyhe6791BZTNIOtW6HTP/WiWvjI5EcUQ79xISo/UP
7AHdGcTjceVAVpZhnWkyGTC519anwUCvYKaZ/N7FQaVU53IpUY2YFA54FHkKa0D9kGQC9NwAJs4o
yqZluYxC/W4NlvtL01z9jV0NRNIb3+MIp6yjszA6CwuxhT0cEa/gnV8v+5AZqRhftnvUsxCEyJHn
bkOOZWyikQvzmA9E+bQYPPmQTbgM42pVztzfBpc6HeLMmt3yPAx7FufVM2WgBRYQtmSG35Rt1mEt
pUaOXI9LUzmjU34SheOcZjBQU/AsxenkU6SUcPHQt6an1ZHntJrJ8vsLzU19ThPwSuTkN3fyWg9h
2LLvWF2D/0heMIlOR1VOmVBFkKH2iVOubSxNBvEoNnLAFK+MUIxOzeeoHfccXDQeQYvJMaT00ITX
HG1JZkBCfY1NxHywgy0HxP7NdJPmS3jtSmkPLgfSwbLnrCHCB4uJkd79dUqNgJfAEaxlrXSNZLww
kenP1srKe6g7LZKae1WckPTFpR4K3pGg5lIBPOJf4FW7ybc3lignLzFLBiU757JjHtfSvmU5ct7A
KkrLRjMHJas57fOfRBFfE0xs/MmidJ6n2DWJT9K6kFjc+b0lhow9ZZaKjSIKHmhM31yIj5b685JL
WommVHKrV3eX4OkP96xHCV/boiui/cEbmzzoPDbjJN29gw98q8D7cxHcp9x0nDWfqn7TUGKW0eEt
0Q9XRPgddPuWTntDIO5cLM5T5o05fSVlm72yu5A7Mq90UI9Z44Mii39rmG3D4Ubm2cEQxdXwFe2E
TWLshc6GuWiox7rTwMppwicy7TQEr90AKdqMKMSuinMYncTXZVQhQpe6JaTmhfE3lSqycvQ4uX1+
7G45XyK7S/o39pQdZawCJdYX+Ugcg8sfTuQXe4weHv2nNl8uHCzoeerNggFUZMSlo+QMjv7mjQzn
Tc10q6v7s7ky++V89XQWU+oTiW0Z71zxkBo2waKf3pzleTGO+KSMNmnB3kHyyigfA7Kbel1RLelJ
Hu40huTWueYQeoh3IB1lOjDRXzRlhnxVmLc5z3x3Hhg0GyvB19GwfdWYqMBfcBQ9Ktg+ni8dL9ho
3ewrwqvkw98TYE9FVSmS6QVtvb+6E2HIzMg4huQ4BT1ZPzw3Ja7VPmJ3IL0iwe74OuiI/dWQ5yBC
Z4a4OlslLrWDSiBx8fWXUPfX2qDyPRG3Ubqa1BJwlLTvwpA8SAGngdUbjiImgCEP3VM2Oj/sufG4
OB97clsvZVYQm2sAQxD8/8yKSTQKxnfDZxqnxDBYzIW21Thl0UuibjV15C/CayBaYgNOfDuYKNPY
hCygeBVJIwd1oglWIvkFJaQpddSKaRACvsTlsMjz5Xn27D9Ynw5xAJQd3Ya+lt+egnIECEzTurqi
/AtzFUsj2RyLWgNDyBRGbZnQbVILnADycsSqoeiNqfkqVKTdR+DOjizxPd3fB0fbmfLPbJ7kmWOP
ajDYn+LG3WJyNOfFahP9cDwsOpLNl1S1yXf3Ayq8fVjsGhINxrr1enhM7ZW8f2GrbcvQCB1tSulb
Hn3K5ougxNSYyJpFoMom0NJ1ZBgWpwu4orRdio3kVDljX2B1+TVj7GXRKGGJNkvMT1wirdlZb/mN
gGR1PiecE3xVdzqHiDKfUuMsYT0WVaputgJsLL5tarqkn3R1xgRaYILQOIt6dnL3Tjex3cq/d5nZ
lfw3DjiqKfxydCeEPKRzry74B3Wxl8Mburcsb560w3smSLKjdTSABMQofwo6wWrJBGLFUhPG0ucK
k09mRz0dCAWzvGH60R02dkO31bLNlKSXqozwZwKaMeBzp6jHfse/BsPBHMyR18FLNxP+Easqtab9
vXFYH4uHpsS6A3ukX9zOkk4dglvJLUd/2eQmeL+9G/ldfHntyEUmiHBHK9lO5NGl4n2o3176qGXg
VPTldzOY7sc2ah+hIvaZhKr+siMxigSGE1SOLT23ql8p5IKckFx2MzP3tahg6634MtefZjesXhrJ
G4329vptHyl1oCFlrmy/b7FSVuVmpZUJfKq6o+Y82fBR8GYuI4kDpMsQal9UeiPSkhx9G5/wx+mi
G4z2U12d8LYn2Zh9rBjK/8K/URWT/z+oLuS6c5qhAmW5JBzyZXXTiMzpu4fABjszq1feorDrNxNb
MKVGNFrgOJEMgYsPpB0qGQ1FTe02Ht2P3JDAziwaBGkd3ADSqOVvqYnFrG5MwA83mwCA/Eg8MNcv
MZnXYtkARWRwv0Hf1AeeV4uMj9A97/A10cgAZ69MrcVx99qURMLO7fzylu2p7K3tLJdh2E+f3EiF
J6G+XYTFKF1atOT1KWTZ0THpDIVysEsveCdk2TLwwPAfj6ZL6f1NpN01ulKj00KpMCYOq0Z2P3uT
PHoggvI6iwmX7DopKKliNfOxK3weh+st59dO8o7BwbNGXsYIoYjuICGU0rGp/gnPMIPPM5NZPob3
bACzI9zwM7KB67hrrte6p+KsEskxEwtolM3toa+GqpLRi/iuYgYxZruBpiTMkZypa8wHjz2VQ+qK
H/sBWf3yLI22+4FwcG8zdFgMtKiVEWPJ6zFOsDmR74LxFjAJ0GiN/KMUeWK8m+tvMzN861O7gV7r
wY5L8lyUUkZmKxmz3hcuEyFY+8PWjw9pZKYjJxswaLB6SOqH7KJCBidCh5tA8OaSUL6i/AQYUeG3
KVZ+w6ZUN4IrUpw8qeVrPDM2N9p1YwRc55q9rTgDXWREm5gAjlLnoER/o8HGnnjZmKXz8ZgXFyvb
mIT4GiJumYxUggd2M0Ok8/2KI9Bx4KPOe3qIQgp1oAO45kCPTq2j4Hc+EkXaYj7ZjfOrl397N8SX
j6gL14iAjc79nSFcMP108joOo61VlOSYJVSG5ANvC8/+qouc526tpZDNexUx+ajGQy/2YeATdj5/
NVJiu8airb16A5GOCfarJTgQqQMEKrZUOocTZwYKHrVz0ujsbi/OiNTOxfj91udFjO/ygbanUcAJ
am1qlgjI28Xmj4rowCqcGb9Av1rwcN2N+VZHm+KuFOaSr4fLoBujgLE0HQj3ScX4yL6lyYex3nRl
V/4aCqorLh7lRgTBXOMoQkB0+hSKaewS7RFYbZjxHV+yO0ad4myA3AveEjyUiN9tJm+JyWgiYq2D
9UjSARi971qBnZ6CuOUUspWEAA47SLD6sKxPCjfW8JS0jbjkEhIHm+XE81+rO65MXQDKbgK6tzRv
XLcwpUhAzDGetXLdJ0NLTSM9niZlkUaIqMn7YgJX4SHjTadXF/YWllsEFnpIfAOPDywnbw1izOVi
NzRnFZMs8qnGu61SudXHKylQMOU4zs9t6hFH59aEyToxgzutGnBJU0dRudZSA6WyJAKKBDtmUQbh
ZmNu8wpjDDW4yd8IIyxVBrsimIY5tV3osdAC3fbRK1y17xWTzACXCPToqtAmYR6jGZC2wjipULvG
4nYaqE+xFJWGxFnGA1vjdlWlvmws2xoxGVUtbqwcr9mCDw8ET6uDo/ZfG5icC/E8onUVkSAabV8A
KXMoLoP3ROa8Uc2lnLUemAIc6NyApibTHjvsuD1wfJLeGN7jCeAqzKIGcNis+WaKgEvnKv/tLa5I
oL/yR1SrKy1iLDhNbaPNuXLE4fH4Q/RCgqE5W7gI1yhZo3ykvE6Luy772cwD2CGNLGnHkiRNwPRJ
C6FSnHYMPmR+30Svjiv0N/ey1rzvm7p20u1sUFUKlE3ElxsVHU/nAqfAYJ6AcYKyZ4P89kX5yIfp
KRzmlnpWJveq0B3ltSm8HfdGizli4D2NwWeuyx4+Ap39cW59/0t9tLYZtXX0O9PhoiCM1wjyfMEx
pWcMsXFzUVnTUqTkLs8wHSTrQi7EfE+kTEBg8nDR1PD8+25NxuG6GLS3M99rshp/PB3wEsG11WMR
Xc8erZoQp14lhioYuQtWhFL47Wz/YcMi/iLvj24neGH3tszwllLsMwxabsDOhsXzpf2vIaktypgj
l+yy6MRvF6pB4TsteEDh9/CSk9OZSz1cySnjmwB7xELycAdnVGYYy0V9quEPdn8uJAL+8dr58cwM
CDuaAvI2WKijEDJZYD6+Z+4Fu3Bl9PwNOErzYj8BZfHc074l0ScVqTEkLBJLdJEwCvjuLSW6mtdT
8Ruzciyg4aDOfBtMcXqojzIBNyHnqGQULJntzbbL77LqrMd1sOEQpUZdQjDLzKPdumQKzEimWuBT
HrST46qsJf87ERNzo1JRXfbLq05epsPr8gS025osIMPHXaH4I7XbTRaugPbvgEXkMlEyf7O66YjQ
Xm6IF/DSd9zoOxONb0fiLS/r45JUtPXNZcwOiWpsM3pokdvHSnR5JKD7sGEbMzGo9zPIUGtHKZcH
xDhTS2Li609x9sZZBfD9cRqtr76R8JJaYKzHpOqelxhyJOuB01RV+aMpsqQxj3rq4Z6YageW7nx3
8orHYH2XYRhU7n//SLVd1eFhmgTbwSUU/ic15tkyRqGDuszq1+3ciq46YQHJAHi0kvj8pMYyAbnm
Yea64h65ulPVn20gFyG4rDaKHmYaa21k4UkS/P6ut9iuYi57s8kB1geuHbS6YF3vgOE4SiWt7eLb
LE0MgIT1cIg0LRlUw5iUgk8Ltjl0q1VwY8ddPMBpTamQKMmpMuqKozxvSOD1K3eJGaIuQnbvg513
ww6wn6XmqrldCuAIJGcyC3y4wG3UlSIiAo/rTjLi7f2gtBRDTzg8nwLCervyLtEypxq1SXGfvG2J
lwmbRBtyHWQEEyUU6cvLjKK3rmYQwywEjwz+NOeg/XSHqTmmBKCH3qoN/bJQklirD78L6aBMwUlr
O0G65drp/ZGlJqysJNf6NE3c5pVHSfhHc5ctTt+hnTPPCBbZQXt7QLPw51Od3tKLl3uspNNYiKZt
OFUNVlI+EjGyprQe7XF1FM3CHX1/ukvKLad5ohKvQRV9F/xqJ8gAuyQHAEKeiUA6qSV4HbRhXMso
hWnEbVMwilFSxUBymtKr1u1cJ8g3OkVmPNyUCforJabdS8SOJxQi0pkh6iUgdI6wPYkVlNPUQ4FC
kJn2ZdJ/unwrGMw/CVrKlU9c4ynxEno9Rf447/bN4WIe5EVCTFV66tPvIwLjdSmeURiJN57L7CqD
CUlGNHtGfQxKt+ES9o5gEfr0P0ZsQNp2XfhSBLfp1zLk6vsQGlx8iVstVHJDN/fasuRWEYK9GV9w
+UWnV3ci3/c1FN4j2Y+N14ZOD03/iuk85e0xIsWucaEv2YO/Sc1EwqXwfNMKb9CkRSMrOwfazxYu
i/yFqs+kSeSk7iLgcE3KKrhVTL/jre//7bhKutkC5L7ctwCHSVHynEjjiwlqICZ8Hry7+55TOX+4
0ZtVqTEtcwbWIqbrTUtT+SIgcdH5U14z1LpXTXbrpIxOEcLsgqV9KOnTTwJ+JfjW2IH26nswBR+3
3gHHUV3Vb1b2pyDvmu5D6L0XsPJhlfwb+Hub7r+2pONNh4zkHnhEv8NNptiTE2DUAFxPDlRuGZLO
dLpRVj/ihXjXDEKuHMWudDL0NfDhyZsVslnQ70mCl3P1zt4/cXmEaZCaFS8Nlbo2DJ3Q35MqGoSK
kv4rCJ8/EZzGDwtU5gVik/DJ5Dyca2FerZW6m5QkQe+Z2oMaVUv3auaYebgbQYC/QvciTbLy48MK
fz9OcJ93d2iPbDu677kKYcKwoLp6siye0XAZ9Gls/2FiCI7CEHGYzgOTNjCsxKC6yCxsj+ymuB3/
0Q+WKMBt6FN9vlYNHqVmu3vNu9WyiVc3T8FkG3lOhRTbcS+l3RAo8ixJWRLf93LketELdaKGnKGJ
ees+i8nsORqgIyi1j73BRq/cMbBvNgnbtpCu+WvoEYpElq1kNyykc3SA7gC3RrJijGiGWC/izOjp
eMENazEQZVWma/+6LRwVb2SyUpZfEQ62i0Eon9wC3O2K95A8J5Om8O+TYanazcnL9oQnzB/m75qY
udw9EBO+KG4Xz6sNNIqxpEIb6DaG+NnV66mOO1Ehj1K7tLpLG4iAxzmVovWlVi7dnHyof2xIwEUx
vBTpTNrAyOAxAQSWSyU+Dl+URWq2RFRIx4uB2pU/BfLh/RchSnOMZza9xs3JBC4O3Gu54p1hMrBY
qrN3imjCA7hTQWmv5dETec+mv0xi7+lKw4eFQQaOTKq1+Uah2XXFFCnhOXQpDP6Aq4O7i4/JaPK6
oVdOfn2fmuCWRsekM5lBjDRLxPOnvpSj6B3EF38GcV2BWs/VPEnYXoOQOMaIlNViFaIl4178XxFY
s07x6uJT19/wWY74CrojIuNfUwdyHeQLrpqT96u1y/k1atry7IT3UgExLUu7N3VOVJprvxFmKGPl
aaymWBd4GLvEykNrLQeGp+MaR6yKHrysdWTI4sQKxCQmKFrBOwoSOPWCft4S5uejkjvPoiQStozz
cj8Vead8qAe8xjiNoxKugvo4h5s1lYLxk56N1aR8rzRcKVonpVMGMZWPF7gxKiA4XFzgqnN/T2IT
AkBwzb1gZr427b6iQkBsHz0Q/TpDhrwNqN+Yg7uipVnrpm4nUJg0qhOLKNhx6YKcspAJ5il5jXX8
G0GYyDz8tKhDS3+hkTbMhjtDNlhMmLGpWjTYlFeoK/jwk+0ury94eCR3g2e0UGyijlBuoGFHX/Sk
RNELRcGCpU+xXB89VcXAcmeDSbV9CZIMUaPUlbtQHu7qOB5sED+wJg4/5b5Si536rAEAPSLJDZKi
ffeI7cq00nGfsYKHftxNLwSXxAIQBDdsyhixWLRVSM/bMUZQ/JlNF6ViTjow07DNxI3n7gmwXQGq
6JlJx68TjZQrxezv083IvzFRcS7atVy+1dBg9tZRpCxvuaIUET8ixLmo5nnL3NPE7/ATNcznQooY
EkIjAkNGGd9YIYXNWHuRgZMHwn31wwcacS5ZDIzpy6bltfNbS41yNVKt7f3OuqERkotzG7iw37y9
/WA7nX0czV7nHSTBzhFeSfr0alSCohxiqKHEgWeDC3vWCNgf+xBfvUGtI4KAkDcY9Aj8tI5l1iy/
n+2nQZHn6Udd3w7kKN0KFO/Y8a03J/9pzdQNhIeS6IkPo8L+psMpbdorL6X8V5SsntGcNHpe8L5I
uPiUQJ2Ebta1NdIaYN9n3ACIboWcbReewgk5RVq69Qf703h+/Y6R073TbAE1maJOg9TMhD6vrWr0
I0HDp6moQlWzgaJeeNgJHpGhW7gz++OIiHJf7usXcGwxIaxh866O1eMSBb52+YhiXlD+YpifK558
BdDyjGLk4iHiw4ntkViwFcZWW2OmVz22aa4NVrBQL8FsyWq4fo3JiST7CL4F/e51Njm95vnpCKJF
IwRO9cqylubnig6MXNtcScuu5qcMy9a4dP+bywKopQZBC4N8XbOcGG5ARilqCoq9Pvmv8tJVlwJa
NPHFCxwwINFgcN7cLfzx0GpKJEjIieDtymmFYWL2B9HRK4kbu561mWISerlciRzZWPFRjNG1nj1a
vJHc6nBtrp8YWjzfYnYFTg9qQs9sapR/5b9m7JQDu1YIcYiiuGkmzu5jP6grw4srghHJcjz2rBJe
mKRgm4+8aG/LPTJxct9ClpazHeSNOubWsLNnOvzoMwtkC5LXpOKGvOQiWEib4h4gXOP24pWLm2t3
TaAJyjCPt4BLu3BwsrYm2CjpcrCwReqrVAg1qe8vcyaeGSvKv1tt1OijZII6ixd+T0a2+6aWKD2j
6n3nTeX8MmEbLQdHUrkHNBsnTttMtVnaajUsApw+YvI+MAKrHzdd4KKYOB57HzvYupxQdYf0Ymdr
1qiyMzcrwLQatubDxym8nm3C26wzzgU+DEH7i0+TUGP2M1nGZbpDkKh5mqBVBHj/rb/8g6SSX/qB
AmZh5NBeSoy2/R/s0c7q8m4wpSa/nT846Mck4IS9tvRB+HCyj51L/W/T9w+eqeGH6clHz7sUCAgX
fOkoUh6RC5QTl/cjcctz9P3iTPpitwZOoTBlRyMIVM4ppv9WvHksz81ohxEFGMLZmNT8W9kL/YD9
tw1dUHlYaIDrsYYeVAvEjY1fiKfLu06zdYrrJEGw6B1JzEv1VDBmRdhTI9n2GaYXvf7c/rwFfvdH
vwTmYk03PvMfuokfVqGdo12XWwAWCBVpIyftpu2pz2DVco//4bTJrju5oigW5kiBdm76x92F9diC
8YZj3bOMoPtbISNklapaqiY4FPTzN6lRaExcWFlBjQUzEAgVSbS37wWj4ZfIK6NaVJzSjRW2EnWL
WVxUxQovZIlZg9NLQMbycFGyWLXOPjqD1S4YjgMgLTMF6qMrzZ+4+44rzN4+VtYQfTDKvRcdsNDz
2ExyVAQr7xQzwS/yWVTK8Ps+BS9t8U0QSD6BcKRUjoJv3sxLuDj/C+VigXyT72UnBul7I24T0ycF
Xm9bCyGMfptBmVfrdcnXpQ1Y5HWoNjAxCIbNDi/zxKnM5G6aQCoQqjGLzJc0xFruPuHtHHVDN6RI
snH8dpk+Qljj2XTQPlpTBKPA8xX29Sf4BQjQF3Xv1uvR6w3p3MH2LMCJCLNGpqdkSQppF8Iq28H3
N2fwm6sN3MNVlAM7CL60AZ98u0cKyyhzT+CWEOFO+bO+bKzae8jkZe4x+SDV0aCs06itU9bPcFCC
sQC17DlI9GSWFsqh8dpTBhwuStVwyfZdiO7jZ63JGNOAcHDhCLLbDruGfrZ0l5t5rMcqq3Lri5Q4
btpO3yNa1fRad2c5k2e+ZVAr7jGpw4oxo8axXMRB5ZmpO/KqjnD8t5tn3LrzvauqfJfHjoJyFApi
Hr3RbAMuCQnSPX/et9CD8jJYvn3g7ALbGICQQfhVjWtTkz0CBu9ST2NOfEtDtvkWYLmgUJvNWAdD
kGKQo7rj+HPuQf2LdJPx0rr+iRG18/GzSRK15dhvn4L522sZimwL5cavsY99gF0bL04C4Fm7wcQh
uALGklD2ess4+tVLLF0Rl7dspbRNDonywiKmeFDKp0IdKlm77Grlq8sglwgeyMoYmIyGXydOiaZ+
yasr384wpqKol6hF/qBI2/3atyQiMhutOmS9LZQaRaA8A9D1wiAMtYlZV/CTeAKozZ3zhNa55Ohe
7D9Dxomb0fs/XeynEbK82iVJ8tGaZt9ZdBZdTJalHksjRIzL9Tx+sQjeo5f11OFQhweE8tjsQzc7
aJdmMID51UsWQFrv0ByyqIMZiUeIB/Ou2oVUCviFDipwgXtAyKIsj7bcBP16jvzawIibulBNDGUP
xNgQb08429E9r+/GUkzrrEX41ymI59mzdVkOIceIoiohAfHfBcuW0t7WutrGAYEgg9IfAJg759eC
fZf7Tza0X2JXj8hAlzr0+fAFD3e3DHaCzY5N143SlDb2jOGjK20Bqips6BY1b2gyK0DK2LNZ98im
SA1vGBIw0uZ52WdhisDuNnMFNzRw6n6qDwcJw0Gsk90OMQQ22RhLA1ITlLXtpKqSJ8ozq59kNELC
Ce9EEFIqeHq8veU4kAL5pXCjhscBI5PMtvGuExTQ2Te1ito7y7BvYNObVmMxvn6jDaEFovA5eyIT
Er/3vrnJr8uloPNmjZeI3gFAgiJNm0fjqtWv6mhIfG9P0PGhrILhorqrkxLcak+db/uIZvhxLu5L
aaPJISf7Lr3Yr83uzbLxPFnCFMinIFXWFVbGvnlLQvzQ6ByoLaxrGo3GauCDor6uzwQzP/QYbdRC
1I8IWccrIX9rvINOMj1L4X6huDyXW+ywbOldYeyMHrm9mi/lr9r2mFUCLbOlZpmx+lXrcPqX8Lih
2i4ZTqwikiU80DYqyoTPhnSiEnoB+wUu1MbuYwGXUrdCtxLUOMJIFnuk1ntCFVJYr4ebrOrUl3AF
opQ9q00l3Pe8MB9Tj8NeIsZVxuG/AeNwlPiniT1Cx+t7hGQaE9f9TZ0thq5BhHQmeBDM4Le9Jktj
0uLYAmppnBaFBg0HaEAVsSHBa/zDLIU96gKt432eqgMN3Uf17DQzTlGyv08FfhOHIhK5DP40bJlF
PE4dElooL8X/hCB9YZRt6wzPuLbw2Wl6JPG1l1+CplhCoJB51R7YfFV8vN7qoRl3WKTVqQizTlzk
y+inwRIIb9LmcrjocjA5FSpfT9D/zDu4U+EM2rKEEt42iYuKwU2Y3yn+ASMdw23kLf/STGEg8Gso
kCHk0IXkmqATv7vq3iCWuquARMwCibgoxzRv3Bm27Xxy818vLGkFwqQAFzYyjpC9dBw6wR5b69an
8sHUnDtizUbV0Y5PGW+r50jktsT1SSM50YYGYdgp1wckDUIyXFjIQ5/6lBFC7cRu2l7AIVlJtRLn
MmtCnihNYc30jKPgb+WGkjw+hBLk4d1URHbvEN4mpOTKDesOTbCIS2aegodfOLSYZyimwuV6bZBR
uxbZ4X1Vz2bOJSQdEU+ckBCULsFWdqLnEwP7SA1NSykNesIZ0ogU5gI2nlJVTRnPER6oFQ8OwzFm
dMqyjeDJCkH3ICKAIx8WQm0z5ddW0+BJZEmaWFsngNS60kyVFjjrJQWt4Zk5W1Kz2HEp7P9yRH18
LurZc49VTiBBjLnBYg8EiUKjVvLnEORd4RSJZL3xdah1od1SdcYzSRhLaoUS6eZmQNySirTtUfOQ
bxvXg3To0UOPCAkj9hVmhaf+gEmTcERV0thG/t6kYgkViKclJCJE/j4y4QJJ5HBUdbE52moaiZnq
AtwSS7v89+rUy/nizkUca+F0nDYiZQnQb6lQhqd642PPL54wN/vOeoeehnqycnSbRVE9StFfKoi8
UKT2fgrklWY7o3um2RnraBmHMXjEPXAdnkrMfnpSUM1qBrhK7BGPnqOsvkflJuX4ImwI9bHesVIR
lqy5uH3afeF+Bmi0CL65GEZ+YnS79TurKjmGg9rJs/scC0UH57n90dCMZ0YwqIEOYVftWTdqEIms
52Rbq3ueHLlcTh/Esh3vEcSjnUNFTZQSgJ391ZzN/mxRUVb4idV9IifQYatWjMzladF6OO5TOCzg
3XKXUnhAd0j0dTK0OB7NL184TnHsDisPTAwq36+lYYSkAno31cm2yM+MJ+2+jukYY6Ed+464jB2k
gW6eBfPhA3xLzlVCA/bW0mAt/stY1FpF8ga4DvXb8eqi2g3qUbtJoRyxsFESDcxJUK/1TDcH0GIt
+TS2sbf5V4XzoVIHqxXEdI54ErGTBRIqqIgv72cPuU+9SoGby7sOeG9r5n/6bqOUgw4b7w5ThGuP
jUXv/AL5OpTdgxcyJy2qhowYKYse8Ds7OOzpozgQZUbDyX/9hb/+hFZkIds/fawtKO+PZ4p7mlIu
VQgekiwfPCiznqiNhIso4HrdWfbJ0/KwT8uFRq7LuixyHPSG+HwJ3UkzOipWRNoM0IdL0MvWJlmm
s+vjJ3gAztooRG0kxt7XrT3PWyfBA9i8PGAfaS0mfbWzdx5v/tduNIUqr5sK51QGsWm3LYrWIToB
TGxrpaVYuKQnSckGL4ACGC3dNMfO7ps56RvcoOTQnMM22uqiz3g+625cmYa03bpyjZiBD22hVeUY
KOQd8Vmrk2tRgg7ruERgw+3d2tG5nBEJdmzX4LAX9B55gMH5tTCCZugPQqs5bfe+pSAeQj6+k9TB
7k/Iaw7NyRdKl2RqD0FKaWAyflF7TjLTFxZ9hj86MeVH+9vlnw4V1cTbPI6Xmytq11BHKgg1Be9I
VM8nekzg+D/5eVB5JUBa60aHKesZaMS61ogNpvdD9Uuoj+1IJ3DMDI0KZHF9hId/KGYNCJrIHHLY
opdfnLy8UGorgVHAd7WUsD9gmHVNkTvCclMlAEf4TSYA4by07E1V1wJwbYy34qc21+A/DRf9dVg7
WxgRDp06MZxYx+fEPR1d9vZZQo+BrqTLYGi//On3PhMIvKavkqEDMALUNB3CdYUJG8tFxh5xA7ov
dps9LKjF4z7+75Zg04w29WL4DvOq0fLE+t2dGxDUUhbH7DhrMaSa5azIAf5JPt6O0yboqBRtpEXf
aWALFgRG71Ry4A3dfw3a5YoPolG55lfyKVTE/83CrV7mgIWXpSOTziP6E/yKKDTDiI6iHSLMojn3
Gt3rTfzcj4Wzxm8Gs9TMKt18DtmH6utuU0cf3Rtnqe7TwJnyzN6tse5MthbcV7agL5bk1cYJTzf2
JfQUfENn3D2FQrjM4gL9BEBF1sf+ACgc4EjbFH+a6v/ln0zgPCcjNQHut+snSAhkANXTTUrFIZrP
+lSKHux5K7o4ZUkTxrR8tMYxzjhz6rWm1kBHEqhqbpX7t/YrS2fhxYHSljInqw7h99AE0gqEAyCE
baxidMjTo5kWNghDL8zAbCry1Rj1xbLvT6aMIXO7e+o9wsAMVZ7Zzk3DznnyAKfqGKKU27JrbW9P
m7YjeSuv6P44vuM7I8/7invvDiEDKKkgeoKy86tc2U48BFvwK6Xh6ZoAiUXYWNcaO9MKceWwfwIU
IeEscugyh36lkpiF1Zee53p/gPKjJ5yex9vYGaJbgjAVqLQpOu1FHHUYaBGt/CH9mB6EayGdJ23G
3zwO1OdEEcf/SXJoprUxzfIqDJfNM3ED7hSTwX5b4H6ttII3C1XT+kLa1JtEriNOtjxnaFiKPCQA
61Zd/VQymLbyof4loqorkkDVfH9nq3+Hsjba9jRACz4dmIW+PQrRhxkdi9u7gXuP4+oRco5HKL1y
YSdLCFMZn3D7nLjrrKfkYlZ3N8mwAMEodOe4pIUXmyDY7zawF00Unk8xN/j4fTUcxOSC4fQjOySm
bqJ6EDdtPLIZGpvevLaIpRIcQ+SfI5R15Rpbn9abMCyHVTZ4HcElV3J2jcbfnGHTY1hotP/yqVWr
pzxnBoDKIyQoe6r7UZtphtpHwmpRsfzZPvoX57DXjYxNzOsZgAonLdsaHdFk7ix5qFflTlrHplWk
EhopSNEuYecqKzDKgNxYuZQKhWvqCZukyhMzTLPJQF0h4jzCy5HAZ5GXMpp/e0t1D0AcnSoehwKL
D7myvAa5Om3pMUPGs6LoiKzFgfIE/vdHLyaQjduWlF+BN21xI0uLoruSa4lDW3YJB3bsMueMoSgA
CcM9+UScG6zjsBIYeJA4vUxav5xtMeRhzrIzF9w5900hvy1chiMc4Rr0JXo3RowFUZssXKYO+C4w
ZoqTiiSjnxalE1qdD2BjL4BLPNcCrjXt12vtYSwq92jdFh0XETuA+hOj7om0d9bjd0OwJJMlwzIo
71JGSJRdQopvJ6OCh1svip8DxNeGK8zRz9UT1eXPCU0j5SJwZQjfLMTurtD87IVbYzyoRix5U4xu
jTbV1PjT5T6YMVwSFC6m1taj2wJSDM6JsM4Xwo3c8JvQclr0YSPkxmm3flGK6M5g95wAH+7agiXA
HX8RR9isvYcVd8pWi2wZN5Eaolc7+UL0JaWyxe19vGaaSDlrLA4ScONQNdh3ZByzGghEq5nWxUgh
3tnOOghnmPi5hxhET/KC6j45Gkf36Ae2kZpshaehNav8X6RpyBV1uXvpPq4U9+HCoi+pEVKxljDz
s92HU9KZ97gGQ7NjAoCU7cynYl6V8jriosBY/dZjesBkeC9Z0hEU9bylFYp4+kcsEF5Us8ubCPZ+
IOljq3lkE/jg3tgMNZ8pT1Wd/ItlB0UBYYLQyFsuKnmQXalAQnChutPPvSEYzuOXHON3npcpljPY
oqxv3anyLTRBZ2wMmhhCyozgYztOvskxzehn2xz1EvzMp7Nf4BpBpMrPN7tiAHEeAy1qknZXppQb
Pu3aqRxIxUBRdhwR5SoVQTuvcSCgnfph63vm+TPFmLCBYd5BPR0jekgHZKXeyl+V5dUy2/70iZbN
4q+O+67vk+6H/SYXTeZa6H7Pfv2jT8BRx5KKD8qlQBo/ktOeyRjFqEgv7k/KQ0Ep9DGksTDkaLhn
iAwpLuR0FV11UEiSkq8BLCBFZey1BrpEvI7zlx6royRMW1ln6M7EVSW6b+NiTR/w2agb/aemDWnJ
kf0tO4bGh3TlBWvTXzrJ8D390N+mMJRWYUA9YCN6A9tkADmm+mCugvTc1t323rwpRhjvEnjO/lvB
xvoqucEFh5/eZeK+vxJbCI0PBOl+ubISGYzpnSVrfaVFnHMyQdNMy+L93m7+MzpPSRcM8JD8C5Vm
l8APo6t0CHSnEHQsbBRpb/sYM97VIKQP8NHxpT+7nz84dDZlKs0FLqnBnl6EKzFPdlsMCw2uqIKR
/6ydxj+5S5BPG2uMy4yu6d/y+CvaUl4m2atjpN7yVrTZWaDaU7/zUo1u3J2w6nwy6qjw53/1x2IA
h65VH4ldAZ/Yw6uLY7d+bYui2xTQHveRBLwQJcHV76wTqGD3waKd8cwjuU5ovItPLMIsy4NcTc4j
uUR9o2elFNMd0SMT1Fe9RQZ48ALFFOeb4lEX75TYKLzankmoYLTLzo2bxECsoxPyeeex3GN0G428
BXrobVlb6vjs+nA9kas3lxqq9qm5WnNVmcfrhN2WmhyLxWrgUIxDtCPnfOR2JG6GptnwYnUYvFIl
8w4y1U/GUvQaisvlgG9anE9n3sP65RGcQh0Jg5N8yYaZT7RFqZgUPQ1SrYVhd6kR6Yi8Umoe/u6j
lv5GOALVkUrYSYa8KAq/D7oaiZUyuFySDiGIKIEevVJt+LHIhkU8JVQp81dbqcE5IjA4k6aVeT6M
tL9s+Jao4nHGeUbqeHn0IKrJruUtlG0q9y0DS5pMN/UzwUYtD90NwPvJ4949skle8dcR23e2Phx6
tV10JKnnBuBpLbM7C3pcyn3spAoqOOyvfikPlKhPMxJDpRmQbpCdWQctKoSowlRfvaGnhlCyE9DB
qZTqE5YzM0ZGtq3dBSrJtqrJzXziR8AQe2ZUn/7oDJeRO3p9PrQ81Xitb2vm+AmptGRZv1RDdDLg
J5Dzslvrf6eAK7INL+N0FcJiSZbNaR3Y4d+JpNq3lcKj4zij7uOLgjnvhpiQML1KWBgeGstH7SED
XCbxBcbZ8T1VZfgAdKM3tPKBHAJNXiypFd22OhSoLqOYpdyL8z6xweUDFCKky710WiuqoJoAJ1GD
5g2Wd1u+pDtEf72L0UlfXf8Lj0FSwYFfIS/ncmgXenE29HprE7iuAVi6BE31/IB+Sjh/C9o1D+m/
olS6AJlpNgJ7R+w+Cg0TvfHsIyqt0S2lGVmB0fg8AOQi7xLExtT6B4rj+ayS8xiQR9ktEzGl8Stk
fR2e1puGW/ZcoeeEG/GCQKPQof1o++/E/jId8bAzfunxHUAvsCLjF7uy5PPAVV/ONv7our7XMON+
EOHRubt0h/3zMFWZEcFJSJWyCSxFfkLiQEowUsme8r2GWQQ2O5/QM110LzXDSuIB5+L/EG+xudHG
tSN4WRSQdK5qc46Rurr86o/kXoCqD0AIVg8JqSA9rs6HgBUZ18oqk1AlJsVyLH7CIB2i6Nez2w72
qoUbGpQqChVZQQssNPdh1Vk0Lzd0WIZ7wYFaltk/xNVqMv097b/ebKMcLxC9tPMIreIq85cjx3ZH
Fzq+QurrjoP/h3pKWCU1TDJBrO4lOqqN8GSFZ+IqvNTO2/SnCoTSfly6mdZCwiwmXraP0yz1/W1K
FuOsIb35mnGQjVRWMfN4N1NU+EPMcmfBQKvL1QwoHkrzazodUDsmcXtve11g2MilqANDttGUm9zK
G+AQK2bEkW5YjREr0zLrBrQBGfGa7c944MV+3fcxWCFMiCtOypV+k9ggYY2AFdFQ9NhyfU0R2aRI
D9kSnm1KxA2469qbwIrGWc2qNuKl7WwJsoZFA2qHPZEbB3h0MKV0iSs9K5N5Byfqyvd1XsGFph8D
bmPcBQF6Ffe4mEv8Zn6PgTBHaFgVHQo6f4YFbXbbpoDlW9BQHy4GYXDxscqeounjgktND7xF1QpR
NNidaU2fYR7yM7Y7c86QX7pJMK26u3iA1+HKBCj/cdpr5BVk2Y666SKPKn9DKFF/UO+deczEjrCe
o/jo68YFMV9EdnJiPGI2B5DMtHjoniwlpi9u6xibiPY828TBX+uXO2JbjoAbRrBboUan2H5tpPaW
rZdUaZ63ywCLUg/C9JOh8HCOEp0+EvvsHOU5ETbDnxmO2xDlKdIbH3nwNWvuJNTlL7VXBFvQ1sbl
Kr6/uB2mP/kdRdBX42cH59ieZMonIvBB8USvsk6d0TpVq2NN62AgVVeh6Q5XgVZxsVbW3PJOMKYZ
GX7bFqUPDDSAI6xEQwV7aAyevfEv1xHIcEp5knsQMf7j7fwKEQxnKBBVBaRtOTufn05P0/51V639
0jrVbnRHi6TqSe+btJu4ELjoLfuzLK1Prod3VFaHLCiMGts0hNKeeuF3SUN23jqYYZUX8XJnEVj/
NbmVN6rS5nxMJ6+aJKRvjL7FvfA59KwxxGQxpMgah5ApzNLv6LgQzhGsW8qO8y7M+ZwtrqTqHyIy
rlmK8iT+5SyQvxEpFdEnt1bqkocOF3HMfC0XIBx2rZ8ZyFDSEgl3nE5dXso84CzAzSVkKaXslbdg
gtVLl+vg9PkZSLEk7nTbQQaQ9YJPDfLhbUfEw0dRfZLjBhupYFNTlYtfRr2rK2v+DHIHQzZe2SBf
2mYXGZHBNALAJXrZsS1DeFdirnsRmWkHgd3naiheJ1npU7AA4uYpthcmtv/tZwt+Izs70IPcGsV4
QaIqIHgN10lRuj5ZumIq8qsYbboqrIxgq8+nbYbve6H0goeXZuqqxiHD4+rEU1F5Zi7IEn8/ewVm
hBI7lgFvKPj5a4ICttkOq1oL+HFHKl6K2uGfWrSJbs3jE6UD/6I9QZW+rHPe1NOshu4CM9z1mK2l
cPuVaMtUXf6FlrOd4e0XKHQU+BzeSTGOOKCmxLG4zHu9UFCdcAVlri0EiOYv7AAB4lFRzcQVVXuv
PuhM/7rpJ31gaBB6aREoixT1J55i/eElCp9xpsvwtA6ugSRC9jprHrfmbkS/3vjPaoSuHBSojG3/
Lb0JJHfqlYKLaqzg5fhYj4W4lYTaz8/XSbmFacBEht4Wd906kaC6O3QlcLvnskpxdUB26VcCU6Lh
vIuzjlHz65UG6HnQLWfrQUQPd489/i30iNuHjRmZFW0RirBBP6UzMyOdYReSAz8QFl10Rj7R4zNK
qDqMFil1fabxk1O0OyJDjWhjIBn8ucfwRFsLzAgD9a8nuPSr1PYwLmyEn7AhO2zs6/KZlj55D8ab
lDM0U6I2n625Y4E6RetaH41jJUURcmv9doQGW9QrUtpQR70tqugfv6OcKzc2KjbXElRBy+aKAN8v
4Mv5TpzwazEkNFvUePQ8eNbDrZv5zLefU3hygKmcMdL/XHR1hxlAqjw2yE6bk/IAPvMHD1Insq2n
TCFupxABFa4WxRc9MSCqXilcK7Dmvr4mrl6jRdDhNwncU5363Zu52Q2IwMR1wUGH1SgZ6SQ8yCPm
pqEQ2QKvLEPbYhbCukj1l5kbgjEarFWIYlLBSumTjtPvo6yeAFUh98deBaiYCx50NH/VlEFcqT1G
/yWS0j7GHYFhpAUQSJLZwrdifPi2XeW0w9xGIlSBBnc3WgYDsUJnr9XeK+IABHz0kXhAvWHevi/A
0z/RYJlSU6e8ggwFAoyTn8YBKBIyijS67GZGE7GtZbgKl+R/0FHuHmX/bhc+U4gDjFF5keTSwSdX
Lkaxe0/XCsWssSYCZ4Dl0Fz7MmjnshyVYbhu9HxAX4Fh+XWGGCpkw/xYpYMfmDOxclSxVMG8RWkB
ItlvKmlV4dOu2RrAaD5AnzXLw33EsDRMKssuV1ifbIdds6RZO3NE1vYMu2k8QLHDSBTLkig2Lyjh
bMLhmeh/Ldws54sD1VG9GuF7/Mm/7Dxehzb2ESHZnklpt7jsLA7rjv7zPXmTxuqTdChVb91T3Sfa
BJbOgRynaKg5rsIk9+Yu+dBAZZuhQx6KEE9iu0YpuqToGJ615FrWLHdQLexOrIFtUAWZWTUO6+T1
xAxbfUQYCYz7914Ktk99JhKPO9vn8AdCdZH27ZAHKwz/UnwnJKCHBdBgWqTUtqcC0+MFu16Did9o
sH/6/oShyNiBDeGstJrnVCz1Xw1WcfYsndNXJKe2rsj4C7Q3DiXIInAEL8A6d5EZuB/qvv5AYv5y
PRfmsE9YEC74vxRfNQnCvnWnApVV6s3xFdOq9zmE2tJGlanSqK5lif6ywkM6YtKVmF6NIAaZo5lm
ucwQVPVmY6FMGic+hJiN/Lnha1hzAfQ5AnTSUigRkRA4vD5cF0yT+21GLMDAS7xDN0scKCRZPzq0
LAdxuu+zQepY2Jvvs53kEqs+t9PhYdKR1uRYe+5Lt8fwVg7Q6CLRkjIDKQhW6dE9Gw9pBct2PHab
R9/V0/mFduW7f+rqNc7gENAA3YFFVWuF6WIwiRX5OCT02PwLbDFAVxQ0rv0h9+Ua/j7I86M9MWpb
CP0Ta1D+WwDV3F8DW2PcvSga6GTooSShi3ZtoMIrvppwyolBdtKJVDNRKPjx0w216sntMBhc+RVz
jo+3UK7FvjeCzXYyMA6+WiCNAudt1BUL3BDtdi9H9jtyvsxERfAMbwo6ipMMN8gX19hA3TjT6sa8
UZQjdGX6Ck+vaHvnmx5eoINJi8G9NI/Rd8asSGL2l1dz2jRElTFD65t+CGBST5qhFtXpUtwDXa9x
C84s5lRxqf2PEvQbcc6G8tw8M/gqGwadBnmHzst+tbD/wbxdyXyMY35QPBMxZ90bGP+Qmsbv5iYg
2Q1P7EXSCCNiZ5GRKhx0GiOPT2VA6UGEcWbTaE+5sV3y78D1ncFfvtrv8JVR9k1vI2MhujZ43MzC
gwtuJBR9CxN5sMmciczCmsJuHRCxPMpa8yMPRZwNlHTj2VCVGlwJLHO7Z0vimcZeMk6+hpJd63e+
tYEanmc+bz5kVxo2X1llfn9cGKxpNydROMo6slUT/+aZpOsXerV/F1yOMDno9AQ6vECF+LBPNkgg
aSaJJvHi1PWaywMk7A+taiLTz9R4RfU8skGQdBSpAkezly4BUC5Bm1zpbrFdraBMHqP/g+7sXuEK
OaCnyiTaP5IRWNhE/uCejh+hbEKXKVd0rC05Et3hIydU3E0u6BgDvoLdCwSH1s3H+nFilt0KcDBe
t8s3iznW+YlE2FBJa+wmz/2ZBpJ2qQl5dJ6Uwr1gFpPfCCRGLdS6yTCB2/enci3K0M6UTgfWQvtX
rql3hWNraTCyaFJpIJE/M/6HLlhJa+5m4MIH3HqmQksjnxBKIa8bOqBB+chIjculWoL2ZSUlXPqQ
Xm+w8vrv+aMrVvp1nyelu+XPEmV7wFtAvj5VqCgKDW7he9XBfuZk1CjR84XON+7Cb46JEmswNEC/
EN2QT8hLrARAkOqk7TbHke5MoF8sdd7lJQytGa28Hr7yElVQBHeKGbetWupQ0ChY8ccyCnMEw8lY
5Qh4SqwwVPuLENBGU0FV5rciTJS+jA505ZOdgRCtNtXtNwAjBne1DMMVN9TKWR6rLI0QEPOR7KnZ
DQvT2ozdVizaZVb5NgGUCftMcnk/fTNIiKnXw2LS26I0Pf7DSPhjlk9bH4XfyXrejnl8Do1hYvSM
yl5+0NuVgQZZHDOPbVvdvp0kNiCdFHpVxTjzUMPvZHLQO323Oquf6ypBoNHgZnPJFTz31LS3EcN7
ohD1B72Wo5YefAvkyRsIwOctkVOUFCtzfjqNyNUKzVrw0mPdm2iocnRKbR75t8GTUJNCIYze61e+
PiqbAg7kv9JqmClpQB1uaPu2lAwu7LvX5HFr3tTzs+dDzhsmuOVINZBF4KmHVjeFN76sqegX80O/
IYxfV7BKMIAIzSS4Q0LfcA2kzarJLslekBSt7NYycI0fXWYBep+PZWjIHK0J4cECrW+AS5agZPfr
Os33Vbq7DQqoBnfHJWv2hH4wxlKVvXG9R9RScuKZkncm4pf3xOdt3c+6EDgUDvOXWFcZXsPiUmrq
F2+EVs9W9Ga25lZa4IQkod/clJ3f/9SaTm925Xleph+VZg4Jo6gb50RmuC6Py58V5IcxBiioaCN6
t7z6PzfWPlKleHHF2Zelw/tYpzGgRiqJgNbZde3C85Q59rxB3LdNyoKa/k8JqQTNDusSjg++QkcT
5SRba9bWWZzBTsTYmlPDj8xQH+/B1BvFFCBv0V/K9onBT8SjnIX/bBDAPCSXZNXYHb0WEo2NSAiP
xQLin8TmZS49vC0N52bF4aOJR/zkJ2dKqJkK3SIlYX8mR9EZAeVYWtcvCqUnD4/MU68zJpn6N7un
Uz4WQeGRpls7RqovQzU5VzW3JtKyxziT1EJ2Qg/16/8ejIv5fE7j7sEJFh+UgkCaWnyX3a2StxRd
lpqevJwP9mM+ED8zpcm5Hq63wgmDcebcnApnmyOHrX9iXYDM2kWzOewRbjX3i0NkbJt7i+6/BPl4
/NOic8veC77kzYYPFgVALFmIlFb4B5c5B3IIBxWSCJmR7rSGqT37cWg32hTs3ilHS6fb6lF/orkG
jcDW7ZR7GGMjoj9QiKCbRg3gQa9wefougU5awS9IUTbffzd7qjPBGSUsAUUMuRDalulhIcpb98wT
FKO3ic29oXGOvLRCck5BlebxiCEGUWozxjPNTfvaKNSvUkpGLd8S90XDrclJ1bWZcnRiJydLXgxf
uYLn1OY6sdB/l11VCHG1Vu32gEHHPo1geWIYlvwQfKOM/di6wstdP0DrVzd7boc2ssk4SLvT2kHQ
YA9ppvCYy4yBYwCz+MR8Z86DV/sYu7k9RdirNuQ1HHrvBJdl0DwZq3gJMsvUwJZC3jrPk0u9xHqR
JWVyEr9ApJLGHIOrpIKx+2iOzWaS0qc8MHBB8ihnsi2rH7/vthC+RKny6iWnEPeAkTCZRYN8eQjH
5lw+l+s9DM6caMHTdyLaE7rIM06VCCSAqjU5sn6TEVrWg1ZbV4rEvHds80PPLlMAvJb9h8VEjLhD
NXaP/9o7U43rDDCifMSeq/tnvquxJukDkhx3yT7GcSQfmMtxgXRC0sFpA/eRoQkS+BMYSSr5KL4w
V6axaPcrmDkZlijJXFCi74WbheubRkxS6NB4ClHAX+VWj6zfplB+Qk1Md0Afoag27eMk6lEMOt/n
/zz5HhQPYeOx5PVCjxI8klW7dXn2vnS+Q/mvKz+uksll6SimFycIg7wLOAxPu6RjvvjPHiTN8FY9
Qn4D2VaIXq2Bes5V4XYh7yMprCNlmATieP5x4+GTH+9Zs42aVANVDTiWNyBTSXwBVP1QyRLSTotN
uSFdoOsBpG0fgWIat9N7cyfDGaqoGBzkYGa+GQoupCFcsIqVBV+t5iPpNHk9iOBzKoKo/BD/pSIf
1LnpImDPZ2RVOjRWPOoFXOFb1SRfKK6yA3D9yOfdzoEIsaWX6oYH+ShaY6GdxeeknHsaZ/Ry2Ca+
1dH2a7TodrIl8Dwey12PPJdoDh/Ds5HljKyo6S2iZ6VYtJzqjmsIfiLbQ1XWo0OdbTwFlY/z1Cof
e+0MgeLViMjaAcPVthwnzaQo653XtIWxitvsfmEVZG5CQkl/LeBD7mAUlc007mCTutd1s71eNAvF
1TY6CHif+k6n/BHgNRHph5h9m/2H83uXsO2N0NLbpi0NFG0Mh0OfqVu78rF5OoHC/DLRMIaHBwRb
a8yY2EEDqlpLBBLULEwWwsYzrRV/TQLe1m/ra/rBVMBOvfsquv1nEut8DkbX5x3+Gefsvsb+6/kg
d5cpIQcvXjy6umVQ+ve/NfgNmu4ym+FeCasO9T3t+m0A9TG6YOCVF3R9h8gXbbnAUaeahL9MYGOo
H8Ox/kBH5qq5B3Ot/ehAeoyp0cR9pTrB6ze0fprovFx0Zit5hYt45FwAUfGgq7MUMrRs1gIwxXhm
gskd4vXBHiotQIXSnnHz/5vMYRaZasMvTIsmjkiU9+ou5FTRNU0sS34eSsi//LvUTU4DzrRendJz
yDESbB6fW8vpJcoR02kEjIlKHaSrVS8P+Uo/sP+R69mVAy16r6eRWiNDSsnWYAhzNGnqE1CXKB9p
CBiEKIEk+XU+3cnPjp57hzcF8QzZomFe1o4nu1lIIgZIhfUzQJXth5gHD8ljfPXmzgpyyaIJRmo4
MqLWoc1rrZh1D2dvI5Q4ocnKDk3giwf3ntwjMg+4+88nWJMbyDh/ZlQO+UEdlQzIgQc/47ngbWvv
EAaizGBRhr8xd6BcpbCdEuxWje9grYClfh5T5MoSS4b/AniC/o52qEWkMM9RAepdHObc2+IeGJEI
FymqM5tS1nSdofL00vFtRa4Ja2NW5lej/dpuecnYFdBte/0Fx7SFln+hJXjsLwJKWV4hkxlrs0To
XVsa6YQCNEZ8+bhYDDgNtWkaKaG4hqLF7uf4i6kq1JnX/prpEzPQyfDOO96FPyHytYfwxa/uovn8
IErKLLqumHaI74loXHJkc5Ro/aJ8joh/XujoalNKATEOOX7LSbn7amp+nvZI1Jlk3rK1E2P8oLm8
DsHrxmAuU4oRdmu0ZtYsZoHzmeSO4T92EmyYvfIc0ItOCC2ylV5S+Bxx6tAjzlFy956Wbru5MPut
GI5U3QEap7fUcHtDHRTrRIk8RRZp4t6+F1RFHtx6sCXfXEDzAqpf5xh4w/9qoZsMWgHn8QQl+qC/
y19+DSalP+ui2K3GWGrNhF+GLQL/jMHSsQhlPYGqvG0tNXA5DczEUtvP5jUopf6sdZ+ExVBE3QUT
Vvm0sFGjxQcKNbzB6E8ZQIbEOmXymtVct0YTMXfPt+7LoouqP1VI0FeKhAAhrPxLXTwbXQ5QI1sL
ykC2n64iWBMsXbkeevq4g55GNA4hLivkS/Uaui549H5Y7DljtWLsviUonGN/v20mZBiwoIFHB5Eh
9tlnkrTTSKN/DY7QcQbaMpgUMi+I601/o8n294zKuLCFG65YoF5G/FEclECo7z0vACL1E5wCsIP8
lVXVf9PajmATYDyF7bkAtdgmFxQh5Xsj0pMJB7SzKRFQu3eGIhv8pFDw8adWKYZkDGhjdVmJuVh1
l6i54tY/vzad2oZCiFGbkbeHpjq5V4HBXh1dmEoVSSsTGjqK2KVCwnwpCuaTECzWAlVoPi7eCwz4
MAwHA4RQhrMqtxYDAtftLu5ndvnyubhqfw/nrwJn0PWxpBV1mKGHw5c3Qc7YROVbXPoi9EeYH6lA
yXGvT5Mwrg2QV2UJKETf2jYCApgRePkNR+X+f+/jQyKeKgAhJIbCD701PQrEnIlsvJQdBr1Zx2Zk
031S1EE1griYNkVm4LtUSOzLOJ7DPFJX55deP7TAowPNpjHj+nVdN/3J7CHRRTSd0KIDGrdEYWRB
KOhWaJO26DBlcsrKuLZIaqdAvqTYDUEEq2ZSj5eGTTJqYXy4FvsTGQQhzjruGg94H/PlI9SD7SUb
PMJ13QwPmVq81RD4zZk/YPgLF9horx00tZs15PuSEm2kydsd0jKm8xB6qmXnSWBXEpDXR3jdxknE
XkFpANrye0L2gVU6a5/wORnCkaBMZSi1rs9byXLx0DbxkVg67yIPcby5S/y9UFXAYkc+PdVQNa6z
LhHINGgsPDajoP/MwgiR01NN4QdCLsSIIR1YQadk2O2/YpbNdIHWqR5xRqsoIv3WJTtRu7KIVX3U
x3MKHsrFOw3302+lA5Epc9UEj0sFUvYMbSDd370au3zbNqGfAvVic+R7lvAY3+Lr6/iMzaZIX6Gk
VxJiexdUeJiWusfh2B3zLKiyY3H9olfC2O9JwUJy6bPWUvihXQz9vTpOwxFjMQ4grnPUfMwDsui4
Xo0zdgm0r0oLlFYNjFYF64hb3Wv6CHkBD7a/YXgXyJdfK+EZU5irCNuZr5k7uzvais/ngQ7xQ52u
kZqAb8dhXVoIi802m2Do5IY/OH39Rv0ca64q+45MFrbdbh+D1lvv6BMhuHrXPdQhxeuk1HWOLUXA
ddYmJJMhEJLv8P/O9WC2VLe12zOTuj78970fxAdiTE1s3o9eOzDQld8WkLllfG91fsh4X9gvoLUD
Mnun4cfA6EELEJmrxz3Q+P9FjaZoisMccTeNO2RKmfpnI93DkXLi1mfJh8bzySkh4cDpTkSB2UpM
gJGg9RXQlAOiaB1V59lr0TpHnjiWLlaxP6hJPyCm5tkuzp++qYYDC8MXiJKUNR198SYPEECL1ej7
6gecVb8+NiRfk3cqn0djAxRrvNLcTkdFefoRriDqmUdpPPfQ2CA4aso1hRUXyuBEaDJyn28rz1xB
ruyhTmJDJ1y8+8fxCTD95rBCxqYZwyp2hW4HCRxEJwXJSZ6a7PVoSFXlZ05csP/9ZRa6nYA1qeMA
Rnv20PE6Vog6ajhKy9FEdz4/qWHkqJVLAFdu9rRIIXOAIvdUdPT0/ubTA26pU3qFrsMmxqrIlSC1
DvxWRhgvCsH4A7zs3EEoxW1OtzkpiRGAXoJMYxS7gx0XHjBfSiKxaC4bdeXe+u6BgWyiAeoTQd4v
XKFmgLPMtHl4H2W5sXE4aFRK529Zlpp3d3BNCcJIWsao7eKPC3Hp81hPs8xx+pjHdGJbFg9VXVvM
nxiZQbarWiP2VBFzRNw5YipOPlWQFzqBs62BSohpJcLIylM/MPnXb6YTNkvxFaNo+3LOyoZ0Pgtu
FmYbW6v2RgMAvTt8zuu4ijY+w3K/3TyHPH4+3RLvZHUIgBRBGBPjcPbXXt+GBeTx8k37LyHlsxtc
jAne5Z+QOcPYxM8v2+P1kyhfEkkQ2P5zlHd6O/8E15DuUwIlhQ7ZZUrXTYS8THhYuhpFdXWlpS8i
Gkx74kp9VO6j1uzic+c2EaVb7FknTyD6GXJaA+dZa7OEVFgqZVkWB7joPpUe4SQRE3pY95etv/2a
7jznGqkF4EmmWpvK1xUCBR4HAX87/BpepzcFn178lK2sJ+kUIdwGeq3QzsgXSOfkMRlsXaWxfjok
W+HHW7wSfjdIEq0Nu5gIbDWNgSLbYxj61jJPzA+fodzWyWxdO4fs9bCsRpdLax15greddNmRk9nv
ElFPL1kqU6qhfTTlCxs1hAbYm+cEjRIy4yOPN39UGJt6njkrmQYdpDc/ZECRnfPvLkx3sJhkjU19
9FBAWdq24qBfPAqb0e2mNxQUC8IBw7e9mSKgWzofThnNqEGXFbnZg7aaRhdDNbnyfEZIpd2f3GC1
JHPAuEGOmTgAmoWaSotKgFyP46/DGoPM2dCVZd/JBmQWvPGXPOo5adjPFuACeyIVoHvXj419Zi9P
N6NP9A/G42qQKyS3Eylr/d9hKo5/Y5pUXAZ8sv3kgu929/czl3DeuIJj+/+aU89T0XDMIYXx0XS0
0/qQ/8NNvqlx+wPY6cGtk/EAR1su3ZkGKo2eBCg6w3+IOx4C0wrHKDCdNB6UvfCLhp9kSuYYwEqs
oY+Bkyid33fY8IejDk0M5HnmJVKnMHuOROmNlwkyJ4oeoszL6n8J2PPi74p8IyijXKDqmpKSRUdm
MUz9JTJQNx6y75jn4Ipqq6mASkSxtCp5SeddK0CP4QvbCH6ZRV8l7NMDo+tU88IFARACv9YnrQ19
hRXGbb9a+0iMZd6UkKcfYtMUStAXROupDIHGZg9SWmeSPw6CukAST+ah74Y7HP53dF7ff+9BtfZ8
8wuiO3vytGNqPYf19XO+5QoEUZEhutizYOr1MhWhN2ayse6agLIseCjoIDE7L+p/qW0yQbCyt2cL
E1FrHEGastDAlNrFKjAPb/D+O2o0rOGxqkmarlT/hUVu14IqUSRJLocQpWMHkpatA8XkAUgGj5He
H0khm3X4cRLUNBWnALUu3zmAtZqU6zi8e65mSMvWjsg2gn2St3zjmbyqCe18ucRey1bJBuIqIM/h
wH0u3PtjhRVxaIGWLX4NRX7IrK3HXzeVpYGXwy7h8GnKmRLg4mvCPIYCqmEcFWgZnnwg4bNbkhpJ
1gBryWq2JpEkC4TF0Va6DLNGXz8n7tXwKmlQll2x69FHxMU+Slyd1kE1CXGgSp0cnk5hTJ+LuvbY
UF4cNLLc4ES42q9vfUx2v7YTEsbnPvEAx5cSHrEq51kKE/AuQ22XvAF2zYsAsbbkV1M8Ww8zfLgR
bXF6dEYi+93CyoUjGVcS09f5L0l2a0jdm/O2q9eC/sE6MY19ISxgXpO2SCFuswtL9VJtn1pCuIwl
Z7/IGF0N2aa5A1c9lbOvrHVJWhRxAgjZN7FYOUhOpELQCvPk5aq8LF0CpEGW6lSjbSS+DPtfcv5x
L56U7unDKEFM7BA/z/cnwN068Q/zQNpRRCzJU+hxAccymYTN6qykGqPZgI0mY3ajc9srVbpyT6Hd
oK/UBjaa5rFqj9DTVJ/OlUo2c577Mqd31AbgfVdy2yrKiiEZwxD6KBpbk3b2kkDuaeLvqZYxI02i
D8uTdVandJjmf6fZbBLtsYod4shpmaeSQ5B4Ecp7TBDPBWi+iBUVREc75sebQtgqW1w3sTLow+PT
NmTZxVqKLGNW9v+sdcwLRGhVpK34ELeyaO8we2YoORAiE4BvUvzIDkkeuW0GLc4+IGfacc1VRzlY
wrmIzKpZwAlBJSnyqRH7KVJGTAsbBvWgnBuSkEYu3wQ5RWjPImsuPjAokmq5HFZ6j3NG6ivD70Bs
jpp9wB1pAvd83gUZVByeVPA+u931ir2vGvY9RguU4aEPZzRNacsOiBnrfyr7Kxrvyda3cm8fMwEq
+Aon3YjnRi37uQvo/iqhBhSlf8/tcUGZFWUcmiUCXwwjnWtGoU87YpHisZe+fQyU7iiLI38mLfJz
8FPsC9fbSBYd2PDSHf9RgCGIo5yQgHsHt9Y/wQIdvjvZc7PLvt5Gsm0nNksTFCynanwQE/3J3Udd
iLd9JZaIS7SFetvICsTvAT4JrQPe01IWYhbkev0FoWxgrqxrkCDHL50eBi/fshya0+U3Zb0o/kwt
wcXkh8d8okEzkamoeqFC0469kjVC8TpETL9Icn8t+wY5AX0QTEBNbpU1/qtmDZjPOqTAs8hWWOHn
EZFYkosejf19zXV3CkfCbRdkSE8NsMZZ4nv6TtWh9Fk9TqaqWyEQZg73S8EwxHBJarKdL/i1fafX
fFINTW88SzKyJv4fbWzAY1PkEq8M/5mipJR6BizdWcTs3ASm/XcUdjkbcj3pR+P0j0jRdfYO/0uM
BNuNao1bb6r6SbfE0irN9u3zgGTvk0lgENgx8FV60CXrzZl6hVWVUhpfD72t45m8QkuU4z9TXDSK
nakks7IkBHzbAzkYx4mXdYT2kEhdJ5eU6Y6wxarSDfvbG+aWvtmAq/TGzh5Q8GNB9svbw4PwYFGT
8oS0grcdzYaB93UnRAXCzE1YuZUnxCp69c8GNHMoQUSWjHkCo+W/iu2J5OsW+/fQCSQFLow8moEN
/IbznvddlZhZJALlRgwxUWJgEKi2QFW/YakIBGKq2KUVHrsW0Fia8JtS01utFTArl1knFuZ0VTAQ
PzzoG6goL4HT2TbeZn2tJBE0D5CMbm+bGjL/chFtGds0CZHvtk4txnn2y0mBnjkuJcnHCH7VGOhE
MNtjCvV0cIRrWa7ZV+zbZZHiTyAbo7z4M6Sziism6MnDaHw/Ykvwp7yuss9ZtF0KNkoOCSbGhQbk
DGgiduWsSuffgzhtB9ef316bnuKUVW2sqeoAZ/USovKO/QRfZdhPBcHNMuyALQTl4fox2IiG7eIV
oAJ/Gl54/Zu+rUZcEPd0MFEK0yQ4llEyyM2WwaOwzgQZcGa8m/zAZMy2qzBtm9cTuORmEpF+V48x
yBSDo05Nlq3XV6FYPE3ll4LGB1pIDDlqTV0vVlXVRHmWIiCTfdQoaTOdaNsQdzzKCRbakhvlqqE8
H1Kk0nKxOAcSMxhwSBemYonVTZlEvI1OTfonSdZF6V+ZqwiRUNjJAv6APJCHGjsOSe1RnTjpXGFV
QNWg88w+5UjPRNfPgQcB9GmHQ+b19DR3Onunrm+YBf03on7iL0SBL60md8dhwNGxbcKUrDT9MZKo
NxK9Flg7XDhtPtdsTSZufll5svMv2z1eW5sP3+eXM1pQBwRGb3HmCj1plncTSFn1yIWTWzOfeNNe
gFG22IFYZCjkpYWBS0yaIge6EegGlYen+CdEvdpT5CKK/h8iLgcn9pQodXED+PELNUo1QSIJX9Jr
WcmJgwAXuX82yEddf/4g8O7pCAxLfy2FcppYj69HBfPdT0syPXqyFhZk4uFEF13yLfg1SyoaQwk+
ojdBejfDPq3/X9hEiIMeIofYZFtPWYzWarYVPvu9LybFhCat0z8m2saV0oDn9loqMCN6AbxBSntE
BDl93Aux4R4T8WO/wnae6eGHiy1Elmiaf4UCVr90mZKGZYGSUi/tL7VfGIX6Erx/w2btXgo9bj60
5aF1emNZdZlv4yKYSgFlozEIhoqcz2+2XL9Of9jXJVZJPld5zNtVt9Btd8xJzvvLvsDoK5R9leRd
fr7z8020xW2QTfm4RDEftjo19fgr7+GTCtZmxJJZqzfXgaYqzvSTfDqDHQ0cdFH6KO6Exq9JLksA
M0gy1iNO7UqIModxdJUXFRRTwMX/+zrbAznrKNiuY6TnWcBkJ0Zj+A5o9OfV/JYQwDewyhXT0c4A
hdWEO9veMZJDB7er1tKhsre/pFiftM2fS/vL+kN5TxXKEbCVCmlOO0udtKG6YUuwAOnfuhpUOkpp
OFPKdd9VTEua4bAuF8aBkdAs/WM12/Zv5x4L9ou7J3QKTym5fmFzOlBLw39ZvIy0Oz76qZyJ31rW
SMrsCFIt86osay94p0Lc2eMqwDUYOJSPbSqqdlkd4q2EL6N++xoQB48aoqbxzKEo7a4YX4wjFVcL
IXwcrKyBz4Z5K3LwZeA8Imao8MfIrtbUcWu4jy0f64EXAeRcf2T4d08KZO2RSwBrVQvtv5fgFZWo
sAF7UyjuQRB0f1Y0Ps+1sSAshGPLaqWDHagKY3lcT4sACBaEOAd3C/kcK2z0Wictd0rfNhjhwlde
v9LnH+012jI3OdhLrlgAEIK+gWYLxDvDik5HlVPjYWGfoYldO4yj2TJo8FirJMrTVPB5lQzcKguX
37TAbOIoKj5252euSm2Houh8rbJ/N7nEr0YhUxaE8BVrW+rDYYqse8ISq9DLvzvZxdUDSZZAACtB
1WQA/m8EhLLRS/6rhXMAegfegNOwwP48ddMatFtjBmwc1RIYiHkmmmGEOo/I4WtGxZOxxs3NYitz
d1WRHQUck41KFzVkoOeK6LbvnPn/PON29m682xQaowCYnga1M1FX2PcOQexcv8XavRAGfCuyyRcu
4daGQaa1te1SkB/TdrvSvEZzisRTh9PBNQGJNIhUm2LNNtFNOUuz5T3LrlMvjUONhB023NeG35D+
QKaGMJWEXmL64PwVYVRxzrIZEP4ZuFMtMYCpvSSZm+qh/1MOvOaD5eHL2xm2LAa+fJVG61XslDXl
IY8HB4dZ7q5gmXKm43LzxBFcUPxdys+Twt3xVBAq4rj8QmE++fAunVH6Ey+3vcQJh5VS+1Ep8Urm
iw4aVNpE4HUPuEcsCwvwmlIiNLUFuI5h0rFMXZ/GX+jHMfmGwvdQkZQ4L7YxycffWpaT/Blc+5dd
qZU39WIz3jU0ctHLYl8RIedj2j109Ny2gaTHk8j0GK0itFSiD//rQQ7AJU2meuiB0i/Zy78Q5vp9
4H5I81ky0UIqxLHzKLLIDd2c9clfHEc8bYU3toCM5UyV3NykUuOThXejpkPNTQJZcoxo2bl0XW/d
r413+DT6DbkIGknX2g7RFB7zDW0qYvlMDXdD0ev4RERgk89wk5ZtYcBid0/BvaGujm/TiNhXjEhD
D1bm/tHduDKpUkNcTcPVlub6Shoqd0hFNG09VusJQmxQ9wzbVceunC+c9s15WAO7YQoICvtIaWmL
84b7E/ykv9gTjyOpX9JolUXnbNKs3WypwAAj82AVTyn7y8i5ppkF5iAG6eF2pImrSVRcCwZOkijC
mgYcA9gKkSelhINr65iCXOSw4x2H/2BlVrS/TIxdaGCJ/yXpqjPcHZ0StIDWXvViqoEvPkc6lDKe
BG7MqqpCpM6IcjRZkFTCCFcO4uZUJvx4VvWV3FdAb8qj+01ii3jMn0xF7us8x9cGaA439KhGI1Z1
eI6tMbHp8tOIeDx0kBG6SrKlHmqvj9gr0H0OxXyB4sFA0CnCJeWCGvOkUuRt2BV31vJKYF1t9ckk
2QUDs5P+YFLs7TkjT2JcKy97WhsWd88f/G9J/S9+CnVGohopGOwxVSKSQrc425IAxNnngqgPRynT
N5nT1qAV42226jc35Hb99SP2LQpqIBYkX7Wyz1W+cLtc846QwIwLbeGGfzGJHYQamgeuLqUgHn15
G5WsZBUxPHcD1kRojR9oOpgY7QdkxGkgBHSpXajroszu6U+9iQIGGv/Eo8v3H6GxpwKNwHdoFy7j
D1pkzrWTEdwLR8xrbmcWZ+EsTaM+DbOclK9JuFSoavNS1jlddLPFbNl54CY7n5NGN1Tnkklcrmp+
9oFFjriMykaq78njmourXpHs1hb6FJSQXWYYdRRbPyzOItbhT23D27fEywfJrlRECb9aCQFVgN6J
uV2QZb5t7pMidI+VHZ1ETzk9kBsWY3s9Bj8v65WMwFiI8ItQPJQe71B/y5MNcCkdUbygbzOizeuI
HFtPuNWlVJ0J4PuNKooox0mHqagI1gzKxRzCdoW1QfXIuVhCQ7f0xx/dFMU8hY3lVMsWDZpnjvd+
nppTNTldJFXOs7mUNtpvWOH3BnGSOQZylY4NpRCpCZO+YXvbaoD1KDuCHC6uvuowis+t7cERyZ0c
2ufpGwucmOgcsP0WJkMAcLbN49Ds7LKGfgekecIJZ3H2ceSpheMe7UEG8j+hAf/BPdyHObYhX+iG
1wmlCFryBvh7wVeXB9RBgnPEDl1QVXoBpVQcLIoPdGPW734eWp/CFT3KGEt8k5UOnzs5S1c4D3Uv
mlQV8MACccOgdAf3pK12lRo60QZo/tc0qkOKawjKRIoaB1I5YSliMM8Gy0yt41dsdx8Tn6YVBj6o
T5TXFDuHFErYNISKM9IF5go9yqkjuPYQA+fdyaWAgld1Z9aca6C+olO+x37d30O7BIghj+h1A2oq
yT2bXMlrVYspNt7u160UWT0bk73GvLqRcypRHy+GnBwYXu4if/uhxzg8xMSOv9OGW0kAcH5d2fiT
Njs555oVaGEqYOV6u2oPdlrFzgo8wh2uKZ5qEoyzzXEHuPy+PDtH7/DGQVXTWeD5KVuiWmyiay+1
43ZHOjcFveAcEz0aVoDyLQAclY99jjEfw6brMDuQjRUs64dnPvZNH9oFDAkZktkFp5XwZT94DIOn
riuzg3l/JpPtxEUOI2D/0tOorC9K+maoL/P7O2aoXWhFUFEGvT+LOD8/doIMDbHv0CAg69dNEGM6
oRfCNxt7bX+i4qTYuXi4CCAmeZeT1nLU07UvqdLJ+FjmM/XtdnPQcHTDEoKBiSWL6wpDr5dOql3j
GxAVLtl0Ir5X7XgrpWIe6AGyf0s1vqw4KxqMpWRerFRAxZ/9B3ryVWRcz9tJbrTT5b/Rb3gDN7YB
1/dgZJP3EB94BXIBNjUVCaEfGVfSrIApDIs0EC0WF3g9RocQ2aHP3wKP0dnZRK12InCXb1y93yXd
fzeUGbcOlRmxusJ6m0Y16TTpuzcGHc65kuISiUKhRw0oQx7EIK0n17i+l9FGnc9f6qf2Dwud035W
MAQwkViaBQ81+H2ZRpPM0t0iiHVnC8Xmbh27KP5ijNX7rvqP6WXYrWCOhzNwCbVoUdTxB4zmqnA+
RxgJrPZ8p5ho0h2QydPIVrSjfE3LvcUB7nXU5LhT1zs/iVQx0M3MzlpAI3ROM2+QOTHkaFMO1lpG
hCFbweD0JXnL0Hs3YJ8zSZ9VA3HvOQUQXI7nNhtN/utYDwqHklcgLva0ZRHCFWZHDDuP70M3S/JL
qzSVJJZ4hppOjYtv6dfnoleJYyGlvKwtX3vlZn+R8daFeiUBfWXC4P4JgpGlPnzT0pTpteNj3nkF
+pXiw9YiESokzarwcT1llIySJkokhO2OYAXdGIHshH4WB49MzAd+bQyC1DPjhIxuLy5fVv8ElKzq
Tz6084lEXd5ysfoKMHUJH0XJZD7W81jJlgShNVbEZ0P3iGVlDYrxIa1vITwKAgjlnXiE6KXpdJxH
ShobCNEat49oJ9T9+WlCHMadDcUQn7muognsbeHngZk0cBs3YIBw0If3ld4wWzYv+TKjgtQ1GLnZ
CpE1m2l0IaRb5VWCz/2Dsh2re3aXt3cvKzaP2XooiE5PaZiRIbx0x1FYucQkXDHOhTMz19/U17ZO
mQGJbeH1EUH8F+TS7uvLp/m90Hh9RQPiDeG4VaodHF6rHtEyZzIrk0+zbJnXdq5wFgM6VKVvrh0y
hDrRg6RSh4qxYOZAv0+PJ2FW7ACUxcU0y8llG7aIkCzdwkOnlGlNPLerQRuLdppLz0e1A6xvcGcf
J6r2ts6aN2G3rYeQTo41EBlMjWrNeWjYWVJWvcUFEVpNhb5vupldcXYLzDA9wwcIQXRyLuJpzD7r
HNhHU4XXcmPWcxkmWoaP/KEvr5LHFyjWuWxhCnDXcvUGAO5fsnspLHakyK28W8zx2CRkDL+zWY3U
gwLCRFmyaSCxnT7WgH1puzqBB3e5X1rmvQqZ/Cv8SWOYpr79CwjvHt/yw+SmuylohMZShokz5N/N
OgMI3nQf57YxFKV7lV6OzUxqe+1+PG64lQIZBtGZZgQwmqnAPxO6kIkAfkdypoG60t6MPlYwJn5C
ylXvlyCP8PJntvkh+PdDSAiz+jOm6S8FOaJUKrDpxJaPZA44LRmwXN2VMMmESdQIC+kHPeXVo/CD
0HgwhOrNT3saEfEpfNnXzESL+G2Wv3atAAPoqOD8cy0Sd7Txjg8IsT/IMfxrSNowVOHAajdpQt8K
dogFZcUUgC7VguVvRrexnUPX3OKavZi1ucCTJaXGE1I9GXTSk8W94YnwDUbFrfGu3IgSGIFvm1C3
VLGm+OOqQeFUs0tlo4gMtikhu5SApKWteTwsGEIAkyCNsUyP+Lk047PtrXcxa9rnR/bZVN94FgWS
b5RZPR/VtsNgXkAKS0+g64kdy1AJrKTpAV8Mc5MARl5MHu3+QHCqjxVTWBotdAxNUUXiqqZ/eY3j
UNcJFJa985hxG3208Uol3Nw/D3Qh8jvdBXKOV/TVWiSlQGsju/x3m2Ywt7P6xXbhmO2a3K/wkPAM
ovB6hU4gNasPxWF3qVmapOrUd+V1s+ovxZmIAl3SfsFJsI36PTd33/oEFR2Ran0FEu9xS6rJS+3V
8NhM6cUH4KD9njPpygs7wm1QE/l4rF/Il/2jyk5zcj0I8wfgS2qNEdjFWxRNInerjpuELEmkbjH5
z8K3uRWxoailalCQup6s2Tc42irFSi4rmShXUw9Fpe+VkeDB2nzYMtXqZX1uWOvmlG5/3079rdDy
uLD47FrOtRmOJlvMDyPXloncX+hN60VDDoSWeWwdkdfwuq2rXr00iouNpUfnyWrX6gCDiLlB1SYE
A43YPT4fKyKCuDaJ30A5eQT251NIYEgQCHxZGRzpcfYrQXdapZHvppm0A3xpnprdp4ChjHQgURNa
KtskF3JTIFBw13lPuTB3L3kD4x5CQSetSw71aav0w3IQhxUB0B28Q7nY21qjrbx9ESy8fqzJMPZx
R7dJr/VKgxvWjLADzdx9mo/CAjYWSkrnxJbHtFfpvoiotu7dtqtqpSVBCtVUV6UdcpHLZ5N2lpxk
+UI6bzf2SgzcTr2K7sPx9p8jYaQ8sFN0Hk4oS55sHY28G/v2OJ6/sd1o7wMJvHBAiZ43QPQfCu4E
yEoWNWXco+PUvGljNVpkUxhOb1lcwivSGHhvqn9NiHxLmMKTNkA49sMnjKMZAFN7axjlMvKbf8AJ
iEndyBqfRNjjqeEjKleSspq6Fm6bNWjJPkGJgkUW4vpQmZ6CiwcpKJwikzuP9A0IphagkOSh3han
yUmx2TsaWqe343OyNrkURoFDwPIZlG+L3H8/JE6lWudt8RnVHNjLhs/ufaO201zzfwY8T8beum6f
2m9FLVkkrbW2Sn+C1cLEhpo6T7f62FFQIAHwlfOqUxElILyGF74f7La9A/G9FHQBgl5eaL/9yJxG
bT5S25Sl39knCNYiWTLi5oFHXRHJ96vwSPvAdKFuoV5BaCoZiKjArH4jmlyRO+pbf8cB3WONMdac
ye7nCsVgWkzaD7RXDi71dRcGf72GS9FnkSyOMTXE6M5bg17dskkyyWfwhmi8SMMSyYIWBFOhglZb
HUHCg6+lxQYj1VgeGipQqat/8IpvXLMyyFR32m1alFvsP9FVm7+kWCWqJlf79uWykxOYUbF1m++2
ThKlfxYtsyGfa6jOUOfzQHSuf2KipQvspdHrVuFnOUX0kfzw+zj/vpRl+We4knkxnV2ap/KE1W1a
SBklTcwyKbXyZofaYQG3TUXR8meVjRtDLju4CVwv9y4vP1mkXL0WhXLSeDemLwQ0TNc4UgHGT0U8
jMHiGKWcmaqcCkHYFnqCuVSWN1wyJz3Ig/fPKLIzPMVDzfzXmyVsQAOSoBVVlqQGC4alw3t0HeeN
acRy4GmmDd/ovyu7vB6NHQ0uprRSjTHSiLuh7jSo5QVeX6IwKd78JKwEM+f2FeZzgHM1ynwyvivo
4sm/vq92m07Pkd+uhHKUzq8G5RhF9TwtypDkHrPLbh0h6eQw8fehUNcL9jOtI4Je3rLiKExBG+pL
2m/ltNDt228LPleScs0pA+Z83rHQOWz1uksCQ/zAYEWmfOnWN9NbcXJP+w8Jc6J1k5oEnEichN6k
fMZYaBlDT0umv2voD7AvxmCm4hPhtr2ryyy+RE1hM2IGFuYWebqwrnihDLf51Cr/WHSl/6BjLG6W
o1JfBqkb0SnzAisifFVSSWmTICA+noJIEpiQi8GcNzzIUt8BFK8duFf9ubNDRq2g73V3W49b1uw1
ZLwrvhGxev/BUtZUMvDdbDWf1EjCKEuxoAYnGwEV4g1/YbKFfCtFj+KTl/o/Riqx7J8YnHPzszcD
VyJV/Nahotd3wZq8xFBAW442Qkn5opil6p2VqEPKtdw5juiPDNgc+kcLtRdOmQmuNblNBceco0cz
i4uIZkMeEKGl16em5p8kDqYzGTCeec7Mp5ZrbpUFIFkcqCFiphfFYx9GSZXnxQ1hEpkRr7qLoktG
NoAo613JNIJWNjDOfeF86NmnOCWDWWduYfKZFTC5t3YVEJwKd6vDAiU4ZzCZCtI3RtP+7Ee/xQCk
kJRFtY38mASoFEcIYXfbFNH28pDoPd5jIOCcJcTc4pc7sLqc8+9UZN20sm2eZAXFnvVp6Ot40KFN
rvVYDK9QMziVYQw9H6nlMSnpS9ja+7p1eirtfGBm/jsxi2c+aRvGlnODpQfWSrukBh2fhvV8rEaS
mZcxij1N85LkXJfdyZtFsZ5t6fAv3O9TVl7m059jPAZmK8UiKpeqEF0hGmYxyvZEaZYw42z6xdcc
xnKdoouvg+kaGtzeTf4Ve4YE/eVBUHwYjXl2+CI7CqoavCe37pbI80bQ50qWElrkD8gtrC+uYo0I
Jq1HA33f1FyY13ycrjnG192u8JOJWzfSiGr8pSU8CYj0oMaMkt04HDWldmgjIXjOhAPW+4z12K8k
tQOY7sVf13dT1aCZJ/pEUH1+jZxQ9m9i+TlCV0hSly/0UZwERz/py3sXk/KRFrUPeoskEKlXz64q
TG8aHoQ+KAR35I4s1MHj6TaSUCd9webQzmjDU6l9EdCtwT86+VunK6zdi7vKbjt73LOTmr2QO3Sb
aAGYzQS+7uEMKyq4qIryQpiPwMop0v4LFHKFy/YTAIoBYYQ3Hon747vo0qT/YYdYlBHsLmuJ8w3h
h5ZxvDqy8rjM8xAzJIE064y3yHEmkv1CDSYqC/u79Ma2hnf6Duf94fbXCre2y0ULNL1Y4LrRbkKj
EGLTgFIZ4ltaueD/7GxHnjAvC6Squ/BTrRuI/zBoV8R12Jd6kOcDvFSm3r0Ga5OU1GO18D2Vyn9p
g4pzjQ+Sy00NPBG4I4YtAqGK4sxeIYgbbKSTb+0prgAOB0/eJLGiiMVohOPZB+zXGoJ9jaksK4RO
K8CtXpeFKm0o/RTpk52DJSjY6S0AXsA4cORZ/jvTpWMMdERpwkZrsza3aSKWSu01M2n3S+j65cBK
fkC9tO1cyL2ApHgd7w90OWjq5NreXiaV2l5UunY1aGemo+DDmJnbDEsGBFLc7QOzEeJx+m9BQ7IM
wISaK5DzxTgMyVO7F1hA5MqSBAz8pQB4BLkUn8lS5ckvJwtXYuV2SdGw301fQyoZkTdKMwDk/feW
efbvxzOe6hAGHaqVrtm0m05zTk6iP++lJSFM94Fr7esD9pCkDYkhyZ4vxhHDk9KHdMBo5QRal988
33ibhyDez0UPADqYgNgBYSh+t6ee4GSvVR7LmMbRiuLy6dV+/6JqMONcxVjRSt/TCVZX3vJUcXuM
uZPSYUPeUTqkbEY3rLqA5rvD78nZU9nNu05WNsB1jy5K5cS711IRqIzTMtacM6cwk8lEYi/Yau+Y
xbCnYrhuso4U4Fi00hGR5h2kOyMs7s9Y2tlsAzOqW/H1epRSNnhceKB9MYY3P260ozvPi4MRCqlH
YkyUcfA/9l9pA2EP5GAOdvjlfdRIVoOcG1hPoNu4URufLEc1qLd1tjBwZl85AGpOcetK6ClQeWvP
/H0jk7h57sfEpFJpXb5FEoVZltLas4MOIdwNIXWdehddQ02GY/pwh8GC+yQrrIv8dzf3ak6i1frq
0LSseAdmcnu9heat8JRK9wV1CoQpehFwOd3BChtclcKLYyeG1Di0rBeblg/ECGdmxXyAlcnRY24l
+AtWFxCKlF3bBETTmJt0Fiz4yhoPXj9qUFcWrSbHWdCUNeyQt/6R5PunPUbKYLjx070v4GGaeJR5
fZgKXi/WNuX1rLyOqHW7QXK6of7J90333GJPt7jRR1wryn3ty/7I2XaOz/gyzuMykNcPrtLqCfHo
8HB0lR/qbqfCoUCi4h7ZIfhXHvsjEYvBl9Ddjn6+9WZbo6OJ8giTg/I4yWqVo9g2WzvkfTaMBo6G
SWvIZZBbgB2271kPBM7Qpw+w6VrNvkY0HI3hcPBuBWFws95d0KW8rSvtPrBv4V+eruoejeKcvxOV
f3+J450+ZeK6jAo7xG8/wtBvr6Ivw7OIo8Si7uAAb0y3MYLrGADTMi+lwEFHrZIsJC1z6tVkepNP
0zxf/qKcLlINlvw09cdU9SRVZsMGbr1KPgw20HEKxXHFgKzgYd52KbYyCwA5oXlfrJq68GI556fX
BlCXSrPaIFjt5qEzQmDLE7w9LjM5444AEC86XyO0nHbHKPB9O7iKYS3YiqLBWKzH5lRpmZ+FD6Mi
dwNkkN2eWjIaIjY8lAACIkjDkwXVIdUX4I8DqtJebEecOobtW0VUP0XXmaSiC5cAwCoeCy+ShTPq
dzCJohjRgkwf2+Nt7uz78QiCnZXxa+8K+u7dfEmB9vmuYP0FTYLzb9TzVSMM/K8611LKJc3ZqmMe
q8AW3uoCi5+m80rtcpcu0Pe5j+fGgZsO0i5+A5sM+GslaQJEJF2d3th6bjVbR2w1AiEi7tsc4cOx
ury9aEVmo6+Jy3qyyEunxi2zzmEpC7rCcl8eV7xee3jq3VkNCpEZajbQhP/WJDBQxQJ6xfuUljT5
8xTyOpNz6X3Yxwt+kwq4kzbhZnE6BwnpjPkkpzZjScd/Dt3DOt4LFRlMmOHrrMZOkZhGNKjQ+ksj
ORokH23Y+4Zr/13xI2huAOFyVjOpxUi/l6sMaFVmjAUBKY064Bs+pLM7DXkkgGM6A2TgBnIOw+wy
7UaJKVmHHl/idVghZAt5VJ+diVVYFjCinnVb7kNLfN62PGg3I9sWHCeAqWwvc2QZBEveJ1iQAX59
V/UHqBKAGcN+h5gwI86CBN5jgNeN4aWqk6aWAliUNI3t/kdJgwGJ/Dtyp+4x/XrYCJ0VEVwQ5DaH
b6tH1nVd7o61vfxqggRwM2XLzpWawHwBYvytNKRY4VHxzIjGxDca5zclv4VBW6mUqUJ/TGNKQpJ/
PtjsKyUgqU8mj8Cwu0X4EqxNmHxSw+klD9JxFSbETVmCCbSGvvFCy+mqmWygyNuLbyXZPddSy5u+
vQld0hrhgMdlZT2CW+RX0PtvRkf/nn1DbsdEVe5agtLpP5VTGcTPPT/OstxDbcc0f8uJPFPC+vn5
3jvCU2duavDszpN7hVhfA2NIFop67pR+bqLTpiEN74+6dEONQrGDVS+OUMq+K6s/VjEZOTwt8kyg
4xDmySMyJDdV/J4jMvchL4DuBx+z0eweSP1nVoXC0kUnH4RXLZ+f3w1sxZgNKJuprXFxXFXRxzom
KePlCWHMmGVCh4Mdw804kDUqH4+/MGtFi7t6Y9rgjevNRaVdXYYWnSaqEtsBcsZCU8AMZb1oqXIO
2eCtRSh6T3l/u1JEkLULtkjdKP5l0F39nLMErt9Pttly/4Ns4GhtYHBUJ9KX9jrJiokfT48pXkKQ
i4tFziG9AGNSyaDDlWcdjHpozme31HNuMPoC+RIZ6r9jEYXzESFMbJ8L9dsyDRvPEPQ1DyCYMIkC
gNahD+xKy5SaFZV2ZEJCSVdzdnsy5XO/U1/kgQk9FS0m7RbEPTDmS4Eu9i5aN3HIYYSBXf1+yYNS
0SYgNWJ00F3JleXaqaZk+V74N7Op8SsyEcAao659gWHGqSijx5l78yimCIWzIiyfPk7YFEEx4xbV
7wt8xzvoGxXSknqvNe4H7yVqIwSy09vottCxMnYL2D3D92VAqGtU3gmv8jXrmE1CAZOkby2R6oS3
WL3/kZFOES52tvRT5CEw+bSFY8YAOOV1sf0Y4lR4B/1qUlC5ifbV3dlnVu5niYNsSuy738StIljR
n9D2WNUUVUDZ9yWBhP/umvi6/jewN60WBm8OJhcjMtIv1PqXMt0P0zs7S/XjFroldw5qOIvrPweW
/Cx16rvN3z86Ycr5Tq9taVEjjnAkMKC3/g8MsYyQA7mDwR7RN6gHCB+X3LlZZKv6NHFfJsvBmMNZ
A1512djy2/7iKAOkGrZjbQ187xF+FAZXoEN/5Xaz++6Ppqz/bp+RM85IRip42EEM7jIacFHLyEhm
muEU79Ctt69RLgrUjGpWNThs4CfYwpz2uF60sJqo3o7geiAF5Vd8wh+3u1cvSoXxYb9Y0LZUGMxY
DaZBKpMLLAdi+ERMOzp8ET/rM9C7ax1sTA/gLiHoAqyHrAuwVv6Py0C7Mu7f8QLjzQW/gA+jaBqI
LhRB1zsGbDDwZLD1NwWZk7nP1CjMYFlLznUUnjpwoNBt0qaSuyKI/4Z3qhgR9InvJ9v+FgK0lboE
12J37projGkhZgTzq3eQJwbP4qJAuD8RgUO51JrIvbM6yIiriktE6Fiavd9HpE7tl+h95uolvElW
X+8tJBwLVBH962yKjRjISln/WjF8+vxOhKfsPoZEBFPYAqxfcF+x8MQLSlgzCkDkjNpRQBlnG8d4
D2pfz0i065ovwtDyDgXVXVbzVXWqD9w58V0ZBt7HTbdwHSWsLli7HWGl5m2qqogdAVatcWIWhpKS
Z7a9LPnlMK5fmoykSpL8K/Y2d0fYCGg7I/AgwvFyo8aPFOsCTJyxBQQhGg3GAeHLvNqs0dzR2Fb4
P69GXM1ZyU9LjhmCB+L2YwCb8IMkszpFWMlVy8aUSa0fGl2CZrEvugmJtq/dVU8TX6Xv08S9qNln
J/0yE5xTwVB0A2zLCX2rhndxsx7zH6URz/JTgWyStWKVwNuqeMp8wQs4zHpw1eoN9keo4p7gTYQM
nawUn+iI2bDtUH5zCf8iY/hi5ujbYgLuGOc2bPmt/nOYo5UbXb8PLB7vKOacDRQYu5k98gDdkhWK
fR0qygUemIRpLbdYj9GQmV9wpVCaKcXFlV/r0SdBk0dVSWoty1Ffk1/RSTIJHmaIllPoa3mkYAxm
oz8c12rObYYteXqtrNXfMinc/uP7xh40eFDuHCmaclxExeT8A+o4lOzFF/W3fgzejB+56B30i/0d
VhjlNBotzq7Qpqz3eoYaXXgN1pGxgCAcd3ZAIuDbjdxMfNzbLTuuFufqF0vERKUM5naxzusPQgT4
uZZBtlh///QoMsYSCbNsHchdJ1SQoXQnpah/RLPkYD7kCvNvLg2uav9z8DrN9HJlnDRmZfz1kJlo
Fxh8KDbvm78O/2hTCvwlyq4zGQIWPYSeURCzW9aC/fag3e72ZOBdBGrFR9PqwwxQEyIEK2fxsbc0
e9ViOjDnHnJd6rmNgAeXli0FdaKyy1fKNQ38iePI4Flgj6N2V4yTxvtLjbXJWJwexsaZEgxWtkjs
Zmnxr/VgrT/BUg7hy5stv/FGJL4KcniQZ6EgAlzz/VCOnskayja/2VQ6KtG/Ed0dA+cDbNXDJV3O
ZLPmMyoQjvA1OgXFwrUhuGC+xCyN54+UV/CmOhmbSL/OvmB7vXApQ8d1DXQhb9YxFP3zcoxflFDB
9+bazG8Xg2qBeMR3guzKz+ZbL3aioh/dsc59pN4zIen+m4X0tRmpJ31hRiLFq00eIn4Hz1w5up6O
eR8P5L/Fx2Tfb0+GwDs0d6W/VjnXTJLAbBLfxn+VwfiU9CpDmIt4wX6b0J7tl+uNn9SiySCV1TVq
ElJd9K36EuWjTPjpQ4DMGBcPV05RE/QdZiKXSFzSAwHhlnoeZmnkJKwPyo5WmVIcOgAbGI0cwq9u
8OWof8UILmSG3lm4E5iIW718ahGPTSmGSBrdH6TkmRyG24DY+fOsyjDS7ZI8Jn3F0KliB1A7p4SN
9Uto3t8NKhonGDfK7tHHWXoGSGvNDjFlSgEkpsKPJD7kCoHHURfJuJT89F+61RNg7auroVZNiKUH
2txHZI50PlyLW3ehavaRrDLySJXz7tN4Ty3XWEwfEGnzlt81SPrBtzWuqfY8zVPhUv9SMEa1gjEV
CtJBBQLGN6gCApiJZjFeCWOumIqbdc/SRdHpSNq2uF5/i0n6DoYjS+pnZouacadosiIZrPmGhtmf
mTeKnRebNCGgGfQTWkRQP1ecb7wRUUR2OFQ5RS64hWqEDW6Hbd9BHmTbXR+wTZzr2DNl2HQMwgj3
RhTaSXWN1f2oKEXlMAr7yUuseCIBkwuqCGWnAsFOgN0bASW66MozbNWSyisVKQJiRGJcqaEILD5+
DfRqgMZgNycg6LYh3/XjGSsVxOeQWSh9XCnb8jsmW2JAWzt3Bj4B1qnzSk1iD0UJ5KbXC+lP4lVj
89yCdXtieU76WECjQzGF3xnEBSzSi7SPc4caNFnCA4pn6ZGr+KrE1yThMBIRiACOjgGvxdJSlefP
Hp8bXluuvkSFpaSYfOT0Y0kbuFVqowpVQiGAvZWYMFjQUy11mzHhd6XBTQ5K7qnhWdZDgG5G9MLH
crci20xlDSpZUgLfAjGtJGkkKouSG2e9akfZotm9CVgI+x5EYdAc9WmaUnI6tUgC6bPaXdFyHxCm
SENY//fNiMdjI8iIYLPlidNsPc7bDW/D7lSeCbKggAjhHv7UNTdS/amTflzB3LWhYbm2xl748y/Q
oiecfPaIsPEWi1L092MK/VWctN/ZLGyHkTaBDp7itH5T04EYbRrL2e0YnLNksEyiyYgNa/L4wHEg
iA5hMJWfGvTg/J2YB9ybyl0ratx5EaV71QOJppk7vvXknEBZTMj2GN2BG6wxSAvPSwxq7Ua6v1dd
mFQbb2ksQXmv+d3TD3hh0N/yEAW0BFZbrJ0+HMydBLgGrN7jaZ3BLo3rRT+R1Wvmq2No1xKHH4gT
6PMeOh6O9jUTri+QMAeCW82jvoXlu9kr6Rt0ttIusIZf7qd6T69BagHT3RNBpPi4YUAkp9g2ggFA
3SJ1bzDLyCc4AV8GUNofJTN185O8ag9C5ezQ2IaMxYNaeg2V4Nksh+Av8vdH5bZTbfIx50Ufl6tD
Xh39z8o4tV4d31coBYy9ojgywWTJuwMZM4sAgv96zISQLy9JEmV2+Hnlv5jq2q5pVknU49f2TV4M
7nsPRI5ecBX+sFPcimdrRJz3L6GA9WkPJww7ttXxjGrXKM2YI8ZM010QBjf/z5oXDT9t5rvbJIk9
Bt7z1QoiA1E60XYMeVDElb2sjNv7/QVu1QqoK52MQVd6Mujf75ErBHJQZ+NhRsozoPFBlv+9bzjQ
lekOQT/hafVhe68UIbfIUjo56hoNKfczUazvHQ+GbT8gO7HVGu7RsyscgjZrACQvCwdNgmpo0jKX
DXpYaC0Ep/AROV8zwW3hG7vLAMsvvisOWbx0Gt+xkTUD/NXooe17c7+o2pT38OV3zpK+v28hCtKg
7ZFq+hg9vilA31NYRcrooqWHPF3B3/kpT5qZoeEfhfFKKuOFICjSWRm1XRxtQZ8CmOa7+XSFM9YY
BuKVj7PjjNOScIduTbiq43/aZtPwQ/EhpZLG/nit3cO2hzKSc6Y1a0F6hpXe9BeY4di0JVzLLsx/
dU54EU1LdzJBxTfjDfma5F/fOoPdH5zyxdGB2jFWF/3oOnwxtFZel14DzqbKaH9wvFpWNLrp0DfR
pVPFmmNLQ1Xj5dpubM1dFwPU1APtDgUmdobT6wbEz/M1BWUvve0E3CVUX6pvYbi8oA7nqTAR9V0y
t3glW3VgsZVS3lEpse+K1khkuA/NK1FjWqY5AxeIzyQwnW8eg7T8av+su31Py9schY8I6AqJcppU
JJXvB/02V81uMpBI5Qk/mMpYBjruW+edbbGaFljX8arpaQDEIBq6/3qWGTbZWK7rKCQVZ+c9gcMu
u27oiKzU4wZ+S0GFLPbIXParlK3LSFA7920KGDHpx6Iia+1gA6SmFiTip1VgTyGziJwedn39YRjB
05i5GWlCOJ2xOaNskrAAqhOuSJ8qLW4mGkitS8p/jsJJldZXJYLmiKhpIyCqKr/h/ltPRCYSYLDD
XqYL1hhnwNM48QwJ1H5Y0KnOqgsU/38iGHo59kpE2d5VCJs7jpPtRzvQwadaXBvoFhmZig2LIa32
jmXbqFCLINmZWUPZjpMyB6YF/jRW+Gc7PhkC1ZJACWz1ddM6D6kyEKtrXmxNOz4rEuqgALeB6Ams
xd0TWkxSmkYPFGBB8y+8YVXn3ruNgWrMDbAqAKSr59Wr6MK1PGNlMKhRbDlk6HXJIQfg3KoJ5Vaq
EAWM/rocnS1td0MBfr2RJB8Lf/n8+FSBk2WsYzYwc/C97dedegtIYFxUnDSh39BqlGsWnCZftdMu
04VKcxYn9flFsjZtd81/7JlvgpvwqxMVtYYfdeo+nDVaby1YAnnSY3HomT0n1vXwn0kyDOw4nR2k
YNfsO6VpDPF28c5hAqbbyQv/uXHfHuBst+cu/ULmPFbb0x+Lo5IhI5RjmfKD+wUC9z+TaozW0T7A
SHQUxUBi6S92rM5qd4b1fo14vODiUZ7hBdFRce3X/ED3Kc8yuiWlO+AtYSat0mVZi1/lytPHx+Ha
qI7n1kAzgUMR5APFc3hVuVpYIVo5EVbFzgfN90Kc0Y1XugpYl/cpgDxlFiPCAFYWmPsxThqzZcpA
2KHFJdWodu5jm8F8H6zubZpYUxusdhhLbhf2JHpX405pI6GUPwCC82L6EIAKjH0yODaeaeTJ4YAo
Lqd1I11/+KfVp4V0W+HWhOBkpeVKv2PJBI42y3liBZSPGhvzOjoDwC5j4kjzHmuqiWnIf8FnjmRg
7KmFDRul0YSr5YLgrzhrhQFs+EQsfS+gte/x33l0aulvWADvao167n8RwuPgXEKLiMaDnzSE2mPM
YZ0OdvrGQbt6WAlx/OqeKMPtuwcjnOxqRzn8hB9hpVI1MVwq3EYgtdVtAO1WPxQyFRgZ4jYvAjSk
+fpwyEmINIatbrI/WwHp3CDnZAASfiXDeZMJbFuAk6ZVS1VdwBAuTJdmWg1JifwwVXhit2JjEToY
2Wpgm6KyQZPBvz27wxSbyCO4N8vdWpBJ2H6Awj+6fyf0xrwtbanGUU7gDXi1HIf6MC9nWM88sUmO
LCX4VzKojntRvesnC7mHGBqXhZdEbsNjju/V3OknYluOyVJhRIUni8x/NWiGekfflrwWYvt+LqZU
TV5iJGy5mXzzkWLOG2LM5b5u8TaAZIO2c8iZUGadATthoLpj2BC39DiliyWCKvDYswuhufy8rV5y
LfO03yDnuTPwPj+8UumZi3CatZSz6xsrBbMBU9dxRnNS5YwzyvDbTVzsXaOQltK1RIegy9pZqrVy
7X5U/LcSCzwlg+fZBoyjsRBkG050tJqL9hVsIGBR9xjDK4bMwAfw3Pf5Iy1KF324EHoacHRwCGMV
938iIMMsPAoLNQx20bwh3vSrkC5J6ha6xwG35SCxL1VBtzhfxunKHFDd52fFy+IemwGjmYWlKCHv
OXxHs1XksdNyohSNRNFh+Vsgw2/QebgUowq4Z01lMV60iVOhJX2/WotnGiZhDpz4FppV3fuqQ2YX
X2sbU2I7R1WsjaMIHmFaax7Eqn9dbircIytR3EvxjscdHBhj4ZMCsz5tbHIM8LzTuddZ8AGp0h8X
rwiIpSE5A6xdeUYM3QnNIDWnd7/qZJHlUlTYV+1ESy66JV5cLbdAbyUiNbtnLRV9BmfR22EumKht
okgWpc8ElYXEkTMUORXzMjM5m9MnclDo0ylDb1XTHy8lGR/nStnSXXaJAC2uBwb0ifjt6fx4MgQz
8DC1cTLONiZpuBWlqL1HmltOfSIbEYt85QVCDcrPTZaNbFWQvtMnnf845gCWUfTcDR3tjn49vXFh
u7UGx5YYY/UpMYy7oF60M5hgs8687ebCOMEyEqalzFQlSMpqnTIIxGGx9KCF0ZcC/LDkB0/o25nn
za0ZKnY0jF/Hq8LuolC47MoINZPi4E76GE4azC70k8pCqNFGTRIIJ5rN3Gx2wX3VQEapU6BkF6DT
Sr3l1N9erXUR0HDTBiorW6xkks3T14vf6yaMniMafPA6cJCzJaQ7Kx22f6dPTMKBJCQE0/cZI98E
YT8Sbf9LHqwIYyQm40qPMt8rtZQlA1TTQYJ1uOBwRbNUz6P55grMa3x+MxnawVMg4Eo4EyiWylkM
Qe6B0ik8WjD8f/z4fLXUXm3d7/e9P7KtTfdNRxV5CoY3FOAaI8aC9eCvuGaawsZd8bu86o9iXj8a
nmaQKtK1nI7otmb6w7MFj+pwHNdsZmK6elf09KiOf9UFoyQCRYfErCJl0A7ChQDv76Cvl0RtaBN7
Fn3VlyNL7MTk/g/RcE0Mvs7EolQYj/n8FPOPXSgg6agoTkP5s+3TwfEa7eA1f23F//NMXPx+P+/6
dv9WCX790tu4zbJDthq7HvEpx22RBxlaQBlxgILbyLNWq5tEGRkLwO0jLYz5PlJ6PWb6VlEJObif
bCPF74EdrdWHVEXYIETiEegsiDagF4G5oNV+JLifxc+i/GaFuaIPld6cEqm48bq4tvsuF551zf0u
MQyQHQmWlvEDUHB0CNccIwuGADFHd814LpCqx9/Gc09DXI/ybl+DL1OHJOWS+wEOgu/Klubn+fEj
RFsHgHFhGvqehHPv2eAFvL19mIH0ulzQnlx1sPE1PcWqw5YJeNViuyBjW3qlLWVMkpdOepuGtXW5
GLktGmxQyMJ/0iJeaXOerdi9O5swVqpcXrHOjVPFgRbhYi13Nn2abVkEiUl9UtiCfqKyUN++sPkP
Af6dEsmwyqMxoUirEX43cXDk+ZHAMANAIbJ2umQ8Msm/OPqDkfObwA56VDNBbT22Zq89S2/5Jmqw
cCk1rV1PF4/znyLIWPzBYDngoAYZX63ChYDOV5GHPZodwGzxOVVUyR5qHU8ATAHhvt2SEq5k24A1
dTvPSFEHDkIpaZAa35A1VUymqSzKVNHahEqyVa+0aF3pqgA6tvVc0R6FLqhO6Yy/S5sGQcaJypW3
ZWZoG1XlfO07cgv5TKCNt1dEOmllUIuiKn2kbfGCHaTEfHVyIQCYNiOX6Jc9eD4HjqzOCyFlWfiW
/VOptfUNiqrOyYUzL1iEg3rdQYtoUKcuYhbBB+QztYbWFiR5qMuPfwwT8Ai0lKOtlCRO1V4iltoq
kouN87xvExQNTLSmloblZ90AFg9MOeVyNDHiBpGWMIGIX+t9029LysfDm+/JfmI+12+uFcWNyAl+
1ERS8Yyr3ONc7UpW5QcilGKPpTSsgScQAkqbSQvZMVuxoHwl0C07AIQecl5+XS+f3i9uO1T5PObZ
cPZHnsVzG+HI8OL31lLIYVhSJNh26Mxd4QfJekPPwiG3OEclcFRvolmQ6br0DSEPmTw/zkH8hj8c
Ze8yYBl5KsdDRY0voOcxVIGgS7uuVd1rQXrEHmt3KCdVTHC/p4Fe3WRGIX8sthGrb6cKaeCduuBs
rnn6PbSjrD7XH533a85/SnajNxsCgahyOLe053GDOYLENJrj9iSuiMdmad9xYzx7z2UNjltIfhM2
+7FxvfmgxBvCss5kpQifKMhC44Z1oucNRGLwIWo58wuOktd2lyi/Igd71TF7hcn86yapn2ZWlWlU
l1BacMPEKxWtm8kK8NGOmW4V+Y6ZCXOhSjCNEfv2+8Sy/iXkYu4csv/5/E6rXp9ewu9CvSdZlTdv
TTL+9oBSlkK+SaCV4IeKwoK8bRgnz7IX5ADZ9d9IyT17zSnKSBZlwiL8XhJCTjGcJq+JBVW3yNM5
AmccucyajB1H9sSFtvte3uBlzGnKNPW4mMzavAILaBWu3PoFk1H9QHsrhFP6PlTDe/WQ8Pq/nr/j
g3XlMS1eg+j5zuarDqjPfQIFpxiilIQg1oz+GkE9s/LEmuRtWMHjS9GNcfZmYeuOx872sTizXkOx
ioLSUWlW3mZcKm+kWBja3G+PsxCmTGZbUY+LHioR7uWL52Ml+aTj5QYE9eTwgfWx1TS4gXqj6D8i
V/4J6/WjvH1Ph/9TwDGD2GwEP/WKVUBm3YWj2T/2Jj5ZLR7HUvxWtlT4ZkdnTThAseRIIVmnkX8C
64uu7U1Xq4Fz5O1oQcc/hnurwa41DJb/Sb/r6U4SS3OeyS8s28auR10Oqg+yG4fMYT6qYU447qky
m65oZr2ny8TkrZdZpGNngtMyQTaKvkBWoazaoClwjLvUtcwlnWoPL+PMkFmAp1rqnEVsgzubdYm4
xquO1O4+qbMwW56Gs2sSUkCgQO5HvJqpFhRsiSNpnvwFVfewYrcYovtvkBzr2dqY26sS2m5PbCbR
NgDr8HBalMLkmGH/Xj8iqSHWY0iCupaqiivHXF4wX3I8GhmfVXodG3yvvYG8+nZ1Ml7loK8V7lyf
LQ2NLMBy7bMR0erEAKbCxv/8kyQUzYrEpd2Y+ShCLuzU/jNrTOvwCgMIVKbkBjRGrexLZ5rhh9w0
HKvNeIoMeygA82wZyWqp+Y/CByxEx8Un1WI3ZxD5enDwcH70giwbpYTh7cPbDZOgy3upn7d6DmU5
bkOJKcQQvKi2OCMVa1EJwb5jxWwhT4Al/BrpSEIGnLnRlNFdTIcWGbCqI+DnO3V5avMPPJD8mtzt
Af64PzQ0zYRrjU2sU1/iRcxXqdYyIZVEgF6DDBzlPH+gCHJY3+38Nbn2lAwsY+HsJr/9TLHkCoMo
DM4IkPlldL8b0H1dSt4BIYhNKaCR+0cYnPWXhwSeWGluTAGLD3wCWw7UJWgAyQUMuB9IMJCuj7RO
bBVZBWKptRiG3Qm9iTIfzd0b7itbnUjy3QYqzcNonK4aUmYqKEcsgoEVMTGCdpWqFExQj8jUVIL1
onMSgNNRNpJRohegb1aaZZt1zrlhC33Cel9be2YSuDE4cdMkgNTpS6IWXQtFKzGLMpGKornrLBdn
SO4NcOmjZCLSRALI64YELk0OJTjPw7r3NcKHMdHQ9StZzWQtok7D8kYGqDyBTJK8Jpo9VheUWvoG
0uZW8PIoq2o6txotwTP+zC9oqaBtboDJhQXtn/m+QolMI2sm9k0/Bhjko6ecq1P6sc08CL1GdDxH
0WburbH3fJ3/qri+hqD2QolPJM1WQwu/sAGcqk8OdR/Uy1FubBbh3FoCYBDDzmdip1JzSJOaPkZN
J4VNN8Ti3mGXae8Gj/IgSejD1aZTQ+OmBD2/vPtIsKqocTuJMwOaCt2azmuYJl5365fbea43t+VP
l/Dg2qWb7ntw/InBjkJCxP6KgOKNdDThsFY/JArvXnFUp6Za+ZzFEi+2WrCTAHuCpdQRSsLm+GYN
/P+7cEsfxJYKsLp7jOr/krweeAyKOEGcM3JzSq/ygWoKWASH3x+DgUIGyiKu6cm2WC2NqJZvXxFF
Ay4MqwipCA1dnu/NxIRq4I1+vW1MiaYGgjuE4XOiSihfrzg5RizTzjgadmcJuZW/RDsnhhi5+ueD
AsZ506lOvkbcVMHuNpakSHgNXrv3hBOhatVJy3VkpEH8ztMyW2gtpGAIbkpNwbthFDL5rB5bmSpA
L5dU5jinmISVSyF62ebX/zBqgueyTLAbkT4ge/lc5N7Mr0M/CYbYONrObmAu87oNnjSz1vbKt3oo
Nj/kxl9oAlFv7j1su7+mRuDLaO1DR6wDE6EZZFTfL4ssGEGqOwpUhdF23c1+JtsUazjVwy/QI93t
TlHVvJupYN4Qqb0cGqtcEseSBLL1v/ri8x+VWA0FNM/e27cFmWLLnqkkSwdqPQr4HZliH/6tlERd
KamphyKLgmGWlRND6BcX6RE8SHe9olsw09jCZZSaQQDTR47JjKd5plwzgrCSuKfdogETywJmhP+i
YvnXM9P/UuHY5KoaJ2YpdDJo5qWVVqtoC/amNoiC45BmzUOIxPbTjowQ1pR9lFE1xAgP5LgdhyEN
BGOZXLNDEDA4mgqNbKV7Ecngr8hK18VZ3c4N0LKjJ9ZrLAk9LXF/WFrEPUNbanV0Deo8uO/48pbV
xHuRYRJSy0Gp25xaCF5EbYT1/P2zRjF+pSSHIIGXDZKgejhppZzJuLwW+CEmJuAcdo1P+71tICsH
KsZd0cvd6hAdJ7C8k0gg9Ing5NRUR3AT/UtQ0r87QNLBsnogc7Mrw7q4I+hNlG1np4waZHAnFgNk
+O0g5ewmepgbbsfiPULrEBjmLHqgMThlhTfkvIfVx3DPowY41IEnFQwLklfpBfLUUUCrtfGt8F68
9R2qI/0toVr9FxFljBpj+oAvNh0yeKTdtwSFBg2eR684WMR3HXw8AfftqJC2CJLIVtdoaAy4tUQd
Kj+jOEohYyBkOIKveDtKMwieQ1jC77TOcTuC1R6N1+gsV12z7AoqyGs49nkl3XzzgXjYt/S8IDt7
lp+nvjdRHF7d5IeJ9LijWF4OvDGBKhFwVMYnUZVCj3MbF7TvKCUG2CWvWazDs4joO+mPv2FzDBME
IgPX5rb9uP6WDsBdcjVa3ejD61CA8Jbd4HyFeYVGt19/7yA29u0lZ8wv4Sa8/sKQyob6GTknMrNY
gEVRbLi6WEMadq4b/EPyoSq8xH5Fq84vd3WQ3k3TtjcroIbCqIiEsP5hWEgbimAj2aHd94X66Ai5
WLkcW/71jpVNu7eRWETRheM9H7ZhnfIAKvaATzSSRM3utoDIt7NkOnGxTpXVdY5iJAZZm3YkZgzN
UJH9AaNG1NZV6/bYXsUEnd0m9QN/UZDRa41eVbbVIR5z1F0aGjyQWLYRTEqgF9+0x8iKM8//yDfZ
XYMPxCW8nkHG9HoF9Pxlgl/C42A3zQ5O1Ewe1WttKu6cjRDbP5xTQftiPwuBlqNRXNM1c6E1xFn1
Nnn6hfBG+CxMJDFbCBSbswLI4tjnIHoq5skBglpgHiXfaI4B6ruqBqr8wD0wfspr09nCrchK3bQx
zARermEXlwoXC/ffNzvcHuzuU95k0gPQtKeBn8x3ukAtQG+iYB54xTyFT5nEfEcWxOV/5Xk4G49q
85bEMv3BSdoNNdu0K46qxU9XCSvEKg8wipB8lxrvKnkRPWsbAFNb847CjZ0HIRqKUIFrhn8tBlNm
XCJtYal5iu1Ya34TUagr5zAaXRjNKL8NOeJcdkVuoKBCuwWrJHlGdHhuIOpgqLto+vS2mFjY/MX+
PoPNaYLbfIE7vgWjVW/OHKMPfhrctkwwDfI/0zFzgFr5fYR+kCLpp5220E94ePbL4QgOEFsukVer
YxukmC13UTXpUKu9A3igScvFspjfWwk3Fu0OTIcGbIA+BjfTaNCgbzW+gwbB5mrdzf9AzqH7oJIW
Vh6A3UlzIsXG7BIR2n0S+H2FFrFOwl73L45CCJJy7D6H+x0xOY93Xg/xrUn77ACPKH8EXLp2M6DM
uuGRsHIytzry5+cpHIKcGMfOs2UNSIC1JXBhe+umV5sstBLPMXy6YQs5hx2szHkGdGbuZ0YaPqQP
ew6d9vpFtLDFbAxiPA7jxoxSP5VDuR2QoailUvMj7ii+ygh/H21N0xZkUa9vdbmWOyEPValKflMq
1N+KDD5OHueE+lNpSh5TYUhpi0wH3faHkPQqTmw8axgKFvoyBa+urvw6LbMsQsLC6ZyWRgbVEUbE
xi2OM4sZtrgnKlJKmygqkuLsk3HcOChsuj1auh6Qp7g/VuGZFoO7UMXFgzjK36/vUOD0wP5LxYsD
LPfb2yotitwbm32b5fe6WFCVBAXMhMdPI5gCynRWcN0hsMGXPPPiZVd8fPPh7qHd0ClE9UC9yN75
JYiJB5NtpZt5b5xvEjpl6Vd39cV/0bInb8RFxTwL3V/xp/xsrRjw1D7UWDff5ebdp5/eaJ7Qx0PY
tTgYIkrqjvzG5HFLPnzZpTxafKe+574JQ8yiLlBwEzMBfxast70PJuLYgyBPyaNbrRDFXzeE57KJ
WaK12EEt2I0AN/x2/jlVd4SVd+E7ASWYq3DZ2E0hm7hrP2iP5LgWBpPnAnmRMNAZ5nRsuqlPAwZJ
F2p5ED6NquSGc3Coqzca6jWr64iYnukMA7zhUE4Ra8NLvxWXRtj7EMwJGtSV0zpywAQIzVcjSzYN
ugBvJGI93BLj6kLp9szfjaTWVhl4M20nDu+KjYfdvYqQRgqdoTMZKtRfLKS9oQynYM5fsqhvRBAS
KLdjsk52BGkNwMW+OVJNxJai5dhULv5RY9KgLWDWHKV5jwTmB93TBo4kDtxWioqzuTsji5HG3wLl
Yg826ivRhsIDBHU7vFwdezQQZtqoyv/NlyxFFnHTPlQ4Ax8bVdw7WKBQUlhmZyn0UYrXifT/IlsO
Yv6H44YdiCPq1yoMkdPHFDjScgxvAypvRhkh8oaCaJwcoZZNmjrHHKhCYdLE13RpDdjK4RqP7XlX
mrmyoqra+Xakd/QvZqb2uZz+V9Eogb2EBUAENcttbZbzNednFNGZugXAB8NSyr8w/4txFfz4KDF5
+qPDB99mBoFjmlzrH6lglPOiR2m85sIsBUJ9H7FHR62AeBubi3KhWsxY6PFbsSH/ULzWh+XFL/XO
+TgizGZ0tIqJ1OCBYSLNz1fJLr4qHm86IPOpn3h1OPUs3u6A982IuuQGuXKUp8yPCMMVmOOZVrtL
Gd9PFWDPl5hIQ2tyrFKaWnEiC0rEyegwUYi+rR6nlMIsfqbEC9sliL3f645325dr0MlYPbejBzx8
gNREE1x8MhJt+lUDZ0wf4BJIRaO/1Oy7p8QcV0L2CCIRp8WcPfWX+/w3aAacM+QN0VIms+Ce1Ltz
ACB/8IFT5+3+v4NnxhWDE3poNB8pZ0KxDjwx6mohGBNdBe+uU2QAxLMZDE2JDofTGJSOBTKezfqv
xYHdCmmA4qHSnyGyShO1ytgeT/3C0bqKmLle8MDN6AGi1FqykWsz4FnIehXTDG0cTvyJ+HpqjQBe
yuAKR4zOhadih9Uew+MOXXbjqvNGa0NErNYZTQWJ+OExttsfpAh3fykKSqkl27mr8Zf2cfw8MX2Z
i2d3haXdKR4OMharJV1UEo3MaWntjaE1H6bq+y10AeXMolDn44SH62Wn3mppKSl0rHd9YcduD8L5
/fmyLhFg6i20gfTxv3agmoASD0XiXQqzTuCWWAlWCAu2VRwSz/MqTPw/a+ozRPkd3j8wmGCg825U
aI3e1emkL+L8f7mErh47xCwzzNmATki4+gZ/3GqEpNmvRsEWGb8+6ceX2+wrrVc8Cxw76nYT5KTs
uyNti1SwTE7MRDrBTQCaJ6LcGVn1oEMjl0KhTsqZW6j6ImFoOb0N+O/z7e6awTTWCEGXTTCiCnX6
ksabdXvaVw3NLLepK8YY+n6a/470k601LoTnQYO3MgVmCuXRy7x0kV0SC5RzEVVFqopcfEms0k4l
FHB8K7wem893AmBH/tZAvOb1t698+F0qUpU2r8iB5681FvbovMbHKiIUKIcAmH6oGLdwOSNwr8wx
X/gXu6MZfZdPMnE2ZuKxeE2hljGIJd+lp+v2YrC8spdTgX6wt7j/QcBvyY3gq2OEBImSR41pjsrN
SJBd4wdlotLWf/VofzzbCYgybUiJpSwEVt6asLInjdDY6a+OTnQ/oFWNucYY38RW20g8mqeadwMo
bP1HYXErEqebvTBoRDp1REsvGGB7Sp7Ahhl8WcScWZQJ5ynMy4AwZAWqw5f05OceWI2/CBdZJqzW
M99XssEiV8NbHlAQ3BSQPFdCyWqMdBh5gayQVKv8IIbJdZ6HTUa02IPsP567nXcA/jqIAMmSGP/Z
6ZNjZgZMB+7XrooCiB7WA7GHmYscyWJ58sMD9Jw1hE4qHui9I7ZHzMmWQuKWNvi0aQphhZ23lC8I
rtezwnFF1KUlsDErlH8OnI1UviwIdw+iRLXW5ZJz/DePvRhIZLrZOduqnnJ57N5MJaERUUYbDO7j
scXVAbQSJMtQI5CAep2NiDBRwqkKsWVB+bTwcKZoBxA+tM2RC8ndFGeXQq2rUqaabpGW6WSjZbBW
+5OojVHfC96jWk4VSG2ct9hwytr6OUsvrg/BgVvFkR7KIJztllpYySNGdmLZs2mVzGo6d27jyXy3
gUacSd9jEeMha6eWbKOWloZQgTaFDkHNSlniDBSkuMGvaa7Nt1GSBx1ClGFN9+aQt4oYcOx0EUXl
tgeL0L2kOZk9hmTtaCpGjHU/MGYvmKuBplWJeAgpegVeeZFAC5zEDGSANwddnC9YmtnNbXEnrCpU
eyEUB07cKS/U2oBnpFShZwZLa0mrE7JmvSLQS/5LMnTrMuQM5Y64bpgS+HXoj4cYhn9Zol+VUUH4
37wAQaWX5rF/mZ1Vua4YXaXkf7YExs6y8h3/FgmvuweqWSVQsOB2WjmngO1gqdJL6Q8Q61bWl62g
5r+VrDe/YbEo0hWPPDxveGZk/n1nP0m4byMpnmxOfvdLJC1KMQWCjzH/sRjs5fGCTB9d5jLrdrd/
xaVKluddPbKvH/GWa3+RIYGt5UudQ1nmPifsqz5/m1zruu8uImwxi21RABbuzhKMiHbWLhgr5Psf
566JyJSysjfCs/eTuGXAVBwL1BpzYDfmmRMObJZ6tmM/2TNmh5uwjD0Kh8yrGqBsrJetwA+tZGyD
Yj453oligO5Uh2q7i+Ju030UTWwS5bZlx2QdFbl1l7t9cVYTlZEyPs64Of6OXeuBR0VSys/iEZI+
ITP7H2DPpDdyVktZuDGrTlMAC+IvFqXXBlUtkalpM2qCm2sLzfdHrY8+9CoVjAD1MtMssmW4nItt
qeXzQqzpD1k9e3qctTh8Cs6lbohYjXGi0IP3HHFm94+O7Qr7siWgPZ1LLFMl4F2303nmVXiHdsIA
YDKmimOt0bmoFMTscfTxjV/dm97qPTbLN41i9ek2hIaT8LU8qHxX/Vf3ZoLoL7ogjIboyAiUIMQK
8tvozwv3W7WnYOkG9eQeJNDDTdPt8TGn19ZgF+RfVX+/QT0Ww4pHgfBHY2DM1fJL22VU2Y7m0INw
Ztzsk56bVsrU/YUZIJ4Mw07xwLuH/4iMs+xguraGC7Oftldn1y67ZJzKb6bSt5TeUHFaYPydR33q
c4D+BTe4szp0xM/AqVGV5YLW7pX7jaVDiYVdFNKGeKWr3DSy8mK1xZP8VJiU3ha0wSsHRHmZn4eD
rwpH/yBk79kMa02qfzeIux2rZyY7HdZy0TG4hFbmRsiYBTr+mtx6olZvKqRISNpRy4/dT0reM1tl
bw+jrtK4Cu7iqC8RXoGbzXeUW59zAuIcxcGqHPdL7SzTK91BYYA/KxNXegPileWP7GFs2lVVaLwl
RLMzc2cK1/t9Ztn0na5TPRX4Fuj1A1KesUfV+n0ppNzCu1792bMUu08Aw9wASpuIsLOCVEIKwiKo
FqUr7zgjDGcD3cgtHUUYaECUlyziPkFi3DLDO2lstMUjyTW587b/ymfJBZre/kC4NkKXb57RHCLG
VcqolqBeTb63EntlXK83A31oPYKv7txzPgAQClD/q6TMJRYzULj37a9J2xGtGzFx5U9nurjHb43g
gGj5TaxYFEoGJHQeG3oDbN8xDJJ7CdvJ1WR7hRpFE/Xe0PCGt8lVqWu6r6LsmLMB3rnz7tXZE8Bz
SG7zIEhb7HVSsueMMdZcUnjkBu4zCiW7HLqzfK3X28XLeaeGOKJNNmu1wdVBfjrLPY1a1UOzGCAu
3XxD/F7hxOAEKdGXjBFhh6UVYW61Dw8WsYzyc5q0vonLq4bqZsQtZuSxBRYzlW17AX5m5dtVmoMI
O8u17WCE/tjLVHCFN0scSRMH42sIoEAeIhaMJ26dGRUu170y5w2v69NPBOCYhZx2t0fPTmh1AdY4
f9ZXEj8gO7TeSmXkg7oms4upAF5mDOT7koJb04MVV+CKKGZX2nxx4QQZLE5JrMyQX4kMJ15TWK4m
zlqEsmXLJ8UhOCpShMxDHLzAkuBV8kkHilSl45lSodt/2RoNNEY3xBVGrhVCYFgtF7yhUbOjGHVq
NENUQ/xkug7dftHsTekZhDbRzMx3328t9oEP0+AXq6FGZ1ngS0XO+BxK8N+BPSZTN9Pt+LuVmiGv
qQN6cWsKPLgNsDMUPUsx2c5j8hxukbuJFp8s+FxDIExg5KHAg0lkqizid+vO4+mcevF/aMxa6iuf
1PUGnX6g8pGzWxrJJZw8xfrev4DBWWEYRYKBzt1BBfXTbdB+z60aY+Mus45rVgnq5WUmEfIU6kn/
Q8HYMuXELPs0Nu/eKS5nRPj5gGU16NZRg+EHw4Dq4F1YufCcJLQaYhzvffgRPzW+pR16zQN6v730
OwyIk96jc1pX2cTLU5NF98PE5J8h2U7i1i3faTCe2ayB6xf9rvGnkLbOKkrKZ9Vw65hxA39RcJGI
b8J0861BJUzWJV3IAYj8pbj3Q+73OQy3JXk1MXxprr9CWM3h8gqzmvRvq/KdtKaZKyL/amaf/Hfw
mlnCt7JgVKDRTC9IsgOL75uiK6RvrlpHbDP+RYUvNd9i3V6aw3sMQ6H8aeBXIR+3KQD4/C4oZ0XH
oJTvWm2T+5XFHioVZd4mr2SrInXboisqdl9T2dRTlwtBOOi3ZhP7Bq1oj9GA7jGRzp3vdLAfIvIO
teQZYrxpYV1gZ8WayaJK4T6wR68HCQ43fBAcyohe04e9f8PlXyr0jm5wI9eAtOGu+NDhphTIF5I8
9mtun77ATtAwSZYsZNQQrOmv5BBLKRoSXEaH+Q53zGl0/c8CDM+R1lBbu1hYRp9UmWb4yj4dytlJ
sFfzR4R5u3oBY1WlU+QjJTi0v4PS+j8qrn7bDZvETH5Ih950OCxFhSAABkSN2zIssxGDwJVdmvx7
4xRPTiCkcrH5wjXOefgXoBGuBKm5rYOeyrkb6ML3svXCfWj6+W2scx++y+jNbi9j57Ht7msTEX5v
cgmPXdVBM30bRUAwOVRldtyAwOW/uT/ZXq2MlfLp7CpccgIHjbicuUgV/WqzmSH0/6lZNqgg7H6C
lZudTqiM6OFPFWi2ISHW6iHBMa+BZIuiMbLRc/v5j8G6BJskRnlHD2TMQKskzoC8nx8Nnbe8Qm4K
So8wcrEkTB6iBeZordaZapiLYd8DiJWtFzyghETUuOhiaUlDZM6AFbcYK/d2u4o1sZBc0mC07BGz
Jonse6eNNSS7brN9YV+ibpoNllv9KOzxKEIgDdHzy3iEDYNr80cgND8o2KWfiyRU9U/nYXv7Gd7E
1huL55+5l+cTbueJfuxIj4j78o11NIAmplRL/V/RpIdHHipI3b+k7Wjo5pnKHK17Rz9EW7IzDgF6
kTwhhURGjH1BiFE7SPaGRATVEICuaD/vmq2UKH661c3gBlZYGFgVz4tskX4yJxCx/dEiQdcltYd3
4Nxb4g0VQiNqcYV6UIPr15nUEfX9PuwpQnkAcympAs5raoZwyLGrlr2f2EZPbZ1ef7RMJ8TuGzZ+
pC06noxGtIcikaF+xODXlIxnPIJDgUv3bUJW2e/pR9VIg1IaRL3dgdCfTfyBKCmzUtZQ9hV3Vglb
E6gvLCSRXWbYsy+thqfXg4JoS1GdVjM4E4AIsfbKBKee6jQ5xQTsfVf++vPCw23O8QulJe39cK4U
qz6zqxPd/3SjmxXlSKqiI8RVV3j/zhGESDx/TSF8vize86HJ+IoMPlU3M6uGMwVZFRqzwXVJ5cYu
67O5d8DJ0ZkiJvEEoVOGT08mK8Jd2RlqUXaVu+e1WN5r47M5NHjuZWyB5jOy5Mhlkv1C6hBzpMA/
VDwTAwxZR8zOVzBacN7KAvC567pJ9Tc9psoYBRy+ZU1Ug1AXIRneKBDja6Cb/2plPWFCPzq+FGyn
KKQaMeTGZKGInHg6zeN8lELq+qRNC26/QpLRvnBboqfbn/lPcUKE/cmcuUTnuhuBSQEnQHRWAZav
4xhUn8NOxLx3hAsxT1W4wXOE9YtYM1HCp5/y4p5Tj1YWe35CzKThQhOfsXv12sP6VtoibD4lhJBy
fb4h+71V8rAh8zmgG1KSsLTAw+6elw9BG4haaZ6s1E9FSWnpS2RCvVRqrfSCNXGe1NrOm0ENVoZE
LclqL6mQm/mL0p7wmXgY0qMWj70CUJsAguPAonFMzggT3PD7YDjsvDQAukH69g0he79Adv2c2Vzu
duw0CwMuw4IAYfDbscu8bPkLplxqPB1wvQvMbN/WpFBfNqO4w47HWF5BN3a8V9doQr2rhoVqEDCt
Aa9G8ttr66pe+3cVeStA4L8U30bo7J7L2gJxJJN/91WPgsEQag/BjrJBTx/ZsomvkQl7M33BO4sY
B/j2INTAL70VfTaTPbw4lqlp9PJInGf2Fi6/tn5QLH1SctuaiLQ2AceWiLzKQ7toWLzfFBnlrVzv
4oJ3qxoa1Kub4Xjxq11QoWk6bVFwsIy+BHBd5c30iNd8lzVHhY/IXtxqtpOsxLsPlX80NTSeUwtU
jj2fCY/eyVeM1qDsdT7vtLxG4oCOCUvCw0ngehZ8h6ywe7Jsej3kaCPkEaJ6u9rC/fZX31IRXYjE
7mJy/iKohPryY3UNpa3DLuqjdtsc8oE4wraeM4t4PR1cdwvGfc13dqrTtDOyTsUjEpQ2jrJll/EV
ZfPfuBc/Xp5Kip0PIYxlsJlOr0DoEX7QAmNlbf3/+cNweWiAe7xrcsr1FfGo/O1scHF4fbAczlr6
rS3gIHdxQQlpAMnEEQiJCAQFeRzehwL055xBV5ZbNpjC7JPLhmJueyrv4k0ajhRYzhvqKK8VD9ae
Yvq519d9QSC3LD6Z5y/AfVcV7Ab/QdatxW2MQFChYfZOgN8GTGQM3JKnUh8OXUultOnvMQG7VepG
hUPTTmavj3gdPBLMejoyHbsZmbieqPxwT/JcCuio7uc5I6Tnu0aNxj1OdF21xJKAO2zT1pGVrsMi
DFW9KQOIylhRo/z275ixZepd/i/4Ar/KPsBhGYpyUI/0YUhl0IUlip8buYYhHIWnGr9CVREdCy1s
7MR9VPXQynerkM7KESqU+iO0n+/mTAs+k3ZMDt4qZwdaxK4JZKFOAjE7OgKuS/+iya8DKEv+pvAd
G7lRZk3fYHYNwUA7ztMeSb+F1PIrUNbAbSxWFyDXW+8hl2lMMfc/fOtdaVB32JuaKm3YB4nxsrHu
n6rjzNV2F4GhdSPkpTSC9U/0vHFiby5F7wuxYLUIM0SGBdOXWQ9pODdvO5AQYRP480Uf+uLchF9T
RWe18X1uz7YGhK2MY/WdBqow3RGlnzEBVLw6vYhtMghbm8jPBFG+26eIl1f1trO1oYuGwHTZkC3M
1F4kMoxqAgfJdAo/j7POsrkvjx6m31dU21EdEMqyemUXK5mGthG3kueJfvdKRYxddwlqxEXAFSsM
ZpseGxJNBjNEwloM1izzxFHl5ObWviI8qzQwFU0GUf3TqEXQjnYK2mUkGHC/Rbqsx7eL+35GEaRX
rBGxJdHFk+WiudfxP5/6pbzn3Q0LUocI+8q7EuCi5n+0r29soBg9W+LV5tPMhDSmbd/c+OXQW64X
J4BHzJHYuoC4GWXZHV1xgokmmE1i7+kr0lCKjT/d6cmTozmtBp3NXkUoiurTl0rQX4gi0zG+Q09b
RGfVAG/aZ7A/iw4jyy+xnhT0HZZs3CxpqP5Qn3Xs09m/N/W+lAsquT8R5QvCOCcpPC5qkAKZIMZ/
sgdUzxV1G8CIAjtvqMLvJnZmW7/2HorfHoYMFeEQ+MhfKNQTFbP5gjTjTum6rcCaD7khM3E4rrwR
14sEo1QwC+ufAzHJMHRpQ6vDxZe0cSJ6Oge8aABg3jvnJimC/8rkbayRhhgJqKriv7ZW1irQwnT4
Rij4BGzUtGHVRjCzwI31bO/6+n9/b5zspDtA7gJCjjwnPWzI/4ACyLSy5FutXAH64np63gRii+KG
pscAvyeHIOcm3PMpNvX8Qx53P+QqDHTzuhjIey1OcVsbljm75fJfTxsZaxlt6wHYJXohCFc8rU3O
zS0CgoufUcmVI9R1V3qS+/cKaHA3jiVzj4NJJlCq3E+o0GMrJCZd79tsSvMhdyB34A7O310YO6xO
TMCCjaJv5arqZJSzohAKnbgzpuOQuUECF4VXreqrn/3bT+GKXYbWWHGtchsqlGSezHj9mhR3y/kU
1bDGkVcBQO0QoMwrcKyk25NSuE/aa0lNvN9aIq6DGJzL9w4Ypj3fA+BNZoZKsCwlJt6FvRs10uFf
lkz7bzXYzqMVpMJNDI9nLaOnpoNZddOWbxktdrrSmwUhXUT94E5Ng5ujLq8D2DxOlGVxuNtXx3oN
Y3TS8nnUnoslaT6vbzQ7/FTy96mWVMvJ8qTGRowVLCMg5Rw2ulXHjW+HPFeQ6NGrJjvtppCUlguN
nCdNE8iE4YYAH7vKR1+hZJqDoLPM3O1LSh20eMDa73U/XqrYz0M9kb1ybYxvR0s2L9jLVLGSzjvs
DpculSjJ24AeZRwlRRw/vE/Bo2UwwENoVDUofasTXeITeOSPMQiwKSXhdevhylTzz9RpNMoUh0zH
kAS95G9JtnXh9E7hufEydK01Whwse4ZxJ+kSQXxSzZ4Y2OC7Vq+wP+NKXCkVjPNOog4IoEiT4dL+
yKY0QpY74RbtcfjbF6c0gCVZ21hNi47NcwIYXpljz/6RqKGZW01M7D9iwjybEUbxxYIdrRwyd6SW
/jzLX0bqzxL71TCouaRe/nOvRIszxD+QWo2Z+Pm2NAeTqN5ZApsbg4HtzJOD8ZLysW9xa6jj7IFd
gAIqQA1D3fXjY4JjbWpN4AnDTnjVmj4VTTQARxlpCQ4dPX4dSYUXip4ZPhB+02nmE+7KFibtS7+v
HXqg10IB4V3e1libyrNEmZE93+q48bImEWVFNk/mEbcWpjNu5qfQYTP0a7cDis0vy5eupGe1+EMw
BtWE5xNR9yHIFvqF3YGOOBDtiQmKt+RXPIAmnKtrLy5zHGZkQUz8VWEGImcBusVm4E8lNXOkjoK9
BZY5162jTvRGCBcJGxNgvr2ySud7tN3JW8DgRmblmnuTLAz/mqRK6/PntWoyDwy4NFe6r6wuL5h4
fqZwh4/hzqFePmeWCghZY2UT75C4bzn1DwZuleZays90TS6h/6m4CkKY1aHviLGe+YHBubm1jfyB
B8fcWIM14DVut67VlHFlzfgDYfPEfB1pxUJ4qWG3/i6VbkwkKIjtil9QD1QucsIyMsHg1h72ua7r
8mrp6Pfdhb5yr/5vjBDB6SZzR5I3EGpfJijCbYeU4je3P4fUFETDIV39lRpHUb3o4CS+vN7ckGMi
qHYO1D74+Yfdef1RJcA7TErklD6xYKf+YQiHj3mTGmKqAtkjidhgVBiiGoUxozob0hpgJ7lyXeoW
UAF7xITbZAv37sFhqEPwTyBtFrqmA2fmQtrddP/hDvyVUF4wPFIZFA9HdzrzUypoUBN/bfCWbtB+
IraOU/3saVEtrEvwRbUJPkc2y9MFokelu3/6JK+kfcj2yc8HYYXSeJZZDEskTgai5UzG+2/CIueo
W78D+BWPQa0BE+b+y0idYN11InwbQxn0MC4Ww2+EZCwGiwpHBj6Aza2pYncLEjA32SMwtyUQsHqz
EWmsgpJ/xItQTfq6zzZELaw0Vaxa/v5D1Y4ucIA1xGhgWom4LTSq5xzslvNMpjRgmaogfcLgwuih
R86AEormImkwtziOdI88IadhWbX+tOOnKuEUxEOMsgqqVt1xuL0/9voRx4GCObzJW/qRU9kPe+wZ
qGOucGSzGpjd6JiWR4d1Xm+QD7udZIg9EDIvqN3CEngw0h+cZYpZ0RjjSyOyczmg8NkAzo2v2bQd
JBBCvEokRYzSaeAKviTmav0t+ElUnjPZ0W6UJsiM/c2vuXmW37rRZ2sGyOw1eIfFxNUuknnTYCG5
BSG8oczU3GK7oYgxYRlbrbkiddH453vJ2ONf7jq/+VyHVFhWdhby5TVyu0jgx6r7/cwuwRWtPMfN
lDLXsIuSQzPbMUoUzNBr0PIhRKGqQlPexDW4sdkhHIaqXuOGWoEEvbxXwQ0bjbHmCKkssgfATruB
Eu2V5wE6af7I1KNI0G1IKEtq8wSJszpNazZ6+ay/BXGKtGuzhyUugMCOQcBm8Ux3/z9l3BEFa7Z4
XBa4Dz7ghpxLcUIRoLkGh72uzkPAnFGqctnJHr5GO4bxmTZ76AAGyDgF3lzkqZG6XgoG5A6+bk5R
jjyHPeMs3nXmD9HJCdh1NgwKhKV/op3bh7ajGK334+v598nBeujQU2qo1joutZjPI4/HwnjPfwl8
5RNN9nAwrKQFX7dveUx805TL9Jl7dP+u4VsSn/hUnwRqGKsd7eU9P4bwe3cDSiKvDfhkP0EZFfei
RbU96c2yunHyVd1F/fHp2+vSIvwPQd9+ksx6A1wZgihITsa4mbjQrrJWsc4lPA0djU8/FPoj4soy
HjwAQWSFTsKN25Cxzz3wxfctTYZfm2vJm6vo5B+AwKrwG6qRdFZOF6+vefFJETKV6Zj1JZ8olCGJ
kMCpCRAA266RPGFnv52Iwfch9BZ1Fgnz1htK2k1eUkF28TXwjfqpWtswLWrgdroS0xeExbgr9Xtv
gvb/pOc3ybFlcUtb9I0kXPnWWWvTslIxIT8XYLwqn2rSEqoJG6wKnQwzWuZS5tPEscheiMmx1UKl
w7Ovao7oMN3Y74SOGAAhY+KUoItlubvUnH++C/p95HUG5zR/AXCeDVZVaO73MDibG1bVTWZWHMcT
KTmgKPUpjV1MzajW9JBaQxV5+PTigxDXdKYajpF1fRYZMQ9QO7u453n9gz4s79mZtsfuaXChk6BP
+zo0aYSzRuh1AtXboPJBnaDcOQRLiAwvRkx7Px404bpNA6K+qgWsxMYiBsHl4ic70k/d70HxPDHL
m2C6pv2N8MtKbvEZ8hDquiHrAQEwChd7suOggMYByihowlLkPfJEdwoclnm74hEZmcLAkvlJQ5C4
vi0PWzYQszYvOciD0A/j58/3iT1wevR7nU9XsyJuSltoOQuYUCF+MhwmGpWDCZBd1Pkq3J+Cei++
edZJfWAw0tp2TSKExeICrW2pU8xJowidZfMqYAWxQgNYHrILLSYhZcHzB+ce4F7/mYtorR4yR0Rb
2ULSgoLUg+iVvTf/i9oOT2zDg7RMlIa5AxKIfxpEpLYorvsfWHEISkdZka/WHi9Sr79NrQjGCRrY
KueTDk3MKLJWf92RoBk3KL1ClnFUzHO7Pipf/U4RgMRXp/7NdBOmpwEgBUhvN8wS6V0lzbQB39tv
FbvXllzcjMwB8R+Nw5kV6Zq+Dw1R1znEwD17rDffcs/AQYV1cHjF5+TM1UoRv0Dn/tmekGeDTCDQ
FnddpVdN/jGWebNB7e1vd3klV771owiOtb94TpQiZtFDxF6cfUXL2IwVr5u7SSQ4dCPW4IWgEU+D
yrE10flHYO5geFVy14OukZ3GRFe7wD5MUJH4TaToh66JYKiz83d1XszrKdNiBZuUQWUuekRgOTTn
GIrJoUYW1mHllklyxqk1WKTawUQOMAoqMASvy2CoD62oEfJMxRm4dhGjpF/meAKjoEFn3SfCb7nY
utZKlfJrLP5FhtWAclDgZgseerLvlI5pE9HdSLC2NFlIAw3jLrkSSdzboXyVR+cFixuuPAKLGjwY
F17924TSdkDngJpKiZQC1Af57urunLB+HLs9/Sh/MeWP2fR3nhE8pbo7u55KHlk9z9tokA9j3xs3
1yOGYTmcKfORdb6KXGzvocJ7it9Zb9pQ/EjXVEXwR08kHyi5bF0dYMIhj+CcDLDpGLzcWyGNkpGD
zxEaqqCiywa0o/Ec1u/3QrQmVb5rL5U9J6f3Mh2TwSnp4Tof/CBEEV44wsdqzq0CAw82W/iEB0h6
dU0io+Vk3au+IIt0IUnz4lQ0CkTH0K2XY9s54YVMFYU15qNJzzGJxoHdzZxUiR8c4ShrVPdd75Xf
CpBIsnqwKESaseeVQgyxpnpTdbO9UVj4OXE/i6wlm+RAkvPlUsAO1UlAmWTXWqLtfWi/gokQ8d+e
qheHXfRXGgD0iLkXILsNDrtzR1/pV5yjjz58PZ3H2afNUIE4NaEET6m+0fEVbFugPqTBmAcrSe0c
hdWZA0veFzbZ5wRD262Bb9UOLoaN4r2DHXiHARqciEeThQgndU5r+PYXqjzHW8BQTisTPCqz2+Cq
GQrstUNGpsx5zeCwxvSYbE7esUSJzaWfGsiNQdweEQ4+ldsC5fbCXhW2eYPOGDK/OM91hyAuurOf
TGqi07c+Cknte01+4GhFumHp065+Zk5YW5OY1hMei8ttLQFy2OLmph/DjT6ShvuzltH+3H70DNSG
53GiO6Z2flSWo/gmpKawVmFAX3La3ofgwSoRgQBTEekSOT7gpay4sDh4IVn8F0pKoG8iPHVzfcJG
DbcJZWcfvJInmZgggJi8Q1bsNxSgEYhn9jz5Bkz9hYwRh3Rj7zscDQsQlTb+y7MH8BSSzW65CI7Z
lu3bIgU2wtJ1RaFrbG2bOMHS3DikXASaWYCR4La7vLSkHnGLpZt7bItLhvUTqmip673nQ7N0AnbM
rpQtm+DlEQVCvc/xN2siHNSwDmsf0hYyAQQwY8p4zWYidotpl0zqnxGB1Nx9KJdUPIpvxALqBiig
L/FN2AZiFUu3/LotT6jM1vDlKCjjhPdOoUTavU7ZvfJnmJHc5M+NIqvq3yunLzBhcNcAVi/S6UXA
8YgnKxn4pY990QR/F3xSiOIOGTG43NLbZR+U9AdmyMiaI+EW/TnJeVVkorhJeEOVtMHet2D/CpKq
SsnBWdWU3mJxwORv7lz158ApPxcZUkyEE87zrkUaHueYEUEsRaw8E+gWF7T3QmXNNGV4aZjzvCz+
XzJcEkiZsBGIVZy/5Q/lX34aTgzzwmVnSeoq7Y4y7dvkM8svzqd35zOajMSICagip9QnzmE7f21K
ZCILwmmLoCNokwMR28Xb7tbR1vEr8xeJ/yRfoyUPUAfeu0mgC2bgxudc/ARYdhMWAkRXmoLI3kiW
oJ3wPDeDXGAgA0G6yoSexJKALvV7CXQzC4tEr2wPM0RK6KMF6OwSc0Lx7XSsgshxvB/3/PU90yFM
mH1r3bOfuwhY14YXhyjMZkS91/8XGhvqBhBCynsMAI6/ErPEA0QA7lD3/d40y6/HFZ6aqGUZXWiT
lPsWiM0tP0ER6RGV9QZoqD52ONKZWD+V5lUNfw7Ciq+Qp7AndpsajBvz5jvScGYR1FN/tM9U8Tkh
Azkss1EVDmCeIvh/DTpScj3BV+hPSv6WO3Y9NIAzhTMzoY92BcJVJO3P9RG6e35Ei9tsW14SbDbn
v4EEsqHVi+6W6HERB0QdRYwawA4yTtu6K2aJGcFOnfkMA+BQNWDWmwzQKTHw2UC0A6O8jcz/CPxn
iaI0KfHFAUr29lluG6ioNwZORtwGwT5hOS447cVcdnexNmLouxvhdkUsgj5Ozg+ndJVekWBMu7iF
FLisT2qupDqK5bdNdRtS8gg4Ow4w2s+Qe+j6tUWh6hOYLTxDGfKvLPJla23dSNlRODpEp9zFnfdt
7/BM46/ivDb5oJ84KDwMymG311NwxDI0ZjxPvMOfB9nkiMbJ6gj6/8efsDOvIDlDNEtZrOQIqK/I
ozXXuT2fmFQr0epqIHbSCu/8EnBKjKmfKwpk6+HKE1fap1IIpf60bfJQX55fuAfa2xIWgwieBIso
UQ/GK07WvoFCwDdES6eh2vJByPo6WwPRG1FDMZzeNLZ6c2UAG9R05t2+dfWlpIrlluWXPQKc6/+Z
Bl+xJ8rC/3QF1n6kKx/a+UoICohV/F4r/JkRrv2c2rUIOIJ4RCf8KOy1hEf0t4X5SKwJJMbD0ssc
3xGh8tTSK0NJd3VKaMEax73Wqy5BqOXMr2eiPlYRZ+LL2lLMpWiX0lIe9gubKrrQpuSPQ0Ofsq8N
r6TYF+HVMhpjA1siBTNFVD+OTW8Dnvv3AsPHJC6qojp9D56wafPnCppdjmvh+HG04Sc5JhLrASJ0
mTS3rVLUlz482/Q81qfdJt9RmpN4dMnKBsVSev18NrNHeYue7sZWXKsfzTsvm/DrOYuApojO9XVj
hZ2TRgiGqKkwXEbMQFO+SfVWi2bqc/pQa8miUzrfiASB9BWg1JANoGBFzfNxaYP+WgVrUJTrj3tZ
x7vgCeqyoKRU+kTRXT5i5ceSIVdOZnT6NHy4LQnhfoP6YZLxlnS8f9S7R8zrBT/yRULN1oXSyIk5
/JrzHeWVf9g8FNdQJybNQtNaYNMPyPa5iwVg2yY6auU9jT/6bbCx7b1c/oFL1IvJDRxvXH91hNgj
aJ/J3DxZndmCUjHYnFFBRaHCMIfhDZE/0b1dtAXY9p5TBm2T9tZ3dz2pWMIy8dwBVxp5BtnFmfko
XPYJzSj1uRsyyUKZTIRBODj6Sge2YFUpLEsGwohESuKdji7UYQWZqCaEL+t8jB3J1aorwJf3yrUv
PbMkDHtQPxKar7+cK57C8zENdo89h0RDPJ86cSq0fqXZuoFI7O4smz6Z6hr5r12JGcpQkqRGfFeL
J8Y1qW8ZGperMMLJPP4+XSklvNwXOpGQTSq9nAIvWDU37dpwXPwn2fSY8+f4DNWgjO0dELEpSxSv
j+hZ7dPzcF20QKut/mtlApmvFpxYLE9X7GuK/LtiomKAv3p0ZEwTqAvFVMlWIOpNZibMgjY7S0Rk
u5B4+xEfx5Alg5tRjAWcmDa2/k/Zo3LC2opIVl1WqKzRxMrFfEwHXjNnX0AVMenCV5UbmsWFjctZ
9XzYQn16bzVJXrwiYcxT6+Rc2MHxDElvOOe6fa9gROGUoUs3Top/JtqpB6lDd6A/IHozlzQfydFy
wqTgTeR919/86woYhg92jzKyPkyw/MghKtaVlaRD7xdscwPhuhHdWeMAO9CWvFQa+ZPp7r0rf4Nz
boOd5l4EEhwIhkxU+IJgSbqAzq515xTYr4lA5KwgN9ZxIYH1TwmDHEpQPr/7TYbqEvRbDW3vjmjM
0KBXYZ03fXO5qVad92lGoA+mecOxCE073Uqa8TL24qN7tdQ/s3Ft2H3n58Ul2Rnj/u5DtQaRiVYo
QWYvpE5Fn6PLyyoi4Etwn6b6/VSXEmZGmI9ovhlRLyzeBmXU92MC7ygFCDLqTZ+i7XOGu1tmPXL6
atvQLqY8ry849SNIJA2MVCY1irulcwgeLscAab7BWGvz/TMtrBI5FNH8h8R68x9CiJCyumb4bRyb
1qmZwEDvbxa1C5ZN1hv6/wBBsHxJZ77vYMjelwO1FzWY3+K95L8hK40sgRKT5wp/grhI+X8w7K1k
TzPmLGEvJdJjbWjl7/jn7Qs7IEcxoGeFmk11rdgtoMFZZ0TsUlCgJZjkKOHL+rE6FK4uvaM8Wo/4
lzjXCo7nINEpnZYPjINB11fKbvWV0HbJN0vdG/z5eqZywIk05ZnNKKa6S7qdH+NLOGxZhT80sosh
oweGJRUU2V6p1EM2OIelftwKWHmDPWs9/fv412+nTSrfA3WXmIBwgGVmjkifJQ3zVUFbp9clY2xv
eDGi7bXrHrNfL36IlIgy8jC77T0bUCK45AeGAwLBS3cfJLV0E00BUa/LpE5WjNKYLzvW8fecSqxc
UoVgJMD6xNir9LHfYCEshS2Quhs8Ga3vzRsSPUNQNq48CowSL7W3im62iMbJu+avRowiFb2dzZef
+Xj788JE5JJDmmG0JL3goBIcU3ygFtSj8Sx+TFEP94TFL4J7kXYFmVL4zMenXSsKamRu4ur3CGPh
lBjfEwIhR0R+x7jFMXn942rGZYDPTEdtSehxKnqqozjKwq8G7qvqBnH+jNkZel4ndFMLUFGamb5Z
aQ4E+eVVglZ2yZWR8iOnpjxREwFSWMjhJirFzUus6QlSr8xZdksOGWHSNllbsXdKxklc8ijjKMy+
fIdaG450adHnOwjGXaRRdIqkBSsWxC9ii7HUqs68Di+PQGaDzzMHs2Hd5fE8APpWeMsh+sjKCXXW
z4gP6+ZtUj6M/IcDruhtEAiM9mwfa9nj6N6AyNTVSnyjsMvGbsbbPZUdmtlm8xPGs9cbecsP6osi
p5dRNSq13jCfYVJN+4JcIBevHlYDwGgCorkmmLQ/rES9TOegN4Q+Uifhzua8myV7kWiPc0dUNgkY
cA7Q78hTopQ16nqZIxRsbaovhx1NMUjVpGXpMCkI0Og+Jp1HiTKgstZ2lOQki8i/BaL71smJdw7g
6hdj/JEq/u3o0ebkoO2+zHwlkkTRfZpCPq0LK6n2/eca+DKSgu/BzVRhJicXVAeqNbPxqNNvfw4X
VSfIsWoKd8ZZEWJzS0FAWbR9uZFv0zyplWSXYclQc0MMU/RxAvoI5xjoi4AwxnqyBaAF1JLsbRu9
p5KahsxiUdfwFh+SZgIkMjoQZLepb7RaWJG8fwYTEzslA74IH7Kd62L5sIcEEgmKPlZJ1y210OyZ
QmUFHbUU0CCT/7j0Qg5gk11oCJq8l1DQZuwF8rXrxQQH20Qz20SjzEuVBZzVJcOnvoYqblvsc97i
lR42Jk/G7mLMF0bohqdwZuGH6VqePtE5vn5mZULkmzqZcdI1DB7F5iArL/Qeia1qg+Dej0Kllp65
4GutTuFOjRehZLGWX1paXR6E28/8E2VIJ1erAbgsj5PvOp0A4R7bEp1YVzHbCDPJmZOfL/D7oMfS
WWhRAkPgW2G/JjUUzKJgETjluZjAZVQhkGhPpMgO2Ktw7jDn/5Q9ZlAW8WaAxKfWYs4BJjqrOpDs
JbukozaFTK0tzuR8K7c6hdjpv3G635F5BW6WGRWGg2OYH4dseFzJL1c7hQxr0Ox3CsHPKEyluVLi
MOijgz/V54i8a/5oBxrT5L8UFprLLz+Ny0KCwIjNdTfLu/WMCk6wsxnGPZYZ/HCGAevPb9hDV6TN
zIM1VFsUfH9sykRSr2XBk7gLhkrw1LkltD9sr6KyaF+J5tqMFWV07fziXIPOiIxkJRIJb2HqAh3n
1jXneDVjhpTvpIokz96NAtcOxqtzJgxAQkjqph6mzHNpQsyyWW4XsC/YfDh1XjgRKscnkZ++D5MJ
rEsUFxvvOTGuLfH+cd7+wZih5mjaLn56maW8roJzxFuDvJsmKumPBoxRfEHdYZJ/NewCF7A9Dqc7
iOrJj/6nCu/9vNNdpGpq2u0D2uSfJ9lFo/sdtbrPdMnH5vBPZQkqHqefWXjS/wdHT3mF74SiUkxj
WEsE2uoL4tctDOtvLgm2qQ7WAPbiPPYq66uYQVoen3eoSOVPTKwcX/fnRMXvZ47mY6KAyTS4fGID
CcVcSKshWZdllLQ9Yr7BxermO5C1/reIkwtcTUR+kLq8FOrvpQkyLAW87aKKtQKWG00wYwjNjeNj
1V1nuV+XD91NO7VOknY5a0nuhF7L7q7waUx2NB9+Hv6/V9sA4O5NRskEk6Foo5LnDbIb4sic61u4
IydRkhCC4eeLHk600e9oRI+m5IdUF02KBk+je2sYkCmDrLot3wcD90jZcUPhDwcrokw0DQ2SRpPB
mv39gqCFlCfLdUH+QmYrrWKz6Vy1I4vzz0uVa8rMB4o1KWaEYGJG3qgCa2yorymrFQeavt5wASjK
onHbZ22sFnsEiSwhNxnnMUmNHzkR/Zstq2ioMvXSHsjT6aB/O6q1D+pfQkUZVjQirWAZ+D8y7eSO
vTqrzuJZBuhPlD5Z7dBBEdOGm4pIkxMGBXPquZYxrgRpKqOqGcv6JFPLaIJugqY7uc3cDCJvQ+mw
RwgxlwQ3DucGxAFGEP1R11DzpHP3e7wWpn5ka4XMyQ6LiWNDMW5in4g5wbwhbQvRLLRckDZ6nJm8
NtnPI2myVG93c2Gu0eB+wDMkTH8qAUqQbmLmNuvDtIrlukQO8sNbuFaO1XoSWar4DTFIfLRPb0XN
ua2TyWIT0UdvhYcIU96qx5Y2FuFqh1yC8LEm+d5DYOKkm0ukiAKJOq+b9FHplVrQsjxjQ0rhfFSw
QH2LB6U5CBV58U34vcPUEZuwIXWuH0cW3EVYnTYmtijJ8xfKpzewflxqj67a0Gn02DT+mk/FAHks
WDuog6AT2Qp+zL6JUNQwPJp80sWhC4Cj9gvQRQ3lIJJd0Sx7WNPGW3gZuHejxP3uCKMbs+1KcCEm
jrZ/a0pPGhTKcdgO0xNEAk0h4vrMpyIku60xwFJ9MGQX7s1nifNS/KUQ5DpeyLPL4NIdsJdpVO7M
/8AjgNWDEp5cD9gwb14W4670pYbrqv23q8OgnZ1zJZTIZX+D6I64ZL8dmAm+r6XhVN5GinQwUQ/a
7puRDdMCQoXajZzA7IKTwImhJUt60zKHCKw6B7Ptrf5pHVDx0qm+ZMlkf4TDs87ZZSqBf1zVh4Os
KC8oeEXM1W9V+cz4KquRxy1nCiTQ+MbFk05k9VgRwvoStEEN01tp4wfdl817FN/qYwzLjQX1JMbV
BdBICyUjAmEjIZHZhA0ZIbLctoGAkH4zMJLjkdQR4ypF5glyPhcIgKgf4B+fASDilClvOs9L023w
lf2D+llwnkUiSjUhJ6g+MjlkYypThU2yuPeAZ2Cma+TIFmTI+ResJfhbheoL+qo7L1Wol80DVRm2
4cJtXVbOYhXnyYM/okhsRkUTTNH159YFSbPiqiiltLOvgYPjNG1Xg+r4pmAnOBzcmI7T8mWYbmir
ab1Fw2qAOMEzilnk7RjqZqAuhXaSu8c192eFkf5FwW0M4kqzOBkapUnIfakcjUSclioXrHY9GLjQ
AxHoL7rW4Az81T/mTEbiRAx0Szsy3Fgzx3/XI2+ELtKGxmGtSW7Xd5Dlrv5qHWSj0rz1hhRjbY1k
yA2tH3qlxZgZjLzS/Et5cv2tzZUo/H+lg+u1UjCfLVooTvYnhFOqEWQALxBYArbhB4MkrgqbC4fp
SucPvS/Otiqacr20+23hKDtKhCwkJzwZflbNQWBdnjPJKJOVPoVLb0NRyzdeUAD5z84KQWHP5bTo
BKFksFlA7ODVNkdXYyVhD5o35e7xYiNTbPFEXu9h7JrfAOKCM2Jki/wS37G887lwmX8gsOTFTGSN
fGEjaZIqXA6RMowuks/icjNIY2iPwwnBfg/5HBerJRMoZ6LgfF3371D26wY5Fy1EtPSsSk1xMrQE
JFYHVl7CJ35/E1VBuogWtDdlyDZsCViz9BRhpDbipfsN2KwohRR6SskZXkUkOOpUfWGr4Bj6KNB1
qlJXnUqgd3ZZ57OhvcbOLPMEUtVOC+yKO9a4W8qd4+u7ki0FYdsDTu2vBJ8RqAyk+nTtkAHU3/pU
/oJVjrKwZ9PNE2+DgTrfpdOOtpLnmzZYxiuurFKHR3anRfJIhapzURSa2OnkUJmbvZQyBuwkaA5H
k1xdd5Un3vm2o2+1kmsVXM3YgI3VsYP8psqMEG6R+2O2HNx5hIbOx9GV1FbC3kxvhL5HbBRavuXY
nZWsqFu1GybyxJ4q7SrZJuyj/8Ieo7B+7axej7EzKtcyTntsuWlFQorGmrvV1znzujIIXRp+WLd6
begTi1NVWd3PUlhU3Gc4zPbhaxwVZ5ZnvtlkAPwxkkNehDSyneb8qQlNGRpksUxtU9XHslnqD8Xw
RWNc6RJxLJIl6aWmlY66+PP5TCA2oCTfJ1G5Df9vnlleGonH6EhaHJO6GBbCxz89xONIsB9Wm4Mt
yYpnyumoWWFG4qBh1PSy+vmHQT8JUYe7307vYDfCp9w24Tb2WBrWZB0cot42JegD+dnER7YpMxGC
ZVM8ix4Z/HgiqAqAd/7GfVzxORbC5U4Bd8zcVGr9aFH901CrELfh0lMPkM7JK+WZRBfK8eZm7R4o
Wk8JZdlODn9GhVO9adhfYJ3wW8TdnZQE1p92HBGNGV6OgsHisZxZbAoe7oCoCPwVQuVGNd8IVlxn
w/KpDuo747ONC7gZTGQrvhdGeD2cgNHfzoF9EpmSpe43tBTI0+oxWKO5z2UJ12s4dLBNrx0ElE8V
Xwilh4bZYbr6xTKmUsgLuD59s6n/yUQAup6PrDhFL5xBuiC+fXmuoPm5eqezBWHfR4+rXOhZJlSx
b7Sz+zLZhWOpY4T6HcyRbZblCOh6QJOU4gTtCw7+Zdj6Mcfkx2rqI6RNjf4e81FowoEjNbhn3Ici
ordz69QRPVj0jcqw6xIEbITvTOBKW4PtLkn5vl4v3Lu2qSZymwA2k5Jiq7itPu3QmXsFt6zjstjX
HgI9niWXhrBO+mut7anhFyHIcQ1+Cw9AjDaMlVt0jLpBo0gJ3dKbPCftyr8zeClrGZyg5xihP4Lg
Fp+sbarLl/AfziV2arzX+STNNOkHmPVUOJjE5Y/awVzezQLTjWJ07LpAi/B089k5MqZj+mdpFGsH
+p38KNAKTJL7tZXmDFQPw4nBME2vXI5y0ixkXJuJBtV2rNd1O1f+74d36Re8GHGQCcEGaznhMoXM
FqOe8nzz83zZo8wlVLfOX85aSmTX5t3O46RurpTC+iMQb1dPWPqSZ1uIs+G5YWsrfapxYgAsvUxm
pypLQEERkEk4Lr82BNjh2KHmxvK4nCP0VP9bnY5xy5+GCUsa80q9U6i9beULb5lJo31DHfUB9q3G
qxfxQoQ0XJbEJ4zmubstokW1Th8lA8aVeLpwIjVAHpRsm04XBLAgGXVf593acsE/fhmt2eRZwyxH
ASYJkAiWw9x1viwrhJomI0vtDD/akfpEI8NEa8juTdwnzHrlNAk6tIWCyNRj6XNBHb141UTgI9BM
oKjfJ1McTJZ2Ie2P2Lw4MYdegZ/6ZJwj8OPSS+MwLbYHc3fiEsyV7KdA84zG3VyAESMKtWBeco5w
DbAArXDLnTyyrAZc4lTMbMVbI6yrsOh3G75ZtwWOm16VokYkRp5fQNYKf+C4pJIFKPprxMx7PY3z
J9INt21Ipl8fFopaQ6L5wWqOF2DMNKmgmaiitsYC+wNxzGEHmEcyu73mj4N1aE+h6xlf0QlhqpVF
BlL4tya9PpfrPZJlDph7N8nRZ5hdytlVpwQXhsigxAKV4AAWGtHQmIaMuufmyg+os1Tk0+lCcOtN
N+twDfWdJ1mjGmBrwN8e8x9Fi4JVSDMUPMif3QmTCWeVld1NvSuV/CS5dneen0Rio7E29OpORi26
Qv91T15uBdv/vJI6TB2XdpX2kD/EY3kYO2OhcN2pM04iSAamsT+ldZczuWef6pLj+9I/z4z/PR0q
xt0kiBMA6fOx1DaMJ96ES3RKd4g5KzHnrSOXlnd0MUeixoe3XVHeSEyP34+U2QMWmnTRgJNqkJho
0wBrZHOjMfKDAyPOxiM/NxLvF4kVls2BLSRTPGXx/pef3dDun11rfD5lz7NEDgKQPEH83uQx1sja
vIiY4XMxOQFuqW8nGOnfloEgErGRreB++x1gxp5vUBR0tIfE4PUUDfu7s3jE2uzGa2TIXfW3eRI0
GkoZ8hbKZSG7gSo9RgGrjqJL+LwIOJrVOnvQh/wQIq8Mh/YkNneM/au6+Vgz+MMfCwp69N0qEXEJ
2T6RXUQMZeWvzGp0WAlLv1XqWuVsr0C1L4o2UcqK/+a2jLDSi+7mBQHIv8pxJ+7IcEe5Mf37/vjg
fePejyAof1R+RsDhiQ8jbBqJ2IB4F+h62INjvQEgkjmhOZ+rbXCoRFzrQrhmN+2cTLqTO/NesZjL
UwIYkcOQlMnV+dDb+yPhHoDv3ffWOJoXO6MDaHe7QHoSdpfHaLgGIVQyMSBLyUdn0rNOS8LQ6rbo
l/TKvll/INBpFsOKinLu6eeTBz94C1bBuBRckuTy0it4izxX9qsdlG5SND2MjIyJhkSzhYML81Ye
6uHB1wQwuAEMJk2RYOJP4SZ6U6uF4wVvjMdGm37ScRg8J3B2eeo64Jm2hpmF+dfg5ql9HaFjGwii
x9HPTDoeqgLzAtI2chHM/E6MBC8sy2LRxGkfHrMiqBQbnpUlpgk2aowkWqwnwkyasN8ZF+vVaYv/
sQIr1fLdbb5eHln7fIU6Xoun9f5wZ072A9qEqGD+oRsAvtoSkgAcfL9tf4TtXXSDMPh2H+Bdn20C
JQlT1Hl2uyDZ4y6a6SRpwVh5RIffMpdGfiN17dmVpSd5tr5jVVGqCzZ3NecLmC0rQGGcN02w9fA8
LPh1KCQr0fCey5DsqTZiP3Gnhwnq9ftmO/5JYfrbi0eFvgH+RzCTR0zPwlP042Yn1qnbp2VxA+3C
7A/pdWLZM0HFiIzMemN6TmyusrghCj2Jt8VPQ0fZkYuBAhxduT0hTe59OmZpBvR6Z2pQs1CtghcV
N4wl8EvP/k9xQz8OCl1K3+g45wNYeSPUCwuyK1TdugkiRoOOhisAuYQyTOI6rFFlMN6ekJPHCFyE
hOhOcxbrVI0OqUEWBhUT70EmIb40EXwG7MSQNLUUZmkdLqgaQ5M6b/hYSPBSCteCWSpfCV786ge3
8snE0cvDZtDnf6Rp6N4HMV7ApoCOLiTOETGVcnpNIqU+4lALHZnDYS8UtnyjYPBIlmTqpxOO/XBc
VKF6hYkc+MXCMEXENIT2IgZMOkznIYmJHNCh4TGbjt8AyNskdccZGQgcXnbtG+I13UULBWmZmfTT
HzxMpsqpq9Fm1eFg2/RHh3F3ZEgnb6U5vEB4o/YTa0+lfJafYZfYrJtsgcfk+356bMd9lUwrlz8Z
8Kg/hOgsL07N9oIfo9bnlQBDmXMu1q+txa+dtlp/9+7B+HEyhno5BBAomVID6i5LAbmydQX5GVZx
YBs4lWJfMvLQ+oVrTH3U1RVOzqdDkwvHDFtCkp6P+Hq5TgwMHgnET3+BRxoQ8ueS1kZJIdIUAd1H
TggtPj4yYCC3X93LYrD++x0rlv6yXzVBaY3oK2YS9OyqCd122rCPULNtgTEjvtErZ7fTN+kEq6z6
AGiVcR22LIOV+V1Nf54mFsQW5zlrdomjxVERkrYKNkpCHbmHdyM5hRoIuYz335KSbI/IX0RruTTC
nBqvQ8F0KkFZfGEsgiVC2M62Dc8eEmaz9784j4uDUkNELUWLOm45G9ClAAqYMfGnEpG5dowShm36
wKWKwD6oiKLi0diCzBuA0rxqZqZufBQfnUWvBTkU2kH2IOZbkNtDQg3DSKLHF9aNtNaQ6kBxu5tx
qK6Fvof9XA9hcDX6TeAggJmOKFxnFWHL5005hioaqj/XwAuC5/emOWismfIYbtM4ihiOAbEvUNhW
HLaepRkQ7xZVzR0nqr5jdFEQBCWI/1tzozFUUm4M9VRL+w6iLz45MjPfsozJOYZrFb6XL40DaDL5
dVR3XUst9J4UyvVLaXXkCBkaJVqQr2ThYX8Q6mlImQ3F0Wemxa2FIWrdEAjjK2rUs3kZXnPk+8Y7
WeKwqWSOjHrrcGjoPRvpjGzvxRMHUYdvKU/HDJrtADG/ONew+1T0dCGJG+dEqfrKfhYJh6yYjlYq
7/LihKIgAJ49nmeAS0boVqFO3bCIpfw6OcyHkAgPGx+kmeqv5elSpuZmOzvSAxxV5VvyeyPnjxQD
InRzel1kD8TT3zY04dj/J8iUwfZLn/I3WCCa+fKzLL+CaoZhxXfUuLLopaZ96k6sIxO2VSlCFcGK
zWznvJjN/tCqOKfhC0IXNJuTvZvcTWv6Ce1oVZcQX4lWd2um5W2Cgwp5muRXSn4dxjoKU2KaJV82
fv690sHPQ6pvIte5482anzsBklxEi4GHECCPxwDqvJvCj7pFwvKyCcUL2Au/4loORrMWBq0sjW0B
SLPNjCW0LzXtjTOvzqTDbRsXk6LiPaq5Tx0+Uj4YNkrmNOqG7j2I2B77rjJSWnG4hTyZv72XHw+M
texumtZZbS0Q5cwZE2l0YKcFCVSaPNdP2rh1cs68Zklklu6C+8DoEyVVIeZbuctY9tLVGqhYJXFT
hZVpmCtGfRK70DfQmMK25CKb7WVMSA0YHdgh0qFNzVGgTrRf6QhN8yEZ4z9iU21B8pXlp256Iu3E
IAhWubLKEIFq9kvlrjJ5LDEJUI08Oh9N5IbLjYZ7XASMQfdO5GKA83lJV9QpEd40RNy1TQ2DWB7Q
taMd7UTe8oNHiHsjI8aheCkkmVlBijShbh9Li7auYjb6eJHWMsFMiGKHFu0S7zKXUW6qKelNLLwc
AksYEWKClbBTw+ZPi42lG7iDqOPOtku00ozJaES4Fga0SPqkaSuVIabRyFsCvY2lcV9XOF39WMVA
MWkrVDuRGTRlDlyIPDFFMrvWGtG52nYcxlhUATxTD0NXFepdLgApBQNeahL/pFbBLXygv8e9jHVf
EiBxLKeqLUqnVfp4mVEuihKU2vB+7x8rpKszoVObtoSc6eOfJOpvOwwlmZhEUjF4iaq7M9EsdHua
eKbn+gMtWt0mtD0cCN43X+IEQCNsktrNQb/OSXi7MnVjWqxgjObebSyA78Ylw88ojL4284qGZ/NT
OeK/1+q0I9ViPAxSvUHmZVcoY6Je2YNFpd8wLHt7hE3GKSyk9Xi7rBnQ9l+oZFtc65FHA+YVq2wY
0an6BMrJ3iiSPP9Y3dOvUJHTnUEG/YXXcQnWmaSvNIlkppkI8a3v8zd0JS7GuwnICBPoKPB4VX/t
31qgTg/TmQZSyOS0Fl00eVyGzhyx70eFWq1/0rct/2uHZas4ZauQ9sP2htWAVZ0gryQFzQ/s5UKk
JKpjgSmYIOA9e63IvcQPL5T3ZqQJ2+8vLjS1ks/D29PQPB10XRxunufuL4kwKgpngTmedWFJO08U
Ldv5Cnc62HyxjVX+Ey0BMtFPW4oTmgqCFG6M1YpbjY9JbCKGV8Ca+feKPtZ/CILvRNcSlCP8esUi
jTVjeyYNH4hLXHNygp3Kk49B+T9aNDrsUcFaQ1AfKkiWS1cTV8HaabWJBE3ejXzHrIRIYpcchbCW
FaX0eS1KA2kR9wRWg587bDnfFfKP+yi9YkHS/I3y1rJhWI4KFvenVFMBsqdGjKVf+g9rBQEQ3IkK
2GYSX+ujhJxYFdG3EbdPmBWwTyGRg0B8hy3oR6QZGyAzM+hJE6o/r6C2sKVlbanu7spQNFUPfxfa
JUMddQCqp+PLw10qrMRz2F0eq7hQ//u0Qh8XUl+AkLtOe9ESJ8SDzsbC3HeWWcGcLLLcpJl/nRML
iFsVhwp3PUDINuPRUaANuwIbgGX7pp1KetCBfTTDppyhQL3mMWisY6HDs4uCCiTKte/g7M77HKZt
ne+10lCez4t4c7upQAfNPnGNacxDrzUtp0qBRUEd5BKqpUdPRcXCzcXtvOVNogeBPt1C2NhSoCPh
l8DURiMNQj2KHokCQ+xhI/rT21DuhI6ympHHj8JdHsbmR4Pe/Rn6v+FQR3R/G/q/qKZUg23T2lDV
mCQZyggTzv/G7fAk221v1PlrKhNUU9hbjgR49yNyaiOVFlWKQ1Nr4e8EqNJFFyQSTkLhg5u7+Ang
/29l+K031iKemejKBDsV5NIL8IExAZvP9EDjskNX8+xZk2YVxn/x5ZL0sFXajmSbnSUBul9q3pfu
mDLfWmjl4Qsv46yyEgVdWjtbWh/lHAEwgJot7vhtKGUab6gjw2olUaPQdJ/sSO7pRmKMBaYitf/K
IlQtLYozMP0/bTpxPAST2KW+kqlBbzVro2XTY/Y5UoraAQue45+/PdUujZJdd4q2TwsJCm8BTGyL
25fpj76kDcnEDDavO7AqeZr8behaqWT6ZUUKCdoFbj8TNvbhIuAcO1qKJKe8bY7jdjmGmeEFloan
4faJdI/ycMRxlPGfyA4Xbw2pCk5oHk3bWs1JmLP/q0YbRYCFhQcFZZboI7LcZPutFcKTD+ey6+XY
xzEnuGDmxBwAaVsjzhXYF7BOSEREqaOb7PRdD4uzpQDkRyb8QggrH6vFU8xb84y3WRu0Adx6WniD
ITCO1AVFVQsOOgJykN86UpnfsxmAM6vAaoH063dPK8oDjqLJIYDR48f8wTTAIlLE70rJbK2qfllG
XE8aZm5cvErpzhMZKvqNCSl7VfJO0c99qj3/Fou3Fv8AQsOMrZ6cRKMLvhTq7sZazyv9pUM2qhxh
FuRoB7S2UwsCU1xdZAnIjq3Lozird9i3ecKEzLFsRwqRsjfRoy50CCCyvZzCxK5XaBug0v0uCazu
Ptq8MzQZOmdVR3GsEIEvGhtQmoeKdzEwVbrvL7fvuyfw5rI9OhaFRE74Ch/BGEGowCW5cxmMd/9h
zcnmnK1tzaEB5G2jRQie2j2qKafax/Py+E8jzelqrxVrbxj5g0DTrYijeYqpu5JybMXbFeBmTKNS
umYFKHoeO5aNM49F0RKCq3ILx89vc3s3ZaDAozwnXeBlRmctH6X5JAZxLXR0ivdf/n89vj09CWrH
qlkqMtUxw/g6JApkNAi9xGiUD7MyDo5qBIi2bHwvDuGnkFNgLeb5gxlbMMf2aiqaylsUngGynrV6
HSI9ohv7LQglLC+DtKZ0BdFebKMfmK4womVhaONr9lqdmG/OcA5BzFbMBSPuqwB4Se8IRGwnWFf+
Kb7fOTfD9SIbz/3+cEEl59F2GcOjN5f0yr06YT0lDSNEWvRRkDWzoeMu5XWj8DZxnfiSO6t9yb4Q
ZYv8YArI/hwB659O2t0n1qFU/YD6AoYvNF8xXQ9AMMnsEurbU6X5d3MgHnkAnzwn4SWARIHGV6iC
+Eth3D5VZMXeYA5OkzCuS/6RiWifoOQHlPjwapKZZlDkE9n3cB5MLdSepyVtATZ0NsbsX/VZcl6R
FQF3/o5TgyJQymSrDATbxkt4X40YkQyQNXuLiQPinPUqZXzao54gTNOdBPcVUOXbgadGSyoa9Mrf
bqm/PtsemTBsGC8b0Vs3OZD1x6czr7mR/8ZfjloXig+zt2/aF9RcVAGDh7Jal/0GTEa4REEn4zKh
YSEuqRzpIfA/2nIIcVKaxbUPLKfhDhqV85yiZXulfxGF+BTVEm9l2hLatYxCoF0Gkj16dDWAJr0g
j8UHVR3wUN4YxcRd3zqUvCtVFRQKwsImD36AA/7AM1YoH4cwJjyMYd0/vsjDZZdqag01RuNQ1a53
+HF0OrzXL2OUkia7OvVIsLsU/9gvpgw2iqWAQmlJKXUktdSFyeGNz2D6fydBa1KBscf2gOBvXcz6
pqj/v0JdzTte0vm48vPsqcQRiyvJyye1M+zlSnymjTXYfI52wJgbhcO/c9NA1GrWKtfo/mb7TKrn
eWQEPhMj0Vss3Oke6Y3U0ZlfAXIpXJR331w/KfZS8PcFXC7Ul8nzKPTNJ+wZeGSf2DnYN6m/K0MA
gEx3MxP4XKNPEz/YsohovUKl2A4sRTQp0iIJidSeIB6xakXWQoJbDX43GekXt/5R8TbHPm8eEqr5
vSF7BzKT0QLyY54i+36ldQKp3L7FnGMU4Hw1uNv7uLh8FiDTC0VrL9QN3ta778J0ybCYeyyu0XLG
tETOMt/8INmXJDW1SqIa8yh0NsZS/M2Y7c62vEvpmcuFqaisq+0pjy5AGJ436fbMJEkPVvGHylCm
GgS8DQtVdKxIVp9JmU9XvyXyDySYXBiHPr9DkWA01FItCi62zTTenUaNfvWU+gWjI/tyQndXvmDs
o+pps0R8V2FGqEvkSGZQHmKDFb9+fI+VziHFB8Pv1nj/KDPB8a8laevV83S5Y7ryU6NtXFDg+aq1
w9Ff7v9TjMOyg0XQh4ElknKjbQ8ARXvOa9UZ+4K+Rvf4dyiTw3Ve6ZPkSpWbXYYPgjWoe5FN86S+
1sMoutLoUJ8irsRK/d39nlC3MRrirp4w0US0IDTxRnt/DeLhBVI9ZlhoNLZrRO+RXapQ2QZMcE1l
Dmwp+O15IMk500e5v50l/FS5vc41leRP+22NlIOXdptpemoEWLgzVXVah21N3KG2IuCoaAJdZz0W
Gm1FSZiGHxNBYniOAKmK5CFFMW4Le/73jiOxcPJIol1KlNkGfZ3P0rM+10F7XJXcjmohuMdG0RBW
tCF6ml92g4SjRGyeNlrscxewGWdR7f/BjiLensHpJ0qdnq8gvP3+JJxXXb/0/Ss978a0yVKtv6aJ
17e8EjbKpAf8wT2lsd+A3Ap7mBoNoz2Cr7gUhQaE05Ff+fKyUFLNW1VkiSQ4/0YyyahStZqwtNb0
U4N3eDCcz9Nr+q+UGIKHF5PHp5pfDjX8o46HuxD4FErGn+ZiVKS4mU+m1IkMAWsxmBZzP9MImMKq
bvv+x1syeAEb9p2SI4w7WuZ2UIzVheNseyYpz+TxpZLal4gFW9oijPked5Sov+u/+Isn0wGoea98
bPysgFczQFttUdOhSRzc/bpZ0q3ha8AvMxseOuKIK56BZe0pvlPEq3Gx4RbI3GlWSb1Bq3vhuUPr
SJBXpSRs4P12S21TRlq5oHVkg4xkdsQO88I1oPbOttLcHQK0i8Zb6Ih4Pm8/mgL1qEtmH6fOp098
lrZxtQb7cHPjEqxAesl6D7vSTHVrWse8JB+BZUt0uVLXHES78jiZxxLKC9Cv10AbOu4VVBn/B+oo
GQ8Sn2n7vbqrLVPIsxdzNmclmKZCEc6cT8BjdJpmHJg1fHDm7cot65RDLywKH3tJnOhd2153XB7z
FLEshWsXzLMDM46t+SDlL5Wx5GCmztvXjuzu1k72Oskq8pugpd5IYS1iwd3c7xZolPqsOnt8jZOt
ZuvPUXVuOB4yQLDKBGzwrofASk/G//ynw9EAc1HhaUK+iAjC2EopZxM4LevW6GSf2pZ1e9AcOf/L
wKufONQUbcavo4Vw5AMlept/+cZ+1/TyFwD4EWPmpRShxeGpTCGokad1TXez5qovzZmYRFEI+w4E
Qdy2QAkr/5aeiUyNELPp555+d8uDY1xeTvodXYw1mL0SUTX2v6oq1skwBJwhywuytgUN8nVQrO1u
j7ppVmEpXSvXZ1nZlsBPqMf4hE2B4wl5ITOfarIlAtipNQIttCcIobGcxQSh+xk9gsVuAKrgWJGE
QPMDnx1H95RIujmmLDuixPWz7wtUtpahlQx7FAu5tuspsIRphNtgdT9UrTuwm+PbhyLbDqT6HsHx
qFQ9qc/VQhP4wwTpU3ViwJiFkO9mcBR/Ru2rpGXizFG2VyqV98c0Ud7AqXTt6OKTuRWHvCmsm8Mb
aN99fiAuKTiMfx0z6Fz84P3SjZAPRZ0ZPGWRPwsApk+6FclO5ftLyfnKlDtNHstK2qFJFLVZDXx+
uvGToSZPIbX/kxOVV3QN8OxbWIQObFn8OFt6zXxzKO3vzAv0QU0KRK8I+pd/WB3zYz3ZI11Z+doD
IbmT/YKOqRIfWInIcRMpeZMDz5QE0nf0o89WVCvI+2k0LgkFbQXnoGLMhQq7HfU/E5qhpPVs3Wx3
K29ozokzXZSldBp/tGOMELN1u0eCrBdPgWWk2en1GFKNheNnvh4uViX6jdLiTcYQ2uNyRXTih8WR
OUhqHZW5BAJRFNyTO0KwBaeUXQn6URQAhGACpiroA+6ul8h0YtWEAfuTz9MFBs0l5XuNGSzKdc2N
+FVR8RJKYrl8d6No/VLMo9dp2WUII0ik3sGBSBcarl/U8P63IJJqNoKulygSca6Gshqpf81YK4Wa
7jmX2YA8J2xFd6QM37komlwxeGxiDlPIC4bF+fJxAVXHhOQUd3QvXA649ZnmPwug8zXD0oK9E/nk
AWXsSpLvYkQU/PP5FZGnHtkPEM+g+obykowS8YWt94oiiFASVBkxC+IYX/9Xl/2HZJ2P+MFlycn2
Q5YnwogshTEJbQyP/0Ap53CtXkzHd0JiYstute30BuOSEqg1KFYpuhAO5N5AOxmoC8WQd046n9Dh
4bl20tz5CSd6usEMma4jaImlaTRyLEjvevQAm6LVJT+rWWm+c2LxYUbD8HmIAEHBnHE4/SKgk2Yk
rCXp8tSLKle/5R8B7gqBRcsxXgF9mQdl5v0O0LubWUw/tZRNKn3p8UQzbqmcrBp+mfGEyaEk5bC3
ST49RWjzJGJ+ESScTjUl1Om6GGF8yj5J36Uob2tOma5F9aJnbRLQqxIZIJ+3g4YCAfbqvTXvVp8h
3hyBG4MmbhpeHOGrCXAlX+Zi0HhDGaNkmJ2fo6uj0jhXXtHUbYlqlq22sa81zaJ/9Ldp6FV9Cbx3
k04wFp99SqvdDhmkiYwUWN46+Hh/ulOM9qLFcRRPIsJd7CHnPsHZnTjqkKeL9alKAcxbn267qL+e
8MjTj9UL+R98yr0rR6qvlVPybHbreDrFwrNzONKMG4RyNXv5OO22ii2J9kCX3T+/D49jyVUikAGm
L4vKNc+tEEL02l6aEcAVM78YabOQSQ1XO1vZgU9u62yHIANlMTVhAVQM4mkvEX4DzCsu0c0AdJZe
py6Lzw7HWzar5SpF916HskTmYDNFGx438yYsB26daHIFx9UNeuqsADGM80VAb/Rts4KjvT4BewIJ
fUrPAJXUof+rcnisDc7HD4ABYgmsIc3hWYTGLoOt9WktgMcPyMrE8vlQFTdK/foQ0osMbaXMD/vb
4xmysCCH7A9iHI1tbDJ3f04Dw5ZgrvUPcZj3AI6cubG0ToCnpzryVbodJeVU0gyWagojTyt77Rg/
nmtsdKXGCVLNacjbib/myrQb0a2fipQFcqMGHopu+lEGV3cyXZ4ICXFba2sR4hkQNTLv8g166SCl
1FvPleft6109v41vv8JeFmzMgpeFRNIm/3IaZCp87zbWfr3CrrzoLvyIhxGXdc4N3VDhuGSeqTqC
mW01s5DSrBJyCezcjF5sveXeZJX8n9wZV3dIWZ401pJlrW9SinOTg5hdyD47Jm4kX6gZXyEQ6HCQ
vgcQ0cYQjYflMk/X6U7g3OvgiISM/Pu8E5/1jFh+kdNNSQIEygiKBiP/VzlIt6KfsxehUYsZi3cN
gzTF5RWuQOzW7RGWa2/VRuKzFXgLF8T1wAkYpbSXzKSnlKUyuZPJGctQfficlApwT0QrV0aXtSac
qUIUoHECp7XWcIIi3ktWVY+2XyXWyDbDwuh1Z8Xqgdq9rcVA6Vq5o+5fNCCMBGB/7dsR94LtYc9h
lt5EpHciklPnvgQUgERK/6IJl86D15YeZUcF2y+IW5jjb6koKLBK6DQoCo/4gcf2DJATKgqlSV4m
2Q8b73aLbSOSgFosGkEAF/w+KA6f2wyKo/12n7TUNZNoshImNJTA+qA/3emcOtyG7Om5/casjEQ1
hpTjjunPWHDq4mOxF8gKsVbpdiNr6QFLIvGIEk7Pfapwf9fXdFi528P9z35uapsArEFTfywkz/nX
Dv+nqW9cxxjpovZa+GoXGS01UNl29XIeBwVXXv8iPc0quwZAs21CvE9je3rgLuMYMWlwoxTDmgEY
haYpn0yheL6qOOX99EWZyYZrRd/Ibh6Ktr48VfRZjfs01TzMcD9u5sKIekNAyvAuE8wHMpzuliiq
iNF7NUn4Gg8jKAGNkd89SaEuDnOl8dTb/N0e6BhpCCYkjwOTfe9LcIKppxFAfdZiSactrKjcDRvs
7SG7cpoHQl9NHTrkmxXxT6maN0Ap5ftl7vKfPL532KCHUb5u67y1qky+gV1ZSgu0f9n5+2l3jSZe
Vrvwjoufb9jvwLYIEls/SyZ1p6jPBcVFRCyrjLe2e7ReSa40Cmf+2d9Hng58fM6veM8Mvvp9AROA
ihgUXENM4mUXDFuTeRNv9muSl2IUjyifyr/EvroI40o7PP5v4QZ7dhJWA3fwrfi7F6lj9ZzpiSrU
LXTXd+i3JbG3dTJDntP5vdV9Odwxb26gPunrjz9aHffmGc40/ahUwS7TUovUKh4I90lf6zm622zA
34not9s1sW9Ym48DLDoFhuwhTwqyz+Hco9bui4l+EDte9CTNE0ra2sudiVCJG6Hk3ydbnnyRx5ZE
G61p6OCvVXQltAFSjUH1tFzUTxiGueH/Pl5fNDZ40JcCjRZwmjz5bgGjmxJOkjTy7V1WLmuHScSP
0KjpIu3dzoHzJ+jANUmKT8PkBm4L0KCMkxL1pZ5fX+3/F5xC4dVeO1Tpnf1eWW29SF8Ea0H4eaPj
eoGofoxA5wFuENwwbL7DnyrLj4SoboKffk2Ju74LRG2RORQbJoXkVUd+L0pnz4Ecl1GHY9X94b9R
oZi6m6hSgzv2h1k0evFbjLYtkSe21p1Vw4WNSz1gPnUzl9thzKDqqkLw4/KZXeAQePnXYMniNt1t
gx0dfP09/D8nklSGUa/9wubM88Lkb0NvUIwDU+jqiE6F73CfXUpHvEzQKPUVOT5wI+1MZc35ffxp
NDnKgJL7vo+cuqi55bZnvHo4LvyKw2hHA5NuiANZN3JlPF43c7tQiXdquC6ITK/slxS6OqG4swBS
6XmGPIjGm4dY9XGv4yaBOieFkbG8wh4z/2/61ql2vuR3sWUaWrE5vLQe1oWHmygJ4el1ZYMQfvsh
CunXzW6SP51XxxwM4YB14tVP3M4pvytJNQe93oONER7NtPSoVAy4MI4SoJL7mz77EXQdD7xelQsl
BeSgzSaxxF/duK+WbTmcWwlXHbPIZcAfyRBMWr7i4/vL1rAc6FL1iRPxltsLaY4TAhi1QXvn8Oyp
SBLIdOU6GBL77vtNgCZ8XLb0/qB607lMr4V0Hw0lgpbg/QzyRkxPsJ4MVDXYd+5vBIDBrS0t/sD1
I7ejKj62EYIf63IpFQHrMycUSCjZxhPYMNRIcBxg8nwzHLtm2Tp7bGeX3kPLKF/9lqRF4PmyyZOF
Wqb32v8rxcDwIwwGsPtzxpDMIfWw7rFd/2fPMA3IMN80TTlrO2AMQQpTedHV0ebc0r6YxafHG/KZ
3leLANiojTeaPnEsH1mWxQ+bqQud4XEqhs0HiahqwFpIJru5i09r2wqHasl0FfOKVzA6sn1ID33l
2MkXKKsqstNH4HMe/hJdm9OIk+Cs/CWQH0mDG6K1esZJ4ihOJz4YtMHyfPE5QD1GG9Xl2veazAPb
/LHQa7cHmyPBkgXvUf7SeZqf0EEJiejHpYqR4/YVim7CBG9mEtaq4w6cOxcmaPDlewVgq/dj6LrT
YSuwFBx6u9E0eUtcWk43x2XwpQEMNTEYIKo7/ZWhAgN5b/uSa6oiRm/qctjNFDXLUTXk3ZeG1nmV
ZOmCPzjkZ4SHC6bx3ENvXJsRXUJAiLaVF5uh9WkQFP8HDX1Ax0qoT6WCUIdC0temdzxM6lSQGmkh
bfekzJ5J15D6FsCfdqoFsAsJFrpOG31wjbc/Hgu8YFo+ZqMdCioSbtBe93C5dSqG7AGTw+Gf7pdp
zLswDQ7g2OBmsNqsgiebfU7qb3bvC9lufapge36+mi8c6fSIpC3cZYBNlJomHpyXmNmiOUj7dtJw
vriVHXvfpuWKYXjl2PpoClqGRGS3aDgLS4kq7dNwxv+f4dPdk49y2+6j0P/Hi8rixgdyB8b+Atta
oAXxi2KZ/t9Ay3NROsvoAX2TIfSUFAH5miO+08Oi9CGo+Tk9OLFrTWrcPNqP2rhVooggDjSblVuR
YGeAWjTn9OVl5k0vWbQwOqNQJuOaE6gvnKtFYiTvmlk2DDDLky0wRZzXk/mTtAOHiaKhwbzPEpK7
R/kj1Q2R7ebRTF14kzYf5UxtKjAxNptp2echgh/As81zDNHRAZkTTW8ViyBKMr5D67+AzaJLgQqj
wHhq3Tt3RRhU2/YTF9tg+0Y6Q+DwanPZIGv9Dx4aIDwxulVsT1FNqTnoqCDruBmrHa+e4KTlsyse
c+IlBsOpFzqYu/t03Rpbx1jGLIYPyfMtpzGw/JDEDVUjbCSBuCup7WcgFp7x9YSIRwRvNYs68Jva
FytHK8+lmBSqkI6vuT/z3WdaBRty9iE0j73KFMq4piJlncjJiOKJ8fQlbxZWY8ExNe56ouoQKfhe
DItmcID460KU9UUpCNhQhA87fLDV6Eu9NOZ+O75VxWXBMu75Wwej0Ui3HVbFmfzcMgPrAzKCij/n
0PGBikQ2HphFLoyYGUne9HmFQKFh9RYOaL0LsMkZmMw8cC9RvTDWiTEm+x6g5szVdTI17mLS5r6v
QfmENMCIXD59OJ1CPCTb3mv4hSm/OfWGjW3wCrv+79tdKv1sCJWPQC5lT1ckZx0CmIFVPaXTXVYx
OKONmh2YYA+RXoDh3eOXRkn0OxF7J47LfA72AacPAn3tDLXePGiOKQRr3onTmWHzWFYm2Vazl+yY
vAScE6dqd3AK6PjQ4ZQkkqhC6+dt96C1rxZasadHLxomtqjq+9VxaFo5zts1/rFlWXPzWjoHq+sl
XOrKpRGI3KrGPKwEopbGV34X1pKEJ3nvXl0RQINL51e4OflehsACzuq3QLY8SwP++r7ZvFo01MTK
KKMNum7deYnxDse5ucRnQ2OS5i69ig1U6KsYfiNYWfKljIY1Wi0aVZIvqsProZVb3j/9fLzRxDa4
eVLEchLzDmID7A6DI4Rx/IYq5L2YW124qSbayFQ+iwWPoQlrWy+5yuVw09/JVU2p9NWp4CsKzW0o
cZeHzoe7ItcP9VwcBOuHrvVpz2M0I8OCVtcEH3HhhehQd00NR7xLVr19+tLCNQPdCHenqHYwfrHh
x84u5GuC+T3WcyAFcVdX90bdb3TDcmnkFxlAhglScpjffb5gfS9BwEqLnM8k+yt+dJu7DkapSc1l
jqjE05AZ0/45Oo0J9CZfUhC6bTJdrZ3w5jlPx9Apdg3DrMT0X7Z75aIsGnjql2idTjQtgFt3xJV8
FcyTT2WUZv/l478E8RU12wvu/TZO2qKPtU0U8e06ftJ9WFV0+Aux9i7FnlETMRDsBHjH7YJsexCO
Sz3pdWGe+YHgGNnImx7ZUPLRjgAo0zBFU1YadCIwN21TfrUsiSB9vIyuFhup4FaY9MWAGaN1XP29
UXImQQya3NGtsgKCz5beE79xoeOtYgjmWodEpsiBuk9iWMnyYWyiQ7wHdqjYK/lC9WM1JymyhFct
xtfvNgBraunLkWtBRGKfOFYc1c5EwyHxGJYXhRdlyrqbwaG0ZysXjok007SC7TFL4Gh3Nl3ftCSg
RezkHYsag+yXmyoeCZN2WxNoG992X1jihi9jxDCZ9BkfEXvBg2j3hr9lEBGAnqtHWmgTuewrnBk0
pnYjIoILAWRyMgE+WYLpqzKXmb7v9ZwUSwkWpWQU84jze4xcm/jTTD/pIcglff5v4ZL9cIUABu2C
8B+cmKR1YsKJ/P8/bktBkZ0olXMCGNWapqMtqhz4vV7PUTmVRvV1xxA4lbKyBmul4DBIplhofpFG
mwVVX2QrkE0HtrMHfDcCrdBA8kgIICJM3q9WAq5cWZgbIMXxtMfkCeE9O2Q7gTOHNmFnumu8tKDw
YgGRJ3RsfFQC965vbH2lWAwd26vRDtmpiytGgN5v8ROg6tK3btF9POb6AW2YJKv6z/Q/KUFYuY8x
qeGnIGVhyCun+9B9Dzm3QRurXW3CUhWtBzr3FzSKjiwrWTlRGNryMaVti0Qvq5lAHYaaWq4Qsih5
0XVU1FXpwKClmCx5BOBgr5yxrJgoPWNxgmHOP07FpFAjy5r3AlZdlPdtZ9W0+3Th70bYbDOCWSlZ
a7LIEgVZpUqsbtOQEIoJ6rsCzMKU4jK7fcp4rqAHuWKHBDIDkN8SBreqMcGsenkTLTqJo43bdHKn
U90RJUM6OKInZ9quVLYLuv/iG1zgJL0BkBGKdRKApVt+/4QvWCX5I4yrl48DQCl5wg7oNWZ9h0/Y
tpHIENIH3w3g0712RMFsFUBNJD1iG85IKCOcusER2lTiuh912uW6806GN1aUvoO9oBnPZneOyLUy
IkMqNJlvKvceCjL3eSJO8hXHy2uQ/54Go2EufxfA5xshBrUBmImmuXn3+v+4RlS2ONHqh17SSE0C
eTvrLlCDaYZjzyiwUIOEaniGPvyFBqDN+bl5AidEecRbwXNLWp7t3zL7D0SMtD86z1lur/xm3uSj
JeR55dt/t9pHV48m5FKdPGyap3NgiEPOBHvJIZ9Rf77OMA/CWs4kdr6v3G6ZTRI+WS9XkV5JN/2h
GMXGKfOBDonBXKohSJGLnO0Ca6sa9UzWSaMumoAq1lMtW5VsMnx0KQgH/grEYolzIz0FzVIwsvfM
3KgnO451s21VSqFsfaX1gFaJkQ2/IJtrHcaPFAA1aE17Dpiv7RK1wb6J0Hg+okmODKTEuj0lY1eq
l8t2jOxwuh6En73Y9pKeemaMD7DOsD+0o1XPM55AVdNOWIQNk4MMjpD/OCKW91qhR1KzHG8+TP6z
S9D4kLyld7qwk7J6MSh6VIxeS4O89BM86AEp0YMt5jJWJ88oCQO5GYHnuLMRrPQ3vmfbu9/hfwyN
7CmmRNaOWGH1c2sVrvTMsHSpPTnCKaaSXPRuhphC/9ZWS8WVO9eHEgEdJBR1eufazppnn91TiUJ9
xgPWq7RT+mKovGGnS8qdSW/fUk/GLV1iq/xM3m5gtU+hBh2amWJFVHP96JDlcRjZuSWgtXAb8ZWB
NuLITUq89k9vE4t9NpqVrtWuYM0TUBQ1D9Dby+MUvuMTVdtKzQXBr/DB+lyVp3g+/IpFzZmKHMsJ
fBRbK+/Uzsb4NyzYe34EHO5iXfR43ryLs0pFndOkIJOfHs+Eg3R6+Q/OhO+/t6qqHxCKH9cQS31v
eBw1Ee0kNODTaTDfG7VBxMyKPsXMr0B2lBhuz+nHWnqgOfC2GKAnZEkPhTyrK+FWZDA9bzTysTs2
hhO+a51VaX/YIPRq87lc8reTwyxazyHV2wHlt4xVesfW14L6glulofcbBa27Y0ESHhBKl/z3Aer5
g0LcCT3BMyj3QIrvSzguHUrMnPWrb+JLpwA/vpvmGFcVTp4gJqRATd1nWcsR0wZnI/23MTacSbqS
X15AavSZHj5qUsWkUF2LrQD/uuHmxMhyIzTVn+00Vu8hXYRQ98xyFlficy2L9zWuhwFTpG8O2unK
KyslCw5av78WOLFQUU0nEEV2uupuZI3GEKN2NkbiWsbjqB3n3hLDGGSuX9tC9Ea37G9OYQ6VCJGs
AKG8+Ps+nNaI9bt7DPPj2diI+vGKUoyDJ6lXm8DrdeNd4vE4LOYEg/os4dVeyEFU1owTY699+Cdg
71KwDTigqz6w6xQd436WAfdDupANM+knx2lxgIQqgeqEOGqKB/Y1Fswr9vv+Nvjw1CNyRCEoC6Ko
tQ9hjlzZLV4XMdhxXt1fMXj0z6+tK8xOvOsx2Ud44I3IVH4RxhznrvkHHqYUpWxaOxErFnIzFp+6
rSR+y42ezamleybfE8B3/q37oeB99i1RxbQIb9WwiffJddxF3lYX9Q6row0ypkF7b2VTSd1j06Bh
6RxRP33rqx9iWoMzBdB46ATbi5uaCNCVQumuel8gx5EdMpo0lrjXQKcocqmMly819/RNqRbLdzWW
dv9MjjWUMU3mJOzs6t4KjzmRSgz4a3b3HfHt1uMWsjnnxsANKmQeqzG0N5ml5r+CLhCAMGwWhlib
hahAT6yqutjSVRKeUCcYYWz6nZ25B4XZPviAOqnXsR2ISWWBAHJJHzhoqtmxyLeT+pmRsmdPU+dr
gVphKgffa3ZzWbVNqmsQsl2yTh6DaAUkci8Bq2P/004FSC8fWX2EYnzQKbX3FebxFZ/6P+j8cSD0
HtzAP5eGXenXqwwgLDWx7ncVCqv7u4jf/Zgo6uy6ArfRfecYiP3/IamO1TxBBp79tV0MFMwjbHUF
gnsdZRR3wSao/3tXujH1aam9IO81q4BSqcM/k5ppFIvcCjnPMXRq+zJMeTYpT3h3Zj6fqvSuZGm7
azTgMUtbg0JcCAuiXIRb6d9PITfBONk2YFqn/pEab5zB7pUktyxUbYGI3QLEya3mbFHIt9ib5FTj
1qbLE/1dDA/eBI2QjyMHBnB/0i8rnMrxxCk9CudpyxAdPM+r4pAcGZwakw8TGnLh36laTjhJOzIW
6hoz4DrxrQE6Qa7r/+cJtb0FS/dhK6A1UNhkxdWmmW6bsdK2aKboQ4SJmWm0vgIssRggvexiTBQx
/V8YEf1QoDGCGdiTzrrVSAuP5YHyT/HqC0LKIv/PR/uMrhi0P/EYL+sOMC6XV3Q/l56RAYx7now1
Xnl63hZhG1LaN+6LgqWObqvS6A2PJKXDXaBlWtFlMNglKrE4319DC3Vlcd5rfJuF0Cxz1L32B9VL
sj4I4WCeLqEgVl69V0PqWu5U6A/DjwfCo/fI2XD/Ka/hilDqdYvKHKO/THlxbKL8RC179ZD4lGZ/
wySFJlSd3UsyAcjMX7M4bFsua4WhIvIsKF4zEPL1G6b/NpbdbRyfMom1UjXlbC7+ZnQtHhSlzBpz
MBNIPGaucSV0Z5K7H54Uhy6rLPmA6kwqIbquCLXOeg2U8CN4g0jT3tCzLNiEJjyauWBFxwRYBvMg
d6jNIoiOQbNvmUTihh1kj2r3wjYZ6pn9Iz0F44/0H2ySoSz6fPpXPNeqdQFc4dqQFKH+l5RdL70J
WBG0zw8rFeNMBB1Gf2xiyqfm6BCU8tMwg09YpxRPvqqESofE+y6lfxiiT2GVq03Dp0176gKLErWc
fQ7nA9bMkSkPABcC1sMwgk93qtlk/AarJR7pE5HdIe8mjTBekCw2OErU7RtILyYkkNo+BQ7fJzvj
ZILmnLlM9rkE9xA1rSJRxNuzT+f0w4o7/B3oDfBe9VC8PkB0zihp/hcG0s/II9R2cgo420EO0YY6
wAed8mKD7y1Jl8jSrxwPfOHY/wmNzKHAj1R6YtMMan6cfxIVVha5vjJRVDjlokJ2LdksGaY8yQQ2
UKSuzpAryMV+CZ8uDO2L9c825FdD0kB8cUl16s+h3BGxTr4quTxup5In0eQv/GcxntuDJSy853Y0
79sdF30krNK42gSj9epuktIwNpkVjB1tHpKuXEIqpIb6BfMcJVYR4AApC3Hxiol0ckQl1QNOY3Un
MjtGGw2VXt7mAd/8DqY5aFMBT5CF1ITuohDGTT3Dj10xfIg0cWpd3AUgdDrU6ZZmMH5fx+ahaybO
DdkXm/TxHAac7qmbWHzMcsum+k8N874LM3TsniWPdaB7KVJSK4JczLutSfaiCbb5dW14QLDHdw6C
8iUXgJbSbHIYeSwb42BM5Lv1P2Ga7qrqs1G4hsZZ01wqHy/ao5mKeNsBVhEd4VxE6aIUG/Sjpuz1
Euw09R0I94V1Va7FA77ZjmrQDqCYeZe9WXbpBf8Vwy851zQotI/HZwosDvuoVmB0dSEstVJ3MitQ
s93nCGKbwcp5ub2cNABvMplF2G7dCTv0CybWTfbpr3PBLPCB/MAiTYWataHeQr/NVjpaiis85ZpG
ESPaZqh1udtj+5ehNbw+yC8FOqkvFqwGnQ2vSL7ISng9sUklonN0jRhzwWmYy0dxW+Vxfso33TsP
7OmvG9upHiRhGH0P19A9gKvEfT1DmFKGpDo6UkqjWkOnEEN0Nw92krH82aEGAfK+u2MRUb91qoE6
TOh8iJeLOKZXjOSbWdGvyvhcQ/U+SbXIn10XmhLFv2V6NKFufYGjS+IXVjc+OmSmBui4aBYdfbBg
gmPcvE8NPG5vWKI92VC8N+CVkL4QauFPdhiDTb93MnrVqBfm/Hug4zg6fWAvpKKt63lypsmQNZho
+UCBHsh9RK/C5nxynnB0i5l2tQd5DU8O854U5QRIAwoU4FZvZi0kSpMLq7trfN42R4hink2IVgbs
W8qUeXq3woz1BsBiIa3oIsIekFz+MuwwvCeP0ZUmWRBXNO7eqicmyeWBivAweWzqrscCavbK15ac
cnWGS/y9Mn2NIKGY/1tZugQdimLbpW8K5xXqjfVIgO6uy2aaxIAiycyKH3bSyX1IAycNh6daVjNx
LRsUknVLUOZi4hiVLyzWJvCLnsr7vtZ1rukvOAyyP7rSqd0085PrgcuzNjpfb4a/z1BM2NLncWn3
GO/2ZwZS0nRDBFbIdDRp9hP5Go4x1ygCmgumsIe0yGaH6RHQXvE6z60FXY0HfSqA1vAKNhr4W5sV
o2RgtKFndO7zhvYydIJFOdiLNorECnmelh/zWVKPRjHwPK04AgYWzpn8nIWKbw65QcyPDYNvbSMN
PZa+p/jXpRU2if49r008trgDOBdxFyzhWEFVd0qZakEgWZeRVkJAuSD+mZbFUnycHRXW40KUaP53
TAWTi6mvRzTSOOBlganDlwypv8a7z0Zs7jScSkpwoZKM+WM9z9tFp0e9ySyvqn8c84PXosuXmk7e
a+g/tapKJZoGWaROGpnMNSgcIYNUz3Ju85cPv+LA9Xy1n9cjyAVk6TB+yoKM45OmLuk4oD3sEr/i
CqURbrN5TaaAZcNI4p7TyZhAnfxyllsX6WEzIPTHh0T0XHlUSl7oUzOkeset7gJcfzXjM89sn9LT
Nw74xzg/874EDoIckqoEtiJbiqX8qgY86/iJMMS3k1mm+67DSE+ytcY/KeJbJOPBR11SG9CrlNcR
uCErGuZ6O4xpqB2fQRmW3RhicZGpK/DcpRoeORO2QuICABYly3UMg60DEpHuFhMB/34jn4dPK1MG
131wZuT8F+jZsY+IWutN+Q/1Jroerct7MArjYgsZ8jwTwnFKvQ+UJ8iWFa8Za5EC81P8xmjXACnO
XxxT1QYMLrzQemefFTJtIqEFkb86R7WNv/5RJuN4reEupr/Ic6YMjLChc93I+rhAzuU4E/fglSz0
Al2qDXHg6kMN2vXmGsoFtfmJbZ9loOUhAK0Tc5T/txTKESXN3LAW6v8USqOXzzRzHF+j3+mjd8Qc
1QU0Y0s4GwCe3HZxNgyyE6ncjTe5hSXbypfhJYZ5CnfNoAH+9XTs8r4NKtZhsrICmJ9vhd9jnPDt
+ufcKRdbb40jWFH7g544oJcaO48xZ0oZ9qcynsdwpHYhihK93RwIRtA5pT0ImB2zz5vQsRrZxrtK
vt3PF6fTAPKccCN0sF/mz5Oxbc0hht5B1BlLLFjdCCuaNdm7LGdNoggXAOim/T+VpM3b+J2m4fzN
Dfw4601BL5O8Az5SnHyPUIx6U6RamWe5DTGmSOURhyNu41w9zbXbRMiIN8UhEUH/Xmm1WSEnCtaW
2levm5Ii9ZMZiWLMKlkUme3Ru8LSSqE15MBvzMypodSR2VuJbXn2am1bxBdYmPJelvovgRRsDjPt
NjFh8BiQisRq7bnbWyI/CCyVTZQguBW9k0qm7mE+NgjjRLb4hj7DePajIIKJAlITWmkpqP9lhu/C
KVy/Kjg0A0dLfyhS5q5Mqr/k7pTj9Y1/s0FYPUD4ol+Nc1VoakvXshD4Wn/nRmnBO3drhLUUl+VG
YjQMcrtf+xyqgG7xvdB/83mUU8W2NnlsrnijkXIN+z0jLi6oLXKNeJPCBWqZy4vPtnrfpBDydR1A
0hYO0p9PJBJFDDkQcxWDPEIDaTm01gp26OzoEKQN3WQNH7k+5qVw06lAgwE1Mft1vaIS33K1EbWz
3oDgbhmnQ7LtDLnSD4KN7vxTdJh8QO/bDRMXU2eukeNi+jfZOqqwNYnuswD0aszL5/lMUk2IqpDH
tdgk6ZIlFO9UxbG31/dHLc7rPY7aAoPL5BTzDgJB1gDCW8f3pXZK+y+8Z+yn6XkaTcqhTb3yn7c3
3Q16jGIAHTAH0VGPOjsutJzwgAr79PHw+CXI0poGuEzyl1FBUHUWugRAHgzeciZHTy6ZuBFFj6iy
eqU0GVhKKug00AfLvAuTxeXF32+bGR5s/vFdpBPOwrxPD3hfPC35YjaYySI5LA0fhCeygKdx0SfK
P+uA9X2GCSBY6UK+ATHauS+AvFMPIlfeicAXki2t7AJ69LAyLerA94ZNmqETKiEPP0w7liZpPHub
zfCnQYCmrJrxOIUrGh24yelhbkfBEX0/DCb27vjV4E28LUT14JYWSn4FaU5KTj0M1SlBfECVxLEl
M2FsoK6PwYvpaR93Cs4lp3rzHvrjm0iVU9lASqFiquE/4X+sKEwbG2dv2yPIFbWb+1BxfND5Gl1L
Y0OYMnyzwFsPQP+HatRDSDMyhHnUicovyLDSK3pf7T4GUkXkJm4gHUZzEgX8LQoH1GgMwU6uVQ30
2lMQgHkCesrxtF3hdWXoP6UMim72F93YrAvzm88YDGZjjRMSt40PxaeVt4nygqZL/Mzx10XEqwX/
7366FW5g1zgwt5lzmDnk7u4ZQ6/976yY2t7LOq+SODw5xkvhUmuJpEcdWEnYqnHATRabHJCDeGsD
5S8d0FSy7HpuC8K15gKzTh7FYrxDatpfFDdtCvrM4pRGm/lVV96pPeGmSWPQysrGeCN9JdsC098k
8p9Gq94NJory/Wuv8suOx+4W9heEmGKCjr84NiVVcuObrUHI8RsmHC9+v+FKZaepYlS2VZ4NIDHq
Ku+GZLlCrK2nvs6K51MYf9+ILSLUpwiWPcOc17l0ReEoVCmOlz/GW120A8rQwCfeU2FzBeU697Ej
9UT98U76DsAfpgtBh8Nc4dg2yBmtEgKYBoNsV436t3d78MZLnuNeYImqygHWA7X4MDUE0T+0YaAn
0yGJtlCbRFryiCqeWfLXkMfCYAp5ro4hWtf86yw+o62S9mfTPr1eS6sMen6aDe+qmRJYQlwjJZ/P
h2W21Nq73/tHN30OGEg7DyH7wSNJ5/7JGN+6P28shwaBptEAl7462DOGZpR65vzVlTNTfj19IVU+
A5z32siROiDlruaTWaw/3YG35LxqKowsxNV7JZWEFR+3ZuEBjGYMyZcJQ/VDo+V+qlPkVHHr2dPY
nPqZCD46ey1BQFp0dIrHqBDlSELrsb9R7pdP9rAScNlmQE19FZv6KRmYPVkhJ37gNe2o3fzVTc8q
LzXKjTCb4dK1m9yMEYnbCmPU8b9VfhTSH51TFf7UIy/0ViwkVmfaJSom1p3pzv1q6E/D/qWTr8qi
lj6wciDT8EdC5mztlJ+OoTAnXEBmRluMbHgoswvSb5KdWpxoXUX38aSjqvme5VUxF6aAsyS88QRf
c88RilbTdDHphYlxd/TmKoPKArA9OY/lKCu77HkEjfyHvKYBbp3aPAp8yX/JSZv6n1+mQdRgP2C8
x8F9GgoEfYaoPf+YDDB16vEhjLSZZVUjwskcZE5zMm3GeyaB9u8A2CgDRBk6MW+TMIPVhuJghDoi
qBKJADc9qKU0j5lL2A7X8WUS+fRcd1h1G2VJsuDO+wnsqu73TcMmHnRO6jGiFSotFYp6mheNtlab
GxMjjt2E3M7ZlYir7C4nmoazL97JJ2bermrK+YhuUUJ+rU27sD+91HJd36PTvkQ/kc7NUWdnLmr7
nI8GyAgX1lCqSt/tQ2nWhYXLOOcelf93J386Rz4Rps2WdcLOBorF8mo57QejNMe8Vi19QG0+H6lD
9QmbdYf7/Etqmt+eWKyaxHBtYE7JJLyggCk9xlhgVu8dhGYMc6uIfWHJI1nlB4TGZ3GZmOth1332
2Po69a4jdW+8idr2iiSd9yQm0Wz0WobXG8hCEluSQEBePRioEG7ktMC/zP2t1twWNaPosu/w2Muv
GU5LqPApkDDGMVoBvDphnyl3bEaD8HzJLIVzVel+WMUiCz2PdZRyIg31KPLQ1+E4pTpVvBsONHtf
GmKkOfv7oJYq61U4h4cz/HThea29vM1G5X1wV6gLHk437jFpa8S4UzKRgS1mk/zB21nobfI57XfN
69iRS644SMJc11L3LpnHw3c17BDPk3w6P27cr49Tdim0TLGeMAUx8heudh5Lw4o34FUXD3CIqIP/
ppc/eh9dKyjOjWJq7f4vDkyelyf39d99XPKl+aFd11uW0TquQkiu4HDjONGCvrfF4cd1pmLojk82
Rwabo3zpXivTme/3jWltYN+Ax8TXrDz4GX55xuOWZdfIRWcGpOoFIICrnFHVCBqOFaiGEk/jwi1D
wFNf01Gv3UQCCHllAkFfV0avv75LBzrK5CCL1DMrgiYJN2YLzsnSr9JLK1Q6sUVXCzEhlqV49Va6
kI+HED3lhAuqnaD17r4YpVOcH6rbfdngtc4OVhKJRueGopWCcY1BdRn4MX6sjFtSsjj70cUAnCqY
GqIM3wI1JKYtcrT7n3lb+g/4OEK0Mmw1hm9VuyMvwr6e7uiSnUFq1Up863KPr7I7OHqjPefSNc1I
kJpq/L876/rRqcMkNcHFtf1KtSRwCxVeyCP3JobaE9hMu7dYZXqZhvR+jpI2tiBkBm+M+9/sFbLJ
6ps9OKJfeb8jqEeEiczHIHcBKMNrBzoaG6OoPXNICD/sLaU4+I63/7bHSi31XzJxCL7Bh7OK8ZNQ
nCwrtt1FOdD9g57g6Jj6hQeK5fQwy/ECQtm3RITEku6WPW5FkQA4ow1jWyZ+gFqO0AWRxjyqdhJh
TrvtyIKduvo8czpJJQwP1DdiAAleXaM21cizn1hbuIXZzqE9EoV8BOSCj6IXeoJu3NyAk/7gNN98
L11vVR1KczFzqG8mpAHnPEnfGfMC2yAISnaj/ICpEPAoJHY00efhT3RkhglVDWaBpt07qD1Zpm/R
u5/cwaWgNh/bvn/4gfUKlDfRHpl5d8IceQhWyZZysBMX+SnxlA9B85Ko6TmQrrxyrajWmC/l4SAi
tMbzeSbdkvGaeHVHFpvcfri/QPLauX4UeTELix32j2WPDT0jtPnFLgtMBpm5tqIL/5exFDrvAyDq
V2PPM58ggayv7h7C8MIMsSPksnxkmWkpR+GGAYQIj2snxuEckxhk6T+H9+M+ZAW9tb8hDEqSjC3R
YE9w60xqxeoAMIhBhMom1QkROazfPNwtbtgEveB3W09XOLpnpbpkSaV/PW9+sciPI4kANvzPjnbG
H5RBvwa38ucuMorW5mP640Mx1SlqhmDXk97Ap5isv7rES2xgOWCIX1CmbKTTSxD2aHOLlLiqx3Lq
1hSGy8Nchg6PYydpDDRjyXQSxCeUBaDYIuNrtwo2vm4+sf3DVxkyH5zRkb8g/QrXFXMWN3kGzA2N
r191jdKxLyRnhR8WAyYBAdCL8BNsGux8bsxb0pAbR1RUVeM3ku2BmcYwtnPsxuZMB0sjA5Y3PgNW
hxfqqJ9btrQ0AffaC3g2G4xhNSIOJjrjmF3HjeGijMFMRw6zjeU598hkY4nUhBRtAp4S1jBrjnHr
0+r3rkivyfxdLEnjrGKdnD0xexQhe627Lsd+VSDQaB7ZdPUTyb158batVlK/Xv2oh2/59GIigrOi
wMkGMzse7KZ+yESTejiNzluOKYY5Y9jpsmTuPacOK6KM1haass+hjLN59+5robZ65VtOB/fS0XXA
RKPyyLzgHBZckXyRwigilRi6UfTeJeAnVhA3m7Qjv9Bbo5gHp6hJfo/RMYh8PI9MS6sVkPeNJz7u
6JId/6NBraMTa+uFyFHoeMigzQXKcZygSVq57Z1p28gbArKwmFxMUc+ksSt7dowJjsQsTetWRIRf
WKKTGqXdJ79tW6BdwgN0IkxG5GrGPfdPpnKDVMnjIjrR0bks2oewzwwyR0HTJfr6njFOXdMf4uwX
jFWKUIJ+DseHqnZzdygMwYPJzsRAyKkSmS0F4hQhlkJYG5qQWPlwf4zAowjfDrWyUQLZUqTTcZnH
sAcw7eUeXF1zf4j180+x/lTBJ7Cmijxf8M56OSyuXf0jD3qYkT0L/AhLID2C0g7SB+VVOUmdX26G
WI/YSaffdBHBRfDXG872tkxpxcTJBYpfZBWqn3TdsNalVnq6BaAzL1QX7n1WaBiwYJclBSH1QlRg
geEVsArrhqjgEnwAqQd/1Zgxx6nr1povMcZ4mnGx3OJTmEPW9LR3vm/vGIFGSmW9biXlHfu7hjs2
wOqq3N65a04jM1lfKniOryfBY0/udmgIKQ6nLYU1fl4mr0Y9qaxeRlCUVUkFVYsV+oF4H1nHN2mX
WLsTHLhIumI1V5q8Fd434zFzPo4ClkGMCe3dMj1G8TEMcvQio8dCKMGhj/tu4o96H0mQFvbwKpM1
BpEbc+FI/pRiRt8B6A4p6IEKxBrqqXKz2Cuz1mVqhVqIWkPvmzUbpw+jfBcGtFm2Dg9Mw62F4nMx
aiS1+dZlnTdD4Eh+NGiJj42LwzOlw4zjIM8kanS1W5a8QL9wV/3451KwgszRHjnxYqYwmVYoQ7Mb
TCaXust2TuyWF4Dcq186dlElhwUwlJEnTl4KorAwAJYwJvyO4Lb8BUg4fT4e8lYg23FXMGJ5dkcj
hVnSghmGEcB/i50j0l4+o5mqR2du1AW1e63QHQF8o0sg8O8X8FGkjJswI5WKIFqK8cvwOIRIwv50
lLyqA4aRO399zHSZS0lLVBMcVP+PHs9RG9kvI3QVbRyVg6UXHLUiGzXjb1uNvwYJz0cTIrDyzn6s
kiKpYQ1S4WyxhKtigyu+jAW3RlDBQ5u1Xx9abwIm8nak/R442M+Z3RDRrVoH+vOdIEhPuOKTIBRX
6WJwmcZdnhfjfCRxUBH/O/cuGv7SiwwHtwG357vcZkciuZcXqojvWw1Gelu5+8ubb6Gr+RfruY8M
XvHWWox0qcxejGnBumg9dsV7BIOElDTpiwFvicu1HeCJkqk+/g2PPpWa/sBRGH73sN/u2hYQoAJ5
BFyT1g0QiOpH+Hvdi2JvfldVQt2xqPTap/G3JThaoWjrPJe7Ys0mqUzDpYepusPPujqIQyhMeJDH
esDuFNkJ8bcF4JZizUdyRRZuw9NDPOhmrSRenL6YR37Kz7yDp2W+0yx0LE/Rc+w1AZ8ado3ZLBh9
1N8uzAdDVJnsymkjZiLKOZjlHuRxIFoZJJvuQd0VGFt4n/s4GdqTTe44cTgLzPbiZSU+7/XQjlx6
7ON50ljHUJAl2HNdOmdPsBaJQlCq7l6Us4vkW76RBXLgeRrti4DGHxPXY8AT7hpBjfwVix2U5NEy
LMl++/e9ADvQ2n7h7txh9Uu46LgGWaQdy8v3lUQoBcgAcG8QaK/wZ+S4NW7Jx9MbHExLjgOXD/UQ
UT9tMGb2YpC9DanQW01Ev9AAIdlaupEwbtlLeWl1rzkOERQAtJYQSXElJlQHk/mmdD9nJrAyJy5h
pLdlKB6923NOu7OvK1SYS9gR0ns73aa0TpBGn3Jr6LhD5R9nyX6WlZ5QLeaShauUYx4nA3J2B7Mo
LILd4jZUPTrDirqSl489PlMgoQFXIlNM8XXhJuWh4PafULdtOfYH6G34ZgkPjsv9XYFY5INZhGbU
FPAdD6zMvMe84tikcufuQRcvcGxA9+7KHSb3JOpBwByj01KtNswTlIeCVjsp6Z2FfTZsNtcLw7IU
iDVPjVbgPOjJ0F5xcuYobU5Tfy+dc0qQu3JKh6y6Z33Z483xAPwz9aq78kiasUVKVo9kXyXVbqDy
DOSs6n5mLJijpEYI52/+jhkaZ6LGRxQ9FUpdzrGQVDWcOtGmEeYGwXVxdO375Ef8vJPmHVUEl1W8
skzfVgT2/MzjJDyX92R7nkVtMhfzRUri9AWfqNukTaC+Rt61QSB3oK7ljJITnvca8Is6Vv7HZ1m1
tJ0oNYN/pSG+FNpgFX2R9FBewHgaItiqnftOUC0brkEle75Q1DqZUidmSjt4rL00mFYHUhDeHZWh
mloJaOt+Z3KEZPnt3U7IYtuMcNslGAEXnJ2dWv5uzSpgl4C2Vag0N+5yTWbW81uvNBoVa7GWOaVI
3d+PzWdNEkHHMdIilGl7oy9q9WYnjY7Jqnbvc8Fph8LCjM0OhNddlXRlMTGMYx9JSP9lqNsP9YBs
wS71jJynISVf7HwWsnaBXSa6rjYj6kl2UYNMCNGStacsqKENZiS6vDpvJp9F4R+jnO/BVVbUUhpd
lans5mgqvpQeDTLtkS/ARnhEKmlTEcoiG8KMPfRYVbEkrBP+gu0NkdChgwkSc+v3u+X9+mWKv74O
0mDszqIjv+2xhPBZ4vfCaNvTDN/6au+1niCexd/1tQCTEzEgqYDGWFOyhJujU3hkFiW44Bh8rx77
5cqZZUo5bm3EFVc9cvP5Y4WfzE5Hg8mPK6AhLTO+RGqL/Oxj2sQXCLReSg6FqI67QRxbH8A4mb69
8m9tqiLCtCmQs/i6/YsVsGoBgzPpTCkZUPyEX5Kx6n8KVj8180h5q8vcgBaRL9p0mBD1s9ikTaYx
NOlCcrZu31tIlWrzkJ3Ou7iOiEQI7uEeCmAKB+vv1virYpC++117T77xKT1uGniEmlcmlYeElHzJ
ZqvrfJNML/TfJ4PPKQwJdp1hEluX/O6bDWsKop888urTdZU11msNpr8uDuJwwtusPPcS1UD0hdvY
itBHoK/Dg7VXP/plPbZEOUGLw1cYSdV5H3qYXspPLKqkH4CB6OWJyHHw3TUlCzyDFDjBluyT1ivM
elFA4DVRnrMuvdaYCAmDCQlNxSh+s6Pn0hLKNpNzTAvDhJHpNalwMaEXoRAcZFM687mci26M5g8D
lSokgPOxJ+2uFn1TEaHl2TiI1D4RByf4DRF1hdUyvm2v8wzmt+NoUhIL3Ke8Wvb3GomJSj2OFVc0
qjDO2iijRkR0dophBr70mkSw64YNvi/eHkAuGtpiX8q84YzbUxtJapb49Hl+hJ1YoSTKvguq3sxW
g3goo1/PihwCqZHi4IZHf3KErIFQ5viT+88fnhKLxMl6Yd5W2Ihc8eZRZQ42h+kLPaIgi0lkF3fj
rPuM5M8BZeii+8qaAeJqlMXQ6lfnfcAS2O7wUhWsMxEp4weN4kqDr1U/+PmoH0DfDPqE7ewHnqZ2
FSEqQscvfC9sotBH0n7lhDdR2BgeB6CMkT3fhf27G5fn76fE2mVYpbetsG/5mwia2Rp8NDdVrKJZ
4phTWl3ZrmXScRGY7XCkoGPCPWQ2ASq4fDoMW4G2LIrQC+prtyWeviwJwn4+jzmpuuwhNP9N+Zfd
w1XXcKBWQ+U1iXyxdkzyw+4J6k0iG8nQ6IrcRYKmIi0nl0bZm3YJHS97eS9IWRjl+ZPXPaBMoFgM
1THEtn0Dh9XEFrWTp5HNWmZpGbic5KSHoPx29Y8mm6ansK1Ue3RE7c0PtRHo+4//hoNZaV2ATHmE
Ip7/dLnw5P3tzJJwMa8P5Eng6AfIeL9w7lqB+kka9d32RSk2A185KI6WgeqrCw9Cp439sNVqX0wX
+OPAiM98buKvOiAkPa0Avk5+mEi5p4d3LB/WrGpyJoo314zoGVwXGaRLcSiNq5F0RwA4jQVGf+hN
L66qmztTvCDEwDQRzMN7aQoJhNgWd9EbIV3C7cV2F8Itdzj683g/i1dOuxZvtv3gjfRvLv2CJixi
eDeQBonFQjHXswctTToeuz3ayo7o3zfgDBGoxfD/fG786SujKV0ASab/nvllYbFus8dX2f/bTY7V
0IbpRDYvEXl8Sg2pFWZpdzFSmuUNbAEAeHMixMwJ0uDJ4DPJWs9WpUbQd2fvtfrs4yyrvXR7s2tg
Yg/jdfg4i95Dnuu2vx8VaHyJfRyE8WvZZ6CS7SXaW+J9PO5LSpHrxlZfjttfQqIVCKGL80hA8XDQ
jQldgSzHLcMB4cMOJ3cySELv08fRnpaxcH31unKfBbI615ifsAzJucyTMezrdWj9gFXdHTSJHmdT
HgGUjmB97MEcmPvqS4zYgOzhYVkZaXmr0k2Auw13PcDWxpdMG4euLI6F9HbO8zm7yPVQVRgRNThh
gmDZHs/h0nQoaSgsu0xzBzQCmEFR4EtL+LsZkOqMoWwp1uN+9VHZrq7kc8HMROEDEOZR0/7lJHwi
Tst9ATlbBQh02pjCXNfpl8H5F4R7kUsgpgqDv6j30GAoLn6qPu02cw0z3sS5z4AAQjjYixGovPyi
52I2/b2yVJLDxLrbJcYG2vyJV0w8LOHvjTuy2/N+Nx9Q0oO3L/BXZWb3uRR+WH1JJ6a4DPj8z1Uk
McOBACVfnQqlLfUpQ09vHToM3QQyj3W6Y046+tjHV/Q7P7082yYG5ph78rMz9kTlHVpS6ls3bNEN
dcPxe5KR8ZsVr32JtsRQ2z1onNlPm33qb4NjD15PdUFLpwkWLvDqEQhwu1AZ1ouH9JApy22B6C3M
QuneW3ZN5BycChjRmU9Dx+NBBddp2VJUbTANE7lt3GPwjYInt0eCSK0ib/REH15sn68dl74HobGZ
yalv83qzfVeYvqthtLnAIMb8OMFARCyW4gTl+3EPoXm75CL6mLyL24o9qCIbD7tptdmu3w+a7nA9
hFSHSFrnY8MtWMHH1S1EJs1566d5DPB1AgtoRtm4hjLFvGxUNYyAkUl+zAJpaRrlkBcFcj8v/A4A
n+T4tso0cuYP9bYVA+hTKXSbBdD30jhVBdhgbKapiqY1ufN+rYbPdocH+Lk2m/BwAt/AQgz+ej73
H8rdhnavom3xoV74dUvsRhagw580AvCZ8a3X6mvRww7q8wyT3mEhlic/2UGApTmxkUjmIXa7RsAp
tUhUT0TD14icz96tTQNzWyRY4fibVP8vfML+uHMG0PQW+wR2XqhO1SNxXlT0jLzPmifEKL7dK7XV
eekFo6BWYoAj+Icpd0L7ClRAvFMnosGgqOIwzj3NwwsDL8e9xGG2BgfN81Nh0dD3WXfLRGdFRb4o
XtfYXHGfykc+43NKMetdlXol6IMIsvLANywASRTeqFUpBF7J5B08GYxKUqdaBIJP29olfc1kX03G
E6zb6RjK0cDZA0Co6I7bknWYigf0H2gQbKpyQKhX0r93knKGvgKnnO8QEP6tHPcaEQfVJ0HeF05Z
Mz1oiBOko97KEYyapyu36AIcTCJjoDLNe3W/paBquEyx/D+M44EV/Rg7L0/s+ptfuWPgy4js8ImS
qFqZzvYrkWd3pVgSLK03O5Ap0F3NO4n+EanvjTPWeHF1YBYIkVX4ZfaZUw7ZXSHbdH/nhqoG+e51
Ady0de6aLmc8ZMfyQA7BWMpIWlA3unCJnRT6X55EGg8Z+Z31D22hZ3CcuvzmoJ4S6x8RKmmWU3fs
okMTZtefmG53LhIbFV1qevSOJkQDk/A/b7kzplimxhSeekFKruYH+5CW6nJHxJ9Cergck592Gz0x
f5k+fjJpNnrlMbgGfDQ6J0RHdcHB7dEIyCNZCelvNWxxNO7klHhlmlOCXssKq/sKSIhxAL6MSkd7
39jrhMPjENI3EXAbUbTpmB4C2ac8Dhdk4sJhzRAhMvIxje5WnaooV5eP1rUt+hBSp5Qu5Juamq2c
m+9pvoFl3vfzO/xNCHfvMZSoiMN3C2Z8ePHaGpJ8uTeJewsvnyu5nHG7JMGDBCndbiOldtFBh3j4
u+zY/ItLyx5cY29l5Qvp9TbGsAyknN32Y5cD/h7ol/cv5OLlpuD+bf/fXlNZDrUfw9xrimCxGe12
c9XXMkeXruXvIfCf/QNUctbxKKD0lYjFAbbIRtKYIEI/mF3B8AB3r8+GRcwJhJCg8Ex0hN4ZsPvW
lo/V6kotRKExgBbNKlPHvbb7lXWkDUMQZHXckW2CJ9FaD12KsHOCkJ6zcQqhQpL2NA5aNdg7hWrw
HF/AXFVo4cJo6w28baM7yxLp1oCGuY3jRzsYyAG1XRx2f3JEjadjZ2nVNsnCKnmCcWC/b6AHprse
OHN42mI/lcmaGNL3rks9mAbfi07MKq92QJbbq2112LtLa4SUAQ+Df8VCH0kJTaOp8U2n/vL6Ac0R
DTFELEDZusZPho0fiiF+sw1CKRdwLhNPQlN58qRSVsYxDDh93eM1wawsx5hVDlNpcu/8WoRWxnKh
a3FPq/3VdGh04dKlcwU2hSXGC/hv5xhZVs8We+gsQhqAB06PDwWI6IdHWKjlFt6DrMFXb1WNgnE8
6Ju5FY3OI9j/oSPH/G1rNPCEREEgyoYPPwz/Qba4IyPi73oVGeqwdFgpBzpj0pFbf+0v9j3mmhi9
kxKyPM1u015iSn8xSbPyB0DyG6W2Yymp1ir+DGGhyrThEMdptNRq1ZWlLMLgZjjXPle/EkpoUuPi
iZVVVW10E8vOl7Zd+Hh/VAFJBPQ4RPSHp17iVBKJTUfdEO5Ee36FptkPC9WOMQ3n9HGjkcoN8Ng5
TmKVNNseKh35tYc4Mf1hn51WrhPMcTYx0kqpPLst6Piditk8OuLgppCfbtqBHL3H3pm7wdvL7VQL
ifDyKuy54zvnB0c4vEYsNbIb2+kbdxkREwR6fwx4msXk9yPtvkAe4PHSOnUseJYybIy22BsrQ1TZ
pPYhsK7fcy3DUW+6IlMtTzsygiHq8zUxnreS7TQQocGnKsiCGGFAuIhJWp30VmPvbRAmOifupfJD
jNMJy68c2yFyHxCtXgnx1YBogwXOB4xNStr3jA7o94r25zoHayRCcRbTKXiD70GIlcB/uXUAyfZb
YPMrAmb9gg9N6owcL8yLtxGww3JIcwwVzW/wH7+/Q3XjRXS4uzejuGY+udg+1I6GlVLOzazsc1+Q
eVJD45ekfXMxWeFH01F8Cjjf5a+rzxTJGPaAL9EFYKlYaF4ZV3H+t5kp/F4pm3u2IR51m0WxNDEZ
uCIE1DU44mqplZ7EepoWOT5sUAdbYu0kE+rDhmN5BWNOCzG96q3McuF87Ws/NCxKkvS6nrwPzsJC
onoy+cp0AXoF+ggoemOA0WYc/lYIMHFjvvx38tFAnCeipbxMnuoE472NWovAG2S9NzxRbPK4pViy
hXXXnaSVcmpzhjxW51tBZMJ6XdRfoDzj/kQ5pW82Z0W6S3TpgwL1U0wqejGNAZUwlO1J1yqYOOD0
0ABdvfzt9+BYJTT/b7WSMWzBxUBL34dhvraKikItCZ8UtvykP0tlt0Gme673f3PFDgAihh2TwRc7
c8Kpp+W3oEVeE7M3/9HFXBowap2ymWtpzVvJjWRymKqC1Bn26/vobImQUtspZnOggq57GqO+VuIl
osvscGRkSFD2h6OajZ+wycMZjpCtYIvCXK5h5yh04SXCZwI5J91FrGDK2g3SJ00CLBqwxo2Wyyo4
PCDC78CwBbxDbrhsFtEG1gK25v5Q/wAuLbaip98LBSU8SRDS7zAsWewxyW54sp4tP+f0SR9iMeAo
t8nJSMDQ+DAjDMoJu5vSLJ6HuGYbS3vdVr2TuvA9q3fG02BdFlF+XrwYZzaBKK5uGAmz/iDItU5u
QVASnB87J+EJvzWn2u9/o+ObhJTFk6Szl4RxH5zShc785q/XHya5zcqn5qYI8pLeSXFyWQyyvIpB
Qb6AssKFWC43IZ6Y/Zu3iwhQZCkD6wMM/frArlc/jGJjJPtmqUBP7uFHqpYBARSR/Mz6y7tbpPgy
QI26zALmpkHTf0QvwgCtJlwHXpvS2ekIiSZZPuglyS/Z/pEPjAOUHtQekWqsmChQWr3V/VL34uZ9
XOVrxfd8xZ39/Ds0GYbqB82Y6xn0C0s/QmlcBUrsG4jFycWMj6qSAbUeEcLj6nISTuYUaz6QGcpo
v202rEBPxmCYdAYmIL5VFJv8OaH1n04QsDvrF78vsNBhI9RS6ZnKOTl6wIn8P/sXkaUzqCVoUWfh
95rLN4jO59TtfLcSlo9ejfq+MckiQlvLk5tvMkYMUNg9ff7+/GJKC8VN72EXmp26Dv2YEeBGJ4V8
mH3wFKmG1Su2VByNWjSia5OGl4EHHbGWwTEfflnCZ6AVnAb++SSyclKvw9Ei3sL+L2Lyi0KESa0j
lkGJp2AlIdb8L2hcYce9oMkbqkyURUgFCV3tN/TNdx8ZiOMkM6xnUb/PQUxQzhjHXXhHEbneamH/
q6nxUyxtQEB4L6KhV6JQzzlLtwEa1fQdZklZqYmw4lmNpeCIoUs+q0zTyjExkWgFsBusLborih3T
HSZ7TdkUqBHsV8vmQiEtanYPzz83RHK+wH3eDDZGBZrLyWLdpOF0mPTcn3R38EYQggjzT9kfTuP/
/JKlp/xDYJz5BTsqJydHastanmX8n3/kzErp+hpgg32Ti3bcVNKR4ZKytlZr++cFFTVmXxnzNYIx
0MIqMz220ZprOJXd93NIM+EdpKm7JLdoeLmhqSqXcalMVcxsSs5+ROLsHQf1BkH32bstV5FKrfXs
8wO+vRyXXCWi92gfq1JrGTCCPCtLia+rf+OUwGnt6siUFLfTYuLPaDFwildYNqZXjQN8UUgyTbUU
RhUtNEqApnml52AjbQCZWDG5p6cqtUuZpc3CT0hsy1I1SqLAcl9JlcOaSeJshTts3NJ3zM/eZKeQ
Pua3cAAvSUB4gqFdB9VwitfYkqEiNnqrnrghjGeOLQQYKE3ML4YEdIEVcVvqm21w6r4Y7M8UyNa8
B4W1H22cK1Z5v04sL2e0F18JMGL3vai/3CgLVjo5Qi9m4X/xce2BMUgnB5GuanwQetneW+gY1Dti
595ZviWvdY5vithWQUyIdIUVr08lv7YSWzWb2didgz8UT4+5+mOdVnfs5R+Dzt+PCAyX2ks3BAT3
dPTO6MWVROmJZH8Jks92wI/x1RYXy9MkrIPRXiT2kvFP4lSZ5PPigKRHKFFYq9gFcpVgRiGrTH8L
iqFhtwy9er6zva17BwcysjlRH7t1OqhhNynxrgcZbfUfoqT1rPdMTkSEocw4sEY/H6wF+TjwFoOh
PTnZdZVew7qWJI+cVsq5UbCU2NZSJk9vg6rNxT7gJuSdrRjw2JBKpUBpTRV6oAsyV+ex+5YVeEKr
r+r25LrkYNgMBPF+wKvdCW/HHRco+GcznfYgKNXRWuyok5f4aW2POKI3EwATc26kaNLmO0nADe50
ivSYxy7/HkTfzRYOCAAikRSsF62oy1Dof6N0BoyysaUyqVzsJPZRovUudxvID2D2W8yxUnbtrR1x
oRQl7uyU62z5qWAf3hRdsLBmMWxy4wPMGDJk5im40J5dTHGYQ/KmNLCBsp1MpWQdAoBpt/EU0fFK
sAs0r/L0TpRuuspB4dabVpgWhiCXBEaoQYnCiwAJ4lOVtN+8jokzF1NRTV5K+2iNup0dTDTB8DZ7
xoj+WSt4kgxpjAnRCrauRa5xJqOkHKf3qOKaXXtkxtnxsnyJlt5ELi7yrq8CwoOWZWed56d+OrYr
tzBCFut3CvQesBqKCiygwIOoY2C1XbYnFIBgvgk4IFHIPQ/00feBnFxpxnGbuts83aTYh7BXvuWQ
UPDu0sUgDzEoXonFpPk6v0MChl+mHSLcMvL2GklvKcdc0/FGs6hyz6/o07BL98TvkiUCSrCeZhMa
qhiobQwKbsUCUq1jnl3YCkwUC+ylVaAD2bEhBQORdAFVB6JX0w7YKCDQzLiTw0Ti+6Q/+N2h2JT+
7pA2UfwwTRsnRB5b1wPqkAkOok0q5wWt5qIKEIzQuKVtQPUzRQ+r5bLIhTHmIbuYyCYJehV4X7dH
ahYXGjw4z81aple+9hKNVcRzwF7w/5O+hYL2u3TDUOvCU+P6+qVm0kOQvN7u5vqp3RDZkLVB5LfM
lm+QYyIUezT7aZ4BWmdcUIUdW/0kSjMZiWVgCKPjDygW+aYJoEZTb1QMFIkTLi6sm6vUmbaWJX0T
w7NrYpKMoKSMuGf7DMoA1Pf6d63gg2MIOzhoNJXVvi8KurBf0RvLgifwhlIXfxA+unqS4SahAA27
8pqAIh2lH27KWFDmsflt5A95ly6n/hvK7GOms9oy6fPmrgLOkIOzOxFd69NFT7nrF6OAFQhM14Z9
4SYv8APtsrHdf3CnovpNmW6mkvxkE1H4FxHwgPBnYLtHeeCqP5pU0AgBqYuTfx5FSRYdydL5P6VZ
VGDoMkqt4rJwt5e0bdqjCqJfmbyVInd5qHZU87X7YbpXx56CGheebeaHL4/MkFh7ZSVW1x0Aek83
fPTM0ObEqNZ+6dx9Nk1fD30G5V800EI9dSs8DXzWSSWYxDiIPQ8h8vJkzHfzo2/kupIcbzm3K1lV
PUXFCaXB844hpPLa/EoQ/yI+X/5HQpHqndRuAEdGijNLO29yvMVPZtNbNFASU60c9xblzak47ULe
y4E1HaOovXIjPDQbIDtrE49k0iPLoaRFFOYIVMC7+vd8OyxlgN0IHPFrnqKPYw4HCwE84YiCHoZF
IN//NWXQeaw5mrrp6+5RcbXTaqmTzhIBvA/+3BV0BUzbiPp2fWHD7A/MwH/HLH1rg7vXNfZVNFOA
7NyH1ShWLWmKKA/LDjgU4PyreTr2ZbY9XiE7WwG4dN3XCcZ/E4V5UEXdHY6iKk7rd2DdnL4D2fBN
PLWPXLll8wnSXKceEgeVAU7vZzQOjaggVCM8f2DL9jJg61h4wEAim6qIyhhBGsnRqyvSai2okuUv
A1qKCk45iFsoQj20bo9VCMeM+TOq9YmpSOUvuM9hmnUoz7PaLJmZaDFk7hZtb1Ys+CxEIxPOuPSL
OeGyvVS/VUtRisNxGkprvtAfBEK+yVFQU85aP8x+M0aJNFyHnhM0bdjRVL+l8rNUvZaD2aC9ayEM
1x2oA5tZaAFvK81CQzaPnpCG1fnYAXOc1CVMn9mJGBtSSrGxtU4Scv+lSscRf0FQUFUmHUqr1oZ9
YdXrv+779iGJ6Eg6wsv/Kpgo2crPHuhgBims7/alFK4M9jroVsIMFm0EWYCY+TjLzvnOEimuAYFe
JhxYv+xUqcbjW0W/k3KvagiY4LQZgR/WhCZ/RB3oMpx7o8E864sGwnra6vWoiZFGbDwMwOlr8Hru
uClHMod6zPeuNTj1/t3NDId7jNT6k2ZV6gZVr4yKOSHAsejXDMMNqMxc/zAaxcsai67P0F0YRpE5
pIE7zL3mLEz0tSPYHwEbs/G5Dr/UTxw/JK/tMQkf4PRoqkN5gD1mw8XZwm1Fyg1tF5ypKVA/xcah
T6knmH71OVoUDeFyrA2K9laFE16B7ipQ/mWAkJbW7o7xSFs9WSl5DOLqZqViFrzoMiVV8+bMvn5T
liRsAKETZYcv8d/cPd3NORuUr4fp3VCpapbX6VKsxNWqO7QQvxEJ4PMS2hUGiTXceZ/4e0K6aMDU
5mpk6oXZKIbSg6a5tfdCONW6B0R/Di/B5dTZGyCeHqN1gsOk9qSOGlCT0xZUxnLrfWGVnXh8x+nK
Vo2FheNOFlyB79W2dms1tPSQTJpRVl4gq9BqanuHMc0PmbPOsVdzX/p4ltWDO9z/lNlN8ugr9ANR
iphI5jHKRbXFxLJ4QXLue0H7kgWkJjyXLTSfvVXiPeqz6Glk0CLxAC537e518kCfHPx+2UspUpiN
kwomcN8MaRFuLeewrwGJa3nSloMPYFmwCHtpG4sb7qKBb4c2LB8q9pEFjhCEHrwgJVlIwTA6406x
tEbAwZSU2u7Nx9IA5omMmwWXaBqJnKaRJwEG54mQLKkZ49eZWvU9JgMeJUQ/+kXlpf21Ct9AO6T7
VHQcoyRSY4YYXql2jcBRlKLuDvz+HUa5Xq6kMhr8aDkzou6QFXuoHAyUe1KUUAcAWBrRhLParhEQ
4qQj/jFiTNWU6y4fWbf/Wp3/5kucJ5Tf6QFafeFG5H9HmNxwB0j4q8dy6xPunZaPYHfe61fcvfuC
1Z5R+wBS3xOpA98FA5oLqdqWuRH/UWzhNvGIh6vbPIpowf7nL0vNORMR/ORg5+iEg/j9NWhs11Ca
y/JZcGEWElzaA5+jHBx7kkSXocTh0T0mVemheubRMuMY5qML0+85lWpNqXXDYCFY3DtdTAOi5LTo
R/T2gLVQljrGPJVix8hSPhfbnWHte2XEeQ5cxgUkNtzo2rbyiWYeVhC6+zfrfbcxsZiKZxBdD8Jo
UJ9aY8ooYHSnrJLPhL1T6MXS6nGgx/K+/zzgj3X+Oq4OlgUA71i6fX96k38SOLVNuquBqlTUQkL7
8aDh6ubGI2bfIAERm4h9A+oH8HuTh9INEFODbfTVHtM3IAPPglXDuh1ipQo7qgJLKwnzmuOlBEXg
Dd6TKXhuRW6e/lDUd2ABqbrwsmRDrtlmkogJHWrzmvYdcIMUlZ+pxBSc6ruzL4vRVDSNhLYgWX0F
LVfWrFMtMu+gDBbc4p8B4+DhFlwLNXUJ92Nuesm1dsNJArgwAn0cJOCJm9TIxc+TF+bDaqGLxSPx
ZVlhXlAeY5C5hOcJpJH0fYRuD3py295eTJt49ixbECAE61ts4DPLuJQE+sjakDEF0S6gsekILwGG
f20WrLfub2FWq+tSjwVAV12q0Ab9W0jMcSxo8Pqt0Yl1akwDmSMwRkyA20fCEPqr3GGGfTE/NlSx
c714oRplFEk4tqoUY1C9r2tuU9abl4MQRIg3/HB1zxRuTIgFF5Du0bB/W9pJkQb5P7FyuNF6Jn7q
2Nb/B+geWUv9hmnyEejoELiYDuNZJJiC+/L1icfJM8lGsazt+lBA1TDfOudRiTJq3VNPdAFpXhw4
ETkKiDkdQdL9/1i8gKLre+OvGdAu+ZWeSTTh/MJ1x7kaB/QugGoI0C4S4D+7dcgUOInPTRY5I5Ek
pYj5HfF4EnbckIb7cFpJfjPv+7uI2a/fmYZjrcmxoovuPFly1pbGjzfjS0FfZltpavOjqluYW5SK
7IpgTmRxcztJSz6JdG7T2e7XfektN1V3A9K5k3BrkV5YTBEq7KVZlVtHIMwsu67ksWavlEY2K4F/
JekLnC9lTJN9k+SfFSOrWFsceyWU3eSas5TBi4toQajBCuB8S9X2135Y4XSHGOkcCaATQtKsfELA
yggEb6uNB11eC4yFs64tAGp5aiyUY792OUmCigdn+Zi3JFUsjP35iANkJytFL5YmksUOY5Zad4nG
vRWnXoaMcEs8bJ3tlGh/fdlamBn6To5YuodCQlE09411Vu2ewNRPtPRmLFASgknx+BKFj0V1dRqe
8v93BrNLqw1WrAdLnA4nbb3tQjnpditicQYGeAv1lcya0tVPN2JXnUNlyAHcxLEZ8UJFN7sD4C6V
hNtddCANM0aQM3MDsGCiM0tllZ9xTU4dGR/zwn9FaMZY5YkTR1+AFGjSfb6Mc3dT5dTA7Y8hHagO
2XE6rWWyiS8Kgmp0lgo10CkPHpyGw3IWFyHlCKClCmmmVI+b7P0jAtT4PNiD4NqMvPSvZDpCZlDm
nts4rFts1kIrnFCR+sCf9iXzLo5wwP/vWBsLLPc7hp+7ccwIizKhlxc2x17sDsmuAX19A8ZXiLMV
xyoTkF2WMfhQHIBd0lcoMgPKsJu01Kb99R3PY7jPeDbAHpA9hPdixJjgADTqaSBftvGX26pDeqBa
d7wjifg7T99ZsqoSNfrry3A+xyGKZZU9PTww2OBTz7p4pexiI4QRToqiq8bzaTjBcrojcRr+uVDh
7g4EMSrRlSRQ9b7a6/5DPPI3pbAM1NBBjIr6cXEbylrTN69It6lZbksjlpLn7hBYzXaK3FMPFIhe
vMuRJhjynmD24yu+ji5vHYzoJPrViIXLn4ngjWocNQGIdTR6bKh4NXz6ZHs+VTWMZ23mgNwtI+Vi
JHs+RmkcbJCbTcmDyDmyJhFflu6h/0RImx1gxAQ9O5q6M055d9WX9KCMcRsQKpXmmHYkU3Hr+8Cg
eOK/nvc+bNiBn5pfGe+4aBXR5OmZddRIq3JG/yXKTBf+r8gsxdx9gc7lwAXVMc12DlLs4MyuQwCz
RJFee3MPyglUghe757qYLFvoKsr+IaWbrzGrEZr6MIVSQKKqL9PfOSxatitWDRkPMYSRr/ov7nes
vIvMWDuTNTsSnUs93WWaXD3MILA+VIAjCZWpe/696JNL5oPSiKPOdZ94oXy0PVqT7HJEz3z3gh+F
RwXva2PB36iPVd2O5MoI+IyRbTXY0uH7pWobs8UH5qkQTz5JZ9Mg/RdiBxRY9ICk2IITVt/mnqMR
DZ4sHf/qJIA1Vs7Uopc7i3kq4u12QkxGF5qkCGJvsiDA4GE8tsDTXU4Ro4ggKkEQCzkFTSax35FS
FB8F4sLzQz+JlRowppD1A3C63xq7x8XKZMRtSAO941RazsjIA9gTL6vfc97Z3ES9do6/d9lnAe20
7rPKYBa7ziozMHzUzQKwDmFdQZtRVy1P8pvHq4tqH5nc8okSBe7S6Nn1mAmYQGQoo4CQ9gSRo9Pk
o73rYcTSQYeuz0wOx99MnPucLZsu4L5rY0M86uG9zLrNnYyvjDrxsuXxoAGsvexfwgxF8DxVMsPH
BMu1r972EJV7cloCRpdFruW3+gHooau6jjZqwCsllpnqLEG0pKKzRwgk+x3mp4mnrIsv4zINVE3G
GKWlhMEVdunNAE4a01qDY1Kh1uFmVhzh7aiZ1STwH0+MvJ4D3mBxp5wp/Ma/gbKp0WOrp9SVkr3I
FOw9AA6Xtig/rfbzKWbLQHZEh/Ofaf9suSQt7XpMV+RxO7fiAMMT3WuHkyqPwf6ha3Vxt+Uv4hxl
EBe0Ek81sVkk9hjMSvRJroVK2ThtWTO3uUZAzHt6SU68k6S7VXQ2qngfI1prSAUHRhDKVY0+ytiv
bS6W5h7cGXX/ShUALsFH1fwnCMkT02XOwfAJl7NJo7UpKWeKraBewwmcpqKLUge4SVUlkyrELTSc
0MBxnC3WI88u+xtkzBqDqkTzNW98dAZAaTxBs2rH88xvdmS5t43McFDR+nCTWt+5pZfWzt7X/QQx
G6sbNhJ0lKp+MhjdS/TsQkQ+aWNFzilP0fi8PZu+r4fUQuU9jeW/THzPAkMCd/hltX3SOACva1ks
hVxxkz3PMUtvcG1V3cj/9c7EN/VXGEOFAlb0rfU0iX69F2T4YJM/LMB0yzq51/b1ezqoXi9qN9JQ
KMMu58cvrr0N3cZKmRTICwHlxiXGyjGUq13iL35+H4KDlnmQRJnm4PxTEWWyoVkvP7KFqcJFnbl6
vPngx+ujDfDbrI+VOxQVFGApMdq62Iur57QOup8raamONM598BvT8ipk3anI659Y5MoJ57TlQm1w
g81B62NhaxTIJyJEzAfuYaLaCaLUlR1LrQCTw7flqrgwzQd6UIGBdy3K/QGYT4tWXZgWDECy1mDH
pJ609s0wh74KccLuJ63z3T8REGrf9lL36fxINsT2ccLx6yPnvuplghY3ffmJlZ+VDo7u3PaL1q6y
vvhHWAm9SiW9JxEz5xYwsA1HbuqkIBVGAFSq0wcMuptFuE2E0KuFAj3cGcqklByFIeOjBP22Gkp2
3UDjvpRjtCgwa6BvF/ZwWk1AtDAVxMDuvBRrH+XhLgBeiDCum7fER4GKUAHmJmVNwsMHGgFt7GBY
X179rpb//AuMgc362wgY+E9DS9KhRH4Hcb6LA4jO1ggdXtGxUJl48zj3I8dz0AypEoxHF3dya8y3
QHP1PpADmNqpRdwkdGp4aBaqIJ+5r4DLeqEzLb7tOMfBUg+uwzwL6vDNWFrO5Z0h2VX7gLdz322U
nbh8ZgDDBRgRNl2UtlgstHzs11Mb341WnTO9aiLLmxdTz2KwZhKWOskGhGwaPIqyhSoE5JCCfBHW
Qmw3hyLfOo/C9COQGVY1a0Ogj2RK+IHY1FeiMuBL/amqlaVbDNkVnJk6m2wXhhmVQp1LZOVx2+1P
b/8DOLR1z/b30EE9PEqM1eYHnwQB3RhpFhnN8wZMM+qk6wOl7QDTMAWQgRmpde24MYMeO9zgxj0t
p0VdlWkQd9RkTdzlHIQlCy9nIfC7SvIjH9mSJTvrHk67IBGX+2OQtWPTFUn6dVsneirOn6VLeM9I
giUSiURcD3FuHYKdUH8WwSQQer1/+nltzyKX9jg+tRRHARCmoRUL+EFT1Ey5jMK9Da4wi/XTYiUc
BQfDvzlIIMA4RKaSNs28qq+40y0RP+PK58m1FxmG3h2egujyu+49X/2pUnz4htVg46MPaHpnAtsZ
Hk0lu577r0IHYDMZ70qyylfg8F6VehNbBO6BcaM+DkcnTa/RmS7ziyl/dkX3kcChFD/lb8z5n52j
u33KmL10KdxXCalWZpvYI6ZLH/g2FwwDExseBl6HAuWvLGmYTFaqGi6LrIfoEeP12r0nBQGkqnl0
R5CojRP+K04G9Xs/tWZev9HK6JZRSchTDLlgUNPLA2uu4ureRq/6XsKcNj/kZ9aq7pQEypqk+P93
9qobOdOERAgjKXAJ9GkoGf0331QawBsry1oesGUgDyFuiHJwSaOGiE2dKw52ijiUnCZpOsqs63mG
W/9PKZmBoLJ9nNlOjK5HbYB6MerG5HiSU+u2sDMRZkIpIlv2LAkoT6WeP5gwRGJ0kqYFePRewVDK
iOmNPwT0KfoMggD1vCECGZRb9b7+TUzXFB1NlaatsrQ7FYUPGpCykUz6x+ZBTMx9NLAyRaEvCijr
D3d4zszju53m82QogUnghk9zODNGWNLg5/8VHHWlLM/P6LCAS7b62bJTpL7MDJt0PKuxgLU3pLog
bqEsN5LWxPffwAaA3pR6Eo1g/nVBeDhOsw/KRvSHSxcQ0tGAl2zIUr3NIJaJft85Kj4szUoshv+q
YZ07WHMf2rHXtHDUqYHL0YiOIHfSwiNee5KdHLgMMXsmc01tgHyEQsFadAZWm0PWW/AvGt4NrwJV
CM8ov0LptXFXYCTwCRKOG3O4HNJDwF1VSQfSrHeuVOe4YxJB0T3PqYl8mji65pUtpNqMnUszxzqa
s/0XIDEg2kx54BtXiw3r03dKyFeMNArI+xtaZo3oAs3km5haMLXz8ae0uOqRjdxzZnKwj4ZLRbRs
eMMjjW9zab6JZOgkZqsPOKKBZFomVN2mk00/Cg9z2jlUUe+mbUdAH0ovVstPImF+Q44FWpQgNANu
BbAH3/aa9/ByGp/K9lzuHkVv0+aAZwVBmAyWpdnmUToKcLHm7aqm1IyKncGS+o/rqLvzbhRAuGif
QpxkMM7KhCL2iOIiYTLasF7xFbl8yGnsqsh57sEytOPpIDKbedsuaxq4pL5pMcnkN48xLEzOo/F9
EtZy4dexdltc0TGjOjH/e9AQqixGVW98nGSl9gpiaJ4VinG0x6EXootlLjdKsT1YHr9Q6ygDPw40
Wzaj2N11emh4Vkl/txDFSBZEvNQyNPpCEdlbZ16uhe7MVKhqJ3R/DsjgKBnH9YlXvE6J6VS/NnaJ
cerCXJYCZhJpBlTjCaWML+faAO8HDL+DBZIBvBCP8Z6esrRcHh9J3aHHxzw4+nuD0Ey1B8/pIxry
twsXaDZrRbCADWbFAYS1XMpLHkHY3824x0I+XLqiyQ/q/kQ5LTiAj3SMlKKFkMOWWuX8Jvj7rHk8
x5mtL21mZ8mdfvUjHcwKbLgrZtH7hxNrHqsTcVVh+yt+/xobg92KQQZkr9Y9DnxlKvOXxH1vNht9
LlyzhC7ACPQO57RoYn/U8l9M31L02G5WPqJPrTYthkPdUDHQleE0Zfmo08a4BpMdH8MQmtUEkmsY
fyln7KqXnfug+uDIJfVk6VbcUHKa7TWQo9Z17QQgKL8YOFVAMGsOzu2jQ2gR3rv2TU2DPuCpUxHj
xm2QcAfiJe+M59GP4k0FX0mIlpWJJYcnR1oLPJVraM7ti/+gEg8caVvt19JCklDqdsR9LKKtmcX0
oDS5t410JZzz3GTi3AWs7PrerB4aU0k2u9/4ZO1x2cq3yGaW5svRYElp1kfK4cLkc93xdy/8mt+f
u1kRNyhuPfvHLXApSoFZV96vnxc92Kf6LzA3qFddffIWeMgbBGshryl9h8i1IAl5QYpspNLoMvSI
aPAbPdgRdh4NRmmvBDRYKQpz3B6Y/bJIpUWRTjHWtEsPLtbg9uZcH4ybTpkI8fsomtQE5uiFHsSk
GPlxtWwA4RH8YRMoX6F4lNImqdODQ3fgJ2WOXzi+NlhgqJpyyBQsXNJEyUF0fq0xzfSoOM/54Ook
i4o1cAChWrrelHCqxfUAvQiwHJw8Hl5iNQR7AOs36qGET8uIr8I4fX5Dg5rJvY7EAGMcDiHecxSC
vpHuuKrKl9VovMSw7iYNB/Oa4+XeBkrFkyQ6pRVhHiK3nAMWtL8Qd6LcUJcu968vjMQ0YlfQUc9r
dRgIX43ROEtbh2bYUrBZVT2y8ZwRohBxU3DkM1p9g/wFnc+Xf4CppK68B1Pg7bu1tGRFYv89103Z
dYnqi+obqHUOwCNcIbtpE39DoIOHXJtDhKpcIQ+lPz38Q28xiT4gPwd3JiEz62ih9hYh5IV77dgv
6Vt4Qbt7ptbBUsfVDTchy1FKBZh+Qwbu84m29ZE06XZhQ6gaqBKWeDoF/L0pADmwScbFzH7pXUFX
cLwWDnHqkK9D13a1Dj+dY2m/ENR1He2C5cvrnALK33H123RusjASxP6n3hb449a+MfX8+S6TMp6B
YpwG4UrMKBu3dLoAuczcJKVSH8FZcNcPSDD1UbiR85jzKdBIP96D7ru3jgwreEpiJkv+f1Rm9Tfs
SeGniyd/ZnYdV8gOi/8z6QpcIfrjEbbr38Xb3648p6AWnD0QsLcy/J6QZnlHJhbzc78v87UIzc3u
IoAl2HoPg1JjNGfZ6KPRLzY1PaGXXgYUKJdQvjQf4SQ1RNdWQeQQL4Sj0gtbJs94Qa2ukAVrkwbw
Wq3VSnhf7HR4LFXdai37WZ9VNAZvTn2skS3fpqZioRLhF6QBzt9kqZFgXZVS+vY8ia0JJkKVjPKp
Gnfni1xA2GYvEmoX7RJMIst+wL1zQzsZgeY9hdM9LAC2P7HLJMHUJed9NNHNCs+aOmtvDluCABaC
66pWXQ77xW+0jYvvukuWsu6m1gomla5H5bSBaMY0O5JIriWe1/a25Uj+b8Xsn5geN5dE5kPtmrHe
nhyx2nKbGA90tzYUexIGGYNq/chouzowFtIeMzfaCVW0nHL3m9Dv6qAi48KOcDFo7H17sknHAlgC
fBySkb0QQpmOPKLrA1rLAqNOzQKQcsj7nOWbkn6mEpDZNk31aBbsbBBtVshsarBh9wxe57Me1Sbm
z/6K5/SI8O418wQI8/WQsNukfkODW8QFrHgBYQu/J8tVJzUGxNRqXF/SMh+xsgHc9JI2w3o8NH+p
8MrX9ADYyieP1rXRYNhjS6Sx3OB+6hCj8HoPHoillx5hGmhzidiCKBHXhxxI9FzvKyCV3QCNoQy8
1H2BVM20mVmgfrUAlpSkhLGz4wIgxNFmo5VPScqAKQwaddntv+RbEeE2QD85V4Q8HyAsHpeCVoh0
oxwsexteuM8OAHduvfVQbg598RxgXXfL4GncFvAcJqcv+XSAWOTRXbeTMVELBpM8pKb4b5EPj6gy
QrW12BTvV6ecKKNTTJOAw2vi3t1ww96UjNfZU6f/eDC9aTdZY8GR833s2lQWXUaT/UhVEqIrvjZO
zn61Etj8mKoQ+2tk6hOPFiUq4jFse2tSM1c5SqKAqqF966GG/ZdD2GfJ/Ed9Xc+Oi4dcW5Cj9sCQ
OHmGThLRoleiCpOm7DyZEyjhcor9CybMwVWdmLSyPTlyGATXEN/d8SsQtii4QQ3IvDWCTRaUcK1X
6ek157VS9C7hPj9ulNiUZj+BcWGm0wxHJHNtsTYtVsL27cDzmHk09iVZwJA7e5g8dtIuzJ1TnF3L
ghm5BnGLTGHpF/2ANlV4PfPONPJE8mgSPRQ56qncksCbqRvIQv8Nu6sQ5tmXGwg4HQCXzIaKacS0
ZrSq7hj7S1yNDgAgUkfWtoRuloHUOvY2BZ7MC44gHGjJdGgvJoOql/1xs7C6UK+EEflencXfQMi9
rR8dEhDop+XMqb8DkWMQenf2ots1U89emCu2/QPfBEqgrDvhbyjk+02Mdz2qAsI4JXSkNJjq8bpS
JsCJsZ7GF2MFTHOmZeRIlZ/rX7iss5c/b4xTfBD5qXJcOO7FmbnjIgN2xlQh0Qxnb58GBBfcldpC
kZNYFEI9MSH7JBprlngbys377UhYmUHrv6Q4QObhbcgM/lZDORp0ksGqG3at0qgnxQXoOrgxUBht
//E6NvBJIu7UZhnxyy4X68watm2kSslaAfq5BASX4h98S7H/uTMNxebxTUqIhI5Y5BaQnVPqWSYQ
3zwP06HdWr+14qwsT0opfTAz6cx3BMD8hH5228QpVEgSEyg5aEoPmCBmgFk2riiSNMXHj/XSgR7f
0t+ifxfO07innhgAZhMB9FN2ySbjhAF3xp7nm0/Zu0xeFWT3cn+9SH3cwkxktxT8chYb9gaqGOOG
hUkwi1aRcJ/slE1Anxn5/8XCC3JgBooeaOA5+npw9DTLYbsdIxY0+lJVUQaLHV6ZmUAkmTmnLVyr
DePgnSEUWKjwm5y3iZMFYkN9jRCvUwR+zpVa8hF4RJ296lQrCMhwqpaSrYhBuwW6S3LO6KKkMBlq
6NSioWoTiAn5OMPqyjDzRqJhZZiublFo0I/0q9up1Ox8E39HyII032MfM1pRQDdZUJ7HXjRQCqUF
U5tBMcIBJlSUJFrEA06MZz2Wuot3YtokJsREVB5NUtOZlwA2/CXkns2UhWh63YLFPxM1a52/ogy0
JvLVXT0UlelS1Gx7KnWUXKq9Op4v5vXQoq0cAJLre8iG98fzGAjAQgFTp43oPvys2HwiYfg/Lp9i
74ImpLRfWEif4JhWua00ZbbhZE5C7VlaSOUJH42BttJmOpaxudTEVKgp1BqiM2nLNTp/L7zfX7Mf
74BUg85WYZbftPA6UAP8DcazQj8PbZ2AOXD2eN7Ghfa0D10Islv1JlQGkt3N1p6JrTi9iWIWpBjH
N3RiTSb/H2ZuoHbl+o6+/7a+jcVNP8cZqONsrlXwPEfHxPRSnKseDsdElGmONx27mfi3zbnvVVq0
bpptWUakE+bqxpNtUEHqlzotmo9Iq8V/nIkFC24rguzplC3CAUrpgYPPQFtVqHHjvUBGb3EOxwk3
XOTaOFAoJ2Py9zydA5jyulmWtq9loqFluckJXc3zh/Ue2Cf4KIjgCEKpCJOYSFBMDiA6uui6yux6
lbVGBifRfd8IQF27GShR4FfUcDqHZ0NirS9GB0Q7rmx1QCQt6pkSEdNWlOMams3zLJjmqZhhVIh2
dXzMci3VrYECOZE48kNolKr81ge02kVgfGuUSLnvR9ZzJwxDxj3liGvEjgy+4rbyer6Qakv1qynu
8n0BwUkZiP4S54z6vDlcwEhLc2k2EhR1DnJXE8L7+F+VeeGGlXZB43xBMcfSE6uEuRtHeX2ZZj0Y
k1r/dbvFm9DOzkPt3seNi1WMrKaYPAPdufblgeNFJqwkvQsYHeQt4aIey3m+H5XZTSXYdHbvex1B
yZJS9EbdmGRgMU0KApqi9Hs7Dr5/Pak4aWOPu3ZqlGj4hDUNYysM7o3+nEbGDZ9AslEZlhViu+px
3+YjS039M/f+f4DbCbouNe/1ksz56/hJSpeqD9ZqDh0iGEgQMT8Ico6naMwf2c5bwbhv23rptQEj
CwTbRPcPTsABuSU8k7SHfnIEy7x+XqLTqK6vt2HILIX7VV1MvT83CQYAUljWXzHbI1epPHMi2p95
Zto5e7i1HDW0WbeqWdI58CheejVmrqDYKod1vPoKgBEWNCdthKm2ba1no7FUeSLOdXIVqixs/KXg
8jX1J+lMJtk0mTmSEvvxK7BjiVEAaolK2MdebxAhrvSzebOrUQv+P6BaKhOLu1JBlDf53NP4LI/8
iW39v4O8BmsIBvWm2ssns0g+xQBImoBj1j0UTuWNCUVnMcH4rT4H7MFQtNgu+SOgH6dywe94P2D8
5aneJqF1elzuYp1ekDiO+q19EZBVGYcxiH+/lQ2g613TrhEGEbqt+GrPtFVZFaGfExtGqwIyHKXc
P1ey1FTZrbOnPS5iN0AeH//8xHxnTLMCJSRq+gumFFXFMhZi4wdvlgjZ4/UnFytDxsC1hoiBXQTC
zamixWxXx9zmJpcp8s3nNdxMH+9JnPS5xcBdgb6Tnt0KUz+IarSi8gKlL7SSimW0i6li4Ww+5etv
gIin7sAXq7NK+/GirWNngyGvv0FKHHEcKgowzf7zJtkDCpJpFJYMh2bLo+MIcm68QicUlTK7yc86
8Ttc9F51WcBEnTqvCWN97jrY/uV6vExdek4vk3a0+ZuOIThzQfd7Xh7caE5UWctXcLK2zjQiJCkA
lk3V90kkNaFq3VjjU150ZClKkXX4CjSpqotS1LQFH0mlp4VL5tb60jk/RMPooRy0qIfVgsupj/RB
1gjfsvEwR2YBqhweipvgJCRiCfuP6dm37romJRGE0vfZITj2/F0vLX2IBERd79fcBex9MDVVPxue
wZjtBllKL1Zv9khNvnmxg/9f/s2rV0qb/iFt1db6hlbuJdjPwyR/XSBrUPGnKfZUgZl/iUx9cgqO
OHBO7Bp9ak/2XBnW7eVUDhhObGRQAm/hn6BAdh4MgSTDRdY1c+NwQeoymYtt5OPX8AVzqBCtqBMR
yGXAnZE+vjdTNwRet/3BZ8J93fpgRynUrw7dwflJ+r0h+lIKtPLjUkkRlaLZU7QUdjC5Nw64jC5V
MDwDDQEbMUdBepLJzj+/UMOuXLkLSJTH6m1cYlc1qjjsa/1eBnuEP+rN40q2fFi/SDc5tTP3mqsb
t8R6btJRz75dkpd1KxmJnCSPBreinqYbFUxDdR8pXV4oDV9LwC4tpTzSmhln27I/JWU3dow6Pojn
NMmkSG+K/pxeEcI5aDjlNZl3EFR9b5JHSt9JeHTgFNt5Z4Y0XlgHixQhh5D+Nku+lNCjF8IF2GEP
NYosYJ6oxteHuIZNK4ZMRzpZggrXZKJvZTeE//eAB/RUjR4ccx7y0KC5xdVTnjRB6rVvHNaln4BI
6uAGJPCsR1P3iAcJr/GSQit5ReuV/o2cAmnhjJgr0gZ8IDy2blGnqJH8SPmhf4nIXIc/RnEDwNNS
3FrhExPmFf+6VkNFOGJC2JHLPLHpWMJfJ99dAJmo7fOTTs5G2VCTOdor9fLMFO0EqfIPGFkWrbvk
dgKE0AUsyVprgTP3Y5nA/sLE2pavrrkGsSYfRk67TKk9LqH1GaoC6D7j6jwPxA+3sb/siQDoy7S+
GE+diCLK7+RFHQKo70vLbw3OqQSwvKu/G0mn8gPz1d6/9N8q9DTRPspqAQXA3eioYz1gR4vdL3wu
CtSxW46HugZSl8rsEt6srEIIMFzIx26mB5RWmnXlH8EDvWsFi/zdXvMhWG/cvRPwECJ6iq4bPNm+
ZZfCoF+LAya2j99GEnZ2tFn3a9zcPgifXl2ziowbPFhY6MaC0FFehvdUrwesSmNKz5vCeAEAm5iT
OqE1nasLpkPWEYSFk38E33jXCs+z9Rt+CXdC0j2PX9TDjs1P93rGbObDfkoGBh8abtxo16/Mot4h
0Ont8CNlo3D2qVuCpQ+MC/PIaRmtslNbvvKx3+PZ9BAcMzaqAIBYmFQ0ciwu8/OS5c/ZWvhD9WAc
yyaWy0znz5KI2RrBMTXiLJiYtZLzv1i1al4Cj7W7Ga+zg0hOukkeMuUzsY94pfyHr2iih+bsCxgo
z7Md/MLX7e4cZzlR7BVGOGqrbB2DCm0Tz81Xm1aEiDpHPZmR8BDuI4vLy0nN8aVlp9gCxUnD7S+o
oDGQmPA3ZMkxRuMIhZQJY87STgWK6txyWqlRbUaS6M4E/97ysphGWabttbqner0gsmdQPMzuHBaD
Z20uM73PlQJPFth6SU+oPFCUlcdMfBWhx7ThQ6Q1+nrE0NT6t46JoUhl/n1Y435MhIuzXajWqpv6
wek4hVFwihv8vZpqVU9p0iMrwqKq4MxQUe+4/KRX1jMEcHdLjpSz9hpnUx7lK1DUChaI/+ONBFNJ
wGki9z+iS3X/zS/d5YFOR/EdWiIQqFi4vHHXxKcUfw1RyVECUn3shBINpnRCo0NltuwgVUYkiEhl
3qYKXV4e5cf9qHvjm6QQLJlGf6LYWvrnxKIClLBQRle6ZEzXOjr2LEAyvSxzKc4vEo2+tZX3Q8sH
tHFRmU2AqfMBLPYACB0PnZF4v4Xi4Ric8xXGHtbRZs1A/+LiEK1NJhJz6D7C94InNpVN/itxFSbD
Lmy0bk0XJxAITsd6qFvyVq1wcZo7jpw2rrijaCNeDk+NzdDIdaJpiEzrEk8jfVXxod6dIRNQsMqu
wSQCvSihONv5LqANpMH3zoB3fn+qyz6R0SUsY1rlu/Z/feIJhjm0CxMqt8tLBpTOszaWkRBk6a1F
Oobe767sIHX6lWH//HOju8GtM9JpjTbnuwV4GZpCfTtiXWCg7RmXM/SFjWOJ26WSlVpqpePacgwu
mGdnAy15n8LMxkZo0gFFSlhzSwEuOIef53XMsT3P2SbY4HwI0YfmVVuaaFzBmDXBzawj2ZfQLqzW
lyiByNuQRIBidDP3TtkC1B+eQWs3kwyAMc+82TGWyOfcog4NA6dJmjQXG8LuOv3JUCcE1E6SMxGv
XFJTr+HwpcSRw2obPq92D3ZrLYV+CWD+JZU+HsBm6lmRHw3cvZH6pMzFLpD7Mhn+A1+VGT7c2vkz
L79ilLJceFZIdfX/ID+4cCxgfiue9h9EutD3/4WZGtukWfacxnphvnPaGmC4YizrQ3CvW+vN6YsK
I2jGhtiOI9//JGjXwY0tQRrfiA3/ogkGXWMW5uITQmAGZdWtmyELoLuCe1f7maZQ61rPkbTBl1Ld
AkalAe1g3gPmhGd5Fu1DdmrYg2rQSUEW/B5Onmup5An1MObwXlCsckEOImV/FcNsj3kXff5IqA6l
VRwaASRq0d3nO63AmiBCpqjK83/hiEowC/m90bKfAPK4msiA286NeYdIBWLyCKWiu7NEDthCVJWG
0OG0BW7ucjLVNxpCUK8qGz0irhteHJvirsUqpc5OG6e2UFnjG5sWmycCvYrbhNp5ovq45UItHa27
UCWUmHvsKbxM85cypOmXHr24J+rYdflb86s1O3GOcPr7xsJXhJVh2bOuQJpTMkAgonNUrZHzSDhh
Y4ZFXbSj1bnWz2uYJqqWMOZfDr0MDPRyHgXtxY0cs7Gd+KMpGQYLG39NBahiMz6nx2GZVEhBOZ2F
HsbLnMxZiSpSoa+NI6a9w8uo1rrd05X8nsp5Xc5ePp+5ta5f6U7Pkr+Ms+i5OKCvvzT0xy6BbZeA
OTPVlQ0a1U43RpwKeRrZP9gp7vOMrUJmR3XqJv4oqL8jKHTV+mZkQ2Y3Msi1oWv9mLtqyvD3X0iZ
GQQh1KiHs1CC6J2/8B27cIofzGWjNzZQmr5KKHqHyykGKZcnskEhLxskbZORwPzU9uTJP4RU4ayu
rMXkKzNFsRIZ63DmfbMdt8ZU8ifwmTaDpLASYAO+nd562pwbPsRLww5GNmPAnx3IRjEwUero5gpR
+VqArTgyjF/l/MTlNB4A6h5stYqnU81zsILD8+XQBtqk2MEVUpEnC7CcNVNoMKxylcOd4p2ODN/L
JECodFe4fLQTWJGcG+OBKTOOA4QwZmqMzngJ7NsiURCULlxHnSdtHEvBdHNGduHldc/dE7mO8a1p
sqG+6+jLIAA6Y6nV01dAuHCx3N53zlJjOEUI/LY8Kc6ykwpnzi7ouuPV2gGSPpaUiGvBIbc1p4FO
1+d1DZLM6VfgOHQ0e9jpdSMuI1BZiwxTm2AeaYSrxOusuK2fIMMBLA/IyU3srM5cH7DEi21C0Zt9
R9z6vurK7tq3Kym5LtIeQQj6uAtjlM1m39UhBUwb+53KqqWOOFhpHc58uV1UlSAx9RppnlWdQhfz
LOvwSce3CjzNtShEoFpvxnYhBVnkZO+j/SrN4UpkiilphKcc5JdSVmTbtzDkM1spC2Jn0egykMX8
nYmp75dZ/U5Gs0B2cBQ9C5OM0rAR8khEm6BDnWk/J+83LJ6J/QDw8s3cAmqE4Utk/RHYkR30EmbP
M5+oK1KomPLr/96afOAMp+eazlaOyED8FPSyURAuKxY784LgMdSgL7xBupfzFtDsSedSalt3dqle
PrpJoAXo1YcSS/J/9Wqo1P+dPPKFuYO1Bz9syJ9kjpaSExugxTTp0PsNCzljh9kq7HOURP7uBKe0
KPUONwMDMDAhh4wh1UsqLErYOc6YEOFM38P/dx+xQw5fd6IEgzEQMn0RjwzbehRLBL0s+OdlbovN
BnJiSjYTRLA6yazBw+uJY1tlID4g/h5DGcK2IeaqHn7I7DTyQky5mDyzTSGQiPX/ZbP9/jf3qx22
3C3edjAy+km7opONal3H0PezTWxaUo3oA7199UXaL3ovfFlON6dqjj/FmHRlAUuOOIolGviXInOG
pcM+lGFMau0SZp4iKKS4Fl9HxjUarAL0UhNibuCK3E34AqHIwgo+WXRmRzQo05AdHE+nXsTTsJrE
dua4gOs2DShvcbK5YygH7hM+i8VocQ+WcXldSKgJJuhFrUn23w7teoqtyIFI/Xg6wooNmz5DC51G
TpNlZgC9RMm5S7op6F/10u2dCqg93WV9kN7OQ9+saY04V7vSXhlBXizRWvd1Jr0eZTqho1ZvJwLK
e/MyMblAFi3Aiz7Cs8DUxfQ9+BhG103/qt9CimvZd/nNXgsFDeTSOnvQhxOlrCZOuzd320LE1GLm
gCBrcprUsL0SYHQcVn2hln46rj7O1QR+Rrsv0l1qFtOVBeAxviy6cvNiL6D1/iSarqWDaUKAUySW
IiKOR4Y4DwOEmi3wKeVus88Xu+v+IlAzUsfYygheLj215Gc1pQtyqx0wQwTWoJe7XQWDWOPjEdaC
wU2Sq2CUqjtvkfz8Dy2iMPAt3AQh+kBYp5E5s+I8YTH6R+AwI0TjvCjU3WDEwm8YaI/ouACBKWBZ
8T4VV1+q+HrijUP/WbzZ89dAbOawIghRVS5feie7EL0Qnatzp1qGjsa7ZvZ3SxCijcfDhVxmlXxY
pqaSWSY0LrxM8/ofyxjZ4zJIIfn/U6FtWxL/oWLWoB8c0oWItf09b/q+lAqRfcSXyhr4bwqwe890
rhtq035sHGglzbpdq4smOnK1eUR0nPKDTX9BZVYPckyQ4cGyuVRc6CsZM0T/Q3/lW6mr46Ami3D1
clV831S0OqKSuhUB9WV5Tdpt4K5rH5pW1kQ/C8Zi4asvevHpdOWaMPgRjCb8K/oGoM3WT6Ob3MP/
5yuJFnnPz1q8YGQySxuoCGtug5WhY91V0R4PIPrmJ5UFuKGBWPDEFEismR2OEbiOi8ylp5OWdiah
P/FcHh2jhfbVJ4welBA4qL07K6ibT1TvEGB4HKCrObztUMc15dpxKWNv/mZ2XtdRQsqwirbrYfJn
+m00UaGgyAK6j/h5t53lCOiwc+6QuycrrxEBGv6IoxTrpVwb3lPB/YklNk4FJ25tSXSc0yZBpy3O
m1hOqEg+h/u/FoP9lzuOsBGYGq4JX0Qs79sOEzeRUFKsa1UNZfiLyMojRXuYx2NJNhPTkTWL+1IE
3h83OuSCE0V3Pu38Xe5WGmtEZ9/NBs3/Pjel5UYey+YW5icyavUcc6SEiqtjBtUisuv9bPlh5eG9
2hqkTNTdcmbzjkzY0i/f6vWN0Pq75badko9q+RclFptRvW7Ur4gBEj6oUQv9f4PdTyg/2qsek3Fm
FTmkdfA1YQKAF6t+fxheAYKIHl4bzQhb/dNSeFjfx6ZCxt1aMeQh2lRO4LYKSOx08m9UX6WBTdWi
4T3kGJD3nSdUetkb5SQ/gsBkuYG1QyFxEJePJE9wRPK9Q9MnsPleH7OgchV8lxyWkQw1Qvg+Qnnj
oqYTjRk1RpMDhQJFpAawQiT/+nVg5CflEZKI0rV3oJeOodvkYhpfVoFACVhg3YLC5MQwZc9dy0Cb
xelMKUpc38E6vvDgyrDjgT5PBKuN3g3Zjs4OaIH2lUxo5C+4+tppc72gnA0Doau+qmGibvh6lkNA
4cnTUMG+F+rKZbbFYi6XTSf5bJQECZ9gwB9mcVHIqmrwwE2OC5Wm9cB5kKX2LJE16T0bRetCZv21
XOztKrfdPfz1VxIv322+RxMUB5XM2TEYvCavAoCXZYiQ2sHY9azIInkVKcBbn5ZdmwNAcgEa+XSm
kQLg+kul03N8Pv1nagZzm7s4/3jBdpR/ruGrLWZiW2QONYL9NZK0fA9DNM+OTr5HHI5McL3vh3+9
Zprqg8FyNuaQmOGVsOBV8hajRm8yVKnrUvBz1T8lZyjhvWs0siAPPLFg59UpzpXugrh3qS9DRJtA
DPl/pSTO/sby2NrdHxjDa0cacru+JH7U6bGFipca+fRUx0InqKnnrt0lNA9naPsntGdVXsC0Y6Oq
b4z8PQ9BXAIr+gBkoF62MbEKIublSDuO4gCcgFXZ1OpNkJEesCB7cayw1Jrdm5sWCOSx9YKgNzfF
xz6OgoROkT+Ppt9y+gdfoguHb9sZuXguY9mNZEWMukjsfz1WTeAOvagTNSJtQf5VkMaAFMe+zn+z
HJ3IS8CO3z1L3tsbl0K/0nI09jfZTapENpQ8+MDiM3L5dr8hk9E7SbNxtppPzhlZbT2184TOtSFX
Fvjby0FydT4fWrmLWdLqM4yjj2jggHNErZUuhlVuewaggLmNcl3a4NWJWuVN2KSZD7WIMlabsh2x
fSy2RNLgeWyJLG7AgoxR5ThfBYD1MnT8CkHx2Q/uC8u+130ZoP4LxexVrEaNqrHi2uNB6Z85Twio
gHQ4JPN//WND4JxEIGdal76I2inihuZ5uOYc+Av7hB3uJJLPKIeS7JzVxPRs94Ikd4I/dfRHvFlt
6fHHr26GeTDAdwEK/qJA9Ogzj40bTmQSONKzBH/TNEI8a/yYQ9oMpvBx8A2mHXLAtqZ+7Z0piuH4
wsdw6sgW4E5zZ8Hdi9q/6ABF8EvKO+/nzloHycHTu0lE2DBUkFCslhNzc0hlzq37HfXb0Uqkl4sG
M97mpuRpKAK+Rb4Il04A/7N4gMvAn+iG3YkW8uWeQoD0Uvqf6iMILLvN66xth4oN6cXFXDljyqEU
NTbTPLbRTvhwXSfACmfrBpmoKaQPDM/O1CFhBSY3hwwfFb1XWY7dXW9yMLx31do9z2hTachJCHEa
m0p5e11jxOpq+BTJyVM7oPSpijP1wW8PX4bSRTGDaFsj/HkuF6G73VL3xahXXN6ajpl3oQxsHdnD
1+A+hTwFgg9T3bQ8ulYm7RBgGkAxS4dkO/m4wBFf6AvGEGdU+tvVGI570DYYw9bw41Yq+hpLdFP4
03wkZmqLMOe7AQkiW0AoZg7uttA3r6ZeuQ5DgnN28wNWt430k1IWYOoe+vObibQXchyOoWPrN0f1
XYrgvX3Wh0MswsL02mcN4F4DIMB5isjxp0C+cpuL7WiIXnNl5xPIt8PwKtml6JNjLcf/cAV65D4i
Ttu0RgVQ9CUBB04Qzmw7UazG0UqyGNGkp/pr509SqRWd5MEXIA2bo9yI3KDeOYKSMACrOpF8sCnT
x61m4JBF6j9HuNs/xkC45m3+0rjUGBtrtakoGAoYT2JTI86x71nWcK00DwTDyzVBL5Oy2esUB+Zo
yrTni6RnXom3nVFgOUC72ijR5DXtF1zevCF2EV7zUPrmIEEby14qBVnP0j/cUcmFyVnNKXi0n3Hj
hm5XMBFnADOZR8ioHmMZbmiHTuDzm3QG4Cp2ufpyehnLAOoWaw7NVpvcg7tp/U/a1oky9594OtMd
x5Ty3p+oefk5oVedjde+lwajbFEtFfkkKfmvJKG6XlXeRlJJhBqujfeaXY5NXN/dmhD3YAkPAYVL
PhlbUIyH+z7ma+adXsyy5iuQXJ2/63qqcJ1agdJq5kzlg13Hxftw+r8scNoJd/FYDm3LgH1uUG59
CZV6Iyjj6yntMon6ieZT6bcJwVDH7HZu5R43XBE8hjBzUu3fHWHO4dXoZ1pYP12xRdi1SAx5xVJG
f4/fgfqNeIQ/q7sl1uNwKdBJ5CMN2MicfgSAP3rjX/lK3nE/DIgbDeevHV1NsFW+A9ExIAjQCES6
hOGXd58tYrxWr7uQWeUCFTKqbV8vr/VarJxQ3i7xpSg+W1aTeM16XGpAISBNUpFQVICxtAaDt5Rt
Fvnp/qxYGj1Mb5es9m4e8vazks/4c7T8jjT3zz6a9Efc0b3K7Jx2Ask+fzlFvJ4748zd2GVIs2KU
m/dDGTNivcml0rDSeL6ADFcC6HcG///Sj7tAotQTyUSBipgqUgsaHunX0XYnf4gwUWbvxaDdBorI
RwJZNkIghfjInkpKSNpGoooLMPe1wi7G+BHpAyRPgyU+rOCxpBZ7xWave5/WLXfp5tlsaVn/7dkW
Iq+VmGaCTsI5EZ0FQ8B11awvIGoDyNK9PFGzcoGAFtXIIWDiBUvPAOUYpn52ZOJaRh7uJKsC+nGb
D+FPjtFfT8J/+a2dNQk1H3WRZt5rqzA515vUG3uEn62j1hOs9NTVZamMMFggGFoEbrtare7ozYgq
V+IJQWNNdMlbP6H/+MImiTzQy4IhUfjq+U11mzpoOj8bTOrhUK1mhlPXZ2HAsJ1vRqQVYuJ2eoZY
ockSAoP/KBH2VxOmr5a9GkwXue+LTQiBQadPiA14a5YhT+/HFkv6e5/m5xM6dcBvT3aEWD+Bquoo
tr4s4A4dKScfMW9YYtSVMyOkymKQ7qA/n6ucjHNpXIVhxcSPZTuqapaUUamRstfPqg+D29+WkFCj
Q4yEy1DhVfnSNAQb3VUPfbWzi+kpzm1BENbrcXgFK0PCGvl8Gabfov3g4CP3rlGFQNMP9d3Jg6e3
GpKHyQcNGiEbw8deezPKxljvzOpcFgge6UhdGPQm3d976eCBa6yLt3r+P17/QYp6X3hOEiF4ieCG
D3HgiEh+b+mr79ezzdqS0r3arP3YEll1wh6354u+zrMmizUAqPRyOJWrqGOrJBhtfrNGiWjOq9j/
Ye4MlscraoA61LlnIJJMnj2HsIapI/zuiagw69j3/KqWI1OHMDKJgS/85pYPWiSyoIiGy0+zXclS
/EJ4I4ErK/rseeq2IwY0dFoy4NGJm8P8i4G/5WOhxT9/utPZWhZkw4MPfP37vReVTG9xAaGLjMcN
gKYXGLZfstlAkyG3nctnVkeH5wo3FPilAw5Of5DhlSVp6zlyzaEmyI+I9A15gyPrWpM5U5oPV8uo
uHfwVdlM89Vmc85vHZP1ezEvalSz4MwlwYuLH0tx4oSxmp28MkHNkikxGR8LLa2ByN3mDzV3w9RL
hRvsP88MVqNzAm7T0c0qvO4JZjePv2QdHNOgMmxfA9ctH1lgghKDMsEZTQqjR+U+FmutEFWEgcyg
uldS+7+P++vGegP37EcFCSTUc6L9EmX4czjr9ma75t4ddoD0tm46SUWaNO+oUpsNymluyFRQttXz
K8q/sqWfhq30sbffRS/UKlCsPTeZOW/lDy9W2aQCa+kXffZhxQ+MEbLpTZ+7rvnCDE2Amy+GrGtX
RYxx3mmYdNepyGxmvHGRLPB5lce3n8FxzRaUy7rguzP1X2PjuZAftWvXtdHrmcsntdYY3vscZJDk
UAjyFFkGGroYrhCgyFU328LKVAlIYUhax2Ve55BHdZ7fa/vwVadywIdKCVwIZQiO/tmKqyAlgRNK
xVSqUTny3QPZTsLd0R5HZQN8wsiCz8cKCpQ/hW3RRvn4vfbJpXodKp+O2Hksr5keN9oGzd+/44gr
OCofgozod88qBquaQvyMuXH3cKVWFLf93v33sQ0XXYBWQ0NI+Y0xB2kY6QSByS2Qs4bMT0CGkveE
oqRDMMPu8MvOkGXpEpIg6kqrT+qw4exN3omobl4MDKg6U228gwDtrSGjOFsoSg15M1v8m/zz5Evn
8E/cuMtpQ3XZ/kXq2m30ToI6omqTNK6REtVatU9CT3dNnbKYIwxFAQ8YiY0mLI3My/LIQxdJT3ZU
46b+n+RRR1usQ6VjyXSi778BEx4PwWSINupwggmPmnFLaC4/zQ/otKKwGTZKRJA4N5v+gps8Nd4K
3TOq2y02TxPyJhjFJbPmuHBjytThVahDDcT7ouQAYVaoFCkn8xFSCDjn/OxDxGtr9xj/4kBkwj4E
a98gBk9KOydINOPS1/LmNS5WtqM83ffxKACCH55A0GLWMEnZH3AXwwQ7fVSCxIlVa57c+Reu72Q/
iN2uL/2OpX52xhRuwUO73nex0bSrh4tLmpkXDU2wSOFGPQHzG6L8B42DBI2Cbo+zFrrkrO5vnLFe
kVoqY5/Xy0kKEi75lI89v1BN7YY3hyBSlzXa3W/U4la4QZt4Tk8HYVxCZhGM1FRCnzpX/EK5kayJ
yxeT8TMbo47KXClp/IRZGz8ZZUHr/DOEaqA+5kf043TgdsfA61+NGTmNBseE4MMTq0pHTC4qdjOu
JMjzRVdBzdETeD1YbfeudcCibI1PoJ+36YLhHtGvZaugIboa35J1oy6piCLdsNSKiycTWpnUVj8b
6J3x5jkXkdR3HFVS3tQDlB212aaNZ5GSecp7XDapPrQc4Wd9QuDhpgkzgbLEWSbNqjTdUu9PzPhW
HaU4mTjn/abrALbfYpWFhKJha8aSdZOfalnIOEJCHTbHF9NwMVZ94HlZ5NxFlFTHcwnfvd6xAObi
gc/wQaGz+RZ58weZAekuS5PpiwdzwGsxQ5bOmrfdVW5C8xiK0nkJUPHsja64N+U9bHucYfncFIDh
gUozwcCynYsaHupLb2RFaBcI1KGqulBdoVJK2xRQIXm9lUh1tQoorUDV+Ywv/mIlx7IP4DXJPOEl
UQK81wlKy7fetF/ZidoXGWLJFxpp19KMIGw+Oc/Zy3mw5n1LZufYwP+oiwlCQPUjGhO1U2yGj7rB
sBc/wdAJDMHEmKVNQBThpZjMOuhWczBMgM9uEh5yDGdh2qGSq/w1OoVkEguTKys2ojETnO9itMGM
RnM5pa2VSdQ2+kjIGA0FOCMXxAz4D//GTGtMAu778E8RwpwRMAYEwOjmo7wqhsBtPiSwgyy0RXx6
zGVZteAEm7zVhThrbCbUthmK/o7iIVtNMYg97ULGKMPQnHWK1/pjWFFErCjOkNmGed1AXmJxP7Oh
gF+hWWJnth8khlNx6E8pUUEA8p5amoRxwj7CrkFgpSoUB73gM8pwvgNK16eJHk+PFyzqWBifIEnB
9YDFnv+Nb9CLymXvQTDvFImHgkrWYinVtS1/PnFYtogqbL6jFnDWCJFXdNPMoNp6DlFurYsBk8kF
JCFKhaiCbvEUjQNNDdGvfHCjWgH+l50Un+u8BqEeT4MQua3DMC1dtKTKjq78YYvol2v+sEZcWtw+
WXAwCybYGg2B9HrvnBl5hRWB1BsNtVeZrilKLJDhaRt+5RU9ZwMpnsMW6zCy6YFQvp4XYF2xs7/z
lh4CAAeJ3mKzrj0kd1bHrsloIA6g1/Omv84XUuyVzJMwlg8/EdJ462j396AN/2WNoVYL8RVGNB3X
CvNjN58no9m/uriL2aom3VW8ZUxkURFg9Gn4lQAqWklJQY0msaUVKg1Fej9QJeE0m5zWMqLCjvgu
z3b1bQN8/NYMcfbkjDp4bUpHZ9w6AnkMZBcXpZx6eQkIhSuWlbl4poGGUwP/vlgILnct34IhGGe/
Z2bpNdFPOsIst7cJjdDxYg37PF+vQW6JKX1rNhdIACOAynKoA+KLEImXHlX+p6na8uq2xQ4nrywz
4IEvyWQs6QDIWSdhRre1pmfZRkmH57aXzSd898Jw6PwvwsMVxO2DiPQBiBcaZ2dtsgqRiW9QR111
1iDKNR+5lD0qlpcz2X50UgeVJ+xWSEacENkDfmwPMcVAEzB51FjLWE49pAOGLB+HHDm4qDI7Siwx
06uiqqQPAb3r/LMr3iOjQhupS2wN1ocRNV0tIyTAVLeiOMCtVlziK/zGLI0aWuNMqFhHJUgm172p
W0beOXJ2YiKlt28X0OHXm00WBoDGbNAcHIr2vqFFuS014OR4IdiWlCexfwhyT6QyHD8QctRmRsSy
3h+NFv17QUu3jH/DVYKC2/sFiRQsDRwJuOlrGNExwnfwqP0JmEukg1dwzTq1OGGAKGuR0tzzNnsP
louGiOwysEparSOVRCrILEFeMuXJdEVYa8nUn4JBDDJCoJGdH+Kym6dBm/qwEZG3LM+i8erIrp2o
bWnx2IZognirMm8Vx2UZuQ1XzeLTnkEpPyqH+YI+pMwqp1SfSFBiu28qSEkJOV/xUGHM7Knj2UR1
rUcBWlWEjGc7WP+OMA3zorxoOQK4WCRuF1e3RJEM4liW0ky2AK62GaSTUXt/LqwhPisfsrJHdsQt
CTS57hd/bWlK4scazE6L5q0n5PkJLTX+qYcoGcrYyryqdsIITq655+iRFWJuMWrsqu6wPjPHES67
OgjhhZ/gXoQOhVfU934M1wkeABG0QTSj6usxwTrfLJH0SX5VnQT3+cjyqCkrKIf9h4+ChapUCVCX
s/lxBBawZ6t8szvhjkedeP5bPXB7p1d8S47bPBXxSatIgiY6R6ryBtMwLpxVhlhLlmyekvPh7duz
aJUdIYwk8RpeZ2deGSz1HcQrPGEffUG7oO3mCWe5JdIJOPDCEeRkw9jV+b7CObm7Tz0/lwaNdtNH
K84ESBcpvHt5ozyQ/74f8By58/e6N3SxSQTWVC6N4gkWw2Ov67+ILYn0/Foox0d7Xnt4N08jdDth
kH0O/xAgJUPVoTVDxWMnbJKZ8LU/dDyOuhkIiQa+nK9b2tJwJ/ZLKjzeF1TBbnT3QhxVKQ5GeY5h
pqpJLPPAlLJeKVzwxrREMqfBMaZHpBh53aVX0o6bmfdbYF64dGkJkwed2zWjFx4hWl1JncTZ7zO5
lukCyNPa7cXLDnouR07YdF1yZfKgCKdFUsgN60mcsJkQpQ/oGj9odTj54554FDoz2Vl2E0VswVGq
dSh7DXvp71rTrwgOk5AplkCruzin2kJ/pKunfYUkSpAt0quazXLmFo3DkGe1GsmOyfwmCllSLxQF
OD0q7HWVqDuio7oU1MMK52+iMQHsQnHmkr+QpFA1s+EXMk9KsM7VKe8aoUR1A51yT5XtBtkOC9ZP
AnU5HRtr/jqjq/le1EYHEZc1N0tSP+LHj8Oif060fKfGF81KwOx+lSJONBg0WYH7GOgwc14039NV
V0D1W3R/kffD7a0eKbY4YgHcKsnnD5F3CdAGSA/id0oHDLgTBo2t2SqgLnURZLxTOlEao5YkhUHn
SHb70T+x2ip/mQBFNBVwNhdNBn31qs7+Lh2otY2lzmRJGYKXpiAqtCIB6Rv01jPoLlA1gv5N/Vum
LVzf6zKjHo8gNb2YvCqFwIBe5hO0UtOrzseICyJ613MhJ9QDT8eHyOtq1wzk8YkkUOiBNw3FAZMy
r4cx+cc+EcGsRpbJ2YGsKnQZy/SbDHucXfuKlbiqSaOI+8YDMU2CJP8swLLRduDb2Kw4ie7Jw3QU
eyZsBWzDIMajc6Ft5w2mlOpM+yuRFgY90AD1/qqn66exdw2JN2+suXRMRB1g19XbEJcFx4JjLRix
c9btH8u0qpxxcOczY+3lj6L7g89q07VINdyU4OJUP+PGYixqt0q/0f82V1jMg+dah2dOdbs1DRhA
dr6icpQYu+2UDxsb2XNs+uLo6P9t2P1/FlHBEporksal2+Aw1NOr8u2740YGxXzSmIMs31TGng0A
x2kWxMjtlYhPGqapok1swFUFRvvy9dQUeGdDaaeiIK499JkT30HaQkUGw5B4wVgWZFEbKZuzki90
TQriQA7UBXpRBN8nezIL1wc3MFIj1TS2XO0oZGjomfw8MRKpHFZPcfD4gDSM5R+MSrm4Z78l5TOe
k97OJofZTVf7MkFgfgwmBrRWEz2C1P2DxNMC8a2g3rqshsnNJ3U6n9rSRlU79z8x/nYASHztgbrq
VutXvefUpa+gvK6BxxsVqMnL3sV92NZVvaaoB0Aa+HeY2NK1hFu/pJS5D3GlVvTZjxp4Mi8R2sYC
1sceVGs9UROCP7lkrNczE3mGMCYF30te87a+W3r1xGnF9DP0J5PjKgxoxkhktS90d2rNu+nZTZmb
c8+OE4+Bn6dYXZ3a3194vH4DqpZ8+iDzLPCruVeIS/F0SHngG9SnEHGRv+jVto8cJkEbP9jDcKzW
LtYmJpMk/rSYueFGmEaseWwnR9h0IsY+qr+NVYZ54MRr3LKbGmpSTPkmyLMAZ4qzrX5y1xTjmgOH
uTkVyffuVp7jYaSVeDbr/J7LnHtSJH4wD2qvp/DYFuBQ1Vb7QxikoxF8GxyB57WPFP/jc0p2ciXe
6dCCJ2mTrkra5RNstHmC5Cd+eCoOxr7toiqYEqhPtI1y13e1AeMXOWFU5hdMImC5neGG2MHlnvCJ
s+W0O1QI8ZFL03+ij1aPZxw7KDEIYWChNlYB9JBOhse5UYlm2B41hT09tqlO1L0EGQmQFbgy+T4E
Z/MPCyIMU27Hs3Utn4DD63N4i489HGo5d4mUSQidYOjEqKC/xhYMhGa6bNaUnCg4wEHDt2xSOZy0
fnoOZdQXl2359+TxjBWxMNl5muk61k6cY1xZgWdWO/vDdEjdTv6H/B4nNJw0lp2V+RYxhuK1NWeh
uUieGqVPs3pxhPr+juDP6KdJp6THMuwSbqWwearvpiajIFLfEVgkNyc+JvX6D9BV+LRJ0fE5ZC4d
d7U208OaUET4vtwoe7cEIyU4wsTE2sL95DQqjmcS5xS6TuvvpyXLtoV8VQz4TieZQjm1B955bGTi
H58TJLsj7WOq6ANEZj/NMk3TORLvuP8NGWSigNYKPaox5SsnAqxQXa2zVWHW5ba+ixGbOdOw8NqM
i5WGauG8ynwfHe4dFFxfHEmJjk9U5wFtAp2TCHV2+fnmWqAvDGUM1I3xLItcnnW/XUQLbkP9zpbL
vxx3WPYSx635OP8U2relnjKMhQ2RxIwyyvup67Mhfck2t7MmyZx1E8zrEHuKsPON1LVzRtw2VbOc
2IL9R3Rp1YTVoM5bDg8zecvEfpsaLpcEKw/o03pjRfBQ164hY8XURu7RnSg4QHWjiDifLesiJYHW
qZ527Ekx+lJnEH98NBte90xnz0lRG3s/Fu0SItsmLyQ13sIchL8QqG3Qg3CBegfX7W6Mfi4G14fd
JgkJFCMncg5s8jQu5C7dLMg0u6DJ0Ommg9ckAAkFQaKAdlGCHg8ccwrQPNdxeNruvCc0bHM/Hcny
CuhUrABPNLMayy4SWNSYwb5awagGH5hOmh72s8vaSsRvMPe2lYQua6nzLTvIykKp8K5GGUsp8SLI
EHEmvZQlzz6LGN9Tp8tv/I6FxAfJqK7LdEURevVuZAcAF1T8Pj/2yf3pZAKoTqrxfzNgRO/JdnH7
PwICHbNR5Fn95m1WkwbgFZtqQ4MgcU/9N6a9hUC1wmAxHI7ldm6O2iPd11tqe8jtRXDx0yGFhjN9
EFLXtGJozTnJr5Rzg92ZqNfQFWzoILl9CMATW3ZMOiJS4gansqu9vwoim8ZSqiWK0akxNVaBryKG
Zx8qxpuymaoah0yH7Q7wmcu5CnFxHmoAPBtCx/r4/83sQqXiU3pFQbPB/jWY19oKwYNOZX0B9NuU
hZsDJhrWLvyuUXdznv33fW2IcrlxRW4Vi9qHZQbFh2tGuQgkBAD9BwlgQ2990DzuQHrDatw5Aj+o
akXXq7bkt92RCbjsz4fhWzwM4920D7CkscSbx3IFZszKMZk2goJz4caeARzYA7xU45vwpAv7D9mg
a0CuYjNvd/GRBMQewvVN7UWS6Mscw/SQP9ez+147+6YpoGoXrIbXEzFfJxqpQKpPiW45XTk/n+C5
oeadGfii3cVkE0A6H/2GXlSGEv4ideDQxFRXUx42ZwQiVB6+dxIwt9ynNDa8izCcyEXWe2hb9sRy
SukIiKbSbPbdokKWiYUWjEPanI7ILjd0DZVvZXe1Y7K1xhhrYCoIqlqGMLIpvBMADlG95kzO7ZDK
Vz8KPn06KtrNb3m6eabWdCGeHg0C5s6+iTHByIIYUyt+LUodhKkrUAxBLh8n+3fsah23STI7cK8h
ndqditOp88mKs6eod9qjeEUDSBztxjf1nWgFxhmRBoCiMvlx4Q/ftnshzqLf/zIA59RmH8ET0xH3
x7B2F7d9z+1PqQdL1AcY6Vc9KVdMjDhMV6kh78MlUi6aCeHQPuMK0BWmVQJqJT0UOj7y8HFwg9As
yNEPQMkQeTHFDUlF5kLDuKW/yzQsJGJ9GRDZirviVGzOtfmePcFPXDnWAI/S0OfXPjPk+e6h2kKv
iym86o+G9je2yZOw6ZmwpdXuNu5fHgY8RWNW2Pb0HKfODlIjnadN/ra8GG+JrmWc8XXpOOvKDZwN
eijUjrry8qO0OTe/j4VdwY5z0ZHUIhNYm4G99j/OfIaCm5cxYyR4pP+ZGP8bK4n1GT18apUPSofm
1PVRUcFoEyNlWWRDRtJL91o7J4R4F/wodpuTYhly92oSxe1o4IO2W6+OH5yYR42OPBlzIvaf9GBj
ORAepa563ZWk6F4g85KvCp3AOkTwD2e2iOOgdTyi59h7UHasG1+aKYaIGMcGCBRELBC3DhuvazYl
CbYDQ31EwTJ/upZPfan1A1UVW315Q7zTVfQ1ug9n7vKXLIRBhHmrS6Gm3JQuvJaEHswOVK3+Kra9
GhJCBBcZBhTsW4m2XPsLGfCNjz2mU5fOwiESuA/hlv27BoBraIBZsMfV3iY6l4akd9UWHfvrbBLF
T53gIVREOfP9b4SqUKPXAWdMVAUctZJUAkRYNInQyIR08ib1pZyxF6LMecUhASGaiai9TFkr87Vs
5G+Vh/oa2PY+HeIq05zUsc5xMqk3hf1/viaLLS0VM87diUsawMbXC9p3ANBxld/Vr6GBWeEa4NfU
DWUgXhLuWEVZAaeXbFdZFR4tjmrxQ2NweWe+P2SfIRUFBi1ImIIhxuLAcgA8yk3IugivEVQZd7kw
Ml9TtjDtdfNP99cMpmYqCTBUdsa1ESLYkgSR3o+2VfYhwjINBDq1sVYgcBbBfhCk/uAZ8mCbD2tk
INf6wqudpquxx+wAd9WRmE1kxvCQvG7BHcAIqliOxowTYfDw4kTWuymBwB96uLKx8QqMaVuT8M08
nGhk2mW7W2dNvKXPEqLV4MFouPgZqDM1mNCE7IxmO/dCIf8fypoTDH/771rnW2zHw8oW5apn3nye
TUmebsRzfWzahpgslpGtfhVAsS6OJieWe+BRvubfyHgGFyAvFJyMUnRptBoRjsddHiJJ/LV+Oooy
VsSV80jtt2ZE+w7CEGYuzvSJixgln4devrNlBjjM+Z0QN2NubrvKZ6l1vwGw2T1pnwsS/VOxmUY+
hk/m+vn5juti9z4fFerV8P1H6JGs8KeZtpLuJQNAAGclFVPMjIJrZbBK4NcMB24kiEPjyNEBLPNH
cxm+CKeP+sBzX5/LFUoAf75w3QBfjfqLIhG4BHUegDo327IOXDez36LjQWg7x71OxiIVtTGoJifw
L2drJuI9IJHUsMgNWXCsmk9Fykb3pKnCYZINfw7cq3LTCKD8lExRzayFfv4ls+/fZ0Whm1Xs1jsJ
55IpSMYh5k2hOdUEUU3e8NXVSJX3V7fju0xkt2pEQXjefkdtsHGZPHrmRxDbmrVtMY5JnGRJ6e6g
/6336c2b0Flgw8qTLdvrMVU794FXehMQ0rLHnbU2neU6DrzQJK+agBL1Gg2BxjtshjyO6RiS2q6m
uNEkv9rXU++ew/lgN8xKzWm3DfRM1t3qbFcJHMLOxjqSzOkrccY3dIjumcOrar4gok9VVZcXovWP
EsEIzT1FDYHBf/nC8o+//jwIeAaETvNSDb4dTp/RjJltpvvqRCiXKhzJN9Wf6q9n93JxAqhvR6M/
hyf4GTud98MfIGyJqB8qFq7AzX23l4bPJ2uPQe3tqdMNAOorJVDSJ44j9zVhLShnsjAp7RjkV4JW
6muntQqFP5d8qS83I9h2zYjFFGhiBjKIyH6sTLSny8Es/rMzsIi3/AYIEgY1QpjsUPVKmBpqIbkA
rscDkCUQa+b7z4IzWw9Q1kR0CezJvp64BIwIe4YeDTbxIAK6TEXSJtD60hGDQ+cHsRfTSqmm9RRh
MkAnjMk79QpBCSE9HAKKiwZ0HpozyLWnpDukI7r9bpubjm0nLzY/8Qa/tQpnBTLZ2ArNt+5DXQyK
4slqjmUW9aOsTUq0DN8ynjv4LqK//SAn+bUpsabJUk/zcG9J6IXFrBvZ2VSIuME/fNyQOgZnK4yc
kp68kr9GYOgLSDzWtphN5sQ1dG00nogPhsTOeOx0r5YG/hVhmzM2Uc5AKKGe1o7mc7As568j32cJ
tWGQj16b7tO7r+cA/LYNuhcVueGWRE1YK6h8VdCRL/8oNa32GGFhpe9iIiKltTNKergV/gUWVngf
5TtHsDSB1sG7mU7l74leHJidJaCLNTcTpou0UTp3Phv9yX5GWPJLUhavQHQGHuEHVsbrY9TCGx9N
3pNJ0tMF1bgD/TwmP7EH2d3bmTFKDBXoyZKWgOo3bfg+ivb2H+W2vhh8ftF3+IOhExhwUtL1Uwde
3rtEG4CVECfcVfqT5ZCtdHtzCwBfWSC8/lyzqjz5xuh+SdkEl8levNW57A3OGnP9nOrh9M8HE5uO
bJh/zNgQxhBlgJGVOJratRFW64JUq42m8bbIQOnP/2BZd4lkErS5mGOk75Gbvrh3Oj/AcFH4P7dT
6QjyWWYE9ikhYZlgZMY7KFhvzrgBVVqbWeN63GMKMnz4lZN77fP7LejK9AObrEK1PZHhinoRIWOg
9Tb+cDCsgX/pA/UcEsGrbNKni8mYOQByiVzOa2wk3vwM1iTVAdWj6n5ZObhyvCbnEP0UXdwq/KJ0
fgFgMEOxZtP1hZLDyir8XfSYutD2GFS/cxWagZVjqmsYOaMTRlVD99w3lTlIswrmP47S5JF/5S3X
wC2+UCrbB1U0ZZB1Yitgul7yW3kLOMX/xEmO+589IIWBiCZ2CMGkM2ffwLYdxYDJyzTHLR+df4jW
oRCpVFGxAbyIAQXl8uf+C6x+2S9uaP6dWcTW1Xx+84fDwezUisfRDI4mf6H5wf38rELrKwlzJ5Tz
fl4znHs/C9LQby52N+mVfrOYvju4WW/bDA7o3Qv1NdNIxlWjiV+GkKDhwvGwFb/rXPuGb67jt2cZ
cSzd1PKOQdhWCystG0zREx7YRUm/kWauU32zjpLN+klgBKSPGY881Vh3VBaqrPBg4nU7rAaN3phI
2XH12jKrHCsFjua88VvS6++M6VO8o9hnbwlRqMUdbqb4GfZgsmjxp6xnQIPKHBlqGhkCKZTwy+lp
oCFrF2QbitYn1J00fs4Kc49yfNkKcHyZwbizYEWpOFhApX084YrSTzmOLkMutkLMBQokJi8KIAc9
bdhPDal6W1lDcLEMbNUrdY+2CLvxHmvYSeJRTEjcTUft4HyFNx31ZrGoxn1GRhdBb+2MdbFbkvUM
GIo2+KoDXIqpcL/zs6Vt1PTX4zemJ+9dvj82FgPpYwK77PPN+f/HtJVp87gupvv6etdbu+Q87LZz
nSRDjdrqMZB6o44pFuw6wDwvA/0shq6/KI2a/3MgrsmL3jksnxYf9Gp64RSY+yA5T56jOUNcE/qF
+fL3FfmkA5wFXzGYUM5vrrlbBBvvuhpDiWwTaQCEtG1wrLehQaxC3UePQVqMVGNpSliIDTf2LF26
B7QE0PUYpyzP5zE7G85p0pTYZ5FZrcSbwQ4loV3yygSPz/Sa7Yw5rVOMv/XO2d3aTj4TRw9qsF0H
0/CJrJYffG2j7AvbQt7nr55WSM5wGxxO3xrdC2aZZm1k4doTs0zd/bPO2S15OOpIqsUe0Ie+QPWq
Rz2O+iR3pbqBIxsWrJ3j9t12I4A6qJ1wBw3uTupXWHXU2TCBHSZVQWyroHauUa8eg9u9KPpwbuuQ
Lw9LciorhequrBiAkkQ5SHUEdhVf6njJ0NmxZm6lZgpRWmMszpJO6GcyHSME1zTqyCoX/c19y0E0
o5IEOsZgUyTs01Wlsk+5T1OJfwmmZSLUjeKgH+52szXB2k3+/swRs04jSaLH5tnMGUd5LmDUDfnj
JgYXkXndpimmIENRtp88GjDgml7CDQ9ljfxSn0EDghpVyJIcn2xkWDjx6TnJBcaF00hL2JefMBdY
4gCzMmsaDrMNahgS2I1ch6mwUnkvRxyXnEdudNYOeCwaE8q0LjX63TS9W0lshwEWbiGbyu+YlfAK
u36F0T5jc0rlh1T1eo/2lzz49jiXfomuv2uQJOoAB2bgqEa18I+EjYxORBR/v+TaDMFlSHXF6Bak
QV0y9E1yOsROhqUtzsSJMV16YhnLldzAQBdvZmzibFWgVlCG96LRGuripF6K9cBweo4uGU4VCEIs
qXnoFR7X6fKZV/dD0Qu7EWtczPYiOn50fn+k3gmtnU30UhNKptfeJJTcNMizvc/HGO0ksK1P/uie
45ZFOEWE5QBAUS7fvGR9/UouU9jcNCFQJZnQ17jCRH4O5T9VfC8BpZ/bUBUa11JLzck87gUh5F1A
6Uh4BXaCksavgwQfCnfJ8ZhCriKEoBWOM7meLmWj2LoZKl9RzsSIMzdY5m4bHIrxOYEMi3S5IdJI
g1o2dscwvNCjqTxGaqMM0hWXuK9bo1/ODFnYN3P23e7WwXmyrpDiUZNyoXPwz2f7JCWuCQqoWLPW
O6lf9IQ/umH7s0pYzovQyv2qab/KRMpGaj4VBwajfNwBwuM4dt7Z6D46jW21xI5Ur1XSu7KjY39m
/B7lTm8FZ4A7Yb7t16V7v5jz/mnUxhrs1KkMIjS104YlaiT258uqT+VlWwPMmwCQ6zg288dJOpyx
//Gs2y4eDUzvwLvETEl+zokvbOrky3GHFR4i/a1/zV6NNbqmnvt43TmBERcaYPK7FMeEWxLxkOFE
Daqky5DQrQsjRA0+N1MIv1BmqIab8fXZ4sLAjZD0Fq9PueDtf5O/4oKXm2oIDE+OqjFTNHdPEEBB
wrxZk4AutIi5cXj1pd5Fjd5YuclXkDgcgp9lzosSO/rogTvDdNPn3seKW+zGFquOpYkmjAeCrj12
qDxNqOSzuvzA/Dtjx4beVYEQCJ+KfEqUrwspm3McO1Z/smqEFzaxVQpHm5AHj6fq4Wl0+mG49xbI
p/HFUuQlWTbWxT/wgxpkq5FTwfutSdQ7oYUbgWfgWnIoEa+c1PVMY2mj959gLFx6/q7KT+V/qUuP
+nSFjVMIxBcD3/PYfyYtT4keIKo+Ue2A+2E9MhVshtrtGQp8vwaiQZDEXdwzhBxsz+J66jMBu2/T
Ra7VNbcssk6kDhF/FABk/5xpT4sQrxCS+JEa3rkg2bCZAR2PzQECypQW/sGVT7/0H7jfgR4EY1RL
zCn3aU4ATwGgHcm3EeY8w7rkFHrqLEayOSruzirV5zbUZIkq/5lg2A0ZnO1ovWpCUDbHtEKaVPkq
DRt4tIufwuWBUSaOVr6pvViowR6KSuXpFFzXaSKsAnrt3AmGkW17REKJ8DcwyqwxfernNgVVoF4m
6/qx8vQ/j/fEEJFL7c8zETIGKCHu87D1wGY+/R9IdF0vjkjNdKCJxEMzbRFTEMhNloE1lrKliyqN
jg+iQjpzIEyu2M08UBBE01XmGKBzY1FrK8Cpb/NMvk36yEuLauJy5yHIJ9ix3qxbasz0ODEcveYC
FjIgw+/VvP4225SMBDuAj4eB02OTpjWnXIerPxvCznE5+V1QZegXYV6SCfdOI0ahRXWwaMMTOl1l
8ZLFP+zeFulib7Fw8uHbxwbbioOla6PxEMy2MKxeb6IHYx6Zd9vXDKWNlm6a2Y3ZqJF4eeG6d5kT
eqDotEvZgjOQBi7I3NUjK2Q2tZ+ftjO2c6UW2dxlh8d64w5dWNSYVgtHtPe/Xna3Tr5wVZjs1/OX
jsBRCQ+y/BL6dRS2lQXww83y7y5ZhG/blhAjO6XN8/UrxP7XO0K73uf4OHoNX0Oc9svN9qnF6Ve2
mF8m58234l5Z1Sts5HuuXm0LIe/1BFxn1H82AX2NYKwakOM2FgUAAdqGrCbkbgCh5fkL4BV+L+oN
EPCNamxbGKGsLDMTFiWid9bhHs70ZkL1vx0XxCrbsMbfWUG//aM5uVWLM2xH9KenzDqN8NNCSmJV
piTyvL4JQzepfOb47+ANbVrOmoWOs+CM5rvUm36phbhUZSXDuSNQE3rCsJPC3DG07B1KTODJYVsU
r8GvQndaD/yM7gKMjpgR7iHoqiFtTEF460rU/q5SrUJyF8XjxIdp3QquDevt42kyczNu2NfN2wiK
qD+2Rm5y8iEFC384R+tyql0iSpezhy3BJ/PVsIofXPpO3/QmaXI4j84VFo4n+x9SCwK3aTV31aBX
2vWm/7/5ho5HvtF7U8D1R22tXM5yZAsbzwi1eU9wiFWIAJVJ6y7vBzAekbUMQCFijQQXc44yHTcb
h5kHsM4Z2NFWaF8GddUEZYx6IuChptpWegiyShCyOb/FgTv7wM7VTQbkk8WxkGe/xcnJg8P+KYyF
H0sKEXmNslbM6keIwHCGlDgtLgz0iOPq7szrmV6upxKg19SMsbBe03r8NczfoyjZQLUSlu7UMakM
RVw2DacmzOIyF+n1bUAGltdbAzRPSOScF00dcPkGyhcMDwxzA9GikB4WwppWOJaPi6O4+H0Vtean
pDZncqGK9d8RHM11j6SUj0KzKdImGHDtMm89MQpu2UTIU0Jjdjdvx3vyEcpXRxTHozHs0EaOqd2I
h1AvZjvddByO7Lbk4RFhrjSbtoMrWMbyIznb3jH0Tiu/ouiAvvf21XST7pgW5acDe9N1REWKMqgg
7DMBunnQ0A525pcaq3y7ZlJK3Oc1HCRnS3Kr/7jAjlto5fR0a+sdTAMRo5WeZpIYeDkV76ujA9Rg
ovL9hmJuJR7FJlcnatioEHIq8h5S09UufYCfzJhe3aHY9nmhq1MOvH79XiZ2BWriKdrspwYRBVV8
YVFIi1Q8UM/J8mZfhadumCqK6ZwfKfU0Wcr/TP2GqW6PvXPJlQknXX51d243sDzbZhFlFHQs9lWX
pRuOZT0HL8mbBGKfEY+FCHlR3nULPfxR/aPhgWgU7/ahBiFtQBWDL0YqWg2+1qPeKc0GlrXFS8D7
0uIEL5waRqBc9Nq/Y37rJ9swzVHoT8a1s1njv8kkjVl8xG3qqdVEoajA21fao26VQR6fsuuh/FRr
JzePjPvl78yK6wXXDDZDhbKsFm7I4ZAclvVEQjETFa9pSphdQwXTA0KHSFzxsqNV3LFyvAHbBGcd
QA3LgSGgQjqbWSIR1Snf9EzlKtx7jMs3ioT4o5VxjKmLrIjqyW4qdom6/nWz4jZlX4iM91HYOcrv
31yd4d87L+KnwzzCOvj7zspReoqQmMD0TuEPceQvS8mk7qQccokZotSSEIya7/A6GzaCKFQxpHpi
oKpvAPmzm+kQuUA9DmHdsz5hOJHjz+V0FiZ7u3bzsJpiQ5y8Yz2uCMfnoNjlXdPh+l879cFWT1sK
YcpAwSiftgouOaoRWzsx8nPjYv6Gg3+g/Rl9AsI7KCKQbCvP5P5jBwgMKj76BxuvmjZ9CeVWYue3
D+NxGmHu1tDAMqwVNkO7r+et/81zSBuyEWqTcXl22TbHRH4+0Et8b5bGi6rduUzayCkHIfWthRWl
gaYFWVvotdVg/X/1ogK9q7OpdD5KHMMmi3MwCbgZpIeM49idHxpYqgIHiFH22C5GLwMR6JGSjHxT
oq8Q3AKLohMP+zVriTC79o74oBVRwt/tWa9isjER1vHC21ElBXTp7rSmbeLKUJ9kdxL6/xRZv85C
zLZBIaeDMJ3XyR8mz713VbN9mGbgnO0kBJMBQOYEvoUayyWrIHKs6CCo5/V+hzcQ5NsRkce4F9mq
jftL2PVDKUa33dBV0uAw/wE+v3hs8FQ3d4cXAfhrBUdm6ZMpKRX/MqqXp9TkDhrN/k2HWW6wZs/v
XCalQiCe8GnhQ6zSKFl/hiZpEpDFHc86k/W0M0T5BxOMl7MdHz87nOL8YQlKuns1FjBuHBEdQ5Bi
ZPQjiyc0tfC5vuP0UJmbuentIR8hAD0O43RuDDlfrHpasg957/qNUpTNh4ErCFZiHD8DR8rcl1tp
1WLEQqSlPKoYE0fz/QzDxZ3tf/VoO2gci1UwO4rQzADp4lXJ+iCCpVf/nxjr2PdRT9KyuQEAoF4i
+3yLJ4B6n8FQn4ctt/EVHKOvdv4Ug/BRBQebyH31jLaflOPDtVz0XNPlPa+TYWc+PDbXMsjKvnMP
BnRaTqgU+rIJcohjcyqDfiWSXV3w2nHU/t49tq89jUaAXP/FFetSk+dN17Uu0KcZS7NcK1Pt9nM4
gR7eg68JLZVCge71KJXeGWYPPIVuSFb+rxM1QtKiwXFRS/vJf7KK2bnVpep0Vwx+k+lbSnn3FmeG
Pv318TD9sDkR44HcKmDxpa8Oc8z6XEJPFuDKkAqfXJ04y/IK9h6kTaGtA8xh7jUzxs86iHKDh6ZT
Pwf9wOYVtF3CZfc2GHCzd2R0o+/cV2pl8MgzNom02YSd2ZCyV/oCML2InjLdSDL3n2SQKvT+YjnQ
rysuK9iJV1N/AY89djDv6VvTQUhTVSKcbznUvkyIBM/NcS8W9q3dJioINH7c+VBvG372VyyEaqeG
YPMjcmhKxi4OkRZFEgA/TXNw57kVhfgvypnonMbbUrf5v5hWJDaJEFNMsHgCBYxRsXgfd3dF5r6M
O+pPm3bhHuhewxmiuOVu/QFO9MgV9peUZ9qZTrc4vG1T5u1sVDjVIgk9lwpRmKi/EYJLSZX+qJkR
tlVZzE53lEM4cthPDZXWPkKl4LPzO+uEvpVZBJJPEekEty4qB49K/xSbvSdOPH+UI7CA/BzbIWGk
Qwhrx1rnWNEOfyZFo94k76dDPA1WryxjBsRbj9ZKN9JhPQjJ7/maG5pGlDAAMeRi2Ukt7eRlVu7T
YybfPiQ5ExipNHuY4/lUDLDiimVgnhrFZBADvCCvVvZvk5liNEvyciB7QWB7QUdYPS6/wEtevGGC
J3k+qISJZdfiDe+vbKklHBH302N1xrX7v3iOkSB48DLazzoukbZ/7yaFWAR84F7QL9utF+6wc0Cd
wwC41NRkFOscIwr7hP+aIEzbdQoLqWl8MybjFEhOBnfJ5nBAyhAEo/vMHFHzawISsDMq6eHk0Zvh
bQxF4lSVexQBNKJ6oBRQP31laRWBPZio8arspOWIGxQKuPMJqJeaJNw3AKAOulmCd4h+NJxBcffQ
Y4vQM4i3icKZmA4aNutvnio4QunPLIyXfxJF3K66XzSPPUea9SSvHKBYxYN3iuFldjtJCWJNe6Lf
TSCEDFI27BGu+KDZuhZolUb4zib/N7/rCWi0FyBzsaxVOLzZqcsIWSnhvEJ0uuiEHAUZCsBNcg8b
QpA/k1RhFwyxsYqzB/q1N/aAw1k39SIB2bsNtBdpO1dcd+u6sd3E8dQot9bp+2AbnDgcLTixHdpk
2/W7KT0YX2R1RDIzy5soD6tRTa94gMushGkXRpaHFEe8j5cPrim42ZuuPXodcqO7XBQvulBI9K2f
+IBAVtmnbrL4qvbcAWHoCmDU2cdS7WbmepBuiaWXCgx9ZgBHe2HZaCJMqWLyZRWFnBabucteQYt3
5pBJVVPU7q64yneE+4DtCz9AxUp8ayjHh6pw7oixCFKWtbvBNuKRHod8GLgwFhuwfatv7WjNHeT2
dbkZ+NX3Oqx2Kr5vaqaszJyPrH9vF9cPdhmgmvP5gpEsyb791C/UAWe7TubotqrhFETfXRiXVR5o
8MDJIUIeejzVHRmBhW3+v+qvwbzPsXPRSX5106EOJORI4JNM6ceb2zmPYE4QB7QAVF6qv/AkQhrH
3iDKKMDeFfBUYTtQsN6GOX0gEUQIWuM+ZEbu/1hbdUPx0Kuqi8eopN1hdAfPQMGOh9jlQsMzsQc4
J2mPjrWm9ZhK+0hwECrub+X+qogb+ZdXf9Unew3wGix2n46iOMyEPh2xmDjqfLEiGBmURQH+ck8I
G/QTpHXkx1sQUS4MfqWqohu6SsAP00o2zSf5t8g63SfAxK6iYN84B8XPoBhfwFXTfl67zRLCOuRI
Yh3Rgv+OjPYjwvvIHEetVgCKbGapNiKiclJl1O9hz8S3Oda/AaE6pUCYpDFgJ2keBB2lzIV0FJU0
5sVy7U0biydn/zT6Q3teqVJq7CehcO4oFMECw/dyYmwuvjilJ24Bv1mA6mlJnGthyamjxNaf1OUU
EwGUZiSH7DqSBeDY6/jhM88tQ0uDg2NJP7CXGztyhRuXOoRmUWJNSTsROY8lprUJikjQRkHVYP1g
xJsM3wFAbL0RFR2for3ypY9gqT9YWknjxHD/oSAjf4TUc/tV1a9/3uPrv3VrWABUdFrb3lU7QcLr
1POcmhG8GIU8zVfjGQ3B4YI04zZj4l7W5136E5C5WABc0VCRqf7JXEtcjxpeXYpP+9/uAHdRS2Bt
L/T4DInSd/Kf5PpBqbfe7EjDc/CHOmfo0utmWgLI8WXkjcGvcpKghQVD5UF9M951m4z8NCRr2K8P
isd6T6h8qwxU1IZg3J7YOZ4wrqarhU3Xxs98H9ShcWiBPJFqcasoXoNya5muaJFNOm5kNmXUNqjO
hMzMRK9l4WeA0zKlVvWVLW8PIRE/3aIw0UqSbVIYHK2a/tOcJ6loMdD4iXYGc3II3Ls32zvLRKB+
dRV9o+qbXSMs53e5m7wNuPwo34oLuogyJ6KvvgiEI8DBlHOA7sdZZfWd98xy4hC+/NolRhtFEMAC
+Wl+xte7ZgGi39azzvOxfuhhdAPj20LicB/tk+s5EirPfZFXg7wVVjbEyD6QaocjTyJHDPnSAeJ0
IrgKJEAoVTUcVyzJyoOOieINQjvjVE1JwAWgkJpObC6DQhEgBdRACcAiw6v+4f6sfkCA+EYonbL3
X6mUjKMd+VVVUuPbBGV0kOotdHfMaDv1NkUaiRvob8wu/KuJpdl6Jpdo/lqccnmFDUOR18JQ/fSU
tue1z+57qSCVZy0OwBV1DnWbIYkBgXOW/BZUymz+h0UaYbojWuAVmjs2IZu6VysJAyvmTVzsPK16
V/wZe+YlXpt5rKGBh7h+IxtI+aZpkxr4kvCb8Mdivb27VrDOI1FX6BA/wGhBbwJBex7LRMaBEEuL
GM2zn2ZU6RxpYNo9FaVV2/iWewS6bo6yeCAjJgCMPf3Xl8kg4b+wZ2MH7GZQOM64OIjgvxMLlY3M
xOwnV26H7xbyFsmubyl6DRiX/DZ0ssBnbzNwVLCzCGFlWHdsfySyBFcDqIBwvCbnLkkarYb4kP0D
/VPBN8fpwvkgSzPg4H/uZMGneWnAk537lnxto8sqgNoLr/fCngVFbiJzcvxMSjg63yH6Tm7RSmgk
zBYsv+LvjB8NpHQ10Dfik3bv8HOoMs+PmygvMDjdStAyeyIPreZsXOKeDRq98UlAOXd2RFx2C3S9
oZvoJY4DzFj+Z3v80UOK4iy2qtZgWEkWPq+QcVKpSn3sB8PkYqBqNvcxwOx/y16SJ6NeeqbnC9CA
a8Sz8mkg7B+vCfL4HNHpg/KqjfWcUAddJk4FP4CsLVDM8nMIfZgwxNqqjv1qDGxTHf0Sdg/xXo5z
HrANgX4NUjXDG1SVBzIJpZBHp5wN/Qz2cAHZe6HB+4nPXUqs/UWA+grFgu+f0Hh8apQ5csPmy6QW
J1qK5og8IwdoXgcPEpdcOCZIsmxChmR9JhkzrzHZ4cz3Ta2M7KPwAz3l7eCAXi3mDDPOuae6/fWN
YU0UyKyA+h5X6TUF3YH6xmmjjcQEnZkR6Jt6ijljJol2ijBTcdhsTrqMzCbCcktHdkt2XPQcye7M
bJW7hnei9DtSLG3Q6XqQb29G4/gr5ecEwqMmBPz69hgctlhxYhZhb4f0f9BD2Jjlgm9ujN7CqTX1
bHwauVfhR3Q1MFTmDsQkuV/Evz3EDRnnXQ8j6pOqrhQxgbR88XUKDNvkLSt3n1ppGrvZH/KDG33h
aTP0P2pYYRc33ofauY4SUsZtz2uF+4LjUP28TLj9Da8N65KCcSm88zhS1Hg3PANOsf9fiYLhdsFD
gGx0Gxb2KkbKOzchsmhpAWr+aF8Vm+YT9Nwj66zrx5nw2wdPtRwboDJq+/5ujGOXifZZwTToTKVh
VUcPzo0YcwYVaexGAZSGknykPS4AMw7uyecieBMSof0Dwe4WzLy+NhxUdtLN4o4O4jggKPTV33qe
kP4cHIsXr2xg33y3cUAZCtVk0EOBAbZm+dPg9FTZ/1QhxRfKuTTJ3pzfDusrsnGFVraSdwDCHB8n
EwleZ42CavdPCDkBxUYOr4acNlVaqxBM2G2Qgbvo3Jn8iTdICZaYD0L3DMQTAoOvqB0naK1Ljbwp
3K4iY4HxFvkj0q8NoRWibOIkgVyXOj8zgEdoRBg32whwsIB1lnuZRDS/8OBHdTgfTJJTYR2jPp0m
OcZwq8fQi6HCtNkr9/xC1KStdNYO1EjCvPxAo55KBqHSp/RB2dPnsMxEPbTwDighMzmX0HRCRTGa
D7wIqjx47idR/qgLVOeDwZYKG1DYKxtVIikyWtlFYaKJl53l8sexrBBuv1uiiLLL5vjZOiWPds4S
WnWqUUucOZER7HSYnwhNhHMvnnsnMfjRpd24QBAgzee2luV+9n95YGOXS+6nqpaFeRraGMSzBMLY
M3KU6hibuI5N/qYDkyOP8tvq3O0tbOrEnOlRApSTzl/32hXUTpJG19/726+gyNV42ifsZ0SRq9m9
ovnZnZQ94FowqR3XXeKoUYSmSzhoMxq1N/i5IC237v0em49RTZQ47Ge37wsd0xGnqC7Ecy8iXKj8
qKQFuABqLiO5QDvv827OJY8S1NNSLt82kOVunX6cxcw7oP23fKPtsrZj1c4vZbusVzSL7rt9TZqy
d9XqmCOAlL8Bt9Nbx5bKxPt4L43McDReIH0x9V+TKssBg8c40RHjLSQFaoiuzERBLiCNJImEFq7p
wHv2FS9QouxnRmdX8NLg4tERZrxLJWcg4nRjYZtXPklwes/aK3lGDgdmbWQtOPffedkmzrgQQlIf
BKNrYlQThF6PbQ7HuArQjGBty1BvRHpFo+oE0ivujNA7IVCOS2hCt5kCM9dNt2nbERxZ5PBcFuNJ
kuThQcpZQMkSYn8s1GVKHzXkd112AAaU0qjPgJVjyOvvBuaBOSNJbvHavd1Fr1psy7WgymW7SVvA
ANTabIcewBN6D1eblxPhWCH2TbmsUf53/NQej5rOfcoG1CNuysjSRFIgbgrSmqeUdPnBL4Wi+8EM
3fHcmbPVy/sNXq1avWMz+gcYJAV7m/I/eJ2HIHLv9scXab1f3YyJgiOcwXYTN577CoROfRJuQdsh
2TiQ86357NlZ8kRF4QHspYlVMLp+Hh3GL29NLrDy04clDcTWSWz8w06cxlYUIne6xQMON6OWpm9y
JokHxdYX2YQ7Ai7CBG0vkeFGcDjswLM7B1x6TL2M0EyQE/MwZaWFVvLmJtUj3qA4OKGsu9lK5cpp
dfICKx24lnGECogTYEj2wSEjN6kP2xRU7afpHr5qXskg5OuJmF+ZwqPuWsphmQgpJhriNkaZp4o8
BdGP0EELUjeyJFgB0Z8UCfJBJ7XN/LWXBNx0G6TGW+9LJaCRzm7LUZSzCEo3PVUjv1mpKDAxBMJI
wrs2y9areHRgU2gZDWAPklrWAJwTHa4l9aXBtkLi9vZdZX+z8yJUoX9NqWoTljhwkKsKVLryCz0I
ozX0TPvf6uMly0kipYFt3qxjdHKFjpoeBzi3F2xotq4ADjNDytYv/tUiOdQS0ksddrl0xVhl01+p
qZWTpZ68UBWLCjW7pJ6IVtpomW8xwizvutNdpb/Nr7gnkVIZd0b6wtXQPBpXStCv6Op6+CnbyOZx
BACvqcVKJz/l0c1WmhnR3RjeN9dQ0EN7U3cThT5MAky6JEodKEoVC0kkLljjWftCi+xIswIXQuyn
Ggbsctj0lTBi4Y7aWuHBh45kkM8G+9sjC3xg86y0ufG+GNgSa/xiQHxTNbclkc0DgJHjYefwV0e8
V5xhCA+rQ5LyuSpeGL+IZgMa7SmPmuhz5h9GrZcZfebi0nx2Krw2ZOGq+3p6kQBFh6BZTLUScXJ8
IcQwnslZo2pRc2DGO6mZovgijyDA0gwHrn4ZuxewoB6cfKsntbAgIPz4O258udy4H/OsNKbkPQ+R
O33PlyjJnoXRYpwXtCKjRvXlPHqMJS/j7CyrLeeubMtVKrXq+Sy1xKB6bMBkHm1Kc2fQSIjlMrz4
D0w/INOR7cdn7dtb+bo3jMsikvFhLCqQOmswelFVgS29dltsGSTcwlsFO5Ls6+aFdzvKj7YWTbrL
+ylfuRAH2o3EJRK9OK0mznJ/9VMu+KC1U7B+yKhDo/odiNQ29/VdnStz8uZ3LpkTzRTd+fGFZWKs
PARdDc9rX7qbqarAmLxH4F5jgJkNCexYRIb3QA+5JStBjMghxHTeIYiTWKizZO38AjVgUpGkLjan
FZlR69sSytfISKqDPRvtumslsj22TmxVHonTObC+TiGN0HN6oeF90HZU1KpJXAvLqB7QXjDFLpSr
cVNHtTqw98XtJZDZ+GXnoaRAtikkphLBgHStkSAe10icVTQ0/UVsXPu3XuoBxuIeaNLAmPn4P38M
m/trOOwOTwwRMR6I2FJ7EsZR7FMjvPVUuh6C3WcaN4/H3dOGUdNQEGv8XEFofK39WAWMGXrPPtpF
UaPxm7XQWdhhNvV18oBPSmm/4QbJ2rLXmV3b/uxlFzl/uSmlsB0HgosKPnH6H2HrMNmgCc8sy3VW
HQaoQR0nQqV0lLIZeneUr+2hxbjuOtbIKlULBWrAaKMZFfjgcxMqkJ7WSkGYf9HzzVlMonsZHs1H
UoJd1jdx6sHCI8JcHGpgFdaPehHhFNQ2Bn4ythqbcauLde+DU6kQQKmRH0JUaI+mlRdAHpXZ6cTt
h2543KSoKdOwVRxaCjuRvUwLtxWpaEkBQWhsZzULGwfJwjgNVPv4cBjqWwuFCUkho6Qx9PxqVGJI
+ykVXHTqzCrl5tjHV3Y/y8OKJSSpqJTvUf4hpH625d4sX2jeJGeIPlyOJovHDfxOGY5CgwaHS7lA
BMyC+aPcjjVKRmq3akazz9EfdELajw0T5NxILJhQ5o7xlPqOkN7W/MudYsYbkGbrx4nww2aXwnkd
gqMPE1wXQ/yW9XK0y0RrJYAtLUe3anXHYuML6kZD/qziz/8Gc4I84da78ZojavWm7qQiKyd4LoLn
XP3xwCQ5paAjaDSoCvvlrLSNuWcpHN9H1GckGaBpQJmCvFhdeh7uKxgNHClOoVOwUpmxUGezJEbW
hMw0LhrKf7klmJX6ht+YgKYfUL4gpny+6hlFRYCf4QNi1EcZu2NQkH64liHP9PAgv6ygPPNlVZA+
dnGJEndjfFMf3xdmnQSxrUbxqlui0z12X+lactaVjLPfrRu32n4yNq9eS5d61rmEFJnVXEXpoiL1
khzEQVYt5txXpdOV9vR6caVF9WcbwcwELkMooHtftBEpcjNJEA6GX/7f1r+PrU8FAL9ohKecFjzt
LqdGj0qkJXaPSMZDCEvLh6ftd9EpPVc/m8qz9Z5eYYHR+2Ah9S0dwmEFdNGG9Y5HOkkQJFykBSoF
GwInEk6fQhJ1ZTXP/rz7arhGDJMDekSAi7thGxjjXjLT5s+eFwpQognv81qpUIqQbjgmcpE6lMU6
akXprqtuT5p3B5x6Zxx+vTL1mOynVi4G3sYxuXYLszaKvmaLN71FknJ0PVJYGX2cCKVatLSM/UOt
6tMaT8H+x9okbUhYU7rXZbAD4gyNf2oQsT1m2x4v0DAynLhZaFG0m43yiqWOPLUVRt36fEnxcDQa
oTMSTQ0aJ48WjMYnIk7o19i1HrYJVqH0vvDC6yc028YnCek9f0Zm62cuL0dJmld1DVZL31lbY3tl
pE/R/GgyORYVcQNCwmZYJfDyjv8B4MycsKjP8XSsMn+Rs9nDWdVCcdcnWoNJSolt0fyVnAOO4b33
Dr7kGVpVhFWpvhuGg5Mb+hDw8lhljui+mRm7GJHuosoyHMZrF5lemS5F/782EN396jJpwNiKpqRJ
7lmHLzE30UnLutY+J9wS/BKlwrAGjo/WeHvk20kNcYgg+2q5s4Yocs1ZXxJblnHDydni+Y9xDR0/
GCkNnOFzQShnzk5wrqlY5g3w5sjgRgJ8jTmeE6v1dCa/hAlEKMdwn5qoR5S2H8UFP2PRaFm8q/Mk
tvFx3DyPTeoDMIMHM44pRqKVL8V2cwPbHJmzuJA3uCc8P+HRs4Unaf4ECw3Omx6GUo/MSPtVEQni
Cl0CH0whI2SjgpISUNOPDEeoJT/03nB3iZYzmCdlF3fmGHn8hHEiTXxJlx1z+fb0/jhGxYiVr1Lp
inupyTjkA1eBhvLCHu6EMsD722NEgwUGnPUuJ/mIO6iPPEXqTtnRmlcZuCIgBg217W8eZNCf9u7I
PHQqLLpk0KmDrbgYeM3hDjJrCUiAeqejZtXS9T3okUNnrL/KpjsRKsaPJ/4j8faITF0LOtVNBM5H
fJbV7NZ0JzHMkukObJaeWb5mgztG5uQ+GeG87RqAX1rFnPxQBSy3J4zX/oNUoS+2hlXBqei6+wej
TSOuQVPjhotoQKP+zFpc4gVC+9Z26KxJg9MI9lCJTwsrD6sSsJAiCfWl8rdGZYDz1RlXJIQG1Vss
396hibQ+KCeChxhcCUOwO0QVkt76peY5Ixhdnqm+Jau7AgWIu3vNhp3KE79jJ+X1/VIdsMBdD+QD
/Ai4nY4BuDULVluhHS5YqJ9b6aBzJlg/mjaY7mrm9z9Mt7BOqXld6wkxK0uFpTpAfrLSEVQqWGzI
lC8xhGyGLIQLamPIVM6P8pKEBPPkzFfmFPP26ZOme0vNRwE4frIbOv/VW0lJRilcC4BXRBTozxcS
rPxIJ6C2C1l4Nzj09NtaVLkPYAgqBt/kFyY+r0LAhWBszMVp9QhhXkYNMW/k6fwyN1wp/YCCbyAr
i9ym/J/GjMt/w88sGCghOZuj4IfJAo42z39CszVP29k8Ti+PwjGSHZJR8E10HpH+FZ9sCui0qPOa
z1c5HGrE+WL0jZM5S277MBEkAtp+xmTFJjJ4uRmrCznIJo9AFHTYiqHz9A+F+uuggsck7vctyGU9
aasv9EjzWq/NSxqsik+56f5i7WSD6q8QbEnC3Roiz8K30W8d/ZID3yf2HD7cygX8hi8vUMwJtQIp
9O1KOySJJ8d1IzZ3SLehcLo37CFGCRiPsB0Ouup/h2bR3skdJaqRXEbon1BqYeFWy6g0adb0f7i5
PLxonMo8L5hgs3Btm0qHwjWw1Ir7BpfMXdxoWVSK0FDWBaE+ZfAZHa1T5yj0no+fOf+sLHW5KY4c
/mcxWCqNukq0w0w6SpQHaQhaME4liYitiARjIOPL22ZNOf1KpqzTrqZPIBVmhpKbunqiE834cltZ
ALoKro4LkLyg+SyAKCi0aAPtXtQgsSXAmwWlioRHoKTVTM5Cpdw7RgfV9mQ7vndogB6fjlvfIY3y
1717PpwmRQikLdiaOlisu+Tm4HGJHbPy7pQ1i4aY0zTF3y7PpIt+KEDm0CHqGgMszbVNGNDdORx2
FvZIwgrMJjRWdRuPjHzsRebh/3+QGtsY8EM6EUdafr84JJGeZBgv77xTPhsYx/xjLbLOfsuf0fkP
y5zZxBRoYtPmAcrDMBHnQpWsCB9OCg+KsFwDMfe2v2pxwzBvB5fzoLPlkjvRsbB/bN3pHYIWMEBd
Cb+dNYi6y4xW2h4SEQ4OG5Pk6xJXqH7mnqan7qQGFNnv7TJ6sMHbSW2I5nsjua9RpxtrjWCZsu3Y
15N5T+eXBbN7ePbMzLLw83aq8hKMd6Oiqu1r50+cd1m/KdG6EizGuiRdKypTMMAx0AFfgPIta5zo
6vr7EQLF9hNNRiURRYbVXAQj5N8VoHJBTAHYB1whDRvnnc0O9bLse4lJn+k3o1YuuWmK2EvUHl7J
DLaEs2pIziGRtMXMgiWilwLc+H4aaRzOX/o4r6cwgBukjy9fSgblB67BIkWBnEU2a6fUOV2RF5a7
QKhjkrSPV2V9qlvAO1lrEdP9NDUnJ+0COcpvwNES4zykkeX9m01xTLr5n9kQiyBu7Js3UrEBmoCl
cvhzUmlIkWtu9o/7qOhKT9duhre3GrKdN6XkONpusxuSn1MmB72sh78fITFzb1ZWsPS9Hyv0e30C
0iZ18CNof2fWUx1DNk/L8GTCu6yA4sIqtp22Yt2xA8T2Y6f4PuEwKONriuRWNEeLostlLW9v3Xdl
Gx9lGAoMcM0cz4pSXcDxYjTu1FJNqSbAM/hz9WPUoE33n8Nu06meIO+leZrlfeTASPuhuj7Httfg
dn6iW7BN0/E4CVAU3HqH9wxJI68lSlOrSF0XOolxyEwSPzz9rHCJxq7bz1/QWNaqCh2EAMspUOuK
xiuU7Kk3N4dThhJ/uHbGvv+2x57CjyejVT5RPW1ntrF+SpaVTuTZGeqvNQ1iQdbNx9XcP1QDcxiP
GjfsUjs7mOEtYYyeSfBUK9cWg0A14Fv6f5s4+0IyfY3jUE23ZcD9x8Z5xqvCwO9plYAG92dwJKY7
iC1dGpiBUqLJQhI5yeEnB6w5/HzHnL24yDYoMdA2kaATAoGy0bipjafI0ZPfliZjKgC5BH3gx9hA
ULE+zfEGNhgTWa4mMZYxl0I9R3Sm4F4vUU5p/AVuFhSR2dT3nUBN6S3FQkcakvJe3phnjcYs19eN
TaIr0x5Bh3/Thf9+0oU+Gio2K38re6sOCAvoWsEKTGL6/659P9CGsxSL0prx/bRlr/0+MD4S1+Lp
9rB1DwnwDqUWo8Ey6nHsmlY38X1eKntghvMGRUQeySxHdm9hO8Hn1tN8SX7Ftv8HQKrdpU/sKnj8
ozEqudmNsJqMTWW6TvjsFnro66DVSiQ9isOG/3pq0600+5dMkgbyH82IHybs3m8xK8iFMUWAljzA
/9/EkklBu+IZIkvrmoEvcPNdq04tTDSodHRcEukM+7d/ppo0kHunf7ZjKmTqGHQIgkjzyWGQBqK7
ansQDkvWuT3sVVNIPkrYMDB6MqYYIOb9JdF7x4e0Szar7tiuaxh/p0u/jCGG3rR2vCXnfAIzcPie
EHvOCTpIz2hhliSxqGPoIGv3UHlOk7YUpcFB/v92JYzyL4VFyWhO/X80DosvaehgswU8xzPHMtB0
v6p+CVI0bOMHe+7j4UnUnk2aNoLzSlaYxBniqpv//wJbhszSQEgDq7itHzXy8HG40VGQHjqwUYi/
nHcgyMghpTsYxt98JBRJzyJhqI3jpLQ9zkYf6ytYVsTpQgC84D492/GdFlr+a2kj6exut0nMIjS9
Z6jMqTuJcbgbEkBY1ofSksJ4Ur/vIEDSQNHbhMxNYfZ088dNndmqXJkJBKpTqlel9Ql8sbEKpQcr
wwQRo+q4erm+1FJ9jUJV/xezM2XcYgEqDcfsDxasgK1Hj9EEW3BBNP94OxYa7ebceG92bzwYm7jo
l7CIB2EyudAK7w81raDe9wKqx4iXLexRATjkal/2PUcUhh/hemKvtUjf7wtl6l0swRJW90hSRbza
fCYbW0cx9J3DiZVvQXNf01vKzgD7pjX8QbwUceo1ExHZifuhN3QqjmpzqHZ86rqr/Ls0Vz3ynMLS
nJF3BiJW7/8qXPsJ6i+/9naNyVujY7A5qv9O/teTmkuOaRnxvNdxuUOqjQKPSGhHKu2vDnNJf15S
wQGPNv7ZXsHAoR+QPtsfACLrgKcC0gkW115Mt0q0wogBPTdSBs96mh50WjBb333Vyc2Qp8PktfXB
7pEV9VWQxIqyvjkDAOOaZLA8zLJ5lkEdOkWixW1gv+gEnTTBloCZWZKwRvRjry+B9BKHcpzBtoXl
2O26EGf7YsVYQZDrVJKs5KKW7R6En325Hq7A5oaMCgVy2zp7bAGfp1ehJ5oMbK8OxvJ1HG/kIJPE
7bsdLTpXJBKfQfw2GYvEI8EF0UKikS/yrjvFd0ra3zplCjhAWbIAUL7jKoe59pT/FagsmCThNWpY
UGsPW8Q+Bo9hXHe2dDmSvfrZXt/CICKp3RWmDeMRETMzf3XLKt9dCuFqkNAWe+Gbm5je3DCt0Imm
EChcs1WpSBaRYuvfS0lTfb7fwmQ5ns0qvd3omrn4DkYZFYTgQIieB6UwcIfUvcwodgAG52CHHr2W
cVvsiPLcc+5W271tbrBYTlLyUtvY9O4aOfYYov+mA/F0leppBorKyAPHv9pqV5IjVJ8OKuxcVlfO
kzIjzIxGt9JmLX44I5l1lpD6XQ/gE3v57a7wIIcGA5R0WkpTb1kKQ/KlHQPOpibAwxkvJeYJjgoe
iPevk4PmA6eYF8ZuvTKcli/9LNwxW2ZVrOZtY+QecW6e6Nfr5E3lKo91RszaY8XUrej9ZkgJFkm5
1/vEYebe6peuoaObl+vzTdu5Z58tVYeq8Px6gWHUAzVbxrOFGJz6zJbnpUx7ilSblTM/7dzvWGKZ
MqP79oS6uC4suuk300ykNH2aLY86k0GFbb5yjLaXs7vgeCXIwsvlDg1uBweWZQ8IQulMEBsAUlTa
+SjvNDiRe+XlZ1QnB+VqH+uj8MK1JCLuEh2GrPVYwiZ4Qbz4aZxUK+zDNlnkTgr6Viy26J+Q3sdj
n1UTgQ94/6ExvItureenHFH1SgdNiIwSz4xzQAwADy356F8CKpzxxd/mSImUIoCvwDry/Wic83+W
22zFoBQrylgCW7ior80nBrqVYjw+BVUe+hWlHwEEcsz3njrEIoGYCyWbkLC1IRl+lSZ0aIFb1W0y
YVDss3SI5OByt/FlIolGUtRTqLmV5sYSpMuO5gFgqjV4a1hpZMQa8oOA8WJF+e1dLNosEiey8IRB
lfIsAc461cTpZxv/XVZXCQp/IDzmffvjBH1sXbWXZSpETleEIx3uep6s8MRNDUnex4LZIrfpj3o7
QZGrx1btYzltdjwQo5a++v4JyS84oRfCAknH7Y7OG03PPyEhE0++tMmSnTXLw4NazeCCqIpxCdmp
QhIHBbo7YU8Xcy+zna5yq/36J5pPXN2gjffI438Gwu7fpgPZ5Kgj5wyx89gVfmv9WT+VRGsQ0ruu
nM8MO5+ob4LSqVhrw9leON/borzUvtoHpR/LyMjVe4ls/FFG7HDFjqxQRlQo49Avs5Ch99AZO0B6
mQud7oT01CDxF6L87ctLLv67vO+p5C7EL/ciCXeeLzzRxFHC/HMSO2ibam49CVhIoqbNnPfNJ/c4
+vMadR7iqQYa9Fvv6zFYpkqWPQyfsqHTe466+VaMssV3Ziscioi844fDlQUIHMHJ6s0qHjsRn5ds
7+p8EQia6iA7okCQl9Xs2HkezOdGjxYD/nJnO+E+WCZE+dUv5K3pNQDwZNbPDPwUhlgW1lEAY9n7
LGtA4RSQKkJ8uugikBWfSL4Lxo4qYuHd8oIN5FEzHN8fMJmCq5RGN+/MsYe7RVUXxm0/ax6lYkqN
WlwaGNBls/Ck7WgOIsuTirEf9k40fNuJWHNVGwqMkrvXyos3r3ysyhjo/UxNi9WgnRdFfr+TkmpK
D9b0qjtQ24y0axsvOwEHvsch4qQ0k59ys0o4blOrUFV/66GCnPV2FkOmw7dF7E1Pg4JcUNFTLybP
+nZ9vwiCJ6Hd22IRhGPajbw8iMXEKQjT+9WY3dAjG9UzGGbM00swr8uOlsdzJNOMknvTvnacFV2Q
yF5GWiDqxgUDDZEuqzbsPvk04d1iXDoTFHHaZkRsa0xy3QxF2/ypKdloyH6noTXF2j5ilvg/P7QG
46okhDYqKJV+IVupk04Vq8QsbT3qaJx07LkZtMoyKhJl2Z6BDUEvSLiaRlcOoJa6eWMqFdFQRckw
UGfhCBzcJDDIYua6oq8slreR1o1TgfQWnP4sEcTfGFLjaZ3PmXfZW23dgBrH5LbmIMbc1ifGjwDP
G/mHIHUZyYXQZ7VlI9PIkLxlnLVYHs6/wG/66tLS/+V9B/0clvYx9HEcWkaHq9DiuJJ+Y2k5h7og
eIKVS2Wv+YtQQMB+q75vWJXc5exVUdWnufkQ/64LRjnPqblxletDwB0dv8b86GVYqy3oUZb4Dl8V
mj9i4tzfPTkckVE1R03MCH1Dw/FVwtEBgCsA/cV3s0ckrV1DIG6w+OTwV+A49yZB2yBN1JOHZxJR
uxCLI3XuwcqjsU56fNhqBpM7vqP/I/n6yJ6NTXERyI4ETztoYMgiaeh8IsYZeZP+C4UbzeCWBc7G
P1furyAnPgTQEwxN8cF7sRPlGbq6j6mGjiS5Nlf4/gS2jY5FrKgjFTdQktEKUEl3CDu/dZw1kaIp
QEA9pEuYHeO0b+ILKbfKG5enmQeqyuAMdxVK6TzjOV7Ef8jZ02Bl50+snEc8fkgg4vg1u/v8VPdh
1Q2jkA3clQ35j8nEbt9Ua5MBWckyONWsUqvRIQQMSGJ+FlAQKJ19wxzlHX6vNwZa0Qc9gPwNJkA1
f97vy4yCwYNAl4pNiJ40aJ5wVeGCU5GNfEwySoAFqX4RLu0cyjZfGH5jkes3F4bDGIi+7+AZ5WFb
2QAOjcQ8vezF3gsH1WQxDfZTuLgOBWj+ZdbXIndXohrriAxXCjAbJ1STYByG27hliWV9h6cklHi1
TyfUAS8aKiJ4169cuM82UsAqToknjLyFSR5q1q+4dwQePl+/HgP2DPKlm0RyUdt9kiYuknCzUFpS
ZjcAc1DmtS59ChZyHrYUm5KeoI7US+SE48j6kAFGTajRZknqcHcO51KoLWbZwf7XxHtqCdz8haag
DDInObb5qtVcTPbIcq+7RnBgk4JrjAOv9msgqBvL83WDNPBpCcLrcHVsWUn9zOxYNsVRJKOcEhrI
MjnPvBdbvK74gE5PbI7DTIEQpBk5o7KJMDWmWeoh+7fV19A5nHaMeoRHLS03fXGUxwtwHiVONkoZ
Ve9ttKZWb3QAgkFkVUQ201q5m4bRopUubS+d1IkSyM4+h4PTzRcTAu9dHLlsS7dkF31YO86VfDgk
ZSUhh5i+y1+buhfC63PEBeQ0poVpymR/ENhBEwbZJ1EQZ+/jUqlE/yVwV7Zk3q6wUA3eMbfWO1Az
i7OP6NUmxp9MesK2YBGF2Tq7YR5bS5ZPaCgB9U4mPPvfOLLibGuf/rEhH/xV5DHr86ma1sg23qC+
NOqA2kRo/LfygS63AYogSzGdZGy02y/hg41QDEz1Z1T7REgiVkEYuev7PXGEkaOB2yf34NQYlN3F
zaLnLiANlUsdDvA63/tl8P5Fqpv+zYAW3+ip8gLZN3ImlMcd3aQZw/b9elkwvqevFkihCLvHULqU
IchPydkNacTNU2GBJRxeg9ZWdZJ940VlqNPdhy2TJw7BDCcu3+hwgY8gIugngIroP2sP7A+bKkR8
2WUy6anZcEyEJgBXqkhr7p68dYP+MbGt4e8ZUfOV3nNggWa0DWFVwoZc69jo0aqnXNo2hc39Drla
PzDWAddEqTgLcRPEvIaFiQ8aqZmeM0gitj/StREbQhS1MRXvI5Q7C96cI4t3CEHrXs8Php4h7TsH
mLGmKRiPgZ70+CWMiLR33JRRMvWLC5toTcMKeUXETipHDPTLg6+qiBx9Y1fSlLduYlhxgeEnmq9D
CF74uVPIxvbrCD7R8vW+1PbL62hvRkdUdPydjFFrIgI6twh3un/zCPFlrLQQUyWLHyZmJTwUqn6o
u5oZrXPmZJSyU0cO/rBLocQKF2jMHZ0VXlo7OhJQdlMXofFk7fCGWpBUm4h3sps1zoFDkYKnDGBI
fbSffiYg/qGJ2guZNNhOuzNk3URfGydwCiircIlY+Bc081QfYVqWxeA8jMQ06PtdiATskM2W99BX
soCow/skpiWhliVBU2Jl2FvaVgJjLm9725lB/4K+gOjha/rItT4YNrHJov+40p+fcCII/vDR0Z/z
xMcEB/ddjl7U/zelScBMkzxDEcXfx+jtF8tFQcT1s+fbChtQr2tbm81EYwdJwhaZXBr4Cj/BspdF
dDVUtDAFUhrS7XEN5SS5+A4lSkvUnMlQ3lNxaAgd7XEU4/lnEB7gbzg+t7zDdZdzWuuLn9A5EnYL
ApKcAv3qK9lgpL7UdJmLPeMnAbRcYx3jjxr/zBsxerMlWfneUxuBY8Y/Ep+TUK6MyK1TjEd/+/zi
ui3yAYT95DY5j6xTOdgrxgfncYL8nlaiWhpsLLGbgXG4xp40w0P8sUZeN4a/izdjdrbc76WE7NBR
cIMAf3qVwz6/rElU5ZEge+vs/46slG2PLHmCZSFIKREKLFAfO16/pSI7lTstQPR0HawYYoSylNq4
jj7e7v8KE5ml1EfYvHjTfUChwZkh4ebJaNLzuAIAsKopxlrygd0WKkbOJxgBrO8DmlslTKTi7sDp
etjpQoy9Y2/W9TsrPSuM0QN0OPirivuWHMDCPz46pL/x83RClM78cCK+Dk1RDn4CFqgyUefWhvpN
d4W6YEidcdpTfqxBRS+yzAvf7hV2rJlUuC5+v0g9nivf5JfC9B5+ZkmL6RHjWvUsEEQ6qj/RdJYA
xxvKSahGe3NF+CPlPRp+/hgf/KXRyfvPMVrggLlwXDwvkoC+cADN7Rft2NE+ZMJna6qMC9jQ46Ec
JdvU4bW0zUUcToFeyK/NkCb6KHRl1Kx7yWisJi8QmAAmKtT7RfnVyn/W3ApL5H1eAdSK5nB6K9hC
cJvBpM6Iao60PDuvlZWWyN+bsQe+h3vt8v94aqxX+3X8/FolAz/QWu1JV7eeRWyLZGLGsqcZdrE5
11DQ1rGhIxk25t8PMWCzUMoa9n8f54LYZa19Wgh56SKsrnImdlzgTqHzkhPkjJmsRSOALzianfwo
NyEIL1BkqgUbMixa0UQr2V2x0bTQNsPFlAK6xAWtx1NWChIV5pMdYZs6hJIBuUT2/WmbPdY4UhSj
B3TcA1cxlq0KI1P0fn9XkIkMJhX1jrMBiemBfQPAusILUMYUf5hJIi/V3ANC129aY+5n0CFBSFRL
FAB2ZWLDOot/oO4azAb57YbVdB+YclwitoaULfG4jG+0URFcgJ+nDEZ1Ar4yebe5YKWBONH4izS+
DI2C0+k1pBl0di9X/sI+Y+gucnqA4c6Bdk7QEwMQM4KztyfiKgNVYzRHWFbsS0/seCTARPN8ppu5
kSVLshF2sdspqjR/yCqlBrTG9Oo9ZKIFftOF2CudETad4itft/vsA/h3q3DO8RrMHvmJmcb3fN7X
OSYfamqrTOV4hfgg0C1AviyxxAvJx9osTUmsQSojQI7VTHJ0KpfBN9IObpzp/6tWR3gO9TQyuZRp
XXNYo5A0c0vY4TMSyZLj279zV0WHl7q559xWJzKI8wrkJALrRJnmhePxmoDnPas2xUoYNcAgb3YX
T5miVEk4g6iXIFt18kGQe7+MIJFeqv465ymo9Qm+d8jn3mmpwSDPz7REkwvwEoo+l6iVdKaRKU24
4qyfgKxgDyuV41MqlROZGnWB5QUcO9kYyk+CI/Wco0D0a6Xo9QKgbAfJSHc1fYLZ4rnR9LZAHEvX
Z/TLImVAf9lsXH1uJIgxfcXYuunfCIV3Mn9WOupiUGAf1X1Ztuq0ldKdfA/Q5Yuyr7lZHkH63ZOv
ilhj5HEMWgfJce9zJcvKVlRcV7Iq4wH8UL5dyqBo7csGMMRm0Yfnl/26q4GvO31jmmWbr7PlrK5H
IBKYttENDEVsdJ6oNel7jGKqAJ44GPe0NdOO+3zvD1akzrK9XHkaFjTCeybAlAqVeKFwqanJtfr6
ywmEOeFNefmI4fHz8aeawnvvl/HC7G83RaDqFAovheGlxIh7kOorCp4u0KyCe9cZv+ihz3iZbqs+
di+Y2vrdH3tAPhnQiNxdY6LWpFLbJNI6BPDEDbEnJAfxS/LL4v7r8Hkx03avAV5Rl+mi/UBUxOL5
IucITLXTSq9MQz+MZvLa4uOJlod77pvqOlzhPgNzK0OeI1r2mCshDEmrylv5mxaoRbFFhg+la6nK
6gatH/bUJV7iazZl9Ef/sgVBXQ1KtMCSeGFpdHV2IW6IEYimaAoXYRijB/aKpkq+Ft2crsU7HZsR
L6WzxkYQgrg51A3SEXWluwOcnJ/dDCk3jE/mXwIW9/vMZ9meKlLFhomr0D2Gdf8tksVe2wVrlFwI
dDd86dV6h44vLKaOuZtdYCORuGCZfEsmYd++c9+oVs0KCvaTYRaXEboqwA5/0gr//BKnEHo1Xl5J
TggM4XQqWaDo7f4PPaf3VFTuywUfxeOo8+WMLmGNynXSPC2PyjI6F3RvEsjooTY/xdtcOIHppACU
i26h0c9izftTCAhsPq2hsuwC8lRWtXN+NEkoZODygyi36yScXWquLt6xgdckRm+YK5pYIFT26NtZ
H/V6XyCjaNNQFYgKNJXHWHkSyfArJb2ogfEl7GyWCpp83G13V8okqoiT9UFW8YNQAvQuaQb9OBgl
vvwprCwaRD2dWBGb6UhkfGal1u/oFjNoOnp4zephgzFBsdPKg0s+AUyDurJbzCVuLKwOlNeJt3xF
mO/D+VSiRuawFt6kjzNBUjn/ODw5XQg44WrzYQe0YcLxuKtUTk4TZSEcfrcvsHZnrDvjtiPHY0Th
Dt471/7Tc/TEu3acx5E+FbOos1w3cpOUHFUbXYMbZUQFrp0a9yEknd36pT5d2WOC6etRrvCdpm7g
yXZRCTQQWewSAfDlGsx/TsC7LDc9IIkrVcz+x1+hwbGIqaX91yT9J6nosyZp1UlNDWwYf0ceQmPJ
jUrfPj0oLIeecQm+gFOCU5OdLlox7sKLnL11V7FPcOC7ml9u+2HuJc+vNyOtWsRJeAW4lE284ZYj
TDm1q6tZQMhIvIT/kAGB8W7wAtXpQH/VfFB2CB2I8Z8d6lgz/huxqpGbV4JJV1JGh0OwR3k+ZiSI
w9kg1g5AVuR+mKX98GNf+uchIvT2F3YYXeV1Vhj89gxB4STuXsxbVPv/P5GcbFrxfgE7y6V6cwLH
2axgRxw385kuZWPRz87UZYmkmseyM4C/276LOoB2gcRiZRC9d+MG7SH1NEiNOcYoVkjH36WL+5pU
CIBq5WNiGiy6aL8GtlTkYcXX/UeGVBbTXSkZCri6IasBOtKIX58ylzSYNqpXzXR7ByGLykBa+QiG
A2y3GnyZM4CdyJni1DXLAVt1aXRHEjfRqSI7j0JriZ7qcZQFb+gapHO+QH90J6RO0kRrITpAdw3T
ILgXVOtced52w1B4lYmEI79CqBYU1Dh/fhSvxeqyGMRpowPvSXLwQfpY3aY4DH2yRrQ3WKTdmBfD
BQPuC5tVioMSN2MfZuP8uN1222Zjxsz3VYHCQFKv/oL1ExVAFjWY47ptNNr/68XrC/VAHqwUDx8w
NUWgElMjQcbUsr+A0u33sU/TGmpX8mjrfvi8vsHEDMykFc8ePV0qIn4Mf5YUjTpP42AQJtt13scd
xsxnSv5/lT+OVERG/2TjFbBHhIkSdIGv4aFfEkG39wowfL8qdefUCtl8TMp9RztzIJgozoqi5le8
mXcv03VJvE6kiurjdUixNHrvSInP5gzoTPZnAM7eZ+V1E1Mq4lYU+aMz+OI+bbwfT4OOOL2Rz+CI
oz9ou+cPwCubRs4c9/p6c2KRxWsMK8NHB6h7QUXN5lM74Ys3ao2iKwJ1hnP4voFPEIcR4Z1iqgMs
hYuwdJAEoVSQ5hVfcThrWqkkzSqOu8ffkxMa3Yd9/4fUjKGWv4L7deZaTazqRVx+WXD5f2gm0xCZ
gqbx4Uzbn6DmGUaFcgf2DYnD3BK+I3JCO3mXZjFf1hmYL12L2oOWAu9uouOeTdWiYJFuRI6gTSsh
QG+VGNKnk6PN5MxR46PSLsQ1jSjw322VpJwSj9pKkH6wJobW81BsWVgw+WR6ThmArT4rHd0Pe2ox
6PLKT7BrUv45NP9E7xM8MQzJ4fRdpUIynUhBK0q90tWmYrdHq0VIuitrwX0mwr6PwXFxGi9nZYa/
yRAYpFm5iKdIkDw+rOeYFZnqhckpvc9ZcCoEFUpqozE2G5ytX5qUTW9fHZskaSwN2RAISprIOfaW
Z9NkPKWR7WBoORiL4lg60t7IBOuqbMsZiJ9ITl1KTSQeb0QSchwwzXTwOUqP3enuQrl9gt7mzObM
LXN7ykNQxKq1Cgkg0gcEjYckC69wtIi8KUWRNxf7OLdN77jlhkpNKW91ttVw00SRxgWE580NSV6O
pmYo2MyMmlfELDBqSfEQZzBKH++BSb68J4hABL+eLduBrEFHqd2OzS/+xHCv7Z58yCayBfHaz5Z2
/G/st0RcqkJl0W2bBg3cTPXSn7DTRRvcHf42UvBc5CQY/AbvjwCW8lv2f2E8KrErPDHGYLA2sBSE
nKelwSrstW6qbOkcRXD9aN2CRI3E6mcFNv4Qy6jogZL5LIdkLoCGEKIRustfyHYSBhsaO8+OFRX1
TTgssQHR0NFIngrKq2ttt80x/3yeQY2avbCdUCTjrTvlBXrVYTcCbxM4gYDO+PLFeKTtXun0BHy8
L75G5hpAcBXTQ3HuIL/JfyKrBWxuYX3maE01HxS2j7Ztd08URcsh8obaBXgDv+3/nxHEbkJdkW78
UdQ3cfgNoaASLpZfmXuSzWAshH5Fp8iJZ2+LDQTwXFq6Wab9JA72KKEnG1rMto166n1hXOCEwT1N
vCvERkrjt/RQ1yK3nTAVzbwSfktWAcLriCC5ENpw58y+32DikF7U+BL/8C0YrvpJJTBjAKzxkz/2
AMRrKzs0TQnXFc/sofhbDVj+cN9EueBKiktSBd4F1Uvy2V3F+qvT9YheZqRBwtP70r0yGEh/IQZq
SgvcgW9pCdkdHfp63uASkifhvIcy9CZHkaGYsxrop+DgYwDhwuV1/kKlkRm9OeRVZ060+jDQmBzJ
ilOe6bcWoVo6f4NTmdgl3wxLJnmTQKmNn8nJzLaaRbMtFRyNiT1XQK+OJIsOj9sRvE0byf2bc9rR
DD7Glmo5es9GeEpxS/QbL7qb6n31yZMZCsgzGLQQmz3HyUGs8s4A8IAewXj8r6Xm67SxAVPL5Dfz
yTdQXdnHyNvaEQ3GceiSMo8XNhHbjjom+mny4bDbQK8R1lXvI4xHbdNT5JtdB3V3FH4FvTlPzg1e
APlTqc5nUMuLqLxKqqstWB606hn7UmLf9ph6/BUKHoenwr93GBOWWMx4ihxxi/QUKA7KGuHYelgO
EioCfjRDlNasbkhe1rwtwnvHDwQaQJ9kgvJ6DO0GsgGoR0yHxJfYanuYXEKzUR9QT06qbE1QMnfA
8haI5PAvQnLm3kV90kGueqC5kAPjNhme+BYXmrIZTpB8rcsXZYvhNop17PaBsj2pwSclOkYWPmNP
uRodjzsTHtmKfZIAGpHWI7FtcrYBg0lwg7aKKoCqixFAQO7kKpwtUdBIOCq05Obi6mNLEMwRu5yu
i+bkLyFpnixMC7pM6ZeHmqpOnt61R6GCpwmwZlWoRNASnUvNpKZYMlZYRbGd8EL38JvfHk3xPyOO
IwXeEtiyNKSla0LwujrbMHTwKtxyUYUatvXPnm0qf6ng7qEZ0WXs34fHui+Z3OQpwoo+qUD0V1Al
ecHzu0+0qSsmsnBnERblHiKFw6mO0QCGIglwBw74QrSYi90m5+Kirv8mEzBH+7YQvtnkVzNquk+R
3qvJPi/mEatUxg9Ph/Z3V7NFrzxtgvz99xEgMo+028BcOxPrN+U2DP8zE9UgSGTLUvFkhRyocVJ5
mP98avrgA52F0VYmLK3SNKkrZtrOxkWn4kOgBGFbIKvu6ciYLcBkQ+LF3GC5TSV1scVa70TNvFzX
e+rLNwn5valmB80ayxDtP3MT7xmOZJyF2zit7FzTgQeL4h9jdtSurv/TPrNwu0p/gSjAq7Ywz/0a
gIQA/Q1wRokKJ0BU7MlANuXvtHYgAMBGiWove8cqhrjRcGSfltRuU0cbLs9pmXIjMHjwL366vfP6
ycTBhUfFBvn2wYXcOLWRd7OT/srbj1HdXKRrltbQieBn+RKjkVACzte/5w+y+kJ83TkgFUNNWGsl
h8GjsJVyWaVjYWDWc4nGSwY5BwUaJPSLfGBmMNQ1PVgOVXtFa9zkLBEq4bJY6jIXq1U0/9Sw8Yxt
ReIEMfpM9q/BfexDFSREqtFl0+YprMqHXviTj2X1cei5IrwxxS8cpAoaUPFduCuwvLAFjq2Zi/X+
Ai8hgaFvyv6mgQrVZcFdiYWhZXzMB2nF3HmuPkxax6FCPqCoujPZVhXTqJYfnScft1Qmhcq0NwYJ
sugXA7iO/FPWqlRzWP6wkN8HTtqrN5TETt1LRjIS5ky4uM82E5arPDit2KV6lzIzBRsay2OAmqUC
U74EaC3lkcDNgq49qdK4TvJbnaQ0wVa3pyBI+j38ESM2vXcsvO5nFZ5Viw2cmTUOKvl3qrzo45A3
pOJ5YzF3isU37B+UmS0f507nztPlPFk+/I8NnnHVLt1T4RlhL5rYB/kv+sBpnu1EY7ZEKbYEahgn
O4No8xoUZ/+nnMdZLpO3Pl08OHHc7PVIlYRKK7xbT3/1zTII+9GXTSDwnbSfbcyUGje+l/Fjtb4t
A/CXPbaYFkDPndr+gaI0OmJYy6TUfLVAgrjAy/z8A0RxEkxfYqexJLLMPrv5qVpYeKIThO1EtVzH
X5uXRZBaOCeR4QP8dtV1ikQt2DzCkojJ2/F+NiIS2FBpyjEeq2W/CsiRdQHoJO/meq4zqfP25spl
ZO3qSLq7HTllh96bGs8NyZ3FydKwgzxT5XEMK1EO1P/yUpRLiTeGx/nIeykCyfmpdvLEudmMLu1S
woibiVeuXmJF2OC/Jj+l9lEIETtpKu9U6wbUNKyXGckNRarJDlEFj6U3khVwnQfsneYBWp5IIan7
7eU2OeDmmwIesaPGFsbL8CmHPPyxLcK0itOqLdz1Dlb4xt79QqigxpqSgECg4r8Jn8UKiHdeJYdP
RrIsK95nJ7gahnh+0/8XtWZcYrwL4CwfxbC2N/sfx329keV/t3cIWXODXQEiN8CfaP6yvm3qBREs
ST8NulBHItX+CZ5lCwQPE1hryqvOI1yVS1LSN1go5Xc0phhWXiF9chlf85ywAImAv9Ug/EAbckCL
s8DsseY9APNoOjys5KV1glnUaCBKyvNvbMscOBnAXeQGKAVXNC8eM5rLg/99SK5NOye9XrVGyVRM
NzMQegwdERQoj1FXbz9gUVNoxzXa9WD/5qKMm5myMaMtOAxYUh2FcoWpBeCPbV1vK+jVsARSD7CU
bQTUHd8DlGD6kB6vvMxYKdiWSjcx0TEjEy/H+s0LVJ9lsJwv8pCXGD5XTQD2KBQEsB0vutIAi9mQ
a4HEw9OiVq+0vqwEiBjygIW9aYRZ3AZa7PQ128V68HeqN4l3WsdEMa/hg/LrXLx5d5QUq/1Py4Al
3lBbKa350qvfqUHmuyjedW7Bh0Gp30rsVlX+RsdPCB6E9DjqAry3rToubB9w2jYdccKyU0i++0DT
sgmgwq+AY66FhCpynVtR19K1C3jQY9907r0X5oeu6OhzV0f73zI5joDXECN7tDCOto3G8motBoDq
hvFuxpQcQLDQD+UT9GMwGCjnBnJe07mdQC8YPgyoO2XVBBkSP0wh9a3hH+D2/0w8TfRHcJiwGHgF
ss3lwYRUcMZciu/0zfamDiRwJva0uGKP5TZCwfAqZocxCNszr/P65P6LdFk8+VZoAn9wqVSQabha
FwuXReP+QVui9398DPeE337FP/ST2Zs6D7I+WRyszg+YtWpAlfRRfZJr9Ruq5wi7VijEDbJu0NM8
oxtIDMLZT4PY11FZp+uR/oUvd5vcD6Yu62kC2s8C7a/OPYdO2nbZSJG0QTLZGcv7VulKoLDYFJhv
UaYdcJNd1+nfIM7AdPkFCeBF+6qTNOoXH4oypOlSd5SZPdE+JgvftJBV0uPZGUYd6feny/O1C7KY
Qbqwtm4eirSufzxqul7YQIUDX2m+ISz98hGasilAiqjZGP9eZ/QtURn9t/bDIQUyoG8SEhVuFsUA
rZhZoN29txq7I844IhOV5x9kg7lbht6ESXPM9jsQlXucxykNNJhkPt+y055IaK9O8bUhqBzHtemI
jDhGZhR0jU3nSdEQm4q6bPmbbbI9auXr1tBxXbdjcg1zsgXuygsKPc8GEgwNdjHIWvjrWVbacBob
OOeq7cavmTrNRnFf+ayapatIDrzki0U373NmMbIo6+wQYTUEwavbW8N8KCmpi1uljvPgaDM/7LVq
2faInCfu+22RbqgHF6twDklISRgz3+5z4/HRkkCRNJjMuIHnPIfQICQhlmIIbeXHadyzILwlAuGp
aOt6uGh3A7Rem7NBwRQT7lpYhMeYhDcVGF4X1BJwi8/lItGXhwLhCt0O2cMPTNVfa35CPFnc8TzN
YBsZu1tPpd+YEivVv8jyy7lBtxZwt8abuHjS8sMDv8aW2t//JaMgkP3kOMi2MiSEaAPTvtYFjN2j
wfnLbmZxNvMEpXxHAMFIdaDaZg/fQn5sHS6JbIgP5hqdDbTlebFnaIRlVD20/v9tisoOlfzBzstN
b5ZP6mf8ZD8oUopEJlcqSt+6Z/85D2JP9nag/h3GJcM7mbV2ZxGk1KvfMt6+Yh8m4lK+FimM/aqZ
fzIlRsG740b0APEPIeiE0T4WdzMUJcoiHtqOOMjLnMlM2vOx1t/S7BWh+TJbmHLKE2duJSG/Nif/
GJwuyEOeLrx3TQV0tmnUQ8fEq/wXis56Yk79psHROag8RVqVnQgh8Dxm1qgKdQtDqAlBRioUlTch
ogbCCi9hat0GNAJ/q7QIgRGruJsHQ9LKBltRMgUVD1dfSsFGzyD4G9SEAndXtNxpm1BSMsjA5u2t
zQfvPrmhKtFl5bC3KJa9IBOt+IRXHHe/PFygVy9Oj1MGw69JcEZN8Fc/jOmaImjyPLNmetZAdlgk
VLASegSE4+H6FGKExszaFOa9iu10b5wKvnuNg8j2V1dG6ZFVNXEPM2tzPtGB3J2Lzxy0jYCSIe1W
uz/xkK+8RaL1bahM+kBZKmZ5b9IbMg2liGW6IiRrhMqxb2yHPIqFyKQB7oC7MPyqY2OzIMXM4TpY
vOjG2AujuqO3kMaUvsS5p43GVbobifqFK5DYj54s2MH1qmxalkMIU16Ol52DJVehgt0wyz6UL9hj
TGw9kOLZ+P/0rsAgOsJSeLaQrKoWZuqjsXteO3pDX7GRUPNoYCx04EVImaxNKPMOaPB3jStHHhLO
BcQ5Ptmr31Y0roLkFR3DsKSBvtHbfk8aTRujeoErgrAu1//3pi+su/rbft9xnofeICCup0HIaEdj
1ij+ubba8NN6QFbgiwITFHrjszptF/K7ESNPOSipW7L5eWJT+RLIvtVZ/uxqWwJkysw0RDE0zGNM
OtuCMYRSj9zIlocwJomqiTxbDT7Z0PJP/7d5xa3L8yymw7jpJAqjIWLP4H3hzmVleJA0mtPOnLx2
62XnwNL/2heo46CnVjzqpgIIy7Xf4qUel5OQPICtWN6kgU7Im9VgxsexYXSvlwLrtKRXoNlc3A+5
ZcK4y57SgTmqD7UtXwsE7uU0Q2n58G7F0IbAfM5SMS9rE9A3+6DyfhnHq4Ol8hkG1nsGNXLGgFqc
GEF7QZYNkv42sXKnoqt7SCfb+1fbboLsTPTJzzGU+5dVLlc503AuBwlzEl0ikvVOBGeogXteX9w9
rAHIMVeP/QeXH5cPBGwmCUgcxL3aoLy0V3Rpy5phLGmadFFM3mP2kM/ySSBpgwD8Nu6rEd6jLMpR
FnQybiiYs0iXilRudyGKM6cd+lDPjJ19XQ9Qw0pc9fzB4OKzKZP1Y1meqf6H7umvBryNuQOwE8jG
MmJsA1dfI6aNp+3W1jQ31qkc3RGvdNWN+SiOcAjtPLYSAxdoCEcJkaPEZw726NQR97Zm7p3Fy0ph
J5W+3mrLegNB44DjS70qXaG3T7m/OD+ggdkiQkjuZb1EK6CJzvK0fRO/YAy6w6AMormMb8xPzOwf
cOkAZpUBf0UFsp78u0Jgs9BPMuLVxdf1YmvCXUqsS7csJt+Ob/wHhAjyYD2TY0Rm6IGSGykZuRmP
unilNui96vkjt6pRREYk+5EZfobDYfmphE/muRj71BgKG3047n1mddion0zIQ67Nrt7iz1QwPajW
SYF+Rb8Qj51O+1Niyep3XAknv53kzdp5BudC4re/j7QKKtBcELRpKaO5g3+raNbgGk86SlOKzeJt
Pf5V/QZtjhIk6ZDEZ8qg4+Gp0NZdVHBZcbeTNDDHaBbYp47pVg3mOxB8+vILLojIRosbfKnj4N6H
kjsQBmtqds8sVggtjfdxm8+cLNSaTQz4eF9b+zHEX2g+8O4jnLZkLI9miMsxseMeogap3tLZQTWW
V/yz9iMSuFTC/n6cUNhf2mv0v90Y9uNhiphR/7L3klKCCHVAEScQDb7f3zRNwvwQfGwL/5EbEQ7y
zQr6/K029rzoLxjxGjX3P28hHOcnuS4aDtKkDiieNWQQf6zg/AfucPEeMsMlPLtPw37zp78GWtIB
7RdWv3+FciLRWTxgfZb5wRnCBLmul5bFOoQ5IOdJNXPc7WkuO1dmwYZIwENt4+hGsbu+FW3Ao37B
7c4eIrW/DYW8eMmVB9EO/+l+3BEbTUuU9BopOaEA0FI2qKqEH3ovwPeD9Y1OGdQXcayjY/DEx1IF
JOpdw+LSDdSF7zkR6kdcJEOYMOIcbdEfwReXLLPyu4OzO1ZmRexN+rCR2Z6gnnr8TpiZRyW9Nw/+
Ts0FJeoe0B3dcPh8c+NXn5m/PRxBStO/350cvrSGAow+Lzmowolcs5kDRtfzWw9SPzvNrACI/+tI
vDPgeg0WZTzvzaZWIUXklDdGJoySZ5mJ81nJlnuMH9kuWgtK0yDcKFMuNPcJ+ZuTkAMptXtct5qG
4FlLZ6Q4PuZU90PofhDlKWUtCw1Q+58L0xPWp0xm/meMx6TsfQi3fHNKxO1BvfUNjWB0MGB7Rfol
c6mHbvuYJoUrxTl8MHAen2oqJQ08OcxdmSBDHLaPA/GBFpujvAN6SJw/lnJVvdU6kwqtRcjgEQXB
3kRX9LZM5CYYOl4eyzV9xD+3LwNfp9FvDGUwcPGrXyQsTgTyNHY7uGAeBk3HOdnHwudu6EmWOjt6
WAgXKG4hymnHb/RyawRe2CtrvAVEL4djsXlsSrIvW+uHwIBT8xi85QV2244VpPebqrnKQ42bNksp
0zwpejGtOQhvcHSM7m0YvLgoka0QYRNkUE6X2ZD2zIdyATPLy1sBNwfCZdEROSMnsXXJ5Dw2Ngs/
UQEKPixav+UhjwLen7wk9+uk68vbGI26CNDSaZdZhkJhAEy9o/AmIWgPItAVmBdpgXfmHVmwQ4Ty
dmpPR6/kVWY3Di7jHAcOWmJFENLeLqvsgwbQYVQnv3qOdHpBNnEmetsuvnZYmevHU4a5a2GgnTOa
QasllMMaUfGZzzAH8Wp8k57LVqeq0YS9+9STJWJsZK4ssHmV4kHjOPACp5kdy14pz5SsLNBoMEkA
rFuH8JdcLmE3UeMCbKCC8J2RWbRyAHRqNCFoKwytvI3+uKMBL9UA/n/I5uZzlCqkbPbBdhfMGhzN
9kxqmUKOu/Y2OGx/hYhD7uDwCx8TJLt4no4lR1z6izdjA1YMxQOb1AzKWxQVR++JJGmbMEc+Y0sn
sxXglAv5/QpeHIRaUWfTumjp5HZ5MAfVuV0XY42BbtVfwhXhFihsuF6bq1bqhDY7xRNfSLp4xjVO
nDPHznJt2G9M9AV0sEICXb9/CHmhrhKLh7lHLR07/CeWnJn48wf2N6QNrjaQLJukzbHcb8rmVsn4
IGdLrVaZUj7xY2omwfpRFGAIILHJEgyo5tQ3DDr/pTThvd20qEhllBxylvvbJpfIfXJlxAHUGkmL
IDO3EYkzUO9kn5v313l2Z4Z+UA+RSzfyUhBi29IizNRaR4n0TcW5DZ2KwL3xxfCn/oWlQiRiUDwP
aIg7IosUGMDvwO94eRBSMDpgjNB4rFavjvaWyLJcc1B25tcDtyqNueoqQ+YElY+y9pPnO8jSIFRY
Yk9PkdVcEdh+FG/AGuWQ0xB7i5jPEx3jXrzh26Pp1sewtcrPy02BtAFcCMjoPyqjqS3+Tl+ViNrh
hjJm3gki8bA2JbNrf5GWZmzyPTwQutWxDjIb3if36B2BvLEzmJxjJOVzef09ujTlEvoGYLXba0uJ
0boRZbUT6LHIHpED6onWEDwRdPLexAimfNbqNRaDRpMOCNosp+mhJ/bmrLBf7i0H09GHOP7SFfkn
as3c7GMG4P28f25KhIiGZ6SjGtGwdAaXXaHhSAcvPF4IdpHlRpoVsfq9RLBFiiWkN7wNXk3Re+il
MatI4Eul7GN49liM5gzZ/weC/vVWmtu2Lc8ZI1+wVv5A5/YekAQEGfaYVPo8Fs+pZ+DfJNcIBp+Z
e0FNYsi6xSp7gKUkIREB5H7tuntMHoNsdbYMiOA/YhR0M4W6MwKKh3uReGc6GCo2K5Pe/PLdn3W5
ECTAyeRrSVtOICmfZvCTWDQ9IRz6i94unakQwMQYALhLbzNNyrDLo6XXX7KV8PVpBFM7RiVwtc2l
zQKHOoevoPQB2XLrkReDACf9u8M890VvMfTtvbSudKsbSL2kriKf9MfPakOFuu5GfccZA/T8TtvA
1kJjjVXIy2jW/NsCLc3pwjHnALi3LGTyMa9rlG9T7n1pDL++NBCzDRFnXyvvyFF52pV/gSrFiEC3
Gvl+q7HfBvefjPLd0fYpAGsBML6j9sThlJ5wTfgXkivJC6rvLfTVkuVRCG56KOFjv9Xdaa/Q3MO/
POrLUTxWXuTS+FS52ta3YmUu1TtFuK4tduMriDCcrggJGq2P+yPnwoas+zvOT614IdZ8vxgoZlaJ
kSP0fXUpCFauQf1DSRJfcKk3IdxVcV42bFu22M20ZXuRDAvMq26YAeNsuUc8FPHmFKSGTZ6+PFT8
LPdjo6ebQO8ODA3sVckPmLu2H5g5TgsGtbG81XYdAO9xLsCrgs4nCjeK91fr7/XtaAcquL6TyHSS
U87nVWCxSM+Bi0rCBBVYV95xxoHLMV7atIswaO314kHXEg8dCHyi8q1DN+Sw93YWI+vr9dRradGN
wNcf3Ceis4EYEHiogZewYWmJ0vhP6TbeL6W5POXXoqBMt+nGTUYDIRRgQWRGYDlDvc8IqxpwZ6P8
3tLI6C2I4DmZJJvHIMEstlGYoy8CZZotxF6O1FvcZS9lAWqgGcLFZd5NkDOyHI/WuBJVa6/Hu8RZ
Y6xUeydTfWV8N8S4oSmyikuKIgbUVSHMRtm3KPS12ac5EeFBn5NY454dsIJ/cFaL2eXE2T02JDkr
fxKy/11hRGgKCHTB5aC+LRNqWU2hlKvoAzNSSWNwe7L5WVgzZPGyO9IFhoefjuppGCKnj3cvCpmR
jfW9uJ3i1oasJvuL3m/HAgk1Ujo2cX8bgJ0Bv50lez/DeYlLwfA2XJGJyaXkxvv6mPPqfQ1oYDyE
dLWNx9Luwk3FZs4ro0RbgqZKs86fHNtapCKSs24vpPLZC0xQUdG9hx7ZEDDo3f9X52lGme7hTpmN
eifTfA8BoAk118J831aTDJnDTOTybMGKl4BUqHLvnD6rbVLfNlCYjyOTn26ZjuxtYRC83986ZlpZ
odEYLTM8ZM1YEv/eUHT2RKocILedQdq2S+cGEBzNAr82uwatEMTpzBDMeA/RxVx7ZFe9Ju2IoK32
nqk5eOmdcX/w4jVWDKrRyDbTAgkCLMuEHe0hVqtt2GLiEE1S7NX1gM0ODF4MY7ZoyO4A+MRPuFW+
RYNZukI0KkF/0nSoeIjZYXkh9l3JndfADICIU9+/Zd+mYRIisOTboC8BYW9/zgMI+jpCDJKJQUG/
faajQMuf4Rf5i+8TIRZTRlzcF2YDzlZrgFj3QIW4URvBxTOpzuI42jXfkNj3iMeW8ddIELH4LQgO
vhrLDk7NRHnaXRVnTmIluRMblqUkOpKkPbWsgCmedFCW136o8gKtATVLai4LmoQW79MKRNWmayMy
VdNxCUYAPtc3vwHePiocuAziZWnqB2Gb8cCa50u7C4bAVJvtNlFIEm1Pg02r7/A6ETO3n8f70G5M
EDq/WpoQe3EEnqmYXF2rpCwL+VWx75sUrR0sKXaaBeH85gF5LrbOkbwNujGq6UDL0rzSAuIiBGGB
1tLh7zDbTZWO6noeB5NIdfPOTgqCIJ3Lb0TcG4dpPNYn6kgf5yj7GVVcWmcq05w3W8Lb19lrTOTV
G4WRNvYR46vGCMWZjvX2U4vPrwMUvRQ/9xH1sJnaBx8NPtXHjLoWUx90jfVpnMFZXHijNgPQ6qL/
czdjAqrQG2fwuioeoySWkNfvFOZ1KMulSA+t5MgbV7kk9Z329AYO/Z3v6iBQs6Jo9JWZT3e6oIIt
Ls4RUDmANorn5W/TuxJ6kKVM+EZiDWOK+bu14L0aHkdkW9kVnA8FE2CwkI+DIohkzWPCoTIOhtE9
77lv/70ArdP7gRXrSbNiFgYwMbBqVIu2CUokE5Cbw7NwmlnJvgowN+lKRSNaEcFQdDO7OYeGyU9I
/IgAcfIQivZus72ec5CyUI2GfxU2EDGrkwG2Ypqxefzo1YRkKl7J1BQ6stEJHnCL9pm6KVYVX7p1
vMJHDg9XUqSE/9fPBDXFHUQu2zUqKzFaoOJjjVNp5lNRasjpwDC90NdhvVDaYQ9b2SH6DDqOQ7yM
7Gu7MqOtM/Un43TaUL7wpZRyBcdCeEGWmmq5q//mPd9RwO1R4Ygg3IKI5i7VgdwWqg9a6gnVvpRD
BlsQj504iRWe0lPxbqov2oFbvl1q6zuzETg7NwoJZxLCkj7dceut8G88DIR8z4qAqfEVwfitclBR
lqRtBGcwy6OUokEr2UrFWRl/VezRH+peq0zuDFZlZn0halSzXFRv44KVyf0x68FO3CB5AoYoW40P
Zxg33bkSbfZIwwoDNo1OepWNjsC7aPH2LQHPrqLCM9a5vm2fSXsqpiwzLZAfmIbOyTuORHHkVdEC
4q7GMDOKmwiopS9vMzAI3uJqlqkYspuIrHSHICMzHd61N0zh6ebitXs1i1OdieT4o6LgbPkDU5me
1V3KtgJzuItzLQfbZygwZkPIgMiaZI0BsrCbWa6uzVcvisXNfRNPxWx3yQcz7ue4yk05NDrTyctd
ulIfoiUc3blyaZrL+pnfROF4YrbDVUMVBdk9DxpOV3ySoJzAJr2XFWxE8ijK69z2FXO6PHZOhNKG
C30DeHdUb+vjuMi04P1QnIArmEhCKrQy5D7qadK0KDKeGIzLNslGXaJU3YhLEK/d3I4U//coTol5
b/TcNVzdqbp7R1iDgf2AvG7Ty3Cs3MMBKe5y1ELLDjuAyl4TIYLe8rC0UOkCrChUGMqT7J4wqdxp
JnEacL6YpxESXmQyYmqt76uhVcd6yfHb74HuMv2jqm7yzvDIcup5dgjJyiQB3RP9Au1NSVZDxnlX
81VS7igB71hphC8CRUcDMvwdUgwkeyZt/ljkn52AxRL0hZNOMtmdIt6K7H3yi6LuTjOnm0KzKLTW
SoNjY15H+B7qCLKkn2jFg06GKrbGmQtk4YXJPR+H1HBGF+/ZnMM5ak2uWqfInYO0XCTYq4Tcu8Fu
dZC/U2KjYZ+O9ZEz9ergQD+41KyFehKBCy8rGKOFUJWdFaAM9QORyNAYPu4ZVcFBAHwdIcxUMlAV
B53003FXJ++WnppZbXWudmBPBkrHnZb1Z9okVIJbXEgFxwR2VCtiX9cin8S/Vyj9INMnfyyvwmZr
JMDGi3ls8ImuX50oyBZlMENC25/YM3RUl0Z2thJfvxH9Px55AD6a0XvbG8d9lhCsSusPQOtFroE0
0NwC1d690rVJMhQvXeGJRUmZihGPL/Tn395Ek+0HaPfsGK8qj9d1LEFCqSDwF6uDY1PlwJpVc3Ui
QWuK4TUBJCDF8Rj24gQaGrs5AG198OA56aybzKcX6/48dPrZMYr/YDq7FEoxV0XlM2j4G5z77y6a
1dQjWEqTbIJAIOinQM8C0I3CbRENhq4JPTWZGLvQHVXXZyG5VE4GygjSQZqY0sDdl8JKIpH6lRGa
a/fdBlNadkNfnK3EJsQTumEoH6NEKIOlpAEb0EKqCPGapaPAlOK+9YWRDKHOyqWQIN0vH1YJMHUc
ukp1ugF50dNs3Dmnc2sh48MLrjjwWsoFDS++RulXlc1uwM+ffXcy6i8PxmIROY0bNMraMEuBOEyq
/KJf4uzMwUE5l9fmJJvQMVLJnbB17HcJ5jDxmi85026n9TxEgELiLJqJ7xVRwj31hURSTtW/7Gy5
WWfzf3skpjn7QmOmAHRaugAE+8FN//F7rbjeGyPmrMnrS/yf1c5Mjt3Et+ejEdB7WXYdtvbP1Vty
K20IFvXB+XyqYL1TcBgZn51FM1pwfsK/9VZ387oeRs5/zVAmAi++Hk6eBeEUe+FOKw9qyULpwld/
eNO771Hgt/4hjL/ryzxfujZieQCMEm/8ouwCw/gvN1V3BPWrWmBN2Rv7illZanPBvxmJXZxOJbbd
x52LJ458YzgKgI6CU4o1mm9AOM0pMHl8v0GP8d5cImK4w1QUWwGHSNyOjfC8oLkDD0T8KF7dX5G6
Qg0ymiF2pjtN3GQKT4aPNVFHApH5ox1AdOwDh2F5z6ZV7Gj2xvePGS9Y+Ro1b2jljoLCSLWZDSTh
ihN8CbEfwGM5V+LKwpE/G/0aafRvFjRrfQZPFyvB8G/mY5o743i4uznGFlYDSdlg07dGzd4mTLrq
m1+D8LiYuCIXYDUsvIcxTQ5OOE7lHOWqA2J0e2meuKfx1NdvegMbyNUYQETbRHR5DKKhHWDqEsV1
TFsj9IW2ddGDvkggLIXuew82+KH6o0JkHH3SjQ9mnEjkvYCE7wqBj5iFs47PC1GGRLtsQ+eMFZEu
SWKg3cLkCbGWs4UNqsDoBnHZnFWKQLuN3QD+mDJuJtR525tI/JiGcgCHRHg9Ubz9v/2C8SayBSOr
f1z6myZk4ZY025/dXkSHnco7orknKwLK4ipFfqzizYxAL94aoXzPz6Zwruf1QpeBe4fAGvekwERp
g2A1dOKlWTsaF83t594FO1JRSvcQc6Uw8n2SfocrFDoEDqqYxcbgekjmTZVDwlu1OBTYOMQpdYXz
MxyZhW15eH7Zwhn5SyEv4kCPbxcMS9Ykc0+WE9bGp4vpHeZisJkbQoobCe0DUeHkdOvRyKJgpzxy
gxkxa6rWpoyx0qOO/FBfq3guMe0hp2kI6wX9P5YTsLYB9lEBz8n2AbYT76Uhoek6+0chdZUvrdAz
BiciBs4mjHPJwlUAKvjvUk/sUi1npr653qPBzIKilop3DOq5/NvkS72IRHBqHhrbBXweBtcLLEgY
m81/h3BF4Ke6zXOoUkv0FO9dmb2KVe5s1ohFU+h4S0bxqgw9I4D0DgVppzzqSCfYjPxUgImHbFfI
0Oteuu6cmewKCtL9mXXXG4rBAPdS3Po89unOI5MM2JwSH/VeUD9S4fF/sBOxKqBzdDkJeGH7WTpN
phTJ38p9KX5Di1URRgp4haonE9NnADrqdeAuZVM6rElmgrYSSl3VTKXSWgW+mqBKyb76J/TiMc5m
MQddF992W15ANHZfKKKJDqa7WCz//uKydtYVErwY23kga5uqS3kGMugKDqupfVGMctIP8L6gdJye
jvoCSgoCx8vlRrDkL8l26MXfG3Gf4AqpUg8BVV2bwtskOw6ekbDcAbe+kFGWcql+wJpC1Yv8YVMd
n+pb60cXUHlPAzH4ihXOpCfH9LSYQo3tNdmpAalNOX9lqlNILmgj+CFpT63Lu19QQas2LtIKRX2O
VVip0VkaALc6ZLHn16ezuKfg+Bf+HA2XTqXjlata7kX+aqM3Hy2WI9jXVBXdk4EUjdfAFEqVW33D
bCIXTUn4gF4RMuYe1AOH2fljqPYuQduDFv8VqgRNMd2Y5yd3I8De24zKQ61oc8JZ0UEUHpoAjU3T
5opt/pzaSAlrLq+1VwetdMbDGnDOlJZJ8UM9hl/tVGPO/9chhZttYdKWUmncCpBu4GvxH3vpud+w
3KpGBE5Og/pdYEgVNJIs3vo6qDVNMNNcep+wunKRFB7dLrZPaQOvr6SlD0qL1TGjt0m9Nn+Y0Ivb
xWloyO17MQU38ZJgJLk89pJOOQmuodQFxlRs7Y+GXZsXiSER5XNOUm2LVj580AJgJ9XxpnWKQmcb
V1O+xhA9S1Z40mSNYniEW1DsOlsbwQdl+pli7G8oq0/KqJaRso8drF9uJkxDl0tVMsHt1SEW79iv
7iimfMBW7ChwMSsgKaiF+XADCmZvBrfgPNGyjxn4r56Rzt+q8cA1TFbBHa/U5pW3GR9R2emIvi4b
8S011/fPdI90OyQm+IgKF/RyOUpIAgpmMQOcLTWKnwUL9hfjlW5PKkqh7ai26XoYDw1CwRwBISdS
Rs5yatPU0zKQVA3crKLnPmN10qOqUdg9LkGmWS0/WEdd2VeoK7E+DPrP73K5W+Iy2qKqOpKMrhzQ
/Pc+o1+OkBYkwDHoCZq6hVLgdqwcMF+LZbOq7vnG6JgD1K8atv8UoU9OqopiVkCqMF19CDnykWty
GsoePjEmx5Feu0/o8gpJRLbdDZsGGQfAvso4vVZ5XcXBmorSRDZ7QWjlslcBomTWMCDOCd/hiQ7U
2+HlEXfexKlyngbxps326IrYOA92t2jYgHpIr4FdN7anQ0WWkL3TocKZb4dnkIscdpT71EAGNHf2
KauL+v/PwSMDBjflYTiaw1Yd0h19i3QqLXosFX9+cQvWG5mGfx4I933CyUSak3UvECDDQ5Ln1eSI
BQDXHz9e9c5L0xgMJNMheZpElqfQUze0nQpE/ZPiI7f6PkecT4yGHIuUTGARCDRK0PoeBWlBK20v
35YRHffcLq1Cp4lQV1KrV5iHJjPv/m0dZnnWpMA3mC9uRgwrN4r7xTNdUSnkvH/HpV63DIPJ7Ho0
MIhlX8ksF8d3GCGMN3BnLNDYb6Vka3Tl+qkHVKOQs79/ttarRYdEAiep/eNSp/RtIFR3ZKz+2bsQ
2FxRIuw/6Y3clEB8mxqzdCciycffOMouQUJdzA8FVk8fKZwzLstQU+HBayY6j3en+8iFCuhhJY8D
nzAmfypE5+6m46JAm4Q5ByH/DqpzisOoa0xhK6wDDTqlmQtJGGGEzUOHbPWB2+9+xmVyTXAf+5FV
RfsqTpbfY5yB6a1VKAlAe07YJFYHGZ8MpXRyB7vt8VJioYg8qkNhCK5GyWMexlfgbDmoEM9xMQ4Y
6GPkA4Z9Y8LAdHt7/NH/nSkYViz2GUzKuGWV5yYHaiLWDf7Ufj0mTe97/5ARWUp6EoD/aOvx00Dz
W5FgBi5dkIPfVjtrCm+AYJeojDxUDV32p9429sCUEvtxqfYvXWElaADAYSP5vK0alxVRn230LAIT
vDCThow3/FjjshBpNsGgnpDUMbFcdns67r9pG4mOQmkx2nW+xaorXD13PH3mtxXB6HPy+pJHD8sj
0lKS6KV6rO3D3Ie0vGFmS3WQNLae3hRE2SlvbC0ocvO67DSdLNozzwaMzospBggpxZ/2VInq5Y1C
qRYwasGnZn6/sz95b890s2skfcwx93jSQEjDG6TSsTl8DAA/Xxk0YGeTHV6ZKf63kCTVSBbEx0gs
lJsL6QFBVWb3WJM99BUC5J8CLjKcXbtRt9GXPRTJtvlsmbenBFKduWhI1x+uRijgXzWl8R1CUvXF
nOmHY+VZJVSueZCZ0f7hdkazqJmwPAYeq6Ndk0grq7NU+NCmxHB8enTMM7I2Ugq8kOt3Ff+qZTzy
jY7GqtxbR5orrGB5fan06ldHXWTdBoQH7LbTPC/0exlGNIk2p8ciYGlzSGdvgwOfjVn+lFmt5JA4
xcfgWjQYfENaUw3w/IVcUTwTCuli3Kz2kSZAiXJ46zMY5n6r0G2ISrmAXwdmvNoac/W2ba9LAVPh
cTI9W8E0sBjgY2HoLPUb+Pv4TjVHXyIXv9wclaoppeyD7XxhjAhvZDsCSBILNzAh4SPcgXj8ioVA
jvJM1dzG8LEjMJksViTgraykzrfrG35kcJ8Oul4vu89NKuGmo2i4NEt7DJCzl9TsGq6g8Bh7gvFs
e/vlWBwxwm0G0HuW59UWhH/j7yquljS3/KzcX63FyfYK+oYVhXw0JQ1utCoBetkgT+Kdx+UeuVSC
BKhfl6PTXLZpybjKywYQCDM+vic3RIcVzgklPhKXWO715PlB2xP8bbhY3FbytDO8QIMp+FNGE8GV
6c7T1wwNkkTYmpsS+ORRh1W8wgH625sOh4IVma40JtKU9cXmg4xsL7a4R1tOS4YazSAS98YdVahM
ZBI24iWxqyXPzZss+EOXmEqCBwYaif46HxgTrDL3Oa7/8kxcnEOH+luIaUCMsrsIhWJul7g5sGF4
Fg2s+B17fMDHgzzX4aj/r8h5a++HoRUa5+vVudQVnNb+OAc+qKxr4O1DaKt5NkENJ3wOSWnGosSL
qTXfhsefzX5xAh2ZFgha1rS4qS50pZPB16W3dl3hbnCrH4v4i3ZM0Slc54j5A/nca1OaPigV9vZy
2edL/S7XiD4CP7+3OBwWXOrDec3pguUaboEeJbspmkPdQxqzrYDulgjRyfn2GFQ8XcH0b9kFFwN7
Rdvvw2YVSsytLCmyauUa4pAXiAuoWBDijiD1qAi/WtDEQVbZBKvFKMjoFHqHffmygFKdoSzBY6L9
1Sk17TC/Ke35JIJR8HHc3A8OyLNycDkvl+coQouZzY9HQCAiQs3rxljSZ8qTlErE6wGScXwXpBkZ
8B22uqy1nuBx37BgCEzFZg98jn0TFdC7391RQpuwwUmi1HgM+nNyiE5iYsg4j68vsFronV6NTPys
NtWV1umB1F0ott1jcETjfbeWB+hL42V8E8fTgPUvVju6dlDBwY2atkmYprjPfXH7lCORA6txX7uP
HDmIej8sAzS3Q/5Q+JmSGQbvnGyCO+c4ltTjwQAvjlPXQUrCya1QVsxRdMcRQqg6MmADq+2TThgp
LukDPXfgNVNxgm574pBNGvph+LClMO7glz1OSkGbUnESIqxdVwU/e3BE7Ppm626zBc2Ry5V7EHhN
Jk2InN6dR2SYsoUhBmHKVfanZmx8tt8FeTRibetN57JsGUbxRncIpH3Fq8E/xCi8q/hkVXB5WG/X
6LDnHMGEYnv+dhXlmXr/qo8+CT7qhLp4So1mBBlM7d8psfBIh7v9uo/6W1MpfG2QHEhjXoGLVBr2
XFjj4W0rMeRlKp6J2HFt1J5vwn/iUHo/yOZfffRv2pXCTrwumSOpgPKnjh1jSJM65lCiFrKIOtrl
wxl9h6yUWPfeiMAgcWS+5udmcxqtTsXosvIxBnZxCkGajNCt03Gx2AbThYGLVWXwMIob4YhZ7wV3
HVVVesDBeWjGeBrrJrfXzGJFAmffAMXcnm1raoaC+y0YZYUCXc1xlGkULetpCZPqd4xTtT6YySYa
1q+XatPBQcWW4yn6SGrsIyhbQ68jE2j2LSQO7sHEQBjfy6YRYc+uwaEfW73n1vbd2nSLc4Hqqm1z
1PciQI/4FbN/ueNZ3zB0sYqVkArYKARMBt8verwBuGmoiYkbqjbMIlnYFD0k0dH8TJ45Soc/hmKl
pMoo4R2QkxDkU0x95tAmBamrgq2R+zHS0U5WHggmJL8hzj6syZslb7/GkU1ApLAKRxwnHoEFP1NF
DMCrQ5fjEPa3+gG17eeriPbInnAtXx/+mNpYqF5vkAI2MpPGl/QrNkdZggs20yScwIZf4pDcz8gh
sBtjyJe8ml3odgJK+7HuA/lhmofxHe7ElybgCHOUrTP7oj42cXBg10xIS9XL8mRL/+Z6Cy06UtlB
yvKDkAZPudio4yvJz6BEfkmKk1mtK8BfiUOTF+Iwp7YEW3SqgBEYkYv1nzYrc7TV4GyWejGkrY5r
0UgBaCzCjz7aJCKxIooVr3Af3VlGmMVsE4JvrejTf93cx+taLieESv2+Rs0+PZpTVrD8Jcy5zmCz
kL/CkAH+ZMIqL4CNpzMpz0THGX028oyHn7A+d7aeTYtEjGgVIkRcpBJW9VVrsn4y1CecygyaAXST
LHs+HpzjNU6ZWaNw5SwUbGZw608eGUb4SW75fWULqj1QR4GyeUvAg3m0roi/jvhzumg413eNV1B1
R4MTo5HAwRhyhlqINtBuXdGJEpy3HmqM15HzCaneWKclr3fKCeMygRXqW4v6OnoHwBeZgMJSkCJy
OasWu6qCq2pRiNcESCwTTz7ch8SPsGrMaEtDokM86AGCLP1++nivD3j0yCRYvkzOz+isUWt2A64E
OGtiTOFS5nrrHgVj/cnN8p1Qfvi6Z+fPRi7LI2cU6+V1Mifkbs6i83r2TbA+jrQ85xQCC2O1xoBP
q1y6C5Sm/E1hVbhaAtyDhoPsNrN46GnethchI+WRle3+nM/rbiUpDQXrrNGKlFLfpqPubLNBFDTq
XMVvX+Pu0WjPz0BkjsK0yfYZo+Vv6LpNKT8bmBL0aznusOlDoLJA4GmhWyivSlL0Ij3A7Qvy6xTF
0L4tzQ+qxocvraEtDg5upv/BuoWvS7HEylBLIpu9KQLjdSMFVvKEjlZ6f2Ln0EAvEVbZgNtZ3Glb
u02GKoAkMOhWnlsD9+mFTsml20M/rLGi1LocG5NCVTwt9OvjWqksSHx3sMe1Gli5mZENv4KfjAIW
Xt3QmoowPyrzGwcG99L+m8bNOtwsJ0j0Q1Hu1Fi+lTk3xgXpuokbJdDvyN0SqItkh6UK9wV7twlv
Df1iFJb7yk7/wLCFUIdL19NObTNL0vNEnsnFQoJ4FhWpSnaseR/s9wOmyMj/NPuPltldnqtsULNA
kPHrvAH1JtDa9yTEzqWgW47ra6LzwrD/z2bdrsjr++DlperVAojA+uCAsoxIZuiuUCLs78bnht7B
RWmMMyifRgCqTwkodC23w+6RNRtkXZgltt53vf576KXRre5tdyXRfqUKs7aDk4nahZpQxK9ytVdJ
vSCJlpLsOMCYK47kQEyo/a3xR9EE2imQL3uPKXTU+OQ6CUB9PlZd3CIvBzST9pul4czEqPSwWL95
bumcHwU1/kXC/Hz2BGbMKxlFPWlL39XHAajGcLvnbTX5FYG6pOOk15hHv+uo1gPVSMegxFmpavWE
nxS0dXfZ3/jyf3MBD+uMrkZ0I9vLviXNyrDADVSzoc89BVQRK8FUncDyG5BKXGX1KTsrDr48Oh+p
TUGyXKKIVEiYIFOsToTRFv8o1Pco9J0/PKkcMmj71MQ3e0MTdqzClJ3AFnpyp3dtyX7tnbYYxao0
It+1jzWB/uNUNSJ/NtPdqyes2rgYQheVfXvUaQUpiXCjm+oM32bMkIphYiWaAcglf9UoZePsJlrg
WbneLzXu8PJ1IEff0U7h4HnHWK/JeR4FGyWhz5WbPOTyNPcIEht6pAilL6+uOHqhYBbzY+8LAmAP
Ey3vuBYTuDiOpR0Rrm81XtDIFD781ASxJpPaUPDdTpDVG3XzS1AK/rTkCBCj9KGgp6yIG4rszsR7
TOvyxcR27qgo34qtIeT7BQRQ2qdVg0t7UtxagIykoorQUkGgMwI6HAWX1DuHMm77kniSTzo7HPTT
BCKZHZOlWE+/o6TsRvNye+TsLiBsUDnMKSFo2A9mbtdMH8wwS0rm5uInMgpPUlvfHlbV5txVaEva
EtCqxCErtwCgXvgy+GsKj215QaVzViRB/ivlMxauSMdaK7KwlxuzTSWbx73h1UZl4xECjnHI+66N
hdgllkhlVaVvOFQCrCA1C7+m7kj2NqOsME1o30uKRHSZ7CQcZHAlKNQGWOERLIJNmFkCcahqVd0Y
jskb94s0JaJNzBKxg1Hgdd/QBuEn3ZpfFZoXsabA5MNdEPLe1jLE51vEU8Juj4cfnxg0ytL5aVsl
WddsG220iNMnCJNvtSPy+yYglTYsc5+u29/3Hxvxja7EoV95GkkAtOHOW9f6OqTOfVZU2eCP7/c3
pqOi88ig80AMECndB4esJwCAJdYpRFBVNMqAVQqzaiNZsSXz+FqUQ5qakkv5z8OcIKhpNDh25XCp
oFiWnD4FaDPZTGNOp/lbnIzFiC2wFXwnvTmIPkL8gG9KETOgTrXK7AG4IvlvxTT6BvN6b8kTrUJN
pE7kTqm1OsBmsaAxS8rO1hwprEP/vSR4wCCAN9FHl3p9rM3SwbaboDhyVdtb8yQo+JK5spLtrS0Y
QdPP3gVZTAJN7WRJuo4N91/WpYWcBeei304vq8qew8tADq+2XPmwhKogDJa1pzDvI6Jvswz7sQDV
isf3Vi4dq4Frb1A22dtxzeJlytRBW0hW+dDMa6h38UuBWoYahyZ/tH1Y1jy3UNRzq/nvU1CnrQto
D2s4f7wfGvk85IMSgvthfmZOJugEaPNFSvr5lVyfjCfOlY8o7m3yay5Q9bC38tePZq0MEtZMY0Uk
lArHoZ84YcrDfj1HX4ls0ApAtR3M9Vc24lfw4yGQ3twlXiB+x1dRDGUElaovzjzVg5r5g/ZbAMgk
RchvZbE7VWn/5yTIFWLCUS6A4CPBfhC9PD0oZvr9e//4jf9B5T720MH+fpm/MOSMkXOBULcyClw7
s/UZdxVe7wifB6d5empdmVXy48G88kkq2o/XbVa8RibJAE32UHHB3F/xFE1c+jnWbrODMVyLgr+G
HAPW79WWBDy4eNqxvGtPXRUiGrG/9PTrAhs7AYx9toZFicyxfubxT7YyVXFx7Ry1fTx6whKwf/jg
GdiOkDkh5EfNvHPKTOqHWiWnIfqzDfa9L4n6mf/95x6hzfGu0m9MIkbgsajOd3Wpgh5FN5akJ7LT
3n/KO3LDAsvNVqznm8AzzmqeMTlVaJziumnRCxlpfc1H4oRtKJSjsFV8PAkd0XLiawuKDQZYm24e
99fdUv3yWPkLMmc9Em/uXgotqgsEPq6HQHpeQOwzPZNIswSrwwE2llqsS1JGdNPQSxFG33TJ9bXz
U9M/2hnAstglfYwdd+HaZC+Y7k1jtpvO/MWQJ9h0pbB/D1EWNGsutf3pgQ850PC1UdipXUAmQxfW
xqQ/ZtCFNbd/q50cn1eqF7JfY84X3y3u3KSXjT8t3EbK3VbvhbbhoI6R73dSg+xjT9ltmdDgmI2I
MjXYSjLWR055G4b1/6FBx5lA6UOaj+hXeqJZwuTAOmBOi2QiTTE5AKJ9J4qKZ3rDxh7C99zCdQ6U
IyVQH8ZR95AwGAPLFm9cepCSgtXyIVvg5rbF9Qofj+pVwgiEtXUL/p6LPci8JByFDcXZnzLh0Nxa
YHhVf1dJzFZNzvQ7P9MTUh8jucibwoR1VCb3MkfQYSe64MttTlJpITjk8Gz2lglVOBPn9hZ2h2Ts
DrjFnl7RzY0wQxJpq0OzcYv57OHHhCb3jEm8H287JK1AOsOC+oY/x6sD5vIK1IIwJgId578hXP0g
HqgeXvnBH6v+AIb243Qg12PK9TZOLlQzMrsVienti39+HY0p3MarglK5xYo3XJtbgdmCquewO+c/
WWno3Gmmhl9urbUKCWU0+DkXN58fWAQMrayp4HyjApWn09KmaUfmscjpt64NzG2r534CzNxUkJ/f
D7AdPngvNOlFxPmdihn2IC8P0mTsn9V0Enl3dA4mOSmwe0kpGI8NBHJ1LIs9putNwownC24qLB/V
pXAt2SwrIhE4pXFgpAV3MnOIeWf9h7flmqb1F0johVfS87x+h4hedUXh41ZyTXs/pPNQ56ECpEIo
waPaP0lPthANHDWfxawiBax/4XhRerfZND5gc5gZiDkZ6LuV+96FR4qv1DtnN51U5HLPC3il6+u/
GYP9oDCQe/kvbeSe6Cd4gBvhZCAek/rx6nNhcX0BjdrNdhdVz2hEkLGY596sB7F/HADt1b09vQgv
+blCffGtnnGJ4TK+KPxk58eDY5tZiAva5jsj3P9HARbtYjLj57JFYitDcOTeHnCc3+3jdFP+LQCd
mREBAG/jWb+l7G0GfmOXCGZigtPyes88cVm/mBbXVNlYesTXJ0Nbdo4BcUZ1A2JR0Opq/Bl6E5C1
SHcr6zua7j7+MgWKo5k8gGud6nrKq6hYpXKMzKagNYrllRYKbyv0QmG2Ky7IjsKWeMFjL1tp2yi6
EZY19dFzhsf21HmSAxW+KJOpq/MlNUEt8Zl2BChjGiapO1pfMNjMLilh6v9npfN5T5P4+arHGs7k
KPEEFvbgk82VY5bhGEl2DJzht/LyLkewWPKzJYDwrpJpj8PwkgGxTXA49EK12gW5KTF1HfmqjNVY
BfbeD4MDe9xucbhY2+BpMqX+ybB08W2ScSpS6J7nQqJo1c6VapQMEsYwadZS/sZHlc5DZiYP+YkE
zfEID7eR3ukCeuX+lgYrjbhgifLKBtJbc8C7hADlphZz+45tc+bIypTiGkbFo6R0e1+0+C0YE2/m
7mx/lqb8fP/VMLqmmctlHx+LwM+CT/AnTSBePC178SND4Q7ZNZKv5RuaLG3uN0HxV7jiX6hUtAAi
A5VtbuXP0SHA4i8nkYd4kKggn1ni7mlPOJAV1YfTX6fiAvf6YIqT2zhTPc4QMug374tUjEE2fuv3
XesijrPR2eqgTI01noH3xQ5NMdN/n0h4imkFbpfZxNyEVDWPC7+DZJ/8IOZYtkWkilCjTuTJrUMJ
tk4Bz9cxquGOC0S/Fszg1OOaQ8or8Tu8TctpC77uEozQJX878E9Hj6iImfpTrXbYUYlz4chTpism
ERFAtZHPoHWEbOXbBCgScEZH72+rGSUFlJe3k+KfCsiy6wMaN4HiRvCqBfACJKtb5iq8a2sddzp/
6XNR7ySmXiACdZ2I3grkQA9/Qx/7FEFDKUIkJfIuS2zE+yV/XJnF2C8EDyYIflFF9LUd39ZiGdck
T4F3loVDA9cS9LtVOsYej9IjhOBCOTg4OLDvOzkWkKZc2EHf5humDKzGmYTxkQJHZMZJszMMzHcx
e8gxtR0G/+ICK1+SY45HaPZ0N4q9H9omKTNoPjJPyr3pKN8Di57fiXAkmVklj5LyY7SgFlLVdfsF
NgKFyCvKsvHN+IBX5+51ozqj13qwDp+yksV3IxHTBUl0/8KFSSK9orizPDKBh0MZftbQMUPdGxeL
LMaaSt8QZ9yYsAaniQh0JyJ4ZES2JmGLbxX2HCgzK7wXWuUwb7Zl6jUh9beHwUtEod/dsK55WSpd
ZUGkxkRuzPtq5J7H7A5hUzsDYNEGOAA+JxmcSUrchpOtJxWY3wR2xywpHLbv5p3Thsb0VG7g0AkS
DyjoFNDFCGcLVETvBjGgAoeO3aTOh3NqzleCDC4IgyYiXE7bUgt5KqDkJiUZyONQbAGbK4g8M+go
tUrcLIPFVszErcboogJLoZCv1RusEj2ZFw3/S1m9+vM0hHtwZNQmcQ6wACCqe5Jz2TUw7fJV/usn
q4V5g6BeqDf5Dfok4ObXA4OAURDokePu3bG1RlJjW5G6CidxAI2BVuKImc018Oxl8DSzWuftolfQ
vnm1Z6+r56A3A9EH99dAcJIu7Ujui26xxBwojbyOBhb6+Q+PjlwInv9m9F71zShS4uj6dsJjpEjx
5Jjerh8b/RV1SKEvkMmLonuNNuwZBYN5o2FsDr0BJnKlZk0DFXlaBy2Rm6MrO5aUMrzLCsofBkSp
Cp5ha9OwQm0wCdZO2ks410nwHlDqakhMkba+xnRuJfoPIffHw9coVUztqJhK5TievbnlQ/2kxiG4
uKGcWuVXhW9d5ohApa+WSz0ntU3e/q6dN42iCNK3rCwp9xiDcqMivg4NSlBjoJAsnHAaNLYvk6ML
nzypA8m/tCL5DJQ7Jb/EiQfDNrMP4ayu1LmBKFkkKcb6+eQZ2gHQFXAQkXcJv5HQiCbrpqGpmtBP
79U3yiUL8qZrPBf05+vVWfFlNhamUtg9Wc4mL1Si9ZUNKEL7ielyQh3cf7joTzZNHKeupNvlJNG2
MF/BELhFBJm4kJMq6c1lUO7huDnFtTbKftJEEa4XaQWNjmHnc4JMr+8VguxlCSX+1Nyhogp3yHXx
TWV8ibhHu2mi7Kv/qPbWErqT6e1kqfFmuNQnWvXxHolNFlgQWR/PTb06SwtkaIhBTcyB0oQFyQJo
xXOEEShEZkoAaqL6n4n7FLpIDxjYCgQT0ZIOzxSi1kDmix4EgEN1+cfKqK2EEmR4c+O2TbfYB/7n
tgW2b3OO7lw5+BZlL2lucEauj4LgdH66rvuIkVD5vqjBDqd6pxR0BR5GQ9xbRf+2Ed+PtSAk4XXf
rgV317zI+3WeodLLttXh7ND+2wyEbpF5C7As4mipfqY2oukB3awIf34AjtUdDHxMKozyUSVlq2Yj
zw4GmYztkYZRZgflw+NPOYOTjjLYpHD38ehtTs25kprHwcSvlGJMnA2K41Miuj/tVZ7NtlGyUjRj
FiRQq3/M6iwNTHab3KD1vMt0l2SQPz7vvhaWohVO/QEd77aUMSPkenOZIWJGmqhzhT9MPInSTcPq
RIvMhOGOvvaAoyNlDyLubeu/vRYP9mDa9yEzComWul/1zzg8Wjv6e4PpOB7rNFeMbjmu/yIHJJ/V
SEaHQ0+zbDlQxny809MPkjJva8ZR7284irmRnWPyd5QOopb1X/WwhBL0daM99rN6DVjh3DWrdFtI
/ZxBd0ru4wIB4pPkfHp4VW98ByOnxFY8h/iMWGe8n9FtXxlC3IGvF3qLi/bq0NxBPdKUCrJtdP6z
2rtvr4L9dQw1c1x1dki5gi/kJMDB49Z8ZCyx4OCM1XiRP/LfUkdCyWnwZyLspCrUU9gM3jP4x3lv
GOoQ8szw93txuUC9xgXfhStWE03dFUkbBqQB9R2/4FdwxCVsNZahb8IIFKHMB8UdxP8Vcwp0JvB0
Rc3ksVsMofYacEIy6/367Pvgy7id1ToDYZnnJM9gcPTwcOcC6HlQ7MWJliJp1LAeUv9wGSRSCLZF
u3POILpe3fE8n29KdszzMDP1tLHHG7kMoC4xNGUaR2SSzjqoS/slV4iLetd9zsfkdFKfuaTvatl5
DqV5h9KDMSVEO/0xvQhTvmKFCCxkJEDz6LR+NkRp2ubyLm/6GB6gm1iuPwLUXljYPmfrNrHKi5Ui
xh3YjqxcUXd1cGS/3GHrfNjr3A1q+mikd4+vTulAZC4g1QdbnHNdckco9TfPocnfbA2ofoUAm/yz
5WfNjrB9ZvQuH33sSkOZdj+NC+/eFh/5LGxXhek4W6lPWkQQgxCucCBurGpYmnU+Le3sm71p0cqQ
PP4hUDLOnB/4jTYEEam97h9gC/v7lLRKhJ1GZYK/ksfKNhkGtlF0Zj5yeyf5eRu8WIQqPwKQyG/0
yVYFZyf0XEeFhx5IqN4MyXwqRBDTinfEE/NTMfmLs5sUgoRhnSsyRjQJM1wNnyB4zrxLtEbGl/64
x3s0XFABLnt6+qqEmXgxyV8uiLpMOA9W+sHK+WIFdYiZP7vMWzevA0AECk+pwHBz69RAPNRGbHpi
IFBgWzxv2RtLc/7YQHOTVd9vXRhVOH7Nh1zZ1tltJx8wHIC9Quyak0nX+S30nbFuMBbxwE/oY+59
ICggpD268f4c/ehVfQwlOqUwmD98pORy0mvF5SHsh/bRbi0G9zFEGEZdc8lrt3QAXmRCUXfBHfpO
8uv2L1ZM0T0Uk61fTag2ZFkabsUlNImqIF2tI+PkCbw7kP9gzFgtyTLQVjB2xnaovMqDcthmJbH1
2xNNk1/lU5SlV7mAI4qU63QGtVamkMfJB9NtguDB32sWsiO5fbAhTDkTiLKCPno6Y01+4NE3HZIf
2g1nnOq7Eefoq1oEe0lyhHxbbvmoX4afGEWfmfMBTQyUw6iLc9EBHUZN9o3OOIT9ADLhEEFu2XYm
tnzekVGc/RdUWv2S5gLeaIq4ituxBdNAr/zitIHKuvn3LEEkV32yPGtSwqLq0RYPFngsc616U0na
cqTnQcf0xFmBiI5RfcxyOdsczdHmjFC/6YRF+7z0IhXNm3WMRsyQlKpaATY652O+QDs6Wpc0CoG9
izZ5c7TEhBU55mwXh1qkKDaE5gijPJpilNfnC17KnJOYP1lE2i/maAfXEqsxRsqLLMAvXsGj/Xb3
Nw4oz/DttNi2ay7H2OZKfAvIMTVV3NmdwLyNsyRoBksBOTyikAHeC0JWpy+oka+17L5Dfqxeb5em
GP65WO5xQCy1zq2frcxk8IY8E9Va/1FvGEN6rXDRwraK+JhHmgREQIr5skXfq0PWTLCq9SXiQIQB
wJTMxo5yqJMciU7S2Lu9lCHfU+VhulMlRfO6Hr9Uy5z+EUTiMKjwGfymKz60XSd3yT4K7LBqF8S6
S5MwkwTIh9+mACOa1+7GnORjsXlqcfYVdfp0aJOkAKVFx2zN4OPj6CFeHx5I1z7GoSANVQGNnnHq
nzmws4CM/MftRBi0iVQoGlTbBUU0wwGZvNqJBGsXOMK+rcvRaT6XG4FzvR5rwP7HjrvywF0ZUCf4
cH/swG8F5q68wy5UrI2USAjSSC9MlQWQ5vrIqm2FZTZMTRL1paRRyWdR8gdlO3za+gwU8SGSlhxE
dlkkyw50OoR8RUDf5OJlNfu6SloERgJEx5+1fUlfX2L7QLqvrL6f6kPwZ9rsP59z85Fb1JwOGyGb
WYMT5P6LU51ic5ASedEQDkj3s4U6R/doJLQJGzBDzwh2580kc1UGULlAo1bqz96/oEAJQq58u6dm
ea5goKBvJBXAxkft10eT9EYnNZ+mAtSQQwpBGux1Gwgwodmi0RzujgXvCLDEntMN2DjK/3ICEC7E
5q+Zu49ofLBxQaChi4WHFgopjSmwb0edRJmr9nTHrW9jHHQiY5QAOXLrqj2PlUUdjkBdAHQSxe4K
WTfiv6aAcV0kSAgnxWI/en+Ob3h9isZLvjXBf0u6ojrNG4SO0pBbikpJ/QsfVpbIlfxtWXPyMIZS
fAmBkF/r/QYawXGcQtzerRpN9CvZ2LfpVESfa0j3AD1WzR+8s4zVwVebOB5tGvmpnddDGPf93EB9
LZ3kc3ald8mL1TC25iO9POd+PYYobJIa57T5P5kxFJ06JEzYjUK9ErLoHKQH92n1otIm6iC3Rb9H
6orSbrxshi/rY5M2efi5OLFvNSpgT7b/mQn8r7zjw109bQE4RM53LL7BjbOaEDh53onhxZ6FIP5b
SFZclUJWGO86XJfmxOe1tZ4PYDIGoXW9Jf0ywzDo+RLZZiTbREmdN6nxq7wfIEb0rFX1KnVYUSWg
2/Bf47d0O/9AIar87+iFurOAgGiGnwCln8yaTvJgN2RhMoPkGevd8Wyo2DwAEjNx7pcxZViZeXZh
LYU7igYVq8Z1b3yxp7vEFWdYl+sFFoOzP3NzOHlPWpxvT+LWECQVrk0kvFT3029+ieZghkyAkHbQ
suH0dcOXsqAqfTApbjFeHzyIHdS9tTHSJru/vowndPnAGKpvQvCs5yD1mAkBpoGOAS+sHFvUuQj8
qOYmxpCmuUIhbCsJouekEucYSZZ5wQ+qDXi0D98D0ITCWP8EDZOVhN0laljxsp4RMOUiBCdTeRyb
wFo/tez3+UcRyKL4zd9ckrvTO2mH8I757qMQ1q0l1sfHo5WUgSBJw+zhQSjjROn8VM4/gE7s5bb2
YUNC27RQJIlVq6v3pJw+ZbUYdroCr80aarER0LDUM08kSdms6xeJV2oUVBSmNPJkBPybLSDTBnv/
XxbaJWGj4ASXCMQc6GfD9L+GAF5cb4hUX18t4QBvCyhonBZEs7qiehHRHx2FDDLs7RUkoCWVEp9S
zuSqSv+4Vt9M9fdAHJjUL1RgDX1SIc6A6F8b84EWwLNV8vlEkqDcHtVxsJDAqKrBeMFf5Z8FNYmA
czXvsxIVm8UAKQ7RG/K8J8djTlLs4qZSrQv2H1mhIFTX40sgXqqraIw7UMEUSloaIzQxb3o2AblN
4Dd9fKIAXU3gm0OUU8VWXkFWcAvI39/fPZRB6WyCzV2E3wuTigvo2Tdl4AL7uXGP0LJhSMiftiNQ
he/l+yu84DQZNukr0h7X3v94PXp6QT3F5xTeBWfWs+ULE3YP6MXcjQKkhVqvhg2OHFDy3E9bTC3/
Fz3OEvV9nKPYuCuFY/C0BHMRMOzPHIHlRMObTgR+evsULiVolgHjqMzyd4foSLcPd6TWlTHQrGpF
Qj/zRR2ycYnu/XFfo5QKkChsWptRK12HOvyepB3g8Nhr8qzxRndQoAqrhs5Yr3UmDw4fgSnUIcOr
jlydZjASAO+JRGwVE9JVeFvH2D85tynDf6LnI6qoE6A0etZDVmXz+anxLuIW1qeM286wgTYSX922
2Kr5tA7xQgJTVsmqbnRmiMUogR34h3W1GhWWBAkYbpMp/SXr7t+TF/PAyFi+mJVHWLlIjsar7QCN
mSmB2aC7EmwIJCWUdwUIX3TN556a7WjK4akxFRXkvatvgIa7ByuK5VhXUrSFVlkiiKxBW3s1jJxw
3lzt+I+gKDEenRI4E+ahEwU2fCjzF5ZeJSp0CBCwtug7SVk9N7mVAmScN3vGQHTm/EOY3Hk/vwHC
NypdTilett09ObMeHRSBZk2rG6JI0IR+vO+0EUgnDDyqSiqoby6Y2bvbVvAsidcEvsgerbe3PJiA
qazPG1pOw4xIMX03F9WPx0CTrrXZM3XmwuUhTqd+NjmhnBHjYOrSduA8WO6cBmqcABgMJvnPu5o3
vRj6sNKayQNGXDBjcKKpYAAUOoLprnb3tzKz0595FA897zFs0KsgE9IMAA39CbLmhvgsAafC4y42
e31WUo816N7BBKNE0gt3QoqlvUEdnmeKzWMI8WE8RsynOna0bp3frg62zpn4zruyYudSBtDumLW4
L+A4lL+TgWPRU2b95wBgEJZlcEy9E0YthHW2Kyh4Uy0d5Rf/VNTWvzgLpldt9NCKm0zJJr+2zeZd
oNp08Wlx2Fw3pXt04tdWgIGX76uZXpyi2OPVA8iuKjy3TQs0MGBh/To8jOnMGqbu0YbhziKtjVHZ
7sE2B/crTwEc5QqBoO/pV/nbYB+lf/ufPJK+Xk6dH2Pde0pGKzevDbce89adwc26Oq93M7dq35zb
NMQV7e6MviUPzBP5d+AkioVphSGSXZJKA/nWrFp7g84n4KLei+zySImO5hPZgrb8h5qFgZPqwROY
Lpzv+n96l6kLrNQIP34tFqLIrV9f98tm4sVej2v6/mrKWhK6r7uPtNPl64OteBoCqKbUk/yutl8V
FWrScQ1iwPyE01cA5M2nORQbjaSuZ1h2H8WuotjHcmoeVks1Apao9TPbsRjblZk93JXI8QbLeH98
3FF2A8pXg7xL7Yf8x7hvQxXEwFQ7ev8QVUSq1IMcgK0Ba/vjtfUdbaUTFdv8dH4GGp6kyJkMA2o7
ZzNaMVGIuQhC7iDaDLSZ3IgwSOYOZW/opLtoSS/pajva4fiO2cjKz/WudAr33w59m106Kvgc7Rn7
zgXT/Y4cAXYRZZf3ozNa0t/gdct3KvkWWDkWgAHMq/ig24MQmUAPoququFeJuUhFy0ze7KKMg7RN
hluJJhUyXM+aoER0zGyLZz7Jfmbt0FAyRGPRUgwPKSb+gHXRhPXSIr6S09SlPG7Uy/vvN1/FF8p0
2mTRORjtCQNIwPIpOtLz3AZKK3p2neUyxfVZDc3/nn2emvlwR6JIWQyGNKx22iLqS/jP2pRK9cAs
TTYrFaHzPSV2tLpeYRLgm2V/upoo3uzWExXiejM5BU/6266igmKXmWxnyxiuLo7cnUalVWfSWQBV
6OIYmp9y8xVsOzSmNIY+ZQHsnOjxzrE/H506TId32QyQqHo8SzYqjpw409cyiXOZ83va1WSxIhxT
9+i85KMSiDI0JuVsp1CqIdwaWbzTN/rScYx1w80BfpYofbvjbhr1W/ipbk0PMLOQtGEIWwsb5zcy
kzca+1vnpn5ckqRZk6rSz3Kp6COM/v+2YDh8Yntzz7QC+FpoWE/es/oCQTxVcMJk4jTaJ96ljNDQ
UWn2jHkj2YAQnRj5KKOeVhA/vuPEM0kajGt/y2iYv45KzbFqeCxJK+wOfYb/TGA7R6c18bg2yyms
Q8tk4A+TjSAYtFmBHI5AbrND3RWwJMiysMv9hvOUPmUdkKVuOcV6/bBjOW2CSFQnkHterQ4E9mjn
np4EKBtio+GUhE166B/4B4IBrdERMOD/Hl9PkzvpraDXXZw6hO2FAqtjfWUpX+HrfNTgKjc2T2Li
BiMc3KaGDWZUBWsWjlzcsTwra77Pl/QBn2yBbe//hn5P+s/WU6NZumZPFROWs8D9oAkAOvJjIu31
XC7ifOpEt9Ut+CxfeeFumUWvG/yiCyAzFa5Wdwx21wldB7bNjQuXz3QhjwaNM78GwGsoZKBR9tv5
0+ZDu97oC91MfCzHBvJeARaZQeYFTkaffWQIceXX3U+RU1Q+BHsZLJTIK9kPQgRCfb8BRYlvfnaN
Q7PbE3alhfx2sv4sdYXvw36pADQ5nOKyqgTkH9k2HHBnBMrfaLFvxtL0kENiMFYIKGxmZp0N/eoW
UR4XdaqAAg+YIiVkugbDg8fo8epQqAW2IBrU+Q08TEh2Xj4Ygp1rlPRX/rvL1MEGru/gbp+MWSgb
dfXmGBc+RmV/cffy7R1KerzVRkJmA0CZs/rHCwM2mZRZkJjRePRMMpYCBkYFjGc9HLHK5/v6dfsS
p3/9cafKDg7PDSJKjNfKZjpVQp0SzOyOHsqjUN+INTChtrJzhgctOQKqPL2QLdjsFlH/qUGyvhEM
DLDGoAHIEZqDSb8J2qY3NQMqH2C2QMapoXD8UKAQgn1WlA2z8ItPB/pMuzwLzZ1vRKnK/lPMEa0X
i1k63XRUAn5Xww/8x4d2VQ3Vb+GNDvvuDpXnoKUIrT8pOZGVjKva/UFPSRsRS4F4s44L18TW9h/8
yAPZVtG/yb1DrksyvxBDcyh1MiIMGDMd6Aj8L+b1CZ76NQuPSFlv/c+sS4AM5Dr/0vFk3/HR6SJ4
ujUbTLF4sM00Z2mcqC5LeXeYcqK2vo9p+kLA+KDLtgQWEK5Dxj+keY4+5KjKoLxG9hrNrISegPRp
yPUJe+PqBT0PYXEyMVtawuMasNKqi1/TBBrkL4nvKZ9ULo7XOepvjtqZx4f1jqaF2hLcHmuSAEeJ
1EmpNiuiN+cPlzMdQJMnGQkCloRyyJ9O6SQCT4jYQ4cp91au+YIKQkHlraNxp0PP45QdRZWpzLIF
spKtK1qwVjx8o2g0UF0ZnMVY2AFTn1FCvDWXSTsCJU01um8srf8DapH7eFnkRD3txrcTvaVTtIV+
ymx0kA1rklabR/O5JxhEfahW8Q/iDa9ZJrmDyBWkwyjfO7dAjh8v+9dG9aZMI+6WS3ajrS162vKT
QQVERadFzLjuZUT9Rfo1IaA5Cn0sKDy1xgWsGqR6jmv3bG0zZ1TyyYUgZWqWyKkeZh8StCJ592oC
wsIQ15RF3SZaR1XE1oBzkbxBUtKesOtailuc6HnDaQEUeaFiJopKX42yq7EuxRxblFq7zz11djD3
u9/u3oPc/veXVEtwOzZIIIcFl7IIS92sa/sbcEe3xDA6uWE6w4gN3DxcRgIV11mbz/BvkYwngjGp
aaeU5Gud7goigbd8E6FAwRcEq85QZ0XVykt7g/a/KDPe0pNaWz42FwoiWroq6MjNHwXdP8yH1BL8
TfWF46T03O/TlDZgj6emPAQ7wj6/BSqs3Arr7/0GqwdYV91JonLadCkOJ0xCthicVbWSMSbIp80T
Cy5riFtGFjo6x1A2gIP1/WnZLUAuiGj4WZ9ZTyWuyecs48xYqAlLeVnxV3eM+lYhcN/EYz8RTral
2xm6Wk0l1QAwtyA1P4CFdDLIGfLJeQFVCAIaQxgL/49neFlVdAE+nYWcXg3GjocVsLo+h7tl21M1
CyqTifoDYpe/F+lic11i/hneDdNTC8jAiU2jN0xYAaTugEpjoJTRosDpFCKcXYs8tktpLUmi217s
Sz7zLLTJ1S/Vq4aQEis+xmULZfhmFfNafXSJWbdBmXIVUcM74+IUwY9ZGJkycZi9hTRsaJeP7VJL
V5gy3dG3YJLKlLcUsuSxHxrCcd4yT5vwdTs7oAOwwphpjfRBGm915hZdRjzYlKrJdle6vVPNlaXC
V3/xRMkGL+B+4K8x4k7+YXvaRzSwbymcPJVM7ErZtXHDMcU+xm7TETCjsc6dBwvj/Iw4Paddctp9
rE/RjwPtNKmynS4hujlvWkt5tOpd36u40kGLSUXQ/1h8Fm8wvwMPEe/KMWBKe50dn0GrpKcHP/i/
4zkFXRCHhK28Po06xDkaN2NAMKbzxWyHKkPUQUNVvOde3zsHkHQs963HW47XOaQAFxiX3Ny+wNh/
elfFULhEMFS6r7/yb1Ljzk9lO1cRySdj0XeApFuMw9DivJ7A2BoIryXvzu7VokfweX9UhbTvOpzc
4WWTEdHQ+Xng3lYyFntwr5G+km/r3arjOToksEO9FwenlQvvLJcYxHI8Qx1w3RcAWT15DXItTVRK
lWkbktHpJN73Vi9gsyt8WRVGE4CdXPEK+pgteRFW2O/KiHW1PrhoKJuNjPc/xjPcr4b3VSR+1ujA
vtd16BEPJ0gS1BaogRdmIDAtcewKcvmcW2FeC0lCzcx88b2o5ew8W4aYEos2jtn+7Vo0jfbBIiNE
7P7WYzhV8401hwgSf8hfCx7+hICuPB99aWfBKSu0SJDw39RB7iFgTMewjO3pUCqVX3Ghy1a6VRN/
fe1x4r21L1ILBGq2sv6SEte0XNr0hDvYvlF0voA3wRmGc5DK2l6NEZn73eL9IymXgp1G196H3W8e
NiqLb6+OM06FC2tyk4IJiXZPsNyjvWMS9yDMi6OzfPoKSzE7Q4yj/NGU929LhRfnh07mHnaJ0/Rb
VuspgLsLj2cBk5VP0xn2QZ40+i/ST2wrgup5gbyRjolfTpziGcTbbC6vtEePVKt68iGpxbxliHdc
isxU6p3d1KKPjvqo0LsKF/uxw3Nz2kj3eqmjIYK5ptkirKReORvnMINfhVkw0u4YT8WeCpOWHKa2
TlC4JnttTIcFOdkU06lrEbVIOc7t6KywosYZHhX/uOl70iq8WFNAeeIFxlgYpGK+qRaA0P5QSfWc
JfpwCOyluttqqc3A7OsqnBcah0KysnpXCWTlD7TKXR5jtQKH6UP4au4CKAcSFZ/CrfY5ag5h1dvS
WAGSCvPUrR2Kl2dnMbDS/b/nmC1dfpFWYlLi1MJzmi9vxp057cvgBOU+P/5TEFc0uc6NjUXvDCwE
Qyp3KGSZZ+uDeTdd6NcJ6cR3sDmGhpiNoK5z11zYgTqZ18E1t1HL+JKRaWBjnxanz1FPgFrfoofQ
paL2yJriGxX7FZ7xfTxzz54uHjnfPytAF6wwJdKeijtzPjVLooYJdyFd13OMNK26Gfoyc7Heg6a5
akuPeaIundrLqU/YuLpaA8kWejtNqnjQ0DVkIXULCjUop1V0hq4olH+zOiqWL2RhIT/J+iutblj+
gQgqABTahHyaykWAPMpVvlU+Q7+X7ISvY1yROkAo5rHdd/3eMrdVCGRo+2X3ReDfMvwOgeu3WL2e
flW+pQYHDuln2eVDqObcAwuzku2IPqnJ+sH/vD8EbpFvo8Az8ZroBQuyw3d+Dx5SmLDBdb4w3Nqj
zpE5OJjOP/l9J2RSuuOx5pz01Friv5OIlWlmoCjoFJcFK/+q0xAOdB51P3HCOZIfqgpN5VXiFeql
ejg4ixwczFfLNjBBF+gOoBis4S6diOp6atHeUjAkhMn47Udl4CWmtOI72z7Rb7rVxkJl0rqmAToE
kClWmw9qXZst1L702YmmWnh3fj3RFgThTskiL/O9EqdJiHtgDiJvlyFxaWGREXFI+DcosDOk5XvM
2LCxl/kZDr2mSYd1MpjJZ5ZdombS/G330MQzk8jH/QKY6BEyLlEkw755/UBpaL1r7OSugBqZH8p8
NsRom9UjqDcTe8f4lCs3ErVg3OWDNapSyOWyi1d87hfWGuqJi9rx/qCq/+20m0j76qKd/A+AZn/R
JKB/jlJ9ULP4ONJVpS1FIa5XrmZKKxeTG4w0C9wZzhhck5LxdRH90CWGpDDSmC/RY7rzS97tbiJO
z9TMHErUBLWsZ0UyXu8NnppKug90qFY6C6Rxgafajmow2o8IqXLjHx2LDMLTzbdwtsZwZPfTYGen
Aq3BVxBsEp1rEe2qS2K++lUAxnU1ARIEHguCVm1ssR7Bn0BTavVYY12Up0qGk9j3x0ThtWEF6P3L
m9QhywCK7SdRbCHvLGUVcqUEa0ZH6DfEZDWgGKZs8bWD179F8vBKbLMAr58F7R6HKH0X80PTv5Zb
GJ3pymJTXZyDzbgz+YPQjfC943dkvGGPFXnIy112S9GOrjuZlNtFk/jJYBI8GYiVev7hVCXrA72W
qcgiGaifoLSCFiU68RN4EQid5YGDNvOZ/KiOo0l5c16/y09R+D9LLJEIxHThklkogNTxwi0QoWce
gbjwQLU44jlJKOFa1U0dj1QjX7l85jOdIS6vH59Fkg3WAXmHCvGkztlYPpcUfRMsnzNM92FeVrgy
jPv4iPETcWSpVrgxv6Ntd5rElOQMqWGpiVz/VIRnKQsAXiu6hnnEPzBcVGx7JiKSnCD5x+Zp8rEm
gCHT8Q8cjWZdmS9HysPlQr0SQeCAf84rm3OCSgL7hIr6wNMasKHngu+Ak2xcXo0TWNppCuSgnPg9
tbB0141shBuOXaBT9XW+m4OYcpqztBauBIebBlC7VXW3DrcMI/Ld0oOcArBRU9TyKwpYI2yU0Dit
YHvQqf6YIM/cn77auLYOyZWCBPc4loDbJZoWGG0dzPiwYqMFR5U1JRuaw1ElTYIzuQJnJbsHIfVt
dWvCZe4VYgZrBwgnCEcNJE7DnXhxMwxVg1LqfTuPXaIVIentVNLEGMEOULKtGmjQUFyl+PmDWgCm
AQ1yQrkDcITgvMHZ8hnwAzJQMFoqyk7kGEpMXJ2LZZL6WbCjnmCZshOF0jlr3TWwmgrzXvDtxPsX
YfuRfKeB6rU6e5fOh7lUDp/omC8io0Q7OUO9cQOkFc4VpiZ8UQ/2KEbeHIoP4spWPldrGe/qVqlO
f5P+/yWXnRZraagsloh1M0YHgGY4q8REM6zYaIlmVgiwlE6vpSLhflwgyy2UL6u/9SV4YwYXkB69
1uFXcOGx8P11EKcYRsBhOYBx/BIevnNOJYZjU+0rUm1b9wUeHZnOSCFZEwJG3AKYT7kIgKGy8VJq
JGGbr4lI9mlAvunDAdw4Pk26tZ8iLTNqV6iRl1baJljUp3PURMNRf4/R21au1v1Ixqyxvyv0J6Cx
auQ+1MWTfUFJ9631uKGoXodIEdbg2WldXF1ICL3n54WqkweJPHVFlPkD24uZKHoQiFyOuRUtyhzj
wcYyo+jfhb44hiof7W23BwZZyOhq8hYmn6xV8eaAvUTA0y1ojUtol5xcllqDiy53JfAQxUWsHL0b
NaNluQYsDEJ2LSjkVPQih6sbkZJv5rV/Mb2gXcUnaThSyYvMhu5KoZ8rwozm8fxDr7BlyB/o88bN
rAx4fPb/tw6mdCGR5MhU6s/lojTrxulwSBqHQEVOA80qaxs+XSjJ3ajB4RuxHKU7RWf/JiielHNJ
9R5cKGrg01wNN4zBR3wCR6hXiShNYZmnXqZA41cf+Hql+6Urgn3ro2zEbvszf6Fqa20e3+HXL591
51gkprCTldw8xGL6zWIUec64lzccYQHp6fgWti74if+chxS5DD3dVrUBVUPteFuGFWAqDPW0uqtP
IMkzUlUOXx6724g/FmfiBFG76aTeX9BRRw6jJYCL1V0BQ8Ux8QlVBu8MxZUeqJgEsdDk2Bbg70BB
ARXHSzF1OelgP2kol8Rj0jAb1cfSvxYmOsts3cmVQ5h1qnQik37+giE0vyStO+LV/19pWbtusA/s
FlSiGD2K7bVfe9ViuSjmP5wBQZfrB3d4ZzlWBNvSzSjokEDTAh0OybOgJYB1G0aNRvFQ/b9syuI5
QB2fFc3lLJQ/4kKfrfmqmYHJcaFyQklvQUR9/zn86K2EKeF6L8lV8tuZRNcjmcDhmHg6l/+ltRIJ
MnM4FMK3TYSozI3spTDYKmS6HM4yz5lMI/ra9hJ7105/MsPy99esNy5azFME17ANqz0Nv5XlXfie
RKEA18/8j4yElEu1S9t5KA7Psp68CWX1z+LrV+t50s3R2h0bZlcbiWqdbONaQDGsM5nR7egc09Dk
y1vQONvrbMG6ITmzgA5SWlKmDwbMjTSyrvuU+FzLUidMjO3hzhZ5GlWskV+Buj4b0Js16NPR7Rnp
kXNqtqMXdtx9mfnDNxrJm2FM+TRBxUUCJ+ze5cjyrOrO/CnKXILrUQvn+F7guwD6WJt/+LtMHqBB
foZLSNol1tPqZePZ7hRxybgwkuHRwqSfv8Zh2A6Voq5wmH0oTUSdX9jwU3XlBwgRRNmuK+aJycIa
10y4KQRoO/CXvptpW3GTN9O3QL0JAfWoZpm9J4VMer8ANisWBK6fm8PUrOTBQjHgZRA0WFuKGABX
FXvZpsm4ZNz4wQ+4x2gHSzaUkQlGZ0+1l5TnF4JksKo8pOfUIAcpz9JRLDSyMX2DApzVYley6WoM
SFUoqzzYpIHLp+ADC1DLQ4HNUQ1/Wdp/R/k2BoMSsqE2NuQbz/AcTEfHAL9+YeCtmYkfdMCofEg4
WHv/Ipee+t4T2ZY6nUXA6q/NBGSXsobD4jrl8jYQGId2V7yDalzEPgus5V1rO9jPnZQzhYAKdujq
UqN0auFGN7UNSEE8InRXkcsU8HFeN7iUxdBxxx4k6FRgjSS3kegqGPZZ+1ZIeBdFYXnW8oQTGJ1b
vDNEt2kfL/plkRNcfsRzT9cSHAyel0lLVlFQgdvg3t8FevuwyS6o4AIXc0nm4MPN2UKwTHx/lN7X
sSYGJiSNXomrIJ6KqwhQPaxiKRtACCsIeEi/I+uAIedu7KYcRqP8q1e+uwWVuJsHsMhc1HQjqEdt
JYGj0ugcE3k9oH/bDkUtticS4ZSixVRsX6RPqDamw++sIMnQyShIrFfbbi+yHvLSv8Oeyxe2XYSp
OCRAuwFnS3vLqYq/lJ4/pryx/pbbifJjEE+PBq5W+rSvu1pN+C74vMYEvw2wbc08m8MZ65RHOX0m
DF3CGboZP8ciMFuUc5lLHPt96wNjY/Y6jNRy7Vls8s/zdVQyIcDNOpz7M1nk0PHiWD6dxvhgUPGY
pVEDiDMMgZ7N8qxJNzCygIxlrHOHZ0aFfKAlxfYj1VKwxVv4B1NBeGTqYbn511ilw1I7+r/2rDVH
QGNef9BRx+4fWNj0yu0lfZ6UDhhtLNxrUBF3kJB7Tp1QqRgvMiUwPanGWnd8sFNINShsnXpOvGAb
UXUr6+QzY6LMNbfSnJTyWM2th72kM/px41ug/uvVyIJPuBQGA/o7FK6G9c4EQZW1A5q4Wh0Oc2ft
2Ua0lI+BtgLOqquZzwePLhYZHdUeIvcseCsjikx64pwnU90poo8RRkdfbxx4gRh6NfbPkgViNA2h
ZnzcjoB6rj4O4oi8hHZXwIrhkT7kEKOwiA/EBtHkpWkWvfdDasHfy7ceGyOcmuRhxkmsBjD2FsFT
GKjgf+pXPCifJtOG1kJMxq7zgO/lFaXpa0HyHEoxu170nC917Y93RIs0TTxAoaQlT77vw/cdPL8p
23bmj1B3f3qlwCXiClddO37QW/VCJuCdfh+zjZzm84GhrdCA6RAqma3J7zeJ20H7yvAQ17lu3Yf2
ekv/jCSs6wmBoWChjN3UpLhWdoda0YDTiecBL5RUZhEvDfQyNqjymhjNWmyiwxh2bm2pNQ+xBGs0
PNslUpV7ZsqnVasqeSpnup4s674Xv6lxvigm0N0Vb4PWySQrQ8HqsXPwgN8uljAUVBfF53kVfogX
z3OOb+mwXMeOzurkKpAJm3vGkaSCkqc6/cvGHkUEOtfw+fkxLco+CjlqPom/lKQJGOfnBXI8wxom
x3603MEktzQgORwTaqzB0y1T8XDWyVoTyaIsx4an3PRDLDl8dRbEF3ZA9TLBkd90+BVrW1JwwKRe
ifaJpFR3hgzZ6PCB3cqyDIEssoqWLaLO0pyag8JvfDJS6JdefwPyS8AUqjIRH2+Z5t21wPCb4qhA
gWZb0+Tlymk7P3rrzjjc61iMLyF6hvFOsVZRCIYR5/jcEZjZIZ8MGoHQuiFX0Lvb3lFhfnsE73Ki
ZXAODBwFkHYjwlTI5j4Q2zXa40rLXKQFNPODG5pazy1mcpS5XLKAyrrRlw3B+w0c6xYOizbo2o4J
76AeDp0K3xy2EMFFJWHR+YuCKVd7eWjznPpfcxIKLKlFGyr49S2Bl2Q4qtYpoIJMBM+Yvw1TgytR
VqI/CNJnHZDr3eCIAw2g/jDIk7oIaiBGFKBBZMdlkz1y9l/3fnnhs7COjxMah+FI2O36FSsbqzxu
XkdxPwlwYHAZfTwvlj8ezmhwHToSe3jZjO5SYs2XhTjgpBZXy3csxBaRZW9JhJlQfg58sBLL+IwB
9S2DK0ZYuTtPJlHZ2DTcZjzQrL48TuOiaQY+PlavcmXBVmrgVeCFmKOWjNGiZzWxkCDlrh7BRaNN
DgtrsLTabt1tftPB/LOvMy5rwAz2Zg739FvaARddeUBKICla14bcOqUUD6U+NnXmzrz3/Ccvecbz
ZkXyMQBsRgceUqNmlZ9soNUSP9LOjOT4eS1GXt3mEpuR72TGHivKK7z7WNUVBnH+nLuu+VkpPP1o
9Nl+8rjxTyvLZhfW32NVZBUY2pLOACv5343aPQOOeoYMuLk1bLLtmLgD7ch+uWOydtpJyz3bBodp
6ytnbAqerEEzGD6j12WBKU5PAK+RiwKT+3S4gYVNg/GnqdglcjiSNs3WAHcNPBp9CCuBP8ZC054Z
AuY+/H5OEBiSfHT/03DWRiilbirjEWdV7s+a0MMAz2DLbZhfMx6vbR20CJXdlDLztcSClBkMzW6p
k7LJDOUaVByXqUS4BeU5nuCmwYY2mmWJgCHDE4vsJQZRlf8gIQQJ7qIJi80Z50AYgw0Y+lsb7Hri
WsU2/JHJ21bl26dkFSTNrqRUVbiGIwsJQghg0FextiUlYDE/RVFH9v45/Pa7UK0+2XOuRgjT/Ntj
I8bJqY7vk4mMAGZK3wDXF2C8zOr+92SMnoWnmmswORL5EoNahjJ99BxAG4cYq+4yPQZMTR/zAyeY
49kQ197u108GstoI8hEXw44neWzKxUyE7b8BSO/r/7tpdm2CpSAURTKjSdMKUuAqFq6ssoisk5gQ
cPJhqBExH90mFLbCBr5rEJ3dLjrHQYDpcxgPfVZRmzjfKFF2B4sBJHTtxKWE+MJ2BfaMwD+DYA0h
bhDYIO/DyjWJlYMoPbHepZLY8rNRlZ1nnf0KCZweUPcsFku0vhY0UJSTFZcl1Gs5KmIOFtuSvCMF
cUlOGj6wAD1rdz/t4r/Ecpxh0MYZoYgfIwce8J5BxpNI3wnmgnXePdnopCav311dXao2MaEK/Wp3
qEavdbq6lH2rfZE4HP+Ud3MmcgHkdv2Gc6iUR41rSaGWCtZo959CedqgvGlkYbSMJyyT10xrlm6e
FohPsF4AD7sZPUlFH4CvM25CjV7V2D7ggA5pKAG0ZBaiWsdxlj3WoKQxSJoJvzXJaGTPkfcWaAXZ
T3bXbzBBqlxkAeiNhS8E51uoIMRpggBLVPAyB/vNHCZLlCcm+P9AyrXjZWHs3bnYadFUoHxCUxZi
CrDu8wv2OfB8GVbIQV9A9T3uQKxzGlYv8gRwwyBfJKfuPV5a9cU6TaAGpAj41nmIfsX2+gx8mU8W
XXW0UiUfh4B+YK6chLrzn7K7hKXj4BMdrq6Q2oosGW6l8VOKwxwOz8MGfwUdyVUGT1OJsP2JJ+cg
1Y1lbvzLsHQjUVoj67F11hTbxDQz+cHYRz1+3F+tVk8RoIptnqqeHcCXHE7ptf70jSo/pFBIsZdi
BErQ/07y7XQX5pT0un8AY2iOK6GxheOGCbPSFlyZMHuPeoQFhUzxOiJR8H9LY4R7i3GdhIPKXuaG
9taeJ5SdgtpkGuBGn5J1/DGryJIamVLvXZ6OgDwhruH8O8Neyv3YGes8L1IIgWwG2kFfmGLy6F4E
grFfwlqoUYwYwSzVMKvl6C+3RvIY9ylfVoUlEuQOcXI0wwZ0P4SKVzwwh52kfXQx88HMxbgxLZG5
N6m6GkQtpzHdGIDJuNQFwjwk9JD8qfk4mUemyiC6uT9pTWYkT379sEy0KujhBZajF/V/88uQgXMF
/ZmMOt98njniaht1NJ6J5m+2NSj7NN/6ItzTlXBdrna5uhOUomUONx7VL1+aoXvk7pt+eLLpN5k8
AIZ05p34orGDpIDk7jcJaOcVlgM/U69hvXe1rqi9v214AB5O9xSgc9DLe3Xr7z5NbzOVUw++Q7YN
/hEv3jpSTz1bDHb7VNd8OK8xKhAYqWlURCaVkj3JZNwSVme/FC2Hxz+OQcJ0UXH0GErffL6zLlom
ahd/hAlyXpTOPQDeswSe6Q1mbqsHC0X2Kpj7FXvEmPiXOI89i8obJoTgx8dn2gKWbOYZSOzEkuVM
6riWhHkg/1FG4Qog5oz9SU8oL8fLuaxN5Jk9ua/EHtXhYZdmmvkZZOftkeaWVhI50bMmI5QrK/RG
gCtQg3Z1fXonyJIFvRDxZf4vdUD7b/CcOyl69OojWoHxm4CeZNGmVS3eFsn0jgjplI2/wCUyF7FL
EiIlnoq/RKxr6pQC3dWZQCKfkTk/5HUExrFItBX8eMp9Buea/GbTOm9dH4I9LwBPtqOF12nYzEr3
BpTD5xdih+S3VACzOuUJ8lxIU4YTMGBir6mF5S4xXBWkokbmy0anyAWurFfqGG/3agyYHaq5G1J0
VCtjQpZPohcRpI1seiKv7mza5QriLm8BOisWlu7bdZUCqf98FgP0JpfhDjUShSBudpya2uydzenv
Y/EUlmflpq2F6Vd3uTC2TSdDdO62NpNcyJb0nEqMcitFL47SOjKkDFHxlJP9+G+/h8jgAPq+28EK
e8bzsfQkFwU7DoY2cTv2td4f7OyzFOGT8eKOiFDvOs2QVtYPeAcTB8OZNszebNxlzhH7m/Gs1ojq
0mw7kEeh1WvsMzQ2fjYrrawRVOIDExzlO68K/1f6nb3mhOLfE79DEn4h0hiTeaT1DGWzZxUwgQGM
h6NxIJlZCAG2rZeNu8VLrJxxu49sNgk/YeiNlIke+rXkOgYv6R34iNYxnr3IGMsPCxpqV6PnJUXw
Z8XI+pSTtFGuTpW7e8JszqugRwNPmP9sKFVoihnvc4CZYGiV+7KtD6bhQA1HKq9W6lT6xQRAAmtD
F12Y8Dfy4i8zPsSk1GdPbjCyYh57tyc9mgs34ho/FylPSSaTSt7pitfwAnCmduNQyflK3Sc8iH8C
JzqbyuJXVuvTAwX1riDAdL/6mG78onHMaC2oa9EZLPZV+noWEP0x4GpWjfeNkusda8MWhua2tAn0
Lne5Ql6wkyF7iD6q7L6qw+T25jARPvLxQ9jaxwMLzjOUSYyZslb4ewISu1V7wBMfMlm9rkrHKvLF
m8Cgh7j2iPxuGsre/dbbnqSm1HnQ0uUege1mUCX92JSkXIGzGa5nY90Yx6+Hn/beloTIi3Np/2fH
liTAD6OA+NB1yQyu7N7vE4g1CDlfKf6cJsPmWBcFDYtMssVzcOU3HHmCfSwsvIg/M4wgxZZ9dYDe
rOX6LmHsSR4lNFzxgsyqgyhap/UG72GZbhLGuKBqelSJetS/Ei8gZB+B97Vnxkr3BHiLfCvzAOdf
Fha2UOhqPg77nzKeTupvPu2/K8h28NhCii2BAyzuEtz0H0RMg81PjC77Ia959OFc5TJUUJ9tfL0+
WSmjWp7ycbK8yQazM+BE8GXT54DBbQjpP7jify4A2fh8dg91J/ls0GTslqvTFfEL04zMWKnleCxp
ntQncoaxruTBwEX0sgOXhlwRdsCVCe+iCS/+BWeVajA3uvRWdKPzIZs3FKSiJbbtLeksaB7TUXB/
FmXOFdm6vzu2rauCqQJ9KEYVHnh6ak/bUDXL7OBV3Okr12zD6qYHC942mC6VMOKtVMh/F1fqc2Sl
k4TONqwEZ3hij/ak30gJwgnHdNaxBbKUYU87RjlqHAMUPxsazOe0SESMD+j6DNE/yZUgGFbaDtQa
dOuoUZ0xBOkx87QaUpIWr4a01HWJXplSccXNvjsU+P0/pMn49uuH6oXmlWpsvC6akfLvEwHu1njs
daJiolpOiNsueoMbDNFWiJUI0NHQVrc4cApW6YokWXtK4AYOoornss2EaDN3ihVw1BI4Xd7DNElJ
QE5yiJyjuYrxPITib48n/qKBCLKkQUqW6OiEIsx5aSHJ2ZwKpwlhW2iJLMiVkb3ORO6PlVQHrc1o
5RlHFfoEqMFvakph/WnN6OROvFodbCKc7Bx5fyO4KWJdpta+2v5I5kjzY0TLzPEk7v/fYT3MTrTd
snSTlkTMWuzBsnAZ6v1Vhh+h/leZlFZM8yyJNKdKTnxFSzfWzNjjP011q/ChOoWHl6hR7o5Dd2w/
9wYMg+dHuv/NbZQvkob+gRGxXD1vPzKHO8EB05AFD2b2JsUWtLxSfh/8HPsZi58JAK77fqBkn2GO
Tq+z+qgwiM5D7xujyPWurOGSQ+yEdvPBxcAPWN0wlS6tQRFpe0cn7AZOUs5Je3FWvo91cLkl1hbY
B19wAPqEMN8AGFfcziN4n62BzClSp8YQWl6pM5UvQHVXszgm0HR8IiqZjHZAAKIueyN2b8EPXxFY
1Faj519GNxASVO+NTLQo3OMINBKjynJ+EQkC/KxMb6ARyyzscfgEOnxp8FLbDMtZ8D0teprjQ/UR
g8K1naC3d1fKHj1Z0okIg83W8sCys1hlqKV5fpoHMf8pHS8ldxBUcno/ALKitPYVtLeQScLnwUMp
ooA4NfSoS93J9PF5l/FeBR0vaRiO+7QYveYTxdQKWDHZElGFS+IoW7HgXo6xNDXoUedzmJIplmpH
oF1fRBIg+rD7Vh5gW6glGVgYT4pagtRrt+AOQBlC98F35qtY8zEaUdnlD7HQYutafz3c0mYcf/N5
b5rjFqJzkOaiycbm3kKmLqzgEgmVqX/hP4M2MCtJPuyVnwX1HvDEMLUE40uZHZdxykgQ3XbJAg5E
Ds2kC8rdrfYn9tmkT3lQFvIq2Y50P77am7ZZfLeOQnQhOSUdSjLZMNl3ikhodaQ0gN1DpnETZFR8
7p3NP2WMLVnKxqa9oD05sUVJjgCYtHkPc61Pb7m5w9LGPYf+Oi3MKIAz3W8ysGhHsSiV3JLvL3Nr
yywwEe+ryyIrdcUg7+zFR4taYFSluaDJ81fdERo6dsTJ/r6LVZBbiwCT6ueLsGIU+QoqTcl4SbOk
XVb2FDuC3M649DUMq6ksxxERa/+vd73EW0nd9iR+CyFhDd/CKPZ+EUmnBbrrI8HJmeyzciuYIV4c
vo/P0IAvKuk6zskkPqx2Rt/oPDd63tnSGyapIAy/jSDpLPMfuGMedFGTgNWFdKKhsS+5aTHlgR4q
1KXvn/FOeyNvFFMLFDWRlN+ifwLTu8YVGY0lYYXmzO/FrxaBGtMzZZiKhHXv7NX/3oAvvS178+eh
tsxmY67Cs0YgVfq5x05CDdLvMj/WrhsRyMmaBoyFi5i6EadKNujfqm8rM6Q2G6nsYA6gUaB/n/fc
VzH3UnBg+/yk5AMPGY10nNnd6B0GYXWPojkwValbFoHHXaxt8343zV2YUpSlSMxwCK/1PShQXw8T
3/fRcd6/i9nvc+ZSy726LQp8joveNUKPvg/2FLlvLS1cFvqhvfw/zNUrso/JIY5LgrYr7eN6YibK
rcAW+j0ac27W6g5Xk4JBi9iCG45XSipcspi6HWaVg9ntsRGsb/+LYtk43UWJSZWUuA36aZ/iSuE3
chNbYxmgFuxnZsyibHrN8dePJ7YRK/fdk5s30xh3Dx53i3XQj2OgneXCYgs0WqqaDG5CMzqQF0v6
fR7bsMiCUr74NY+W332qF1jqHid8FoRqyDxE+BuXdwUYdk0/uu8Q9FNZbRenDQCFNpmboe2D8V2+
Q2ZW3nFPDqKds8ZfjdRrKQnnm/FAGYM0jtlr/GGRRZcrhSsMDACaig4zBi54MDX3B74m9OA71alv
Psv+QWPHDV+Q8WUqNHSyb0ugFbhSaD5ujKM6aovWz4P6RMpPo//h0anYieoyfbNs3w+8CSQqDEPz
ZMKhFZBciBg5+vOEIJTNQC4I+FOsYtctKlmovG0uh/vjRyZdGv5mRlVgmoLZJhI0R1lwp+pLlnVI
1x9BHLgAHb2jHOS+jpxatXZEbTghMFhXUtwIQEkOtn/c1fbPuDLWSovgK2n5EmxDhoA5xi8LGrxl
6indkOVV3QIhPl/bCC7QnwK5Pb9kwxy8mko/cR4htPxZ+tpFoVqk5M39VHFTD3BmQeuTq6aity2C
r0+90ZRvD4/GHNK94q2xcSf69ThuaFteLt0fDDzf0CT0FBOf0UzB96p7HUPXIo3We2RrynxxQDzi
GtT8nuFC6EH2SRvjbIcCR9lsPruSjOUBsQXNd8BVNRAL7fqzPvzXIaaPbGQTe8wTWIutfynr7ROt
T5OOTIG9YCTqcUfKixRtQsCvjPdpAk6o/tZDhoTU+m7Zz2TX6H3zSTToV5GzE2RT3XSkxbwqNg45
TeEJtvZfMqHYdGgBO6fOb4zH1793DzHF0xflCE5v4FvA8KSMfFoltq0IUqm+Bj7wDtHmFrSJMFnN
L52tBVMwCRBzpYiQSI0BB7P6QGyaVeqp9k5AqgMY94KKQRQEU1mqlMrjMxY1q6CPD2muodPoSDu7
L8/pxmfgSARalFj87HpkmuTTHlZNN0HOIMUVaZkYRbw9AwXViw9Kz4voXIp2bzmSckCmTM8wgakJ
wjdNsfoz3TqzszsKNUiFPrh8Dnm8McB4t4udRWGbFvOgbPsH/Gwste1xKLXWDhthZf7UHMY4yx+4
t4x924dahYcnTJHMYB6pGPQrI1lmPWvqGy/DbNBIbT55orJ1Axi+1QKG1te9aujY6lWK9A9iBXDG
RbTCFJKMvEcyIFC22yKQ6fVJEqj8cewFzgwh4SZrnD+toHY9F/IwHh/V5fsYfdinFZ4n3m4p2n0I
xO/Mn0JONInwkKriPaoHM3PPkvC9VkDCn0/PxtoeqYrtbT7MTnNdDFxw/6ASZbiSzf6kL6826vqI
zDoUyeTdlOlt8Krjf62ZCABRN3cr8rd8nvMJ8ZpZgZPEkVjbBA3qHFcJD7zKV+WYvnAHg5QEsrXS
xOt6Eoh5WH16jklTOMDbSXagTI7j3OMg+f503PZLXw/6k7oIu0ZTT2x6LT0eCIGIuNQootvWZrKD
K5S9kRKNUFfAhFEg4sbHLiZCcoEEehERWcem6Q7tslKG5qhowzc0gQa6b9vhSllld07Vmw/QnT77
cwYM9MyEdNqd6aFEpJkak+XQ0VcWn+yncr4FJvr5GXaHdn0rfx0RiBUe4oOkzPRkZYxWK0maM41z
++YZr3zvHZErITuD3EoJBBUD6ovqBdSI7FxSHZzVt5XfyIJ+PiRvlQRfw/cjQk5shRpPZvV8oMQv
f+4PhQSL67vSYkVO28HI0r6wugXFkDLuXPtx6F1NgWT8VFwVGXXBUYPbxnNHLB6YNoxNOBuZAUjb
Kf9sfCtb/jmyZd65IJx5Eq4xlySypL+ga6SVnN7zvtxAftFTFO5FVk3jmOukjGVPuJd1mV8WCMZd
6J50D3X6qP7eE4C4DeiVuM9S5t4W5KuA+Vuobt8tLP0sPNHooxqA0QbboNdOGXhAH3EHAAvaagdj
clyqv3niZYT7Mf7iQB6+KMm6/k2n7PfT5f9fUuKwdShXx1yDLRsUJzRD3Pu+XG5cuCT7Vkga0dYS
aoqvx58nf0g07CNA8yycBOi43IyqICoHyab1+tXCVGOtRHd5agmCXaYJyjdLMPO+bSUyVgRYa+d6
d4Si/Dylgb5ujqAQ2JZkdRAk5LWzQc0CbQaUSfzLnIlXxKMNpq5hpOn0s3OyWfZoDuAWt0df5ZYU
z7D5nC6YoPasef/4vBq3On/D7ckPnjwXE7/+xus8zUq/Pp8lSyzZ8mBa3l05I+0UnyAarkJAKZo0
Ny3MFgp1vBlTUQ1EsCogF8XyUGLn2CdzPKFUM2Egz/E8UU0la477tZcUuCQT0LwVV/47pwMDnEFx
uR392Mdh4SWZBwIpS1GV8yZYhlZHYygxnomHzrdUphuNt1tzCaikf75BktBymgn7AXFbOAqTqx0i
DxLQzeGYZccTsJpzRllPJ+5PkqWDTHFw7RK4d2+6JtxXnW4mbSrPdiqs8QuNGuwBS3oy8wHlR1C3
/UIvEG2cupp5piqbEsQMFWejljzpupJpp3vKbZdMpwwrG5yAktKaaChboa/4xgAt1qCq2+cjtSVQ
HHtAceBhT2+CTHGcC0a8wpQq4jvwQvIQC2j6gj+Abi97iquv42hKywo7PJTc8iv6JKELHf5JaKsD
5xcEDQ0l8enthY4FTGKQ42saA5+Svj4iY9yhdk1ccBgYViPHfTjZdaISYv4tsK1tGNoVeMxXYlk1
c2kGR9RQdA05DPQr/4oWTziSLrIVgDohelwhUeObMR+BUHaECE6SGdAPzn8GCGXWMQxXvvv2dcrq
rDdoNqf4qeOTa2ACO+O/GyTLjuRISZ4ZHIt6Oie82LyhqpYlyxrsEl8fVoaezORaRApPXo2AStID
0NSG5HYkgmjVBZH/x/eAEvmRGYTCpLdQuJDhjS3DR6e3kZR+s1TfyFcrvhn9sEchOSgst8l7bVEi
4hq8tylqh26pOk2NwF3M/9QQF9rPOOiVs77kTvosX5dM7EKO61uew9y10Xr6hywXbJfzAnLJC4ao
nMV5uyWxito+neVm7b6dSOsmlprXClsafQH2jyKYDyHNYJWl0ly+2SrDuP0Ei4G+24YJA4NKofIx
PosIY8RLTcr/5TEIG/Ju+RXf+KREil11BgGGA7ZQvAEChDhv5p7R8JB0FQrmBeBRGUOQ02JSz26g
qF/I6M6AE2o7wAUjHw8AhWTnwLG8xfkkvEdkC+xDzaVHI+/Y6mphmESGwPbs/qo0XA1oFvYHh/34
PMEw88aSKXYX0SMTBTAVWqL8IRHeMYGmu6MVZ3+eZSJlBXOPHyA0vR/r7tAxHZxc9dzLBxb2NkHp
VS6hHGqukykE0LIfs2KMbA2KHhnIoY6dmiUWDPQYknxzxnOnklxET1h0cwrcJyf/L/wEkbesmt6Q
li94665acqy+zOViCzkFtH19IOJdNDFHDKj//dFEUFUe/R959Hu0HGTmUSamwq2NkFvaeo7ZE+TH
6RLeTb7LnTbiK753hfLGv2SmvlprgLgAKFFxgFxF+yLhUf2GiVvo4yri5mvtv1WW03apiP4eYj5u
3hgchksOGUTkQ7rhU/1xLe8vRsewkfgIhu/qlwq4d9omvmAoyY8lGrEjJHcXLBYCf7qQ5OWG30qq
5hpf0nt/2s8SoM1cU8FtKzupcxoYwwrgiF/EGNneUiYlm0MfhcN0J0WM6V9twWpG9xVtCRB5uIZr
qH1VvS+AT1QVwNR1+MU95m25979hl3pV20GIrWz9VQE50x4mQD7OOR4SJXM2uZ1/fIjfeW6FTgFk
/gg8AvVZXNMCeeHMk5frxAAeFF4B7TtNvTc/FcJdZJstgWra5a6gJUvmWga//yDwplhq3Qwz2Y1+
lGaWtLRk1Oy+cXIwpEVqyI6f2G+Rb8ar3O3FkhD0We8yhqTw9fYhC9VrmPNYPcBIAtXADP1kg8Ws
iigOWmhnn6P7zYjofnosL5QtBwud4qCb87AmkxaV3Dw4JnhaS5VQj/JAbNARc6Fo5w4ddJx8NP7m
cCI9b3YSiHyKdCWekS8kF0yeEZ3wRUKIibJ+BJdYkREyNDcbjc+oxTgOd50G9asnaLQv2RuzUESq
8pypKD1txrfrhHq6ADITd7oh4kVCpnJK2qFu+mBxMOqC+KbNMAaRbxqks3MmBzBCsOcCssKOOKe5
AsJr64DJJvfw87wnDjTL//0TETBL2PAYoNQGX01GT8Jof1qAuOUgBdgg9oGP84rOiUfmOJDsaZOW
29eaFPZQcXZLt7TNHYJx2xvEsNG9v65Gp5mYiDPxuZ9ha6mQuI2bnocSSAiRxXVywcIneFMpQVQP
qc0iEnmWDNI4D9u9bOigNpcfXKa8G9ZaM0SpJwWdVSQpZt30znqBDxdSjBNPtnwCk/hDYg12VOpX
fdN/PMQTqh1zrJAIUC84hXvLw8SjjeCsTTYg8hC5jRErLoTTQ1xpCyS1hjlygnnPLemIeua11mKs
ZD3UoyiFQijbq1/Xdd6FKsVpUbwmdUb1rPRym0PIge5VypF7m6Mf2zUdJCZLSGYxKFM52zOaZ31b
o6Gngf/0lFleNyMI9ggC76S/jZHM0xkLkJFgbMu9wI2MJpA1YfyftNtZxkzFh7pXKz3zdumQMBNC
bv4FIkMYxaRdQwtTb+lIEyD324Nyg3CBQFHYOKr7qXo+o/nTUatoLvNMATTKUVDN8I9fhKOQYff8
xEXRBr8Hi5DfDnwXO9F6MshprsXBUANWFhDuImwyQQS2BWNtxes33YjdAfhrVFysnbx/f4WzJbBJ
BfVM5g4NviXgKd/Ns0M3fWkPjtkzo0urqIf3V/eijEoU+uAtSWz5K4vykn6YQaDLq4ty8ZnVbZ09
CJfbdTI8At8yAUI4bnQaoV1h5FM+t7sY7Jp6sR4qGJ/i/a4/7i6eIM/LxlNqjmweI036cvdaMW5y
kHa+1kuTqcTj6wvOpP5h2cGLFHrcoZQRcIswIbB0ArW9F9oDV2fNR0DCwcxtYc+kS1xDyZv4js1J
eBhilYiCveyYBUnxEjFZZGu1DQzu3fKeKdmFW+QeWKHIvh/zAo5PNqo9QJpHXGHgsadY0HTKSGgt
9ExM1ChL3sqXJbbPVCYOJ/o5zRNBSGD5yoyN9pGd0lauY7dcnLATyKWIPKLQdMKpQG+hVtLXj0vR
5f+6s3RU90fEeW3FKv1/sYBj+j6QsWEXc6PXbo+7WCw9HHg5VJua7RWiKRYVQc4RHoFyp2os+Rw+
2CfTwFhKleMP5LBb9DMAAy78IbJhyPvYAGGK7cxYbOBDb1Tbb8aaXtHl0s7OrhjO5bGP/cvRHzXC
LPTShGxNMWIp+EMDiibr9ncuccz8B5XIiYTITBCoojpJkqcC30PJbfaiHMihBxHt62+UzzP9/wpS
t77deI020+6L1ISyj4jsniJL+aZaNmj9y0aGSwy90ZubYw7zTF9lY7ybbPit2mK9D9sXR9xJNe8y
Vu6V5ngxaY3+zOLP3tJK4j22fQLfr1dD7zMxfBcy4qEzREoDXOBeklK+MKerJ6hLhIsdSBxiHdIR
XJlnSukfbtlqBaaMi7weB/rM8qF7bGaQl8PVB/i9jEZVEFJvLVWtfvM5ZxwrydjSPA83Z3OyGF66
fc+4uuiQ8CMObBDZ9RSEaQB2jfTR7v0ED8d2X7mdXbBrwGiykEZzwEx7DXcLQsAV4SV1z3kTCXWl
5pS8Wfhs0ZXwlLjCSvwsZmO7G7p/L+FGlDzzkbq6hnmi2ev/zJ6DadQUSkG07CTi7tqihPf6fxDB
DQg4tdmfYSTSkswDht2g6Nz2KOzr3yB1pnmkl9w+dbXLH9qgDygUvp8ATOvyKRl0ZYRBSiePe6rK
Hq0/gZ86k6kgUCwnzOID0slOi9rJWRVls2ayyfRyQyozSLgkvLMljAFfEG73CVwyj3aTwYiU4qPs
D4B6b2fCaobFb/C8KeWNUlkuO+KTZau21ZdlJg0Rx6iAGTUp5aL7ULdxzjahBJ1OMX4SygHw0cZ9
wqgov9UNICgnZOB0TCE0tN6XDItya3yqgRcgm6nOkJ6brSgGWZ1BvvO2N0NzHhe327WZ0Q02PCMq
P4UNON6vzT/W+gFOZfLZG6mB58mbBNRUNF4qn146zbR9z0fnF8mUw4scnB3mHWT0KEjk8/ghE1Eh
6GAsl4Q+f9+/lGeL/4iK7AKC9e3iKJJuneyOHSGun/UJiteWurar0LQJPJCStZurPeSea13X+ObQ
cf8jtqM9QVORLfQggRnV7a8952SKmjowZ8wSByeDXAABTdIhlcCIE9ngc82X6Z9x2KNNoFm9G+Lr
Ch4akUTkTQsW0E0svsFRkZyQ5EVm6BLoiNhqH6xGc++hjyWSu6GuWmQmS/sU/OUhl3kzokQ1JYym
yQ6dp13mYeA/Ecw4GYTUsQSKKhHjZ+BIGd9Pyl3ugEkuo3DwahD1wVXZrT698alL5DZtQvRR1h9j
jfxcjCm6TUyp35AVwu2veC74Kw8uogxEupzdtlCYFpVelu7kc/juEKjUJ5xr7BtwFyLBa2T6MPO5
0nAZECwBgFyYzJK5+USYyW9U6cl2L6WqmvQUXdH0Uf9uX/icpQwRA+OCmbH1rfYjaSXv/woP0Iz3
NNJ8kp8HzcsUsKXxyfBSGp2iNLPQVDzrrScnJAwJibuYC+lJvcx7IdTLVB3YUn99nb8AbHg1GmTg
9va16nvOr3lgI+bU9se11IGjb1k2IAhwjqQqHolc+xNHIDgfFcKYzMJW4s9zM9zC8bEzSryZ5iZW
XZMtU5bwgfvqvJZlyeGyfXnhNCsL5gdyz28FNS3xwUlKb3T86L4chKrVIYjWSHcqsS/roFtVhXY4
QbMkhZAN1zUlTfas3QGz/KfIr3e/0n40OPVHN01g+SSQQvwJaXg+qKmYlc/oL6rn1DPZhbUaXs93
RiUTOumeauStoSRMch82Dx/fhgQtWd4CU5GW714Rbggcm9vPxqhOF8c3Vr7EnL8YwGrMYN2QkPuq
J0wPFT5eT1MOaQxk0CtORFOvPFeD/80av0pEUwHF7kUzyhkk2wtkT8sRKxTWS7qMXST/uue3Lblu
KyVl38Xr4487Ah5RKPBtuWzlxxrKbfQSw9SKF5Vx9e9QM4w+ePirNfl3eeDhv0OM3NtBAV35CoWY
HmQorfPzTZsmHK00B42OgLDil+7DY8eLPUg7i10qbrsoKSDsc7pjdamQtPVop3uf2Qj4XntHwwx1
DjIf4s94j5KdKdUzXDoCoQFu+rC5iD4bD1ZFBqKZVuemlm583eyvY71IFURQAWtx8n5By7JkkCJL
T4gF5qKk29fPTb22AFC/7gTEgPKWKk1xTMWKfBWHfaXU+xQvBUktgWbgi5byY2rgm0qK0Hu96zD/
FVH0SIzNJPNd3oDeUIK24P3BVrJXT4EeLStruam1R9VF3Sz5HnJ3o6MxF2Z0saafuhYR8pZO7Dvm
pb1+2ivlcxTVBHecrcMsF7/59zxBFQjnODXvBtoKS4JoTdJWd4AkuWNXCgyTNNVHo4fTEOsamAM+
mmE5maDT/wBWN1q82QLzyZjJiZTr40p614filNqPEGfGbL18LK55p4IBaN33ll5WK+Hd5hRnYx03
NVogb5/oY+kPcuU9/abWxbPYBxnwjs9ptTt3S6saJv9yOAs5rHq01Yk75KuHlbOgHk/aWu5pdyor
fnRueW+gdlRZ/CWAn+Ri8/YoI3m53izUgIfHL5OMrcLTiesf0BloL18WTtADw6TJrpAlrQTQ8dIo
LZgLF0Jb1/wUEBwtEGg1y/CvkJDzuDdnfelZk+NTRKG9LWWdwYZsBqLhGXN1ruihIRu4SQ/eF6YY
7vF/2mgst6USk2QU36URHvnOkvOz2VMs6Aaxo7krBNqsCa78yz5MKwDEMDxBbeObiTIAiDaZb5cc
qsMtFg6vcC/9YeDYdAurx8zAFkeCeIf8FJZLSE9F06+Ups8qe2Eh2/6gF94SYwgWwmrYsM5fevHx
PX5vX4PT0fEmb0k9EGP2HU3ESt1OY98v1UCrVheik/T9odOjXup5On1wy23UxB8Mp7TW9Ef9K0WI
imgnWPReVXh26LjWG+nYKnbnTvXrCjySTVCMDBBCr0PBDloy+ZISCR1p0xh28WHzvDn5VFcRuIYA
HwJBwVbYhjBes08m8dM2g5Gma4q1UXGYrkcQ0sJoh6B2+MBVITfpfJZ0MgUqOfJW3n16SNy1esz7
I+OrvQQzDHCysbn55q+j3EHHYfOmq6WqXByUfXX5RUcJXPfuBpgGFiQwLD8oIvUOi5klmmQmetUe
4KIWsAnakhoZRqVkQGOlFLkqS66I308zKRdOiHUbIcIE9ztdS6ZZd998WL/OmQn6b/s/EMaT4YY5
lMW/nkiuDZO+jmbQFfaevqB4ufKkjDEohJYW1rlJd5mMdA/S3V3mCzm3t2JKnaIZOc2g/rgYCpR7
3g4VqU0YOd7p+PpCU/4lYXK2mmaWuuImQ1YEQzqzeGMSssKZbl3T0GBtgzta5eJVHjVQ72Vt73ti
0NjIWFRrDgoMu56Q7KZ6M1n7+miArb3lAZr23Sh+Pi7MRBJoKEOEy0qLeuZaq4s3kvrZdbluZVWc
auMr9bBpWhhvJpGQbdsOElWk+Pwe4CqMdTRRJCCdMbftWVLsxTfcKG2JSrinSU+dG4qP2gpSt1BJ
WsWkYUkBu+tae4tLP5qkZseZ4WkAlWkNLFY4M710xlBOxHyH7i2VgPRB0yEGGCIUcw8fhdk0U89T
fEpqmOjzxS7piA+vKNg0mPKX46VqNRs/dih2dH42awsVAcReJYVexAphUwpzfrLhQKdT3oJ2ueZl
9iY8Dw2BnoO1HmThf1+6rulFAme8HMx5GP/zIFip6YzB+u94jgvdfKBGfdAiWvM87ay4srEqoJDE
WzMPCRTJkq0RYYlwfz/8ufmrJNik0kuqxKE3+uDLsPptLRusV07CkLWf0u3PvuwvKNQmt2NsNslU
B98AN5tr45bf+TAI23oz0PoIL55KhfKd3YZvAbzi96Sd7iWZ7DHl4k9t4VKuBT5PIMADfENdOQ98
Ic9NiMNXGWc1rcc7X98stAhxXFxd7YYL6saHr2eKyhgKaWYf9v8eR/qPFhde6AQVFZzZkm/NKj+F
3goCE0lnnUx74AFc0N6+GkhNHo//bQet54EDU6kaFCOOg38RXHSoXEaMmG5BKEdpv16OA3MNPDZ4
RzchrL/7vjRB07y+hS0JAUdrl2y9xNHv0/SZ1Yj4y5ZZ6tDt3Rtl5Zv42Czp/vrXVbeq3H42TW0A
51EtaMLYGzsoGC8CFa19gXqEtBuZWMt/T9MP5r33DmTYcv52HaPjYGUeV4vm0pHURLGYBbAsM5po
MEA8FEkVLOVeBZIys+eK3BElD90GHTfWiPPAz7/TfWAH+7Te1+d6yFHxdOmTEk8PTB9ZIyPrgoPR
seVP1PLG3MbHuXAFmo7I91qw9jFIGy6OGTt3Kks93FMn8ncpOcpeNWN4chGRE5M++gZsnzMtGL+9
aDgzulCQQbkQfchXErPeRPrqSFOOYibB2uQDYgkhsF8o0gF8SpMI7i+XoWmQKMPEZOCNE1gnpUpa
AOwAnfpANvYnVlnNt4Vln8s5MwvC5dDQ772UMLfMGQQoMoxHbgMwoPuHeNMxrh3ZQTaDZt2S4Op4
hN4kdrQ9UXcE6wfBIZzdlgzBedRs0CvOQBrbPFjTp13Be3lTw6hO6qS7USJBVdbnr6fBElEfcRD3
MWkNXEfiKSHMR6oDs2UbeyNXGY6DQ6AUWpVfLuO7cu5pB7FPECHN+Vrjwoi0rEaGQlgmOdyQVUoV
Kq07CMKvrFqE2FGQ0cErI8ti0tqKc5PlJXuKwZedyOPxnbq/cYIwggZTyzrWOENuk1dsqUJnFjzt
r1NnYhJLMJtTFfrgwWYeop39pmZ5SgKVM0D28YoNDDFRfWCfmyZ8MchXG4RWV7uQFTCshWYDXu5d
ZPkgn2tL3Y4sizjGuhsD2Odi4PJlYDTRMSybEtTgHNb3p4dHf2/cfW5qbXEHAWVRuF9vxA/lmB5E
72RgxaXAJC+uCpOuRYX3LYKFFnhB0nboxEoBVAe0ZNYDj79lApK5JZ3tCtSVBbosz8ETFUZFmnEv
MgaQkAk/IU9RTl9UxZHPlnXRxzeoQGlVUqWjCSZkb05vrdoLPChGc7Oq5HRwLFxwCGRRETebcxxx
65quW4TRnxNTuz4rllKHOiqA2Yogcwe6eH9caViGVMNt6qvpnaUuleqfZy3qDe9p9egmnxK43Kbj
IzcFHdqqHPmYIDkmE7Gz9ZRdHW793mwR29twfjIGR1Ccb922d2iXdK9iJg6hIaaqomW34IJtF6E7
FBqbDD1KWpkdEgyqPSljH0N/2n+YFnT1BPxtQGtAy6vg93N29cxHAoSOcIDhLRj2kejPCNhhk9k2
4To1td6fHat91UebDR/SCJA3YJ9X/QEaFuuE9ZSqno4FAuG5rPya713PkaCabR1Bvpcpl4QWI7Cy
hlfQP8e9vM3ReZxO1ZzlZCAjzyUhq0O8kJdjAaVfnHBATms2Ud4SPJ9bYsDQkgSYTR9EC9kJmE2p
DQmovdk3BGii+3wBRv3XEFdlPmOV5/4noupJspG34Mo60ASh8GLvHTHcnQF3V+jM9vo8xSkv79U7
4MW3dYBn7Y5Ia68qH0vZRxk3DUfeSDMm+BVgtaQ0oiF2wgIXrsYCZs3YE/LL7UDk4FJ0Ry7Wt/Wh
n7b025Xf3+hrhjkwhrBMVJisoL3fyBBjzVM4sKJcxuuOdwhRSHM2zlPucrcAord5qjty5/WGzuWc
0cumj3fL8gBe23Qg2hALXyPSOTR5/7+gja4lTTK8R2SGg82fyaUgjNecSPgT50+OfUyoPMurMXl1
9UCs15BZcTxqBrbCWZESkx05Q+57hQKM3FfACUNLuO7Ku2aNaNkoFLnAMebaEXLSx3UEgFtPhAf5
/wvIQJhYwmx6hAsj9WMF2srK2WZyE2Dwg8GQpWrnd1vnNDN7AzM6G0zDaM/J2Apw3oHl+cmfUSkg
/AqnnjqXibRm1q+wsNeMfADL2p9XQTG27aJt7FYlDpBlw4yvjX3C+O8Vo580b6rQpnORB/7N8y8F
bYy1nL+E1Lg/o1dnMKCq3pYU6GWo12N5Ejcw2/mGV6jpf1oDmQpL6rXIUgnpg7HYPFpIsDhbkfeW
YMHGi7nXXkf8RiL7PiUIQVCQBg834biQKzAvj8oui3uGrDykQZTk+jcISMj87ff9DXuxtnJaXz8s
5ZFHUNbEtUOfy7GxpPOOwCwJGLjOsHFI3H4Mt4BOAFCzefiOr9pSHWuV8oCuUtL/nluOBZQd/Mr2
Y4Sd/+Zs/Tqf1PR2Rw+BemkVMFQSNCt9CujOIn1sdzWv4j19EIWID2sIN9w5GQ5yiN5KnnMMb4qN
Hd/PAUnwpgndBTN2iWSHjkBwGE9S7fbUHY2VWX1WKqNqtg4uqgjsKl09pc9UvTYn/MC+F7pZY5aF
oZ1lPDp9WwP+Xffb75eg2fZJqovCt5iY9VJNVp1BvJ6E7cytZ+1RU4kdWoOMbbZH2vsSmwXYyHbI
YdZm9RL6uuXmM3gi1YzbnICWLaRQG0ZhZOHbwSoXs6UvTo8i2SBtFMOAN8BUzYIZaA+Y8cO2+avB
LkAaXsRmp7ivN1dNba5Yz8LYD6vQ1qlZif8mfvbAOavfZ4U92c4OHmOL+qUV9hcPdJhiGYwTbW28
becJGJ1ZVqUY/7eO6fnYbBuR+2ks8Cs9eBO4csOf6VnN+Z6fHIQu+S+rjVPVnbz4xXRVCnRKaGRH
xW8WIkvPkqltSgxZwJiVvcTMLBqxVFBgGwzykFdFT9hRautaH4UYKkdw9A6847kISACYp3U5ME4A
CvkDZe7qArUgOnzBfa0cap8MR6ZVRkzS0ATKPX0oo1CmZvS90AbFvFglGBtIZ2H+9297po/qq4DR
SsTAr9uNti7NFiZwQQJvXLVvAMDVmrNIXcl5RFtMXfStyHUbN9FkMXBsAmo0ptEO7tM7PkKcrSP+
i6nh3d2U/HWPZnfay/VT6gROEFBcoWDEIKFHPFak5OtwCAZ7TBzlMrhdO7UlXnvRlf4YZFTgGubJ
DukZT0whis6YLuIq2S4pOn4hlKBcv3PhJQNVAFPAy3iNWCc5jywTaUae98Ivfnn026sBassua2DB
oM32maw2QSNzUyci35fUCmpkCnNX2fF0XbZocYycN7iJwIM3SdtRmpHoXFWarBGSYBztVJn6jxDQ
Y7bauXW9JGotOHZNTlublsP4yC4wV3F+SZyWyp5MMIHQ4aAKHN6M3HRpVsNsHb7Qx1QF6u5K3dRH
ECnJHIdebpsdX0WVDCQsAyRHOhPhqHfWmt7goi1MoNIV0n9JbrrGxmzG5QknlQRQPO6krKwS202b
vhtH62RY2j40eLaI27CVLgcUCElvnVFORya0YkRWjdqgQxdHP3rxpZ61hX7hWZCs/yGdY5j4gsE+
ucNiCSLwo4tgkdU1s9H5CjS7SL/2PECLh66mKiqiRoIZSR6mGwvw8yIIFiKjjwfSdd5jba/bkXTn
qm3qJPOeUjF+WDCwdxIC2ByLZ9YKEGAG0zFZ4YdvoC2vxK+pppxkLp41zW3N8YO1U+YJovdczmuV
3yVLsvc8wxrHGpQwXlu6Ug/fJp99ajtRzA4fBIEXxluq8Z62CnrZg2z/gY4hRlXk9d7I+kB/xdtI
uT8gZB6ybqzFrO1MYlT//tE023lWl/YC+fbPMLdxv97dP7dfbPFe8fBXEAYeZMkycuE9eRhZUSlX
MxldPx5BExe6Hyq+nMWtjEwj86prfZsY5FvIaGCEnGpT9Ehs52q1XH2Xuerd/AEWhkxhGgM7JBEd
27iI/5Hi+96wKF+200LyAP7wh/R2nnAvxSsggcpUAxufZdjHYdWH4gS0YxHtztOLays/pN8Kt8ro
wvrvgn5Oh2GuglN4K+0AFSKtWk/JzyA7gXkl5YxE47YQrDCP5WxnNwl11Z7InkoH1SeU4llVRWNY
YpV/t8auyXGL8c+iTgDWRyokGIfF3dfrKqpOXAs7P1cOKixGjQz56HbIM4jlropzEBJSlDYoQdjj
9wzxZ4qUFS+9WRU2YCn/X9mqW/b54sRGnx8DBzMBnPGCJFk13iN4mlJdGjGZmOMrWm3dTSZg0BX1
feS2WTMlZY465fQ1O3VptSgZhYhhVSwf3PPVh0Rmt900OX+WP9bIOADPT/118s4w2Nf+eIS6azXl
UVFqGMmvOogn8Y6pgT6qgKCDCbV10NZi5+yDPSS4DgB61M1bTYg3cOuYzpT3Xjn+PXG5n890LkNc
d5l/+KIUv8OStd/RZXshPFLbsXzyNc4JOqdySJadeFX690gOqCre3wPobp/kRNGc689M3WxapPrf
2jeKMmvn8O/kHSVK3jniy/PAjSksez7llzEj0kkhN2sQZ/tyrE2YQL7YYK+jBMYqRy5hQP33dcLt
24c+Ipdt07yMXytBaY+dFyP76MAvq1FR420ipobG09TBYyJyKSlBFz3lU0IB1q2rrusoxW04vmr8
hh5f9SxJGw5JfJCLL25gtlIb6DgKUm9cQMa2Ty8RGDHSHgYpQIZc6xf19+3RaFCfa8i/1VYGC5cV
xb2QQOLQzo91xWl2VHxUCLjwQE/cmimPNXlNXxAEg4o6F1g2BKLOJeS7JEsad3P7q3GS6+Mi7SQk
ItFs4FVjwifl9u2xcuW/nsT7yA6RisbLVbC4puSdcOyOy5glpeQh9m54dy1180BJHanGbfWkO5L7
ptNJ3XFkHcp7fXiGyiYClkFqVg8gqMONW19WEwMNY+lsLG5AdTZ06RJyF8vJVTThQhy/ILpi3d5i
S+Vp8gf1tUrKAdWV0uvTLBnUKkunqtQNb/L+xdV0lvM2G0n7ZNQ+wN/m0jB8Y+Q6AxfuJp1IqTWJ
auszoELaFSOUGSGf9yGNu23X7PU9O0PuPE8rUNKs313l8vNt0aZsK7aQBemNmSIS8sAD8LqvHalX
ukW0ERv38Gt3z6QBOY9CDf5D2sbgs8Z6mi8xv2/DzID93lel5y/arLWMeZsYVdP0U0TDI1SBN87j
ztDuZwdpgWKP0Y1vxy5z5ZP/Exscxv2HZ2eWo/ZTT/wNrzKmHISBAGL46QQIVObZGsaSxZtpA4gR
aU/cRLy7Z4ez97hP7//67zZ+DZUst7GuKS7b9Xai55UFzeHWE5vpRSjt5sSMWZB89IRUdYiudICs
bqaw1FYOaDH7Q4XtMfsDQLua6xGnZBhzF9VnZvxrTJtZRRPPyEKI4Mo4Cvgo3HbIPUFCCpoypCeT
xppCoqIsef8G9YlT6Yc/vzYO7dp/+7xrUzrQajdO5AL7DtOv1kGQ4+H1vfOlce4z57HqkAGF70u1
TKPlJner9ndUPcXUIqF1vK1XborRJlDAMw2gBpTaHw2LOUTqeGh4oYdRcJUiOvC9L1PcXjkJm0JD
7Ns9l42WlU4Mf+MHI/57LnaGh6GDaeiDwLDDSM/xc17+kPTjLDKz0W4iX6EyRi1KrD9QFtEz9oiv
fqO1DkK/9bJFPQfZfdq5r9uz5bWOE5ezvEHllMPSB866ibUWwLn96iCAAxXsrNuwg782SJoi++z4
r7Z9KVPt2qw9lbWFmKZZjOHUJHzlV3wgiAd984C1S6n2iucixLN9oNhInF6uz/O8+X8XY0u8d8Wy
LjPfonS0p9xXYn5NvQ1ITJbJHVpM7w9l1SKXfkpR7WSyfTe8LgZFOPqn0P9gNBtpGyP4kpVzuMww
8xS/jAvzPVNnkOTnP4iOeX/PtslGccucdm86UvdDqBFL8p/fZmkElYuypvD78VvLziMfrpg7nxcf
Ngn6fbbNlD8Mw20Jj2VoYMAgX3+NTwNGM+FIqdieDkN5l2pr80713vMNSBdhjBES05N4RMgoQtN1
kDQ6TLN5+eKz4yGsd+ohYBvCksMqMmi4vA1CGOePz68xs0I0a3rfjZBhjAbIsjV5LpsjdhyQxAU5
uJBOYU3F7TeAcZ/NQ1unOinJOKMGw85b6xQvV7PIey1FjpRWrZ6/nsZXWup+g2NnsfMKPBgJ76MF
61y2Jh1eU+UbcdnF5VyenKJT+GUUidFvU1sTAf1Ejbpa4Lo2BBHx/tIsC3Xe6zhN6j0rbtxLv6Ot
ZQ/hvaAZmt0iBbXBObWq47Ox9SM3J1RTE8MohPKYb/CWY2Bh7PDs+TYmAf9hVQcT8+nTUsyHNNjA
BmQ7KqAJHQ0YyxMiPTrEo+8MRjFAos5ihAV8mMZe2uVuJUgeHyv6dWfQfZgNc+LhDyfr8HXB5IU8
glj+ThDJ+lBhXeIu2AFHaN5GES5Gj+GTZ4aQfFonWv4iJDoXgOBxGoMKSZKbMgrJY27vP8/Cc2PY
TQRWlIRht0t0XD24OHu0suVWOX8ZI6YOTQ3iGf1NqwubbeRxW1Xd+ptGW0YfI14nIYyP+X/jBNDD
S6Z1/Z2wVz2SZLZKNwE4beOVnH6COlGYmSS0DKWHLG8rC/ythEFC67lJubDteWg6h1kUc7OHKBg0
MSnfrt5nf9gEo2OjEAvygwBmdhW2+6uGeFx4pZD7c+dEmtOv1ZPhv+wIDwLANEA02G2OE8/ZflvQ
WNj3dEUBR5bC/9VJnKT5tC8moS/2cPGYmnIsPSfdV3mGTlwA78syRBHB435CgorADx3wwBqmXn00
zA86Ubz2jWn+5br8AF+L0iqcCDPtb+H/IluN5qhhDUe8ufsyK/sxLVAQ/QsZ8glJPMifoIFXUmLn
LYcwMT6Ga2qTGBl9CcB3l24VssWnUaxoA9jR7j3SRhxN4F0F96yW8pxgG3pxFJPlAgWqoQ8T1e8p
/Tn91KVjQJ8RIg6qA2cstZO5WM+bFzqQ7GM96MHGQJGaKERnaUGZhV3XoBZBTUIJEgcxps8TN+7x
mxYB84tgcqG5Z/VW3PzYOFapH8v9yoMplGcmFnBc4+3PtcM20kKdoKdZPQEQH6O+3DfYIDLD/28P
T9e47DxCdHMLcKSxrJS5ezTolxWGaFyGPbAoiPX2rjQ0KlnQlTy2PiH77rUE2NbIh/7hyStrmkDQ
ZkjTUhY4l5/Zs3pDqSATbTFIBvVV59Taibr6A+Lt4/hKaFGN2o3d8jUKalvZ21X8kYaG4pzk7jnN
89YGeHX6V7c7GTX9htzQvfHhCEpdzQouKMhIMhc94yDgZmt1/So+tm5hIpXOWb6N9Qs8Xk6esCJh
ka4dWtzvDWyfokqo62lXVH+7XTvxHfeuCZf855uJ0cS8ORmtWnjOMGInQU6s/nSWVyikK/H3ywnF
6SkI28esydFKRGFY7gg3neMufrEuaby3HCKR/RwA3n0kA650ss0xHNHEeM7xU3+y8fq5M3eIN4Es
08mq+MsTdaot35ZjhIJpU1ijs1GbHPWS9h7aPo1iTYrVrq3C9EUxn+si/TzLEW5j44eTGSYfu/BI
5tlsARpglFcQ4ryYQ66JRcOKjvhk5XG++1nqxcJVHGpAAo40i0MBPu+8RDMMdo25jIXhyq4L60kc
uNGlqTQqUfmz0DUOWguVEuxksMlLqM0Kr3Z0a2PaLkxv2xiilMeTwXobRE35N+IxEIw3zrhuLP/f
9yemKUdUVOHlTisZcrX2bmtfDLaPmvXtk8tQZolW96JsvOYMHFRY4zHjjxfJ9JMEhxdnnY35W/We
C/Ar8c7Pz/lCHWkQRor6JiTYM8M/RNiMyruClj8D0Q0M1YASgFqri4MG+TaS/X4qarlFkl3JVM0S
icbCrcWnnWwtup1WnoCiLDRotdoaUvIu2EcCo3tYqwq0xQYvqtIAGhacCzbCTlfC7AULb5dsM7fB
1cgQMLrRpN+VmVOhbSqmb9Wn8UIE7FMsjf7UogUx0BCW0M6+n3GsfOnUZHrqkieQhBaSoXsgBmeB
f4at3aoltL77NurLqrI5r+deQY7tt59+VSrG/+KDtChpLI+QHC340ZgGMNN8FbmnuECEk4vlFuMG
gW0EmnGp+pY86fX1SfUqW7uhLyw1/OjowSwO3F3yP++E/bNC2Oi778/ikLnfuCyfId5HjvBf+7tz
VIeI4zaRoJsF+yppSGLII02TDGC2VosZCQQW1nnqLF1Ka6LC1ROZf2388o312QQZSnpS8WpejJa+
lun/bY05MOIciYsvBRWpIrnDClXsU5CiqTSmGZuEjIcZ9vWh15STlCWQqvwD+ZGUl3pq/0DCsJ4v
jK//C3UfeLEv0e0qeS3e90ySnoweoRcgLN12jYHa8fhIVzsXYHydNoX8vqxkA8mJqEJbaxOjy0mg
H2EhK+wX77W0xLHoPB4ns7ZGSZbxVtm+EKaPKUwBTyZ2gOXDlo7wtvRsFtbbZhNwdORIsv7d/7L0
GhrStU+NkfcKSQNVKGKcf9FwElCF4owR7RYqcZ0Bn7ABGix3NQvCr9AdHqKaF4sUfPP1CtGPSIMq
HVpY1fQs0P6BUG5fcxsSv/oiZjVsoJOBpKLKAMH0YmSM6FLQZe8gtCXA2ADfr1WdBiMYA/xebORI
utU94hMgMVbMiCC887TjQShch7fkXhsMwKEZSDXfbLubNasZYvmlV3iIXidRItgzFOaxHH3FAA97
dqs0nSXdqVC+bWSHKZmJMSCDLlhoc8CVtzuhNkKcU0FHdNnsczuYIz33u4EJRtC9jL9BnraMrjdg
QBf3O/30gLzWXAoeH6UKvtlgfc8xq80aSDp330QDei7Nf9bsPm/jnD4zKUF4061wWozowAePN/cM
S9KrsnQxjPQjaNfBqu2rSodwG2oDUFbJPL3OeN47XrFNZrFM42+SFw68OpVIM0rWIzh3dbaXYFGt
wHQeT5EbBAfQQpMjh9jhilu9aaxwlsHVYltfLfLi61AvNcvP5BNbh9P8rqxPBODpml25hoPU/98K
mHTqvuaeBpoc8W9/641ftgB8Lk8P43gKXjESugk1rt1id19Ktz3cG1taMoZwg0qxxMfXNwb06SB0
LFi2JcVDM9mHZQbRCCMjAFrTwBBQlT3k4EuoU488mCgfX0ZmGz6cDaqPmcnSqiCd+jQOX58TDy88
d5EwzNH0he8GFgVKeYQNs1FzS8FfkFptaFDe51SOTNyBkiaxjfoeexv6r42OyIkLYwmZS7tJkbZs
9M0yK+nommxnlFw38aavh/U1ERKwVWLzmjehbSAT6AJqxeqPmWny8cg6cSXWD8ASfSh0qYyaFN3D
1LlXjr8QpMbIdk1+kGrU3868zc4fTT9zx15jh/8wh6tunqLpJv8ifwIq7yqiHltcZaD1mmfg3jl4
rAB2t0BveaifHDlYxp5TqFo22YA/JSBYrIw98Xb+MPMHo32HIwPtan65k4eSd985ZR0cs6HHeR0e
keYjxdgtRA3Txn6OyV1EEe2PYO021RUF83k7qgZxbaOs6qCOxXzSJz0GPrexWmyC1Qres1XsIqg6
0g5Rf8ce82XOcrepu3YaRu/J4vQq3ZWE1EMlHSzQAe9DgTLNFQ8MqHp8G9rhf34TEeTQFGquuM9I
b7/ioQV6FCTVUm7O592WLmLoTxXaOgt/FVxx8a0tut1u2XE52bpiFcbEMEkD/oGbuOehVXlnZS8X
7AQ+WpUt7rHy96s8arxwW8ugbQ6MJ2NvyV5yqSm8v7Vxka6gtF9nOzCRx79jQ5O5ciUOCXr4Lp25
ZtoKDJqRW9jEeu/RKJfwbf/oVkebgzllr44qwoFzzA3biC7sUYd+kK1kanpK+42i66s8VTeTaNnj
eT4MGlvx/PWlJiY87E0OOKnkfFX7jiyBkNYBzd08hymN4HyaGsRrHIoyLCexdyMWjNodSQboKGXa
wRNDd5o5BFbHTRbMaspX3GJv1cnFJnLX5y3SmIUivpnjEOcncOiYc4dPIwbeOZ3xWlvUu9jRffgV
138QvWvmN4ULsvh+9BjrytejPVQDd4auY5KKKQmY2S5LvRflT2k0g1usCcg2tSKYZ1M+GN2ZQH0D
zzfRLPTeBTISTXxWJSajfBCTaUI0RLdTo4tsb/ZtQSchmXUc8itXTPCr5TrTk2R9HVyJBgHF+f87
bBPPgB0pdk78pnozNAfPJy+cF9n58Svt2mRXX/JBai88rzv1BUtzeCfxLhKxpHPzapCBfFkBqipU
OeWEb0goR86sPqkZ8vpA0aCXP8Um7BZiirG5bm//GJEVDkRoSiElzSgyCGpmS3Qqj22mp9LRXtAk
AwbN2Kf4Ne0R48KSEoGSx0LDk+1Y4kDIwK/OI/nJjWRHME+POJLI1s9/QPZ9e2xx3EsF3ldjqGKi
Rrzx8q7q/Ohwf06KbYx+dhUJALI1kR6uR3Pdkl5rmizl6t6G9I2/DfOSko6aGWllozCyWEoPaSSl
L0CBUxCgMWL5uyuSFJ3OmAQmmx94GlWRUORL0D/acu5Zip1oCtNux3+cmj3tT4up+CjCaUEvUzIg
Lbw7M+EB/Gh7wZgKABTu5NCt5JvLwfwSPr99MU9dtSNzZy9s3oAxldseVQ4tw0bQ5JsNIDlJqSqX
P6Vak36lL7Sixe55VXAYrS60UgmcPnQ0fjXL4RaI3jJuQS7xa6XFKlk1tDRhTfnc6175Tsoj29Bf
kB7LNXKRk4sFlEoJlDImZu7I/+PWebchGQgbieHC93kDufpm8f52ye3U4/sLP7mqCD58Z8L+rcWn
1y1BOg31ZLEempPUiTMltYFMcFGgqqTgb4kQLWN03hRVuZr+Zfz930KdTJ0jLQnfgRfBfwBKZ8ow
Z/A2lnvS8UGgcmxNaX9ll4F/7ktH3DW4QYquwTJx0MBSG0LdrfX8hI2YyH405uXAbmRnoja5/+S+
4YZuKjXgWwj+4FLOuBSUbi5F4KItGxSbX1j5OdKQiAnj0tfQNOdGsLBCClg6LJzPruCCHxnQ9fhq
2Obl4eog4dschqNYdMPahs+dwL7TYYmDUKhYCmTy+iVWt3kpld5L3BOxnKoU+VeWLxN5gJNCSOu8
OKyvFvf4wpQ277wRCulVbI4lJLtc0KlJnR2e2+7L6eB8+ep+gwWzxttxl26pr5eakMH+WYXrVT82
MLK/bsuTjyXWn9K9POtCm422huxrCmuY5Zkj3zSVUrLA7GXSIJBJRjclympUsdMcpA2BecBruiCS
8Xt8j7UNCwV+mttWBs2TfkbNc8sALunFgYqrVnwPgt0ea0KRVJkp5a0FkGJ8fAE9A4L49Uf8EzQF
HoicKT4WBRNtohAeMoSXZZso/eHe+o2x3P/PoVoUxwfUP8NTC15U0p6zowctLRM5znIVQTqPfZsI
V+wChmtGxY14O5ls7WSXJhPZS0qmQXaH9fqhW8f/9ucoHj+LJWDI0YBF8wL/Zk1u2ZqdfL/h//ee
ClaoVNw2iE2ikGfbH3CELOuGoj6jrKrysY5TKzVVqjaZ6iEI4o/br3ZXyoROCeBQMexGN3QXvYfW
PIiKDBhVMmy46U0yi/2IEMFmI1ATrQvWP//zI7Lk6FHj18jN7wXr70er2MmHNAXHfgV9cnHSQiRd
w+c+IXrzBWXt8h4lhwFvg9wQj09iMvhXifAJtIz1L4eWDmYuhMIMkOHs7e95lJ3XjFB9w1VsIYSh
Oj2Dn9CtCyQUanhxsUCRlkMnnqANH0ft0MCLHLZ1H8bhsS9W9HiVP0eKNSJHzkMgvULi1bI4Jc6S
IpY5NDfBAp57/XmA7QuimrgL4jCjd9oQncY2uIlf3NGj9xr3HiwKV2Fo5YWuHQniG5fgrusIEZ+5
ReR8Esde4doqCVjcZxXzHHRkgzD16NhaSMkrGOz44JyQWsayJriOtLqTm7hcidyR0zYvhz13fvpL
ouYuJqQnKDDu1aAFv4mIB3v4U1d2Rzx5vAtdqufMtlrksJrTN9lOL1iEWyR/h1KL7AGFUUUjUHR6
xuYk2TzZhxH6rhFIv48VCmeGKpr1c207kdjPbizsbaEYJQJMpj4SGONgtDt5s2Emy7oR1xpBaUNO
7P3G7x2ofo6Z3AmHsGYXmCjH1DaO/IpQPG3Yzb6ZJ+K44pZNnQ8VmlVXs4lV5PXL7ngwcnCSWqmZ
MN5Yq1E9sKuHpKxlPbQZM0vfG1lkqURG6//kfb4op0KWl2H0BJcV9vxvFNP65yO0yUUxvEBGmBpq
lV9AYA6b/wqvrg/eAiLWgWOX/eIzMO8HNmrt/O9CyG4GNb+SRDmEUj2DW7ltEI6kRZod5NL9hbdO
Y5x09mWtj6kMB3zVVvxxnBWdjBfHKkjlNNxgdp3M0lrUI/zBlyG6KViFVYNlBXqgx4ThrMwHsvO3
q1kgh5tk+NgGzgBnWT1G5Quag9at1GH7uCSsp1J68r/YkDPWgs8CKPplHWFUq6RE6w9MvYtOzeYJ
hsQIn/cbd2MI7WPXJewWK1O54QOqs4hyCKwl57IVtz1bFyfq5OZVQ1y+91uErcVScmZ48Y9dOdnk
hCzMATLVGANJCfwfkBubGDXLo6UVa+IYguIMOA6VMldiV1+ABqlbPniI+r7kmukQ1t1Cg+LzxI01
J6S2PfmkKjlNU+7r3T/1hx1kSnwGfaI1YKMdqRSjKUn+BxE6OF9Z4uEn1jTdWlURpWmssdyz6I3K
n2N9PyR/F3WQOq3Ui3Pe1OTugx9JXREsSsUNk7AKARDongl8Oa4Nopq6MSwCoLfEi6YEW0vVgVyf
j3yPfP9VPukpiwSNKg9boOs7sI81J4gsLJWNW/kGqfqxLMHIFTDuTMUYM1yPyBViJPjjpXwtSmhN
o0RhtBd1zowhdIIqa3mIrRIItKW47+yen9gYJgecL1Sf09nLZr3KKce4LWo7EHHr6IuYdeWZcby2
/QaD8s7CJx9mk2tT0fx+1TLYn24fHh4K7oNrH3xREzV8zCaOwwhFj7t3eCSbO406/GRc9wY2Rv8h
qBt4gmwufV+CalcX84M/LIO/17s+Zct+0yJdbKmXiwJrDBEBrRgsZfH6KcY++T2J/xFpz7d8ntN6
wzOBuw5EjH84kQShr8nZy7pELGFELOMNXVUAI7h8Yyr/DqN0lVtnDtzgGG+09VoZoJUVXYAVh6p3
NMKqLw4jxdwFJ1r+eXKMnisE8cSXxUUYC92TNXFXPPPS2QSVl5TYZVm8rF73q8ROw9MrFYpci9xL
zgIoTjOKaopJirWiBpRoTEwRQ8GG7V48n5RM59R4FPXUgHsfpZPq7Xr2E96+joxYL5zwggYZwyit
F2l4N2x4TUUAbtXJBQsf7Dx+TE22KRcRcJ8DL85+ZDGz8iPwUefiF22H0Zry0CD0DUZQcWS9MTOe
TZTp1j5P6MrGsBd8RAqWG4Jh15HljyhAn0uA0xP7DfhcHgUZ+BsMEBwSJVPpQZaEkbaajK/9ignP
ANJN0goShIcODajoYtyniAVRCVKkFg+fpn3owuI3j6wIHMSxqaiarjS6n0cgOV9vQ5QXgMDtljkd
Ynd4WZfQITQCmSsSSGarpKKHkWg6dYV6ihig8i7g5IRg/dH+Ll69bUUFaFVgpa/NB2Db6I7wFryo
1XFLrPlmkn2QlS0K8n/qW3CbNFnZfJl+cJEtvDm/zPwu4CJWTaddzjVYgJ9c18kJqUHwqFZ9stM9
fRCqV2jMVlGuOioUg6xH2Bnv8dxIMYYed47VeEknKkZn2+PqbhU1juxRY9PmPeEvv+ahzdd6EpDV
aTj2GOiA/yfB7CnH/BAJwb07/fxjmN5TmK3y7Rnh08jTVP3zO5bg0cvCBYo2qTDGerCmhZ78/hTQ
rnAzQAEHA4q3RmSCtjGdmIO5YaqB5Bd9XOon45y3RfLdtcjaJ7xurbMZYD4h9t+gQdMKvfO90qlw
TjDkDWLNtZKoNZGT/TrHQSdx6RguRDmKk6/lQA/+h1nKVYYmDT59fuHjOir5GAsBFcKlW7Fr3fK0
docr7hWxDfVRv/rNTVL6kRrB5lDu7H19iZpb8mqz1CT0/k9eAdSt8wGsvGM0uAlnDB0iJSVzywj7
K2w8VPnXrM+pxaqPvZ8r3sPO7AJb7IvW2ZEuVUCvZwwPagt3jL4y4OQXtGtBMNCCP8bbc/BJUnzw
D8GKbCqCp3pcmJiTIA7SC2gvOECRz72De921FME2XNkafPKgSBTbbTUTdp6SNMmxHPn2FYC0EtVO
TDSgkP3B1fpFi4yL4wVA4sEd3L/uV5V/Ruekc34gIHQg99/xFyARMOFgyn+41vCKN4qddINUgNwC
Q/1eltOxbvSvsh1MenfOc9RftX0j04ROOhe/Kdv2ye6j4LbD8aa9t1H4/p2huT/LyCq/HYcsAxvL
3efxAFGRdQ7dRQFHj5FXjjeeKllWrnuQa8zqeC4nJa7pCUp0XIefNJTUaWzustP44/SDjb7ybM6p
vNbvOJJFyjqAdAGHzSSQ4mwLd8LcLHVgyxReGJiIKhXAWcQNpLS9amkEQmmJf7jDWYAyxOuvFtLK
GnJUx16D8RgljI15lgtUOfHaYkxpuLk5EgEvzSxnIBVHbHkaziqGrEPwo8PKQxXpAR/lCTRmH4Tu
cyKmVOgdxShkrESQSkDAj9r5BpS6Q801Pg9h0oS2TmlPr3qQ/Y4m4UZ4MWSUmTPhFnxbR8JF9eX1
jBefgJbmjGV1B4Sy88TrtuecKeYaMf9YHdOBrHlH4B0vFhAGN3slvYmiE99Fod0w0+hJ/bPbYzTz
BFqNfWAhXbVbiQHvl/Vs3JJJWahjgIAj2l9HR1n1zYbXucDnD/WBPtBYcj/VR+OBBqmTqBFW53p+
0Abddd3iRm/jqhvKj1RVnvPn9hPf/LK7rzWW4B2IpEu701WB/8V3Uy5/2pfOdt6czMwHOuaKooy8
4LvX9l6nKrfKIkncoKosjaKxrzYmaudh8lSsQeED0pgYGuAmey+7Omh4gCOZWt3whlAHahkWvp1X
MKJhkUvNSqTAZwaR2bJzkJ3XDGKjTRdewkEZ/fJNQlArxYrKbryTiPx+a/sstp2ZsRDmr/4yvvlr
DLMIs/UkT1p9zuBHCBUFTTwRA4XBurMSgZNfXxGshMlJZBxSKcAHBfIM7mQOWqDgTxQNAjHPGOil
bguz8YhQJYxnCmE4T6R0lSAZk/sNogCAHV69LIDmweIU9f84YrACOalk5Q3B6N/sxRDitaoD8cbe
R+/dSPKH0MUdK4PHOWwtn7dcVN/X2VX89hT5wDwIlNAOGka2HJZUQkdceBDfWKkRgzImbgynRWIt
pQfsp4BdWKI3eL+wtPTkc49Rx0gSaUJuIIhgTj+Tv2MfoslLb9dNWKgR9EzuQTYpxihZV4Bg7M6d
kjj3Y1MBIjYki/SXG8Alu3JOdWStPA0NZyC8BZTWcx47YpQVPS/HuJqFSo+0ZqhoCWMyTq9DeWSE
VMtQLGGMHAAvK8JVYzL+891MCmZs9U+y3wHzv79J9Uzo2FwCPDVOYAjZTjRCXRK/xylpvzAFm50k
s75uj8e0UhQYQuRJmrvpNUkoATihoe5SVX+Ad5/T7C5aiE1M5rqcgddgSo8UXquXuCAX9p8/MUn/
TD3CZUQUeaKGiRn1pqm8X20YeK9a1L3AibIIkqrx4lIUgaop1YmGsqLEaZIZhi//AMmI0Xcdmm/B
XPF7P5WBwu3nwYC28nnChQdUgcC9WzndfKP856YiNKnf2JIKgi4F7qbXBjG/UJcy+w1IZ/ZKYBoj
FOw60GxBnEZvUXhiXywKpamJqzG/G3ZtI4T3RjKOik2m9e0QwCcLh96Czye416W2XtDHWHFBODTW
cztQoqo0LPHjo00IY/BP2EBaqI8sPAPGBt818m9uIrWsXHmhQJftuWfJU+9WKbp+CD2haF+fQLeU
IyB69Gi0e9ez0FilcauqMOrpJl0x5ggIJi7x90YLOcl8eX5LtdPDdEIOfFSqgEqH4Fx/ht3/Tca2
JTIrxHVJsWSAfuTI8ChVE4OwVMP4HAnm+gwpYDiTdZVunusGeT/0327n2OevTaddqmPh/HXRkKZT
RgQuUJCqzV5xgzaoAS/3xZu2+j3hLsfS03g4XcIUOvFaIWE9Hs1GVPvCnIWnoviMoT6nwAuW2E0S
QuAIFKs8b2e+6TxJESL0ISSe6AQzdRHWEbuW3zAhfyNeAQEyzsxemrd+sfpWfkpxEehO/HaYExNN
lY4cmuS2y2sLbfxuuhW+gCVEa6Ev4B1CYXHEEotSimWyrDsJJEqDZ9oZ+YR1F+oh8qly7VFMog+a
N+aDBXLkSa53LdByncvSQ7c8laLC4jbD6qyTQvL7Skva9eMMAvBljpwpjRMt483JvdI/vFZV8/N2
kwINa6WjKgeI7pjJQdiHIdfhHE8ldR3ITIJ4Dgm58TA9j1W1XjpHGFomnrnyI76K/VTXXlQ38Swv
igP0AVVmOclzs+kzq/cA5gm8WJusbiOAAEQbQZh1U2c52eu/BoNKLZ5BPUARDjsg33AKMYBrLDPW
g/BWtyCzHM0DGgfy5c8xUHRKSru1PvTY8XlH23lcqHQwpIHRIp28Pm88lpBnC+kyam+0w+HxX0i5
zN+T/70QeN8++sU4ym/W8Kp5ChMf6ETNcdajCiWLZzS7eR1tnD6xklULp8MxfjwM+8d4HI08BrJV
UXd7uT/OQfXlXYLrgCBKXSJ7XW6olvNxvEvrLtrKrQ5zVPw76v9wOaNUg32sMqJofLly8Ci3RKTZ
UiuIDiIkb5Ak2b6AdoIc8Z4yFPLzxDfC0sBTnP4XNgIZlhTKakHgSQsQYVxVKs7B+dvWtWwqP8Qq
yYPaIClnAhSDs4YLo6pF+96ACzfcS/oi9xxtlglh8Zh1P09/FVXrw7rW4zlCOgGk0ELi/zlhMtoG
46jnivH6NUegFVAU29j98JrCXeeqN4sFrG2Z+p3c/voHgInetFsVLNvVyygiKKDgCsAS5WDcibmt
nei8/lLhFc6Li7MdU3JCWf+GiZ5J385CoycUNPeJJyf4Sh6qcOA2BcjJKvdtYWU0tsjkqEhfmDDN
Fy0uEZDefAr2wNBRxEy645JhxsYcyUpazFnOI6TNJfB3oT16L5k4Zb2Pha9AGu27ML+SOOhgKief
ymBmVd3zrW9WDi/CL137AQKxiXUo/crjiyhESNfh+qY/xQMwrMRPdJPZ8yRd5VpHgMHK6CV5ddE2
nHXOWiUprOHVNO/lLtjJwnQ6fb7ol9wNSeyWbrW0ci8SPhZu7oZc4DaJS3OKSS7tG9DXfqCjUvT+
gnHOJIhRjw1ZCAQlDjHDpoidDM41Uc6NruP8tPLYrY/kiJUMvZcz9WBl0Vx1j34N6bGx4sHflwZD
V4Zm1+rh5OgKWtbBRJVrSqNqwCvNrBFLL9zWFqrYsOr1c9CwQMgNcSCN0tFEmTIEdvBsAmdsFcJ/
9iBQ+y6QlSF0S6XACRFmTHuh5MxBo07X+UtI45KHe51zeqszuKOq8qy2k6PfKhAcDpEXVVEKH7zj
poS1Lyoh1o50vUYKxNyqUHGc31taWVC+X/0sRm+hJbYjgZ5HYAdRp52MrTFoldVvZgMmejqIYtgo
sWNsd5ALWu690R1pQQ7tf12imMlYJDT9nFskvYtXM2n4MWiGXjIA3Yrf3jM31On5kuBNFx9NF7GI
SUp9Mp1M8FvBUoHv3hWXwCUs0/r5FViaEk0VazQVv4gsf3Y0dEHYCn6We66y/wwASCyFWfUfmllK
JboYPYxyw3zhQf/GwPBxvrh/Rb2HIg+4SS2dfJv0dhvokeTdO1IzLeF3vUMyfwIriMpE5NizDx37
faDqxwd3n4sEg9/Abn+0SCya85+v5UBNB3BFGyKyqEXBuR19T4QutODupySZiuX0K1onfQc8WxUD
QATptM9fuq2eA4jg7pP9D9f0eT9osBp57Ekhwz88CqQXwtOLXeFlVleNpaaxwQlVdFhBlEd28jf0
G9b4hITNNEgzOw6jXOo1Oss9vJEitPIIVZiEvuj7tYYREpfNwfbxll+CuFr1+qvUTdmkX5miF2tA
++uaLoCDT8ZSBSG9iyWbj8bBhohBe6xnchTjWz4AO1lCDOB43RpVrrdhOv4/J5eFZbHsxUENc41z
vwqvmFao/k/pQJTVvcZVn95J469T1FvyHCimxkzMADisk7Z4FRiOjZisX+ENyhXI33Xu3eDq4lBN
bLgFDVQi4Nb46fwiCUJm/kiXHUDD1PEVSOLH2LaTv+NJUnm+3+CxRpD5l8w0l/w5lBGk1tWQdQkf
zP8BB9cn3YhRr3jKm5kVzLB7elc8lPKyZJ6wDy+zHjNPsU/mim5xLOAtx28SNh/kGW987jV1wS58
Iu0GlI0wnls+If/dGdiMP3J1LKFqN1lB79y6QPX97HOw7fiWEx9LbeKkL+AChhPGCtxJf1LT92cW
j/ZK/5C8cKuepI1u0Okul/e9MMCarND6EaW7jZyIUNYa2MmKPtDal/bj19VFZfPk7ZTrsPpHHDW1
7K2u9dyIhQcYYmzjbi3bN5PQ+5tWH09nPuHhT7tt5tK9vGYpKEtSq+WYbZFJuAdky3uzLGB+C+m+
iEseAZTIpIDKqBbW4tPnUu3zqGEB9kkjUhsVTtBfeYjJUltKgQnkzee72GB5oWjRaZwBOa333LpP
9Qc/56Xp+MbSHjmP+Q+Oe4e+PVRB6w6fV4FeIRxEuE/4uz0PALZYTkvZZxziokTOqlq3i9VyznsE
d3X5iF1X1sgTyD1oQ6iVImMtQi2O2YOquQjbNKG9UILV5UjaOrCL+txsMCVjtygAoui404Ns/laJ
+RAaIt+FSvYfTF2DepZTL4ngWaxWWZMup2rhzGNrw9X08SZ1wyhoinsNb1VkFLJo+f8bIkmIfcuw
r9kWTVPh1/BeN1uvg0tswMwRdiiDLMGbB/QwZJVy4A7r5/zsASBMXBOW/l84w4IOzTpv9uqdMtHE
TIpuV9Rh54xj9yUsj2FeIE88hc1F2skHQp4Mk7v89BLxGoCBDl1l87Zuylpq/Ins+CROpHwittDA
9IO65TBRjfPvXQPkBWKXKlvr6bgpLX90pgG2SVPS+6ugGJ1DA5PoQrbx9tRzzIVvrE4o+UI3vdIc
wmeAH5mKiCYDJXWHQkguaRgMAvNa23f1UludXVI51Gql9nB99qvnh2EX7HxXoSpJDY9LX9aCoP1w
XBgMs6S0ykFKdKRz6Tsy0b/A/6ywLwhtlBoll+jB7e5jNKMXWu55LNKJCA8L9/7yQ3yD/fg1CVTe
gwmDxqS5v5MCxac3KQOQO/5NY4DJf/XsgKOpeQCnRoNoRw7hATLBaZy50OqWTdWLqiIN42sW/y3o
nM5IiL2kTu0+wZ41i//aEfA7asYMMDHXJJmCTlsaN1Vz7ZzTPmQUrJF6GW7Lenbm2o0aw9Ff7z1k
+GmCS1UdLswgC9WeQsgbNLGOh/eiUY8bmT3ADrd8/OziolJ/fDqUPUcwAcfwbLuCnxksdiI0KFba
ShBsu26tszKKhK/4HZXwiDrGg4m6LQtthUpMkLm/MeD2FVvuYzQmztHgjWkoQPQ6m0StNaXYPGbf
V88xhJxphyC1V+NKeKkcWnY7kaE81DigxtJmdr8T/wgJs/wISo/vpVddBy6dG17CCNZVvmC48Ree
Iyc1PPZuGFoE28ibKf+/ynkCyLsCdOuRBbxY7c5ja6PQX3m6JBTVS4mnaOx04uNPIX1co0Cil6yE
EmP4Ps59j9zie5OirdMcFYPmrBeeZOcauBBpkpA1aMQxEErVkk/6/C44V9Jq+IiOQxxe9POKBswM
zX5DwLs28pib4BxNhVk9Vt+NuMjVf7lg+l3Uf9gOyprlR6WHrahFW8h76OnH/G+HbElWN2mG3d25
pg8k3E53+3NGsKcUVf4KfEIRJbzjLuasOXTwmpY8Q9VCrtPrNwEcS7yScmC3uMPZh2nTJn4MT7bs
2x4ArgUrtN+maZ13wTP0fNXX3mZb+LN4zuWhfYw5BYodB0iPBVx0L+3RnDaWu+ihFYUGeYhv7JxF
DkBWm7Ew3lwoiGP3O+IGkLQu1stfPD9RwCKjEd0thEhPu8ivgeOIMJ1mq4IU4T0jCoxcZ3oTnnZu
eOGl1Dps8iQGIe2FALPzun8H9c8lVT2UBgJ/uz8nHpfPe0C+0enGbRYlHpObiVJ93ReXlEvjBWMC
ehPbAZV1OwN3FZSU+hN01jZGV35O0QUa5+6DFuqirCICGepxM0l1I37mnm7V0kAz9FkEwqvHEYQ8
PDGPfeLR3RS7iIZH7neYvifkojCDihVUKqqDA0W69/l5cc/+fprEwd4c2X0CCohiz4zU8cqpIYrA
RDjYnHD9rufsv/LMAv9H1lGxPNKQu6enmxTskIwbEPh0Nm04m3ug2bVmnjL4zdxVtchCGHGGsfp5
jlu8fLdQLOjTun4ilXTOl0q757WU3S/sZ2G/ZX1/OtK/xHMqEhrruk5bZA6lPscK2HmQKqw85z6E
mJ0I5X3grHJvtxM/1IpFfyNQz8EIQRk1NcAZuW3IPuFLWQR5wl6pCVGthVmTCFnKuV4z5wCrMZfp
Wi2cDxhNefpxX6v9rPXOFKh4PEt4bI1oMG6NE5HFUGIk9R0vcInlxQpqT7tX9ISs0D3S4hZcUJbL
Ugsm1j28tRYD/cOPLq+YoaeQ6t1sii6et3YLIFkWxIzxzIpqiAooAWmfv0iKRhRrGeQnC43thFOh
+fPcB2AGLmviP59pdG+MkD3pr+5O0HfdlpVefVLT1uo7NnWRvnDyEC0N5NvKv4ucE4dDI847cDFP
fnkYjvrkkA0sbok5u1rIXJn+r0TQYoX+HhCxXn93vG2ZB7CUNBoLiQxpXE05ZfL2R1pN3HWofaLL
bNMQrH97YnfjT1cqJtziPqt4lumlCJWiIJ6RuE+fPbCuontfKikglemNYrwYMDTu5py40O2NruXJ
ppCYbPBz0FzbpmyEyX8ECRSprcBzxql2dtHTu3cY6BySD3WqDJl4soHbPrDkUAC6H887Crlj/gYW
C5E4gMX+vxdNXtqo2toN0KDdtUbsvifYY5j6UICkBDQAZwZv58vzhig6vwbfiWwlvSR+JH2Q0Dpb
cl210VTr5xAuK4SXyXu0pdi7/1nWVvcyS6ymfVjmvHLJSx2KjjcsFLEuCWRmMxxc1mhPzMpT3qLv
0LXf4GyNzW23n7+vexY5M/+9rUT84l4kViGEtgjzzlvOTCNbelBwivz1YYYdpSucZE23Qf583SZn
nhdfq+lDEd+UDZdZGfCxdJnenfAHGHjNfCNWWfhQI4KkRA7CVYkbcbcUmSnbL8zXJGSvPiqECHKr
lYD8XlZYDl/aoK02EQcIR9g+Etgmj1OHNgSII1IA+9p1v8B4K2jzrH5eb3+vawz9DKFoZo9ViRSg
bp1/GRHJErjJBQ91sEB7Qa4qgOCCcmTl6psTdMuLfGdHnZt71GI0XmmaUVA5ieEVqteaCZtB23P8
f0VGujIe5CAYWsJiitJkKgogw3bMsNeD1PB+6Qmf1EhOq8iZOINoWe4I1SbAbaabvDJncrMsJ7tO
iJyl6gX32vobtmC9mcvVCi8+yj8Fb8Br7DNLu3w87e57dEVG6ThYDyu3ZXYHio1e+xTRVH0hZSus
oZTsbRFM+53BIDNM7rvbRhMPkBrMJen5u8twFAICoFIVzkHUMLcz9mrgxxcWOf2z7+MdZQO/NolG
+P5hRAI9G9JoCTC7cClsFnc0Bj5TQEw+heSiP3LZfjC14gM+RHJ5vtQQjaTgTz8hbxXlFhYv8zZY
6wBM++gDHsBTulb94KXKfCFWzFg8+5YrfZGo3pfuzHAe6wRosAmA2AfdW+2r7S2d/+IkAs4dT3zs
+jKbEI5wsxkvc7fhT3QPPMEasWgcOBWdGOWDtGZHXOG9NrQ/AHSRSKe+lgE1S/NolFns6A94/Umu
b4bqlVjX5Sk2K7i3Gb96jokDu6v7Noi9paOJMoMRVjZ7IUhvNbGd0CKS25iSP0VzLycY8HL7Nwf8
bU3886c+z4yzjzmc7vt3XWrFZtPVgKTfY7yk098UK9O3ImRaHeQzsYE38G/dgTHalDxToEpv4ocs
y6AgRMBbjCeXI2WKxrhP9aHvtjU0W50cHUeCXcVrxRxzCwuPE4ZykgQGX94RwAH8P5SDCwuLLC0V
/5bmDGeXQiYJKI0VS0b52irF7+2eUDM2AQnWhZRZKODjWp/zjoG8ZLukl4y70SKVH0+24BauAPxN
UsitN/ONlVgwTONOxOdDPzzxGmgegESqLNyZaBsp5Z2ouqMRjlk0n54M5sIPnAajgavOw7qhcIMq
iQk3QJjI8MaW4/G+wQt3oW+eLDXcfJG0iUaP8gO7RM//PnUO+MHURKciAfHMLM3i8B0QG9fMANoF
n2nKCdEX+uwfi7vTHwq4+hQiV79gAhJkXIu/ZgVO6AhTN30BGo59WsWcS7q/oekLvcm/wkeC9Zlb
038Tjb6W3ZeaHC2nxTOe3d+SQ5ZoU2WATq0m08BNirLmUlbz0sjF5rFLa9s8d5mG8mV/ixWsRHKJ
DJu7p3enCWeyslIoyoE4zhnByV4hZpBW9AcmczWUet9Yey+AH/qhz3cNjIc3k67SS52bB4Dgj21+
66RqzwCEUX1+MM/cJO9u1rZDucFpH4BzNyK4dnkyRTl2612+a265I7ABXvfxdTNXxjnE2em/8rvY
vNjI7x8TS75ZJVNMYg5pX9R8mjkaIWs16gVBjnh21EN1w/8MPsfW6ZYdVwyjMTAR+ZZQwvtn+FDt
fQE0mna4u5/4PYwQb0ZEYxrW8++7bjSo3h47s72ULizchVudpCpdQzaMW7LJBjJE4+vZ/dkf5Nrg
qBsPs80m4lQWBwNEFXdMYLyx1WoHYBjIVj3ptXqTJY8D944tedwvodd/7vbUMzTNgMozLPnzyYWV
dn61eE/DrRwfOaqOVE5uHKc+TOFBlSKmsPA3rRD8uv6vjFeT1yvqnVTfLzJdZXtTxVOxX1RpIbpN
TzVmwuTfvRQRO/kpd6PG9cMnP3ZCWbBfVZGvoHbIipMvU6FcB+2/k7wOUhzG4NC/9D7YIXxU9E9u
RrKoHRpsQTfcIfXapJWpGViZS3YZqmfbiPw49ZO3cEy+3aU1Uhhp/mMr0UDFlbyhFqheXM/0VWjl
qUuwAwkxDMisjmTKSE31i5qEQKq8MiC8WTwZzvUgkr7+pBhJgQqb4r0Js4Jx6OIjF46iqc1BbC5j
zk5NRkGL44ljWPkSd33MxXYXIXKfDpeGy9TcKugbq2DQBqjWmdsQfzMvy5U5GiEcu4WBwZfim9Nb
9hPVVNriJaRU2d7gAWRGZqcHKadFf3cwJS0jLMD71yPWYBdwksyQezjRBuGuuLbMwn/YPEp5y+ed
XLaaPu/30lWx1kM4zP3O/tmSgp4PL+skUgPJHmbTMNt6AUqqPs/mk5isDUtJgXYJjCwfiqKrjVYf
B9PJeK9C1RQY+4Cy+/EM+wYk5cjnis0+gVKeIDEN6wf7DsxCnWekQDm0fHf/mGJuXmxDw2dLqZDX
O0vhN4JLibCYCSBQAhBgG4N8u+dPAnAKjifIdkegstvVCrF7+vR5ykC3GbUU2ns2Ov3i/Jvw7888
CufcQbBKqTZMsKakGOf11IGuNssp0rRau6kQ3LwlJqDa0JL6xQPstMKCwkeNiQ+LB4bik1MU3RD2
AbiN7NNRZ/VLadQmCQ5vGpT3WJL84ApV3lRQxYF6GltLcDrSu9Tk6NhNIavustpVYbxmJlRgUuIQ
CR2TiK0AA3fzSwwqGTpWHiSvRxq9q4HVlKoTE385YXRdhR+pWTo18vWtTjw8Yi4BrzsxHB8x2ygp
ESYMWMUcB5HAAu7MlC+cil7zM2pnSmuWMjPdxh9Xhk/EuuASWnxUpbPKwa1v8ayHu2sDjIauqLsT
D3GtG928q2tDQm0yEFo9/oXru+9gOO5hbGsyOqfzYvzHbG+m0LQ9Lr4R/YowqjKU65G3yv4I7sW7
emNZEgue5owgDpogYyBpje+N+LLcBCtN9m6w4OSyZgUfcFIRdfuc/9P2NJzh3EqBNK/EPwq60NXx
pex8M4nFQaUDjx9VvD0jhn8hCxkFHC7tq9tG0+ojbUDERfha3tFkVMWqmKZMtzwkNKOuhaP+Q23U
Izju//KgJEimPLRldCPIijqnd6fIgJJDTVzBkFZJRyhlggG+xYsnduGYgUp+Auim9J70AjS5Khnu
ebtqH+ITBE7Dpxs8Fz+Y1p2FhCmK4adCqeSN9yWq4X9DOUu/7loVQh7OJH3l0NrqOPVo1/+RRh+m
bhtzrZVcWNoxyJ6aV8woT1tA3/PP+g83juPu+J5Ju0eTqabKp5coqvmDyl4TJ/m39kVgvp2DtLEe
RNAA6KpRXpCwFwJy7vIOIOOJb78LUUpacusaKHrkjOx5nwAmA23JE1Kn9H6YFXDQvCeucC/LcCAd
vvFSUPTRSBWzNHWTtvVGvX9mHW3W1sPJRnEX3w1JPt+KMYS3VRCcrbfijArZuHSo8y39GfpxzcNH
9qp/Wm7Kqs0CPg/dnW7tFJXhW/vpSo3Uw1u1L7N0h6u3w27xCcA3CSAf8ghxrydm3VBhfB8GFLa4
5u4hHxEtBrwONn1gQms0Xo2PVJ36fV9+2vP/bNyHdIc/oEHh9LzIO6oLEg1DZV2MxU/VP5pUONfs
tNsoD0C/AUNIHhOTDwvmBg27di64OEyN1WfNp124gKKQHqyj7/TCOVgf4Dr5dJvVPQFpsbMVsUXm
cjLKbgTG2+Tnw3sfDOkOKUqCb8PFrfRFvqAOrIRKNeDxxVHWT4XKSPv5MYOihd3iBqW448rIchFB
9LuMD1pP3yNuFaSqc/RmHK/evSzpF18lj5eZa3xRA0zjgn0PmpUJCck3ww3JYFJMS+oivIiOHk3z
0hDWFAntkmbefoD67EoMYwBguXNaqdKyNk9OfzyvbcH0cwXBK1yOpSdbahpt4lZLPJEus9qNz6QW
EKidsOs7ydRSHe4+AB4TsWNaYy9naJWJ0iC1fr88cct0vXt1qCYyfmjBmLMJu4m9EqQaPXgXRhQ6
OUrjjRIv3ilJMmwusbw1sfxfB8U9RSa/eol/L1RsgAGfe7MG7PRYMOTMNa0NNh122sfoV52p+tbz
n31EsxImIpf8azPlXw70ydJROPODM1pX4lruzBLzwHjxwM9XDh0x/zEgsLQyD0zdbavUUFWMEEfr
WdgH0piHa1ZnrdQ0vd/zgdE/GYBaeynajWauFQOGtwIeBYohEEI5NKY9jHsYSGbmQRa2oB6hRtaO
DJfKUZ39cLxDs3FxjCGkqfgdtSEj1ln4sQBkKfa241jn5UEOOcalo/D4xkIRXrgK/39kcp0pp1eS
JsLCN89We6O/2Z1Z2mX0a12RRVk61mV7Qy8shrx426V7ib8R11yWorCFLarYxYg1UytKR3slHHG4
V+o+EHMHF8yzezbTAYCbM1bKz2J10kDf8FmFyFT5qB49p9z0QaZ++K/5hX17OhuD4RqZrEaUjGtb
qw6B2ge7bSzbbnXN7KPX9n/Cgp+wIB1rNUZdA90Z+13yhm/HCcbQEPZZfnlomtSFZxkWHK2OPwSL
juUW/gfc4+0H0xBB8hxm4UJC83+8zNsv9PVOcj4YxLTFccfulYGa+0H1puy90hVQ3gxlpsT5+gJ1
qM9qBGyfa2bKpJ4SJG6f9sh/6jLKNKFeeXtcKseVW67btxfXJAy8cMuDXb0iQ7j1Pky47dPTTCz4
cLuu5Pcx+FnmzdulHQVpugvceIjT2C5ll5WL4WGupOSBaOQ4We4zHTAAlYxMhmcyLtvhae9iszSU
LTffwYflGtILCzKFSUzeg63IehBvlgWnD+7CfAGIBaUGPi0ByFf4a/Lri81g1ziYe5wDMURhRLt8
J9azezinPKUXKvyJPZJov9PsZQHIZI/QYcP3UMkmMAJM559NpZ0ESyurxw4TWImm1R42GIVrVN3R
Mfz338gr4leaKCkr7d2bWc2oH5hec8rdY2uhQ15d4c3rTs6YrwFUVLCDeHXlTcyntGn9j/c3bJn+
tSrFcbGmikhw/u5Xv3RL2NtTNSTWHqOTnUuE11XmpmbP+zmgGnckWUuhZFpfPHVixalwltX8Dj4q
VOozdBKNoXyBX1sQDI8e3phMVCSunq8ZzeEGoWoChM/YHQ/DRa5CEOQHgg44tHrixZPfGxiHBFhu
ZXG1QcYz9MsVO3+Y+m/dRLf1+ApQfyAr5oOW9NbQz4e/9xGZpJ7wUTk2tepNWi8lJPDklkol0MRT
V4rrrAh9ENfrit5W5N8hEb6PXUbpJ78R/68bKA6HDm9XCeW0ucX7U+2vmnLGjglhC3G720g+Z1Sm
OBg2nlPG1cXJXJGF4Oj6cuH/V8EZZOQ8MWtenzaql8tTVU6DR01kk1VNsIoMFP98R5wao9Hw1nKV
qxX+kyD248KoGI0smhoHyW6xI9FLEf6VJu0R8MXS8etRRqMJ/1I5+6luRqHyxOKzq8PKl7GtLZTt
An4cC7ixdd/wFozw184nAkBNj606fEVjlU1R1tlciJzX1edQvuON693VEsPaTWr0k/tmBr9vKVsE
/jWWq2JMav7BgRRV57shSHv16JExzPH1iPMa7HzrEzMzZkwPggKUYAtcK4d06MOj4nk9X5AVlIan
6YtLk3ookH5vjmRax3MEhruzaUz3L+mOMWr8HF4X7qf/j2460CwtOGayjleF61hNVR+R9rmODZuy
BrboTbcDcvpLyZCIo5QRfJgRQG1tyv8HPilDj2eQS7hIp2NgVScujm/ZXr7dsgagb8tHpeVwMNpj
GH7Ovr3n3tcpFYmzf++ZVUKqLMJjgY67sBsXJXqVKQANvraCZjwNqb7dFtUjbkEkPAwAk+2V8jFo
Rn7ni68Ib2QIMhaGzQ8n8/mIhL0bYZHp7RdbNbx4ub620l6dCCFrP4ztggYkZmSTHDBQs23uwV0P
8rwcAhNvPlQ11ln5I5vvNOJDim9UoBqCixHNG/jk8CjXg4MVJWV6Kv55hF47iDcexHc0QmHb0t7k
/MyizS0WYW7MuVWAnr1fRGKY+T28uPliiRHm8jY9kMZTvdrRWFyb/53sM96L5oi6J1yv+Lv6tA6j
7v3bQ+tRS3Y+k+rExR0/LZqBrBSL8+HCKYgZg5guZXZAG8wz2zUF+LNzKyvkr3AN2UdF0beJ/Hey
evPZPTifEwSU/ZD1GZQIX5Yo54YYfqGhKaVQjP9W0qHNLFzwgJa5ahpOyjhBhypvwVsVmUSnKxdp
MpqQVeGRpLUcqJN/Hsbvk9/PZTZppm0kKmj6PcEBIa3fqBM8rAp3u4poE38v7hQl0YLtttXfeYV8
P0VOaBA+N1rtpPAozUkafyP8/XKecNM1VXTSceu9H0Z+VTuaexea95RtoHFT0FVtIjUIWy26MKT8
mlc3Bx7vhP0xfaM3ZomBOUKKPAUPZjQPVkgjZKKkirXtvJmzncvJaVs9e8I6o96n4kP0FIlY59s6
2e1ABIqSsgEnsaDRK9/AD7m8TemePY6RtcMGKBUIYR9SySM59h45/miL4xlJKJLXLx+a3MsesdTm
9uFphMwgjJWu9XJ02Unz4BEJDeHF4lpOXo41PH6dkdNcwOSwXnKTqAgV8mwsQXnTdUUCheOy/krb
DmpXg0et12TcS9D02A+m4Pg3ka6RnpcWypBeNybx4sWaXSjmExv1AaM87tdSF3PetZVaxuLT8FSn
vhJUQy7ALqPqPVdn94kSJC7X8ZKt6Du1HRpUx027LwV3tNjCOq/xvgy9px5yeOmZoO/Y4WY+rGpE
JVKpBF36peO/kek7tB2P08d3CsN2vx9JERlO7zbGgHQxM9j2BZ66F1FfOKa91BeMtBSQMEM1U1jJ
zkG4TR/Y8PGfq/t9Tinh1QNAgC92XxwKSDyoaDAa2et3p51WEu3z8b3+EmPfVJu3RWHo9MaPjKRs
FXwaEBHJjGyAjeckWS81tNupHTW1Zo3EfsSMMumJV5tBEncIqiUku1Au8t4EOJGsdimKIxF94TUh
LOulN1eYwNSxP/6Q3torO1hRHaDhAym/9QvYDidwiHqIhEhr+bkmiQpGQo8B/RsWT8PIG6+cBKUU
LfOxGj4MZWpGR1tSDPRpVjTDsAZl8s0LXg6FAy9DPPMvj7Fqd7Lk1dB/TcRHas03UCfrJ4ny8AEE
J4vDmm19i6gZb/1f/p6YQ1ElCVU+ACfQYnOBkdfWBKgIHRRku2Z0trrC/yJ67F2sfzE7nRjZDqPE
Ze6BCsEzheBYFqYDrn9jOQ19XW1vBXDMZiJv054LDZ3yojnkin4C7QHDQAjrzUGVyjeimOY9CSuk
HRjXD3250kKD1zwvdSEbdeO2r3FXbu3BqvDB1+13PHcTkFvGfui9K6KIdQQp/MAUEEeibJrrtSYo
1+prPJeifimQGlymniFnnZW281/xRqnhI5q8PjVQTYG9xRNrDAeLhlep7BKGLC9j5/xnszKU0riR
fT2aOgANM1jD5qxyvV8D2GD2vPqP/1HFwfvBdUjOyEsnJipTVCqpkp5geFXXtcJ6DtdS2FaNUrdO
nVUyg8AzVJbnj+twa4Y45qc71rwKbC7DOqzRNrMuqP5Z51dsYj9KfHvi9zJOnqZ9xBD/lX/XThm2
4RSszVLtdnbK1dCkBw4PhsQe+N7+U5mPjuQ4UuP74OTTMgeSWmXAHMoOu9Pd9nYUYasQM8x1SG29
K15HOVWtPDxMbnmNkXzIQ0TbCUXEox4D1U3KnfwyPBTpuoKCSeRFrdnGLsG4BHwB+QkRVcH3fkEd
hLPRuV6EkhK33eFzWvlB+ALpJBB2Mb00VFd95En4iHO9ijX2AZkxFSIJKsj/WynsGoaD6zlBytN+
663CMIGhQVERSd84WEY23qiESBAcEiPT2gvb8SFHIbJvCUvUL092gQYqyoS0XOds3Lh8iFQRKNyN
SiWC1UlCzidv4M2DHyjjkBQ+oLxlrqD1IB7KAL7gs/+rC5pRBusFzNG5KG1jqpbYt4KyGE7Wl1WH
9lnEcmLtK4t2pLjHuzDo+1FtwwsCTT5vakHZuRVCHYeVQ0+HZ3I4UpZJ1BRb8P+6L5kiL90umXMo
str1+WafJUggieoRgPMXEIjMDhGDwH11JJ9BalKt+OaZf+E8Tw56Fup2qE9onTuXuRM9ZSAtykPS
0YDNqWNG+eOsB4YqTL2WP/rjBohOnmAQ/oBpWjASSqHgozg+9hBYcjFb4GfJ7gmoYH/RF8SUMEJM
U4Z3tbuqifU0aOuanJLZeKabafxoOTWTdMm+DKggp+VcwLf3ihR6HeqSxuhzGmfPn25seUbvh9zv
P2eZZHsupSsYY/wGirlXUQD3YErAFxuK6naVEhOqXhEAQB29RYiChcFSfRbqn8Q882qjkaDUn8Ju
yTdqjWLmrVJeqYq+ayNYaRjYJ72hPJd5Nti4o4L3FJoTW115G7bWh9F/rJzwpdIqEltf8ih6DY4g
zPySiZA2XuUVoKZ7rijCDmAbmGoIH6oqDjODUTDBmp5sNi6gNT94sT1K7xIf2JYStflKmtQe/4ks
aPWOo9adSkyIJ2glII9pFQP92c/aNaxyPV8Ofc3LKyz2HL2C1UyafbSs8im+wKntCxNL4ryvKOKx
nrlqp8IMZCvs1bDYAne2VuJZAgGJOKkhvQ0KggdhHlqlkznEs61kRBCMGQAb97p9hnLaI9WZkZig
ZsICRZNJ40+LNqLM8wP7p5UlT/G5SVTD2oa1JEWMXmbfmLJP2y3GJsEvK9JjivpMP2t6aS3jz3m0
rbHuYI4EGBFv4PYZH/E6ec7sHU7fGLIKJZgOstDXK1/C5/k4j9QnpVV+D04X/1ytD1NhbF2ULGpS
opRj10vtJD1mt9cEtkemHiioR3VebSm2Uqjx4C0u1F0vanCVJuFbx4dE14v+d4RnRbhWiy/K7ar1
2CgPV4WFolWDU3xRUdyjOql4WD2e3ReQ0SdpD3+1D9H/8YNcegOYduvVt8CbXzqebp7NZV2rNtao
J7CZ0/kpP7ylCMQEzR01gAMw4chKiSIRnMOMukTB1zpWVBIyD0ato/SETMi9qjQds448GdBEk6p/
PSeqzsYDOr2HaKZIY35S1H/eyRka4ZHLokkALwlN/Mhd53COgkPCckI/TCsNlC33xa9RLoaiibfa
+trF8SgQePEejm+pPXv/teN5qWPf+jMbAXqUF+vyg8X58XufU35iJVRRyAmTR6Et9pyDClTycrMc
ZEfXKhCjoakFM/jwPIJCGDXXDPBiD7SdrbGBQfwkZOU436ayn7Jy/pAQ4R++rGz9MoxFuBlbR9cs
aM/tqe4pVf8a+HRJhT38FAQsbyEw0jBkDOD2GbYPd3crF4U2qQF/wRlm1PxKS0XMOCqOCbMNjgHq
wAG61Nwr9SnGZNNU4fOeNnBT9Yfd86kLUE4Pu0reM8Cl54l75la8xsYAktX9Li+xgewHfIEAZtZ5
cE0ioGv8Sj4YjNv+83BH0ZJaJ0UypwwhG7TBMoldTI7HOfyEr9B/d61liGmicLOwApZP+4UI8+RA
+z7EGwUoMQkBnejusE3+d1L0Hj5HXjXTDsvjkwzjQ+STjs8H2hNXfIyCmutlDyNq3PYFwdsEYIo9
bBLp+pXf3NfwZVQ9M2H5xiym22Q1ENXo54sFLT63AOwljfEe5MqBdO9q+KdaKumBTeC5mNNiJgRA
ITeJQQtJ7hwFkPeY6u6PJOPlMjxlsQ3zaRncs0IJnnp6J6rAPWs0a+JPLrdoVmwz3Oxke0mM5nWM
TynRGV0s+N+bU8wTZnAdBZVOlBnjHxrlZv0vscb0h9rvMZ7K9qKWzTrtWVAQkhFy1ySxtV4aMMQX
1xYS21iIiFFNzHC7+MBFrvvKtkcoopPWcau6hQXxy2PvClbRw4+q/K2TNrg/qdUwZs79vx9+aCyj
Ni8//YU13zW0Iq5y18yl6F5nTqo0dCdZnnEnOAB5I+ALhjIgUZxhapu+4FLP5S8/ibsPMdLTCaWv
nc0FB8w6jJn3Xdp+jDZHuYzKXmgbP6WjzTMVVGWDx2W0zYLkErP6Aa4QkxfYbO8rkGH43CvksCJA
t6NFqn8kT7NhZCdigzSdpuAZeOWcH46ezVuTyVPPFCPmKP1BN/zzUAgQbLN68R85AfAGRdM6wPYg
pgvZUfacBXC/jlh3Y76WfKn4DmPHdhIpy3zN9NiMmqkLX/JD07KuYa3Kh2BkExgGtJsNhdP9ZBEl
RqX8Ej7dfEmo62NYQu7dvKzNZdcPxc88QOfmWqhjzisvQn86I8kSdIClMeLsgOP8Xl1s+ApZASuq
jIpsVA1M1Nr0y/2FNitoM2Vlx2vVJREXkliWhxsHU9QhjN6UpgF2s32bdmqGaB3Xd8ptdyY2RJ2c
qXm3IYZ2X3MVQ/GKbr9+vtoWVIEjwFFUmLuKvCY3s8UtMEiHg1JPHQqzOax65OgHgIK+MM0Aqy2a
1j7lC/5lpStvS5PKXT+xUSl67Nf8GCfcnTzwfV7QF0kGTGYSKD1RtXra5rtH6h5P9/E8PGf8DbA5
o1tUFvp/AKp+foMWhFfKdjg6S9cOl+IMNwiGRSIVDfUi8nPHMP/zElNdQSontc1nxTXZiPD6Zjfb
dudlBBt/SyCBiBMCGsMVmJnm7El9mRCNn1GNaZWoZ8OKnkI2y+bvt1Ss2EQdjcZFgP7mT0Res+qn
yivHOUu2BYnKfFHrNRwPaGgXJInOBTujbqbE7XD3jvfJai/ciwfTFt2JFdNxzQ5b1EjkVqZYQLQn
BVSYgdvI42HLDaHUlZmEejpS75tq3yvfBhJgonlRuLlmU9F5BicsxQFuROZwehB3glypMyX0I+7z
y1Lh4S1cnYk73IYU4fX1lnbo6upax1TLKfx1yinwHdoQao7pWWtAE/mhBE2rLkPQboUA+LW3upci
UXPDM8f2DR5tqLhgD8q/+tk9VAr5upJVinBTRdK9RMIreEInwL3oOyHdKLaiBPa9ZcThneuC6vOj
8J99V2IzZ9pp6KiRQOGxes+zb+1YVeApVlUJBiolVLAfCeFEuQ9uLWziOskcGVn/0MfCtCQwy8JU
su86oWEonBc8X6Cswmvz3nFF0Oj8kIrYvcUW/Ocz7mpnsFMzkFnKta7bml16LyKSmLs5yetleT7i
qc7A0FWXUIGJt0BeHkkdRG5kRTKJCAgv1Fr9wsK7n1JTN2LFGscPLCV1ZK8nBAy9tZVgYYgkC8/G
xkGHG7omfYjhNKXvGsPlrHBSQ9wm+0U0ZXqDanC+xwzfCF2Niz3M1GYXkcj9nwH5m8ltqvmHKha4
9wsGzUFAmhoj+Ik/Xkh5+5Nui/b3hG67m/cS/yArvD+GNK4IdaiWrDUigovQrMaFjD2SNEEGCF6R
XLSr5XGzKhj1oT6xO84zhF2VsRwyK/69ZB2gsECYCM16NbKb3pjjLJ4le1i+asPmF9E1XuIA9N+d
+kTiGMTlr3R1gx5Rhv6N/AvfI52yasVM+kQ0G4v08w774oh3uSAxKFJrF5QPikNIQr0gcTqHHh04
Vr+SHE7cTvECkRSl3vbNpPSYalhHye7+7SLTzTRyCv/s7IrKYUUc4HRpUyC/Yms6maVzDzx8+xUD
h2yRlDRX5TvITisO41lWwuHPC4roQGzJun/yo5W6pe85T+AntoZcZlpx1cMLlLKR7lyz7QiTdSLv
jcmKzuDiirdbiKiPeYotswlMeI1FAnBFUJrel3AykzQchksgv1tDzeu5pp/KdSOYj6iVgcIdmB5V
bqAlmu0mpJCvIMr5UogUaRqtpYmzjg5WIruR+/zTpALVRnFwJIciTrndDzBuZqoMCwYUdbS/Ebl+
sCqAz7f76qykwJmFHOzCydD0wW5veALEPY6rYHxwNX5FgIytjvAn5Psjo28Y/rsCzhpe3az4fYH0
QfzVGY5NiwWJjJFyCYh6iKCfFv1mqJinzaQYmtr3l+mCYxqdlWbFBVwEEp0l2POq7JLfFSBViE3g
LyjSzx8yvAEh/JcuAdAXrhYSI9J4W3SJVxYahSIGm8NCVHU9lxM3qxHx4AYLmZ/DOCSF0NpkHpI/
0LL2CYWoOQbcXcOf25Ek/vyLTO7/mIwKS23cFniX+F3BpgjDZt+OLO7mpp5tzt5znJ+3kJJIjHh7
4fXWpoRXAXDjfja242tmSMsPQMoTomMQVMZK66ohw7ljmXsz4pyhBJk33JBQ0Ug8hqiTy6WLOu0C
wRsDNL5ubBM67XTD88bgVT/AnZbf/jcrkjcu/f643S75tnr9aCF41MQd8+Wqjn1YkuJn0NeYR7IY
PGgl/G4KwII2nrBM0eZqxkEDlVRDSCsYWQga/J5UjpDFa8IakSrRA5GCX5ulYabagFVT0NILncad
K4DpQ9zN+Tmmr2LrP8+uus4mQp6rmaO2pnK/i1VukoymopOwGB4iogXW20RrANUsA63nG1CTvFmK
z0hpMJUBjGTffEq7sRi/4JebA94/n01rdmNnQHNru7KdOV0uoz0PXyxRynwJ5InawK1lYU63bfII
daGr+vjfFYDP/aqEuip9GBfFbCBItrhEljt7e9diebOfNP1Ae/nuom2H06C2GhwfyvLun/wlvdXR
XbTz7JPnCTyfhFNbkK6GNHVHUEOQA0/7xGeOf9jALH5I2MNUbAl2Tef+y2zW02eO+pZ7OIf9770/
NNVoE/OT0U0aithnMcFLB5HAouUjpWX3QT5whkeQklUVeXr/GP5AA8KRjybsIuxKR/0fzTct0Chl
8i4rvwMZOrR4nxdQq0v3AYsiQuqZX1oehHKJDHFfb4VWJ01l+ajQoOqPG6gNvkpgsAyqWkhnB21b
b8tuztfENqLd9aFtorszMzRldIJroUNnwVtCJrxwS3KelIH6C2tgjcaG+ojU1Trjq13eRKlFyJR0
TNPOUVCcqk5k3z3JcSS1Mosv71lDiQQb6dYqv6rQPQpatNKOBrVi1B7+zrSCGUKItyypKQ7ZjMZI
+xWEoCcZtMPuzy++fKDncAmRLU/1gh+JRZJNtQe8BRt3sSP52kaPIRgyNHLQHiModI/OsL8uts+H
/ax9KUUyoV3EDmhXhmDqfH+vmtOJMGOrg7pDF8+bVWMmWOKMbZ0MZCo+k16FuYdH+Eg44mOq7Sjv
o75n8mBsAkyYqk5dE/3YNP3nBj/V1FYtqbO8IVY2+4iaYWmVN4MJUjlEXXVmClkiaXaYejMas8dt
ULV+uYO5Hy1caKsfecoBEx78BRBB4irgt8J0i3LnD5OAaT1wfO86fukSKQL9Bl0Ay5VfLclcVB7f
K3iYvfHc5SoAo17IU7kWNjpeE+himz4joAFm94FoIeEAlTmix7+LJAUdtiBVmQh8B+muQ5b1KwkN
4ob703vKHoLa5Opj7S1McLaGJtBQpP71kL02hdPdvPFOJOtnO3N0A763DE0ecR+OGpZiOf2s6EVj
KOC8cRTB5VGaJKA+ZnjcIqMYv4ACS+9AseMN1RC3biSA6ue3Mk7DByi84oTB7fbk6AG3kadIdTNp
Nhpz9qfFgvVMAXT9CreUW3aTI6Or2ar60cXi+0ccR0VZOwRUoHgM+8hTrDOcWZKbGNAQxT04+ygu
olxV0DGfqpTpNmQ9+/NSLfJ0+/JzhAZjmEUfmgvSGVQylhbRbRCpb8nC3LGv8NITiJR4X13yFrIh
QPLAWv12Wq6qV5FkMMQSZws6mppvqbKyn3veplovKJByIP+8kWWUOkhiqevEvCzy8hmCaPR9Tapv
oa7+s7eDrFSKhz+bRZkSKhsNn1yIvFrh39v7p35Kt4X22CMdcYP3k6kW62LuXxs9W9nDZeVbNc3M
YbjwSC6XJk8VVE8Or20KVJEMPyToJ1WvZdYLDPxZEEtiGLA1HqZfc+bkO8V2SoALq5b0yVE5CXz7
pH3d1gObd69lBiM6GoMGbtbdLYRKjEDM3GLH1XvpY+HbffWFSGinV8qjMuGNudbO8FRAZuz1r11l
KyuyOmuQFB+qIgIW8oRj0KWzqb8UrRG5+qqT+AIxr6PyBCqy9wCLxpgMj9ONZvfJWI8Y4XXxN5Wl
k5Cj4FyQzB0A8ZiXwaqZvLqKdxf9FyFTnRiNtBf3leW7/+XGB31s5bSeFUqN8qVdDt0sJS3YRieK
Ih+X/ZdDj+5kdV6YOVgihymsRxK0InX4KHJV1AGsxAfKJ7gh5g7yxvGU8L1nAgdQMZzgOGqFEQW4
xdgOE7P/d7KC8bTLf6DuS0VNZY5ptV3Rinpy5K5/WgFpjbMwkrka/ZuClt4k4DyGJjtMXxgc+yRa
7X6x+YLk+nGBdOZZGAaPT8so9d3Y0QnpC3sW3wgaxOPB/m80xn+p3A453fiV3oZxKFhpWi/qEXsF
KiZTvzBSPvDe98bs6X+bvzsn5+hbAxyC7OeJL7hYpx2FY+YZF973u8xHn68ePXuCmWpADr8jPBt3
xRcCT5rqQTuzz9siWZVqwSiHKDaBG/2pl0X5aCfKp+o4tdiEn97VaD8CR+RJ6X4la+5EJrj6i499
Yvob5I4qHm5AlYsM+/TjC6r8cYA7b1z8rX/ct67N7ZrnA1p5L9E9x1gaR69FT5iXCV+WnTm2xIrN
BWDdh3s1mxi43TUmJrJ//9Oxg85idh7uZmdZxRC1hihmCkNQ2mOxlzhKLiuusSLhuF4fAexbdnKW
Zu1m6BNbSN09DuJ11KK4ZJDDLkSj+NlmrTgzYGiUr8klOGutEul59tdp/u+mdlX2vCI6lrK7MRwN
Wt8PPkY8mUmlD4b+oPXDyaYDwKDVTfpnc++s5CMHFy+HSXSOcNFr84hBeMOyg060auX8k/VtqFV4
53R2g2WSluZ746i0zbC89n1YljK+x0eBEPzMe6Xk1lgFPSwuMDYWm1NXg1HzrbM+wMuwMweTgF25
a4KEsfTlfMXPd9LpxvufrcDAImWBKAJ1pZpbWgPP+HA46HrWNlE78PD/ptOk3HkLwfeBNDYk2Deq
TcdtF9pVhevlWniOI+ogysMM/8T2Xl+ePcHS6+38D2ENwRAlsXQWdtWhrO1H9BtCeBTzM0Eh3Xm7
9AIzW68ENQmEAbtf5xDUhqUW/6dRsiKuqlcoROZnQ15xu85M3A7YMrFn10fi/4tn9HmDBlaa2AAE
emRdikbCQMlNtHtXDEM/9FrsnSCBfU6OSDeKQZnPZbie+9/fHu+Ec6GHVqOzijmHEkLTGJTwMVi5
iL2p/1m5Jo/abEjJ1YdiBKRQd1MSM9nGS4g0eBquRFJeDGxTVMCN5Yl6VwQSreFzBHWbMAfzmPQZ
1hXOtZsWuQtJihW5FZ0aTY2gaWznwOtd1PgYPRDYOCwx9r05zZilMqlGM7bNxjP923vfwPiQJra+
YJHIDkkMOdAHXponazPQL/2Oq7Q1b6QHx+yg3+KauNZHwBf6bAD09pJgayyi33GNrWlkSVha3xYV
LQglCFVNKT4hGWZTxB1K2Ht0VRiZPBljGmvJuaCKTgPViGX8l5LZKkpCvI7pLbNT8ZCJy8UEYHiQ
jhdFBGaGAjaCFH6unxzFkZfrc94edHVaPEitE5WjyfuXgNfWos7EvnjO0WI7uObk2auWS01JPJkj
XPfrzNFISyoqKEOAhpLfvsMa0tXxVJk4Ic8J77V7WARbWF0J8LYQnA+PJ5rWJ2wA7jCfm0FwejsG
KLcmlz418CJbuPpGxxbO/kl9sATqq1we6La4Edu2VQgYtEpF4Z+1oCx8cUUZoO+l4keIb6eKuUed
ASZDDcFW7qLrK1FbCxCxpD1N3VuIyJtE06l4uBMHrCIGK6Ri7C8rKzKtfRLyOtH1z96UwPDZIynw
kN7R4HcWlyVxAHzVxvk+7Ev0VFtp1ekHSwHJySli57VhgHOKOml16BTafNtw4hio+lVC9Ve2g4ce
6am7ubWvfb41UYQWLy0I4va2CXgdFu7d4P3xqJoVNDzMSdN5LdKXdfumy7bcjqwPgonGXfBZlFy4
8iiOLmFQqNUcpP41pe3DpiSumR6QtzWZBcK0TFsiHUnCkeymoWiJR8aTRn+UXmxIx61bJINGcMzc
zhKofnSmtFe1MNyqOHTHzrpbat0GBo5NhUvTAdZrihjgXfh0dT+MVjlk4qkCyaW0VwjbB1BuSAnZ
FBnDvm8CkLihlAMUqc95VtViwruBIf52r572Ux0oOieaBHYTJh39rOr8wLNOaPC+fPle0TVHx2ve
Kk1c0VuGq2EqzlmxEuamAT7LGBj/0d56RDzEBprr6CX56Xh3rmlVwKpACQAii8xPmlUw2kLfagJJ
q/Uli93iLloNZfPcmNfpG52BHfsr2UYdyka4RNS4eMpFLmcOWE38zcnNzNfagOBzToi1KZQyn7KV
1ogn1VC1sQKG0gV87lxiOCOJGi2nsxEXwVxyRGuPrMmRApdyqn1PCkwzf1PUsF+sv+g8Aead+JF4
Og8JBOyKLsrS6TlTpp473vRcv/N80FDwSl4JdOj8UzbzQocMN6R0RykTIEb1ukLkTjZCbEr1HBEs
OIeoUdjaK6T1gXAoUmM63xf+Lar55xsZPy2uHGv/XK9NAk8sS6JkjunSrw6H+8WqHXRJyqRQy0RT
nGcO0hJ++1OTYba/vBMEjC+arwPDqDq8a4o2gGuHsSJZZ+q6yZp5x9zA6v/leaK39DDJAbLyb4P5
x12VAMHZBxAjp7wYxk8mcwYJgga5X62EOXg19X7RlsrBq1vsPpX+mzb1jhsTOHF/pT9HSru3b0a/
1ELyKfiI9eXrpEQPK3n6ov7pPkBgloqCZLFRBqwL7EXwLqsOAc+oREQsnte3iZ65zC8rbdcvgxHT
imsf85PoM6bGxrRToaZerRvCtYonQ8/oj0PjqBBgECDUNbebT0jdJzJ39ZdhzpeaxejyeUaVvvSe
a+g/BJbRi/wN8GrGHsbwy9Zki/j/29CU6sToJuR7KSgp1fK/l45Z5KWjs47iGMG9mJfmwy7w1I5Z
iWbmRrgc0RJmPKbxcAdwV4ABJ8TMKiT8ud3cNY6AZPpFTRg3NVsgOORbsrHcGBFQw8B8s23ZPgdp
TBIOMkxwSbmoTTwWvaBGP8uGYs6uiX8tyXQ4FJjbuAestOyJOy56ZN18Cr3piyNXoAgb39LBwbHP
7NvkH0s9YyON8tFiXq9YhY+kB6+iQARvACvl6OuyD9f9A50ekDgNdCWnNIYSoYGg6VVsKxTvAc7D
cZ3mQwKpGsN+FliI3TKhXQdpvaXIbT4KCVxQ1mtMbRxRm+Y0xDNsvp2I0xr5FIxqcfgm1ttc9VQW
D+oxsgR7GDkIbGe8VYJwaY27A+NVRmthtjeQmqJecDvyfs8F48sP+DdJeqQzhq6xpkfV8AUC2P10
6MJ6fjtOXLvw4lboHm/jV+M4Vqqy39Aug+U4AgexuU5s0X/dx/Kep5+WAjIutpw6PvVtZzXT7vqK
NvjYnS+xe0IESIKs+iCZPD2bB4+Nen7XiQ0lG13AhSV0iAis+GRXikMnzzCWwp7THYMW7vKFHave
Qbvek/uQxY/V9RJ34VLpT9RfvRhpwiY3QJpa4O+PynbtKxsixJlXqdZ57dNLRnt82mUsAzX1QjHq
FnnqRwjd+1BznOB9n0Kz2PBVN8vCjt56T98VvNYNVS+oMLnhNOX7TEWZ8zTL4GYaL+t3I6TLKtlL
rfRxcEGuUUyWVbzc4owaPl4F6fxDFJrXPehDoJt/zAN8QbHh91keKK+6I36TdpXtDl3m12kdfyOy
k/GTdQnQjkSnqGa+fEDgIIjBKcFgHGkqf6NA7g2i1f8Ck61RsMGSVbB2GMfsjFtT3jzD9Xm7xkF6
ImOKnuw4frMgk8scVoC2N1cQW/fFs2QT5ohWDClzEhM8lJGi7ZajHSi0KV1Ofja2FBJeWupiS//c
3jGCUZ4Wn4hxWSHcxlsdTaexhmOuu0Y9Op6o7Qr2UOIdKpGfT/8KQY0KsMSaJ+KYoz1CmB/mddcO
MenqgwE4Lc0bLVnTc7gulVfyGQPs5awcUN/L07nYCQp5oVxZi7QfzZcon9QG7GqLGHF2LSOu8EXd
qsEyCCcb8p+ONV7X88X/8HXjGixFb+L641F/IlF12g+xsQB4/zF7BWVf/1L8ERNcNjGODl3rbms+
raJlggn0kwRIgOPJuPedMeTMxWTfGgeRnx35efMJDu69z/wPQlsXgvro/ZiCEtfF3ZYzBk5ZL9c7
Qg8Z0zf70XR7w9SQ3pWCWnbx3bppmnXWFrpMrvaVz7eTqisuS/xxna2xxpuidzoLMpU4q81mgMkZ
+rTjSN6w0o6+Lzy9gad9S0OYmX560ggK6ZSIf2z8Ojz8RHIBmAxykRRY1y6OpnFd4I81udHDMCzS
++36ohLy8EAVw6UDNLIDnuQkEZnLsWaFDzo8tpvVHj/sboQog2VExHv6Y4kf446J1geu5LqunHtF
nStOrIKMF+6MZoQ+y5tnlfy1LjL5RJqUf0DbXQA/yX0NVZlLfy7BlxoGP1CKSJZf7VvxNYaHc4rn
V9iDJaR0jyBlAFVJlHGlcwZltko4KNimasyDBrkMeKdOgRPHauxtjAMVo/tXvD8j3tyPnHkHrppE
ff6bKVI2hCRFeXOI49DTN4bdgP5HEn2+qnA0KcSv4zeXyYYsgPr+MZ6Sb7TCl2kyZYmSeX83fNKu
GL+bnjl89Z2PSauaPsDlaino9pfFVo2HPb0IETlO3iVOtD7PF1+QV2RKZxjV815aeGa3dHVyp5bT
Rj2fPF2+IQazBYg7xnqrZUyFX84vaNSBnWqLvHPWQsehEYb/7FAmf+98g/6xzHkwBje1LI5JZAbn
MxOxEThh0OyebCeXSQygOB5Ps+bBfQ8fDrEEK8Ite7tNxLQzHoiygiyKnmt1ha5iae4N8CPAsvEZ
aUS735PhOLX6HvZXVwzZ5qkYdKJ33lBUIkI7N9lLONH2Ih+cl0KktvrKBzK7arq/Z9MNwo85idTw
L+a2exLfcm0sDzrOsESXCDkD48QL8EgApEo+LWEqiE800i4cCEEs4a+7VXE0FK61gpBJ968N86QO
fhmK8BRN9PIT7iWn2S94LrSVfqejEzVdDSgV3N+P5kGanmp+8cabdmwd0P+ffgO5rlLTcgJ4xSk6
1jvCY9GDGAgYuZ/uPwx+4FTbhiBkygDNKgJpa/H4ZbRz+dMi0acQAckKpPyOIRO/z6B/6IeX6+BN
eAvCU/H801WDGdIVJlPLmho3rRFC8XGfLyW4pe2XjKQNexILmh/bqgdS/Tvgqjgl6UaLhyE2kg2c
d9x1jG/iaZcYee9O61xwu579GrCUO4FyxjrRv+/dwFsWlJSLTea/luZgP3FyXNwLsaOjacqVSlOQ
Kqtbj75jLq6c4UTOzYTuMZDtbTbHCvFOlWrsO/R1gv1fEsrdsIi3ZYcSAe6mndUYnZUJ/LrwmFfV
Lkd/JurAmBFjPItARvE8hVbH5hnyarHF74Xplvn/vGNbPVrL/qmQAvg6nqmx9m1vio0LmIUiyXYX
PyJwgHSBX9ReW3yh+Xa/Q4EHTka6dfk6JaVLiP0BQAHprKmrycpNcjDRnPySakhPL52NWG2PE1xf
pcYPSVmhzvZyPia4Vhs7CNkTK44hJpqRbWOACq5H7aouQhkMf1FL6mOtwwEUXPJdaG0T+guy+8i3
tdaF6whmKFJm/5SHBIoNIPvTKbfzUoTM47GuU86cQOPSFHsiND3aL+eAurxoXNajwDNN4ioqIzmu
+CO1DORxJv6kS13uKSNPpIlumd960cV73/W0Lzx2iDuq6t2KwK8jSOKNhs4H9Z1+RlMxW9v+fxgC
j1BS42Qz1Ow79auxnkzL5rOviPzXfrMEP+dPHKjr1fH63xB9admxNjA6L81SR3j/J34fUKZL7qIg
3SVR3YZzUGj4oF0xgMjp40PNHcbj2Oua+iXJvXCzUuhmI7cpcYl8zd14GeyldJTVoPNoT0faYGoT
Uo3C52HjCRcTsxEl6oX0/inIW/Jpx1vRa5XFbr86xps+jrKMK3WCUUVD0dzMlcfnrn7k8U+ckZwm
dfZOQrRFF2SvytMZbtcnWHFIkGI0DFCSvfIjHmZyBQvc+31Xr8djgmcIXrwN9H55I1AwnBG77eYF
ujjRlfO5tAebtJGRbd9iaKgCQC+38PyVpHox7s72rROjtyWuq/OIUjrEtz60rRLUDY85kD38j2GS
Lb+5XrcvjoeUELEFM68Bln4bGT/l66yb4iMY0IIwhe26hgiAtmD0myqoPZ+UqPru5vsj0FCkGdVu
KhdYI455DXQU85vRVxMFULfhlNnTOWO0B9mwzQvvIwDjK+7i+BC7QRqgOUWsaRZfXkSrBcsBTJ00
T3yhcbBeBxuUAFwVZJR4VCsuAZKUh2Dnw3y3D/vw/++Fr3MthIKUyiNxyyOLRHpneoQMLvocl3ef
4sehQlqi1o8kg/s44CJ6FutFK/RpLBYWIdfcgO5oqfBnJMlaApnYeRVPuIP4s8DWIVQyoHQh6iFJ
yK2BbA21O9+cEm73fiLcSC+Lt6MC5+6NwiZwvyh57H6rUTlYuSWku6pbH169CDMANfH1ypGjU/D9
kAN6F4vyXFzODXKZpgXgd2KLQJiI+kZCDoirbYlQqOW13i5oHZkNW0Jhj9eRSEoT7BNhph4dVxkl
jkxvcpxXCG5VjncDpv50IGydSy6CxBed6y6BqA5/a4N1EQoKH+EsqQ6EqslfVdtUbhQexxS4GIAy
vfDE9RgU9T9d89lm/OIbO0jhgjUIL46ZQCJ6rbwKjxtTf0Yq6o4kBq094ykh4Z1ZB9eVQewaWgIF
SkhdNnNCSwWcr1W2rnDCnFVfogWggcAP1esJY8HORUgC5FVhhLs0lNi77B8rkzv4uFctZAWqhAls
LZZqpPHfpZe9czHg437n9V0aDNqjxLHRyH4z98i9weNSD1GK5gCA9CSVwbeQluuoNYzeeOtpbGDI
R/rsOGKUbxtPkAYt2a9+dBYvugnImAtR6ONmt0nWIqNcHsW0m7lD+HoBb+0GWOTXqdHGBpPASpZI
LYbjdh8Vk/DKXmnd9uOcvHG6Bc8oH5QUHxZJsBSh4TDYHwkk9pMIAaI9wg2+hvcE/NTJYu1mXMUn
fZLgj6LA18+babk0a/JJAWuEPB+K6Zs8X6YBrQMohLt3YYXQPzmGlhuCOF69GE5upG8aBVWp38Ox
Y83rnmj49NpO2sq1NZq9lfkCHkG22T3f36KVb0qYyP8q/JsIu9RytwF3p7yZ2P/SC0HlfE3e+kqI
WUtFSMSZHWQ4ImvGFRgL/0nja7p1bY1rbYkBboRKToGwyHcUgrBgD/VBnE+WL8PN0k8ojUHWK0/y
GEOcm5Zp2QAJAxUIbu27uBu7q3gOrX5wp/ao10xP3BF6soztku5MulKkK+iV/Rg6UeztqPLIWjWA
0bl/n8/4DkwcusvCoz6vrmp6+iYCiA/Uz49RUf70nRFouMNV0hjssM4FQrbcyLTt8wMOQO31Dmwf
UZ7TyrWGPKzWN0QGI6wigKN2mUfHM6b34USi7ShPQ9n9Ixz+TMyN1i+jSphGciDkuTtR0fployaV
rgm1Eh7o1QWai8BoIcSwhVR9hY/BiBpfjDQote9AP5xKlDmOLHO/Qrsi2gS+eHC9Ro8+H7lNShsr
t9fPjvayFhjuQZSit72BFnUMB+pXTYUEGcVrd1TfmGUgNfoTAhdXI385sk+XDrP/1HHEKfbwvAR2
008R3gVi5nUq/yS2GKr4sSkfxy8WnAiBCqOO0BF1YPUUcdybIxAQy5R2Au6jXuVOV4c1NWyp3Q8g
6m5KC+e3F3DrKqf4+exBtQMH3k5sFkmDHyWZK6gCtB1ph4XuX+ocl7WGOmqahb0ggbyNy+TqNvCr
RTDc9Y+89DA1L3Wk465+b4j+e5TozC9d8Svl7u6H84AHECSI8WvJ8cFGwmytJaM/kow0mTpDK2dv
+3TatcUKlUzQwFYUjMiAM+KcI5w1yK1cJ5uUp1r1JX58ZAGffNeAHEnSGocXHzG34M0mpBX+glEG
382VpEU3gYJrMVu52PLhQrj+GfCuUQU9foWq58jfAd6fi57SZR3bdouYyP2hcjgtzQfZmqUPWEmf
pC37ZVrMilbPRlNPUh/eswVKdYzDyaIFdZ2AExeelF6wBPeY7d7Wvg2EYEXirrXZsXwZswQrDIIv
LK/e5PJY4O8/GyXRE9z5WsNVZIerap61q2C4kBaJAoN8/bcmt93H1V5JChS5bu+wdEtzjxjX9oEI
7Bg141d1U2xkvVWwhsD1x7DpYiQXau5zg64ptSZJJ+uE2RqjwVDwdDYwWWPJFh07WeOp62BXpCQW
6jilyfBJvO904PumZzUHs/gj2qvMw4xcNyWZGLObCIdfl9ho4H/avz8ODySiM3svqIjki/Vu/Uad
+CxZbeCQ1+qgj/KMKvWcxCX2+RN6P1cM7Yc/t57XvdgCA7agOCZYZz6ZffXwY60lcjd5YY3EvIZl
zu1kc0oQoIehoXpWbfJzuCjVJvAfcGc6w+1eJhTvNRVOHGbK+B7jFbFwad0naJj5IYcQ/iliZ5vA
j0+QWZY6wBL41E6lg08sWMHcFcXAV0lZ5iCAn6zACyQCQ0EwqCQkzd4hl3cXqB5qHgQGfBJ+L7wf
Vi4qxKolA+MRVlN16MXm1t654BdtZW5Rd8OqKNh4e7/vajUJdiobHkdAo2efmAdH6DE5hWM//Txz
zy0GqWRyCP60zV0pmLmdYR/xReJ2mFDR2vZyWgThLGPbpfwhqgiMw+yhZlafJ1ShKoa7C48WCKR5
DYlqgnsWc2mBC5kFfNmfhqW/5+wlBvh0U5bbQ839UmtHx2aAWIqY8hxZXjrjLECiHcTC7JJWTQUA
gIWtE9AiosbKfZDrLCJQotaofABU7TqveKJsvDUuRgHGC0lS/9NYyNAOY743Z3V5dfm446aDv8JN
NLqs+u3vHFy+IIOzYs6oAcKjzCH87Z+MBVYpcSfIdHQpFnA3BRI1tRR8iW2lEVuC6/SixIvymqnX
a9dIJJwpuVtDayeSrY+FPBgbJccQ2JmmU0EibiptSAsXfBvsay+33DeU+3szA9jTv06o6Pu/ABGZ
LBh6BlcXyUkBwc+iEFtM9EZycgV4LHcji8/MauAgM7nr09H0fAzjv5R1gzZCs8TKTouZg35i6Ac4
xf+Qcq8rGrYs4Coc7cc8B5QvmVG4eA9T7miLfFT/QarSsVt3mIYWgL0fd7as+o5ag6GhuxOVaEUN
X5zNN1aMZwZ+z2Def5c4f/MHbYVw40rsMSP6TY5RbDxZtaKwret9BL82rWoxVaPnEn2kLRzOjQU5
kn5+nTLgrH8ezTjm1oJqNzUPJFSM+WbPPPL6yXH5nlmN5HFOZfd6RqEsMwlitxS0ScqaLuLTW5yA
TIT+cAbLU7ec/CzVPJj12uEXLudaKIa9uChpw0T4C+k1Jfx2cJLrSuAr3yYnV0/gYXkR/w5gmYo0
rbYKrcyFoM8FWpcP2gpSoG0qGTmf6NhlcIojQa25uDBc9mfPrEFU6NBkFR+CaG2cnwoDuADqUrRH
4WVWhzRfxNH9DhdgBuVaYxiBeeDecS8aD9zUVELZMFOoaJovGrQNUzI8yJgMSQtwQMJC6igCZNw2
QCJWHgTkVYgeUySd3TDfgek2rUQ6Z3+Geml3cnhfWcTE2oWFGiNLet0uiuH9znUuUbByg/EcQrhG
y1QO9OnYyn3OevsL6MyORwJDf0o9J02W9trdIzntij8qtdaZVBsn0UL4pUfEx9liCL3e2En/Kr3/
GSqW9enhJc+L65a4Kn1wldqBZT9P8ZaVTBHC03GEheV88x6Ix2XLP9Y8Eeu7W+wKrwsAVoojU2wi
Y48hk/oTfs6/GTCkXE8kus/rEJJaVFJ+9asikhDTTaRbMKoHvRtr2ytIms56Q3ZHOj+k3LA9/Skl
9es7p5UOdC5xvrWAiiT4l+2ghG+w5AItwdlEnMG5TM1gy7tBPXkyA+l+U67Gwv1hx9QGXdb7SDuB
mFfZS3szmU0kl5BfW0NyJFauQt5qV2ym6UyK0hI6PYpkeqYdK7cY4qKN5E7+KLYfG04+SoWdtn1Z
+XgNJMlqoRhfNh+/eg9jc3eGeRDLtpAhrK5RRaN1MnNpyZ2VuYI1Wte4phpokH3Q9OFwF5XI0FPV
ZkoY1PERjH2/Lb1aX2FrJndqY52s4lRHcNFJzIhWrJatOhZHzftT2/Tj1SIVKzmWBiXk0bWteLH/
XhyakgmrqLMVgDN3qaXkxZHqEv1nyLBXnvrb7gzaBPpon7kf6s5qD3v7gg+/Lsm11EWFZ0JaR66Z
jlsT7WghhmmrFBR6Rb4GB0qxnp0IsuzFhQ1cGoXz5MOff0o9yxVQAkfRB+ajFMnj9ROdbKNH5F8l
Tc004VNWIGT9xDnpLyDzOgGIjRoIPwV3eR0FTZUJWRyRdsiYeEFZ2sCYDKu7M0Hgk9Vk0ILziKWe
/hxe+Vb2KqK9zjxvC8F2ba9k1q0vuaeNQ6OwvRgt2Cd1Rtyd1ko6dOR2V48ge4n2FV5/PhtvCC92
AN2vTpII2CChl6HXDsL6Zn7a2IhQUv5tBiiKiidBecjCVa+ynHr2TBG26KNaJ5Td2ILPtIsywrWM
zY+VKG0a625ciTKoGd1SPNRfIBa66K2sQXTVlH8UuWcQbYlUdalFen18vgy0K9HIDV8hd4OFOKb0
gKuZTNRVOAm1RbDeuCLiZ+PzubOH5QyohyXgJEB5verJKOGECSiGny8YmCGxY5n/+o9qCE+5D+wv
NfACjqPX2KQV1p7jON7JuozGJuz4Dh+3ry3N8lHiddnJLmHYX/4Y0TIUDMeN8Z7d+vjD/RAfVZPi
7VdcxAVZt82YpyaUkDF7vOT6DCHHwDpLNrI9BqXrdwQCd106U3XXlcJb37lHvARzjeUZl+0CB4sC
piJZUh27GhprgsEsdZ9Y8UoRLT2IT1tSS964MiHkjWqka+6BJah9obk6xDr6zsfLi78iQ5VkNjko
oEHs+yCHkotQauqDeLInl+e470vigpTyf0VRx1/OnQ47KkKoKaT3WUEyCdhy6epNgSwyqRplVqVJ
h3YOwvhUCOk0m1PeCzf8GtI/lxG6BDXxduQJ2j56uEOD/jtOnyF6f5rZ/aB20JoQTlXDykYX/vTU
LBNrT79qoF5S2tj80xRkM2uDCDS1EHSLzrdmqPoBmf0IK4c/y116EPReIFYG4M68HflkZzOQcZfP
kkmG/C0Jmzmw6/Nd128sBS+rSTSsb8qPQEMPzcsprn+5WvVfs5QYEbXpeGcugHflZ2qKcg3+DLJR
3pS1E8l1NJoSuJ/r7IWwR7AfKBT8eWVz5VojkiA2gcWtRP5wVEaizg200L7zUfKuVe8B5MURea9K
Sy0fKuz3+YmiYqlRC3MhPXkSdMxnx6MwmFDzspkDdq3ehomAi0UnTjhtqIVwMF9JUtih6L5yKFp8
5GxP4gILKdi8TC83m4sT3Z10LmqysmbOBYUTLySMnOzb9OhP7reWGrhZ8xSYm0IRZ+trU3b4sHeN
/KDNW7iIXS7yKp1/9h92vxg7YiYHicYH6HQE1Qw4qJbrnOCPMFs+6BN3gFC93uQfly3hh0jkDhWA
LUxsQ6sMJlgSCig0K5xOmHszml98FB0aceu2xgqghYKha6J4/io5vaACTJuDK/jbV/BjB9fopIs2
pT0sQnr6XdM1/lThWBrDu38lz39fZxikCZMoSwVvOZX4Hfwix2rzy8fh21aGD2p3tSCUmoCWOi2b
1myyYXsTIDdZmbbeddrWuTFzJYUZ7/k14lx8N07VMmnkVnf4HNLd66XFGxYyNCNia1SQNadOHX2h
/N3xmLtUVBDyw5z9qqWMtNJu7ceJkeXw41m8f8hLaKAV0zOO5tdNdfMzQ4LS+n7T2xwz1JeZrOMq
Ws7Mxo1Jp2nG5ituP3Ti+PcVlH7AepcVJkYubx7SIfYMTM3rVwod6y8+cEq1uyH90y7u7AwliPiU
+b0goVdMP709uPExhqE5b4dsJBqaym7RmS5z25iXoksfYlcdXpR7ub/kHtciaKphDCmhijiTHAdN
dC7WJTY15cCOGne5xvijPo51+wAov1CfKCOn2G0C9OzRPyuvxaioWiMs+/M+nzrF9uT4RAVaaSIy
xNVyAgTYzKPPZRl3jDXOfbH4XrBCN3y6pYnoItedtZ5aa11XtgU4ojnLd7dvai0lVgwTGw9R+3N4
eAR8a80+xEtZUQtlPHg7/pbYZq2be+68rdVEX0VI6GQjJzt23gF41BWSX2jEsEfOL+5yBNy1Q0Bx
DR+FDdw31hRbsd1UczI3fvOsXfrEdbKZmyA7hOkJ9Nil/IcKaAx+HozFYf74GJXZ6neoi1xMfqqV
au6UGThp+ahWHhtqRBnn3TkicerlWuLDX/eEIOotCCwTXZVqfmEnNpWGGQFpZJNu87PiiVIV7Fj1
ZiOqL2SlYwteeuHfNj8JUFSHAK+39+MAPwlX5Nhtyhkw13h191lPQdGeD95sIIyBNY78AJ54AZa+
ekg2B/i0nCZaGVGHRiu8cXGrioFQYkJd4AmGe4Cbr9zzSxuKqUrHFYpnITR42xmk9zWtVBQqlvzI
+jom5Ra3D/lR3JiXZiliXwYcD4WSE22JK4bhpZSqc81crbCAD5kzfE7YSE2orf9agAhgu0b8FjlC
zEZ39iAU66r9s4DcFyi8kpXOKfysSKD75mrHg2hsKvwsFpJCYk14KWpQiKyspChsIpcL8W6QTy1M
1boowElxu5idVjMTKtWkMeSYvu0Jbd4sHURakyK3vXVdSuUcxNwFahDQoFEAVeP9T0CDZ/fi3xEi
UCxvgw7VSXZI1c5Je68Sp5hYvgX9D+04IW/rq8H/bUB2Xvz7Ca+gvOrs2M27ignG0IaqF0mOJS6v
rwhnwipKvE33LoPdAbB0RCku73hUAMdojumqKvcCaU4lU4cL82iYYSZxKrMySVV+4tfVmXqgZd/z
3x2QhvvwFOgRvFbC9TjBBiqj24ZS8RQlQFtQMiUFfNaDRLoNVa4McraM1EjT0d2oGg4VkYpCJrmc
0r7Wx8F5T4d9JecANdngFEa3EsN7Mp9OWCMkMtcfUYT2CHYXWjkvARmOVnclqw80VB1FgKMRZZkX
iig05kzjk/15OeOnUTN0d99Wswkng4Ecdrw35heoNuLqabKrpmJm9yBL1gDTNik4OhcZqrTrAuxu
XC3jixfW/eYzp8eHsKeyqoqWsIHzurgJOFa0tT8lSwnsikNsYegtJMM5XjB5z2/VykEavY6bsK04
tEAfCW0QFSSz6cFkj4nSkBVZP870H3IDKPesFd1nNaZnCOPbWDHmCPSyqscJ+K5OM0uuAte2DXqj
igGOCU8RbE+q61Medl6Wdd4WBT5xkOSDunMWxEEVfkg4MOx6uAMwacPlJIDROxujDAplfCW4Ow/B
vjK1HrkLg+E71/l8eYPMDEGCfFQ51rcHbC6leaubyOjoTthLMiM6fP9dZuc6jB+5+lRjNdlPvmCy
r7kl7giQd5FpBhcZ0DT3+M3eWDuSwQCbL8UT21KCTVwLNg0/xEnaQx2TtEn2hxxR7ii6oWLFsjC4
vrAJDUYzj4KUy2Xoc3k7MckAC0Vwd0Hbm4CwgvlxgCDgXyZaY+iyunw4ukVvyCG/mXsCqIDMOInG
thhUkER+dOpkEKVIiogFnfDC8Zg4bAv4pUr5HITG9xA6hoo8PcbvNCwzI8Dcs2KviPwwIjir+mZo
rYdQDIzSyTS8LmVzNymFJFhixpAqbpp6o7OiY6a2p+SFlGssX12XWCrSsZRkUcnvirsUL/Mu2rSk
F1A4572Lf9aMuzaXgsbrH/R/2KX3BKi42UjL5zZ5yu4dUrtQxcqOBVhBWI30oqaJRirAIGDk6OqF
hrZTBN+WFqfhpJ4b38Z8pKPyTRru1LN+L4+uaw3NG6VOMHn0gKf5y8y2u88z512nC9yHjm9Sb7km
S8AonJ6HNW+jvMGhFd0UarOzLpbebEL18dQd14c+zp3/dC1E7PVt0Yv5D8P14CiuN2eSLE9lSG/E
9eA840v5GFM0jJSp3nyoRKJJZEe3DLKaTAL04DwIOYrKcABdvaeGmHoaRuNKm9mTY0zuvZjL/jam
HZmMOKjiFgORRmIsp8CHJBBKkQ2xqw+a06jxvtCArl5CQz+2peE1DP4foaFsstoGYZQjEHYU9ZrE
5guo3zhBuYGHRfyM0/LK8/O+5SzuMIbPu2ARPHCAZ9l0pOXJnfS98UtnDSi3DXR4gxd/xDuxdENq
AaYqvC1D55UF7/M83SkoPJLMKvUYak03mb4XpFLQe+shHAAxHtPrYwC+y9meECwZ/qVt0+QgHgVi
DnvBlvJdrYmnjl2gazQwrrvYv/61lEhZ/hK3XlctN4pxxLRuIirpyu9NzkcSZBozlORCAGcFiown
C75ilY6KuoGv/k+359HhqsprOsM2Z0nt+HkKvqPO6WetW+NeN4U4Yv8c25c93j4NJzawLc3Ma6bP
wpBM6CoyBzxtYCjIv94BC/o+Yr1RTYwj6zuxwTKO6yIMb0k9jRxpxU/WpZpxfmoI+gNE0mva5nNo
hPBa8dM6jDZRGGO1RFH6kwXcXnxDEHq7D9jPAl07Ek3T2bMo/YIo4HzUm7xCCOJzLUaLGWB8GRfy
brEITWjIxDka83DRm/RRmBY0CbBJeMX5S9PLOzdekM0LoM9X26swxkzRD/Dsfql6qoF6KpQmvizO
fW86f+GmAzHXTkGNw3mhMayAvhXd7UxBhZyaoX/C7XCcDar/i6t/5T0Me5K7ejMhyq9vZevTFnIT
17pRx5gc6Xn7iHeXZiv31CEiXsIWE1R0CafPLgkQSRW6E6teh7u8csoqpF8l5aBw+m8I1FssAKjG
DKnTJAG66qD9uFjOJ50lydM0lfGR8Rvso/iJ+7oUFornS4aHOHOEo7m4G8kevWMc6ttZzbjci4fs
s5Js9+wFfx2oVaWotkIiWfcA6kRjw8eMGicjAROl6wL6kIQm5rMk3Gc26Md9+qnzyUrSuNpmBdyo
lszFL3Rn8HyeJrJb+qkc8PROpcKSVXIk2Xh9JBEnpNDVypdLZc9RTzIwI9g1XFXfNV/UFlZeNcj6
Hrws83X1ySJLl3tzhApQDlRoZjcZQSzEvGsN6HwpizAWgUWX6OngpGg0Beb+idvpO5keV+3PkQtB
g+g+VnM8BBaCTPyMr00MTIpe35NBtOTB07vbPZMZMv9kRqPF0hV58cMBvocr1ph88b6/Wbh6eFxd
3y7XVurZPSq5k75uFuDXBvoNWXgaVkUytv9bFvDELQGaUwUOUHf18qJxFjqWT2q58IHnND01udfq
S7BoezusH2B6Co87Ptv/cuZka89whmQ9FdJRLBAoD1v82WC7HwTRq2d9ebU+tPrhn3Cmqo3/yHNi
xy43WnKHJ2WVp2EM2IvZ4k8dzzSyVA6elyU6ZSaM49/b49s90dghRtAnIQaJi/IJ966DV0kbp6R4
VVIg+cx8RwYY1xHViisiKwTEMvsm5vl7WblLbTzkN8GOo4YXgrkYkEOP+NaPBfY11AUrkw2rcTIY
2A+Ah2pCg66LUc3hYKrhj0kY4G7ZYKUgr48hEWWSe/InqWqWlXZciBKMGFALwWccqhz2rADS6l64
d43fB64VBfyBuJBJnETXRBP2a5cNJL/23LUnUVHYpuhSIsmOUkYIxjM0GPXbPiG477i9v2ktzOk9
2Ve5TBSCF6JwZaaD3QnkLXQYrcPV6hkX5ncdml7WeOudACV+wRYMFRFdFiAbU6apNsFNmOfy29NV
tqWLViHbKXFQYn4RvS2v5ICz1G9+d6cKcyLpmzvQL+IzJS5Z7E2qlGOYcx9K1fDTsOrTKvN0t/ij
UuiwNVmsWUBE9PccoWc11lwWC5ngG0vBaKRkh/qVCD8YCeK14qoxtAqIJDZDVMGhClgFpTgkx3qR
hjHAyiEI7VgFyZAong85L+2NDzZu8cex3AChC7Gu2qgEdm1+ObI6CV5B94nUAuh9AYc+GLtzGVe8
/+0QpuR6e1e6tl6t2sCbCGdWk/mBwu3D8FhD/iiE/59T6eWDSoE9hpaRdHfA0FgijF8P2I8D7g5L
+UrHugdy+gGOq5PnxTnJqaYFHuhfFL14RaTxQxF+vLmasbWsypaIS1/kiW3sj7Plhz8ao7kSquL9
nAnG9wPGf1A47Uo0eL4c3YvmYSH5aS2Rs+ZII+BIz/Nuli7X9JS4vB5i8+OXlLFtxm31m2Gk72sv
yDXFmclSwb7XZrKPDaxqZSETKgm9syFa+1NKhgzr7tsl0dGOCMIEcGOlb4zhnI0U969mxaUxMQ/h
uNtzIFTYUYYmbQ7fS78vCh2gQscqsBa5LI/u6f24tUCm5BRtXjlYjWa5+xdUzosGp3GsddGTC0kZ
KPJhNZPCpueOsHGukz2z16CeJTbQm9oZBfaHw5895cPI3ODgiFMUY/+RkTzJBP+8ZG8N7iUYd3X/
RHVSykXI/mF1QY/LFyKk7xQLGuQjsVmQB31rhJhlh1x2aPhnVlrvZVGRHsPqRDs8w+yesmFCms7C
6ycoXAAHR2fOyqVmpRzZTf35Hxf18AbFozXtUeypT9NFXaiBA/wl+OJwgcTf9UZfMeIARPqR2n4N
bdpeSXxYs3UoiClRgX2DK23nILQJn973VPouATF2EiJMcIL3ZulSdhjfNc2V9X9eF50jR1Nk96/n
MfJU86PB68HE/7wVHAm6Mljz0XV+H8GLBlwm0fMD9pGngYqoMjKhTWqBVDMFeCDXf0GJ7vHooIoh
3bUCFEq0e4VqIN55kEYDungEpj1Ls+Q7hvagauHYNtAzee8a2M4f2RTaSjS6Srl69vtShes2WAyy
UkZEjTu9ZOrifEWkpWGyE/2AvJT8CHwcy6ZCuj4leYWX45DekLNiMLRL3LYbKF6ONZ03BHRyRL/4
AJM5DVIYUAkZ7mgnwYXhBzwpCsYQ23ss91CAND4tte7cVD5huPkBQY520JAyBL/pJYIl/Jfo/VaE
76Vgnbh1UVo4o+ZNG3ET/VvrN9r7+MxSx9hZyyxPWjBRXPqNZB0vlMj0qVZVc8Ia3YDz0KZeuY1i
UKmd1YoyjLTRqfCL0HNFpRaC4CJ2BZk6R3z0GevpsLvbOD7TCy770addtX1p15UHDMKllAacv2bu
iWy+e/97SlIzLD/PA80OpI9YaQjLumndu8nTsBdos+WTgMyF5DC6m7aZmhdfzTvxZLar3KPeMsXy
m4XzuYQGSTt78CaJwVEK6imX84L4xHj8u7/AkkjTiiEYRFsoog60fdIZ9YK+FkX2LzEt41d3guEF
4g/b4kwhHZTD/+n0rS6InHCvcsWFpweuLh7gxw6QfZ2zvA2IpXGJoct7kL/g2W3RdqBG9XL1RA0w
WIYs1VWgzvk8LX3thvGAThQOWS9/YFM8E0IvyDzAhPB+8mJpflkPZSfF5NBDSRNAPK7982HCkZ7N
6gAiF5GlntumpWPm4jIGoX9RiLB3rgnhm3D8rfcCbtBzSl6OUyBiBS4OTZ5al8S5dL2LgDgNzB2n
grdp7FExH7IsCZ357UGy+1UB3ntndVf8cb7gKf5X47CKl2qWBJqXUwi8fKilSf6BmwEuajbD7ADn
slKwyQqFDEaNypnbzV6WqkfI+7tuln8YZxY4aKFQAVu6pgZBqC8rvcsb5pT73HTCtpB2vFKA3Ewg
fVO6Oqm8fW3npegEJaxbyCc+PCOCK5ANUoVQ4WiG1jP1A9NfzvRHeILC8s+uqgJqX/yLoTyTndEt
d0is1KwHt26oS0KQSU2joQORPqH85im1x3G8hXhJ+Y58O+3VKfHvb9dRkn+oLT8G9Jf6PjXYFwsW
iK0vqWv1Z8jvsb+gn/mtWV/O2mI9Rb212keCRbgDaCHvQG8EDp5b0ewzQfINoeBX6rrzGb/LaN5z
AKsm162dsiCQCaFuJKXWg2gdS4+g1Fiv8Enyjf1hro/OmGYQ/QBKWmW1ehoJ0erds5NWclDGM8hy
rKw4UKLR4hwKaNqbfIRN0se0hAlZ1TVHp2fMsAtM3ATXnqvDNWCz2f50ASBbvc7vYiIuHQsxwc4j
RwO1z2vZIqZvMpxWoXgll954UpPETDeldjFrhxPuFyzfRzaQ6keXV4vX88ouL8fsdxIbU5Hmiitp
phRGp88v73TN+Lq59E2KFCNkdWbyHLe8qy91EjxEpQ+9CcEOFs39iBL0Rx0ZKB6NX3facBmD1t4f
kW+6XmSTMnAMKqS3jXDSTc298QI4FCS3iy2qH2yw7PaPObvH4oUpf+ugcXpS+WDF5FI6Ig0OBpnU
CTMSP+HPWvlbGeMmOK4ND8U+XiKuXDtBGfgpbSACa8rDmcHRtSxb68d/JeJ5CeyYw6bcPYnKwBVX
dcLGhuBd2yk/B8xjtd+ql1+XrQvOUZoVX8qu3w9t/3S9k5iZBAB0ufEEavPlASG8dNs4Gga6ifP3
5n6Rs3zRDqXIs4NPUqidbb+WY1GznAq6rZ15ZmorF6W3DVspThC1NY6z57/lpEiqpDVAbgBDSX3B
HYCk9aLezCXIky7ohMkqDyfPz3LvbgoQEssn+1ocpc3o/LMbOg1dvLcq4yBTlI5y/ypX4WX9xmOG
EAqnwLHZjrg9x5G1q1CsGCWmcAVc9tDDmdkjw70Odr59HnOq9yTkblqj+ehwtKNQbtYZIMunFmkc
/vItMIe/Ck32f5g7XumGXpPcLjLvzBbYp3A7HuQREEYoC5f+8rzPcPSvcYLrm03RcPPnRpszaNzi
OIfGofapqNk94x8682WOSMysmTpl7LHFG/abZNbSu0/1MdMsXvC9mkTHRxbF1g3OUFpGvNdERtqU
RDCLTqhKjuuD8sdL9eNHzNemxBF1yP4th8ecdJC0NnoNGkntPTwDtu7YBxnbjIolHxU7BR/Kpp0z
N1lsct0Nc7jXCb5IyvTvRkgPcE6U+nnozP9hUtP3aXwdnSpUXp7RoKMrzsEoZtlDeeGUY01632sS
Mi2y3DIeTdsvDYuJ7nakazCpFR7+GDyez+wZ+/NJxG4m8jBUCG5M3O4HKG1jjL/UyyXLh7PU1YH0
h58xUyUpKL/wKIzgl8RhnrmGxsFn6X9QhDxDPNhbFNZ98vdDsQBmDsTA46dUk8uVMqbpBGfPocCe
kmcGaj9l878Jj7EPc0941SD6ETjPeaTGEgtjku/7lw1IJqUmp0wnLKJM6vxhL9PI8bgUzF/acTFJ
jVKQc95qsqJgXgXnMiqnUg9GCbAAnGPedSfIfyuiQIGnfskVILuabNsAkWWJ7Q0ihNBYk+gcbIK4
d3KQHuoyWqSemkLl1sreKjZGcPALcYSmzjmNzhCiJZI2/gXT+bFs5RUuxJJtOSj6uMAXuEyitcVj
BMWnPzeMH2GoY6i7mzRI2ccRWrBRVd91n17b5sFk/qZohYpa2Y9aY4ioi3sbHFdAm1Qb6mnE73rY
94IqqKukIEm0RmO3IpWRnAS9tF1msQW3ywuIWDHDRAwPXvn0FVzWAYXFJJhswN/lLBb2Qt9AVTaf
18MubYGPNXxp0OP3stYozAkJQOm6LQTxsTyUVWWpGMVeHwG955zZMj6lcqJMYzZukOx4b4gjDrzG
FtJk0lg7gqbZTBwo67tMh+7QUi1rUO2YIrKplehx1yxYWeuZRyor717NywytEKzg4NtVrVUobMVN
bhnjQ/G8fgy+MBfqrytWGGlHJ5iZ8xVP6Fk3FTRKTv4B02zHi6Dfld6Y99Ga2dIBtfIKNJdsKOth
NhnSnPpnkOKk51EhcnKoiH0OV0/vO9SpK7qATjD5Vzr/hcJHAYEIPQZlQ2iGMLs5bbtPBrAdCPOf
wz83bZ3GaN8PriBAvyqJMfGH/RI6kRjPFdEKrQNXq6UgTidifU+JTrgNf4gJUXBrw18aBUCloq7b
O068hT/5jN2wPfTD30/o2KMXa5cR7vLAhb2GypWjOwgAXwsV0c7KzldK3Qm8L4JOpXsB6rRkg3xi
r7Nh03rKI8r7x0fHF2WKgk389mgWhj72gX12jTdaMxFvODLfJplLzN3AGnh45wSmQ+t/XCsnCWyO
OhalQZLocx9f+DdWyPsdCgbyrWAc9zRPtUqXFfapzcBw4WwfZW8dWSYLkbHARCjgr3lHFUaHthwY
laLxyN/7MIaQRo6pPMuGjVOGSd9mGFEhOFfVbO6p5MTc/I20NWoDI5eYNesVJBgrh3gb3xdQoC+E
ybLcrQo5JaACy1uxcmYxQVY51gNU8TPfRU64TrSZAaJXLzjPAgxGMOWDOOIDom7kcKZnRBD+i2Ki
jV4rqpJGQ2TwOs8Slq2jeLXHmwpiE8TNcLFMQnLVan6hKWhMVxE9cQGBvja1jv1x7fYUbc2AYquF
KOST119/HOnvVrHcbIZE2YfNCrlp2hnmrTzke9twi91WWspGOG/FnqFuw7yVwu3K5gKVU54fiJi3
cy56wBtuUSn4gfE+8xiG8IJV3NdxHgTk3eWQO7/qsMs/GstZEPlADpIZoO5ggcIa/UuF/v5RicNc
y7uUubLb73zaUY8wsUQ6/tFDze7S2YWsKEXNDK5LINfrS47Oe9mzYKAsy9R1YMSfIdZTFQ9oa04H
vNx0mRzjom+HyPCGZMpXJC1+IAfaWlHua1Rg6fg6HinapFuO8+VZOPeYZFJAJhAxqH9//QYgMnUj
LwXC9j9ffh+tbt9fV8DyEjIOoiud8d4L/jOnF5Q+VuWtqSXMk4Yw7BYkII1RPtImih+u4lwJl/aa
tSXzq6vzla/wVSl79RkyEYgnfRLsmBX1DeLZ3TWO8ttEJuAZzFO6JlyuxxiB0x3k2CQBPGeoyiXV
MoHxbOUbIMJnm4FmXc29NTME7NDbA85RwTzos+nXZeKc2LfqBr9Rgik2PTsD7GtMh84304M/Rvix
mr/8l3ZAEWRqKtJ6sUVAivW/7fcbTdJYlILZ+XDm8jkOkLTx/NtFbbo0oNKwfuCojvzJp62fu0GT
TU6PtkUvysk6lRWGYchTu/z+GzVxAG6QKcMZFl9gPXVRtNjJ0YDIHmSk1SXp00gEFbMJuwT0HXCr
FRvio2yR7vaCTHfKfz5AHtmoKE9JsesjtU/Biubyim7tQZIOe/ihRXekI9ncE365TYl30l9/oMg0
/C1C7gIrQGF1iZJFyANEeLXvlPQtkPFs3XU9L5RRWLNiPap7wQdvavVo0RYEGM0tkTh3NQo4PKDw
HLfJgGJprXKXsIhEa9RlX8VILuYkAnH7EhiEuWA8D+8AE0vXYi6pWzB7ajtwvh0JzZvY39Ca5J1J
N7OUujv9gRnVrQev0zh3dKcprmEmR2rcR6T9ImW3Wm/8nWm9urAduOisJA+KLL1qX3GZnN8k5zlo
IlzkDxHt50NQjM5Ow6VD4UywOfiMtxRwqjECKsgVudHH9Y60aTuIuXO/zEDB/8161DTXb5wXj/y3
EPIoJLVXuTYq03HyKLL+nX0aqLDwrYFuq/slO5pVtSutedkgfgyZBZx9Kk8z5Vmj5azyv/oxwwLe
m1CjXEXlklsxCfWmkTllR8XzIJmqTkoigZ7dTcXudEDggni8UyERHLb4cCtFbPvK3RL2Tfxr4Foq
ORgf/cuyVUA4e01VnsQh1f3biXDtfrahX9xFnKtB68vUiTqKlnDn3ol4EueQAIaeK8gGxPnpe5zq
7Xjw7WxOC1r0QdSazSgV52EcIhsI31APRcfLj6d8L+Vu8pFXhCuY/shWo9bxZRZgWOFYSWmfWk0E
20mHoVupRbweA7Eqx4iFPCpVxQtgOayqIa8Zz3BzcedrWby6rLbU8hdhm0TcCRobsq3HIghb8+Kz
74pN2xyvOm0abmarwQSykYli4RCS1ZNePBTQBaFJyu34t8HIUmKb7LM9TEilCJKw6e7geAERjH7G
2jmoRSkBA2VrkEIFKAi1BUOwrtgnlc0r1W+Mr2WccPoF5h+EYohnFJboncpiNuc+oc+aomt4bcLI
o2YM/yCXjzIhw1bvlPMTHXfJeq5WhW0GNuanKGdM601fFGQ230Rvr7B+jJzhhwwcGfFI4BLtah5q
YcuVUapGfDTi6nnVQnb+Hp5znJar1gQOKYBp/cLCATYWcRxk6viTgcxEJOh2KO+3rXj/yiYbO5v6
gVeSNkL284j0Zh2Kx7TpaHBG/SYdKIpAW63WfJGmRH55L1wilbZT+hEeyMxKxvV07yAA+/oYitk8
FMzyBzAC+cDWC+2hEE+b0o5UP9d25Gp9MWbHIP5atPhd+V+uwwQY97E4ddyZuCmwestuGLIhR0QJ
PqQwk9MuWozRfYwk7yLSIh6d6UoJ3SPT3525xjdv3SADSHDMlYfX6aXitwAcp+06zmWhkTvhYC4i
+YpO4BDv6Ef4xf6zwGjsTepbvdnVPZbSbBwkrLA6Sk1pLfHhWUdGLYg52nnRLw+UApvH8iuMUxvO
KfFWV42vZrn4jkThRZBJdkiIlKRZ9SRJaQWPm/zmrmrEL5zXtpNqx2XlACSo02UPi0Yaehc4v+zO
9y83AnTFCGZdIhmG2P5lsItINYqy1fZZNOuiaik+mBrMbWFowieKsrMd/Wa+EX2xs3lg5/nILDdU
FRuUpxyn/qhc2rPpMxl7GC44ouUWRmK5NgHPZQtzyQFxTX8bRsCaya/EWrP+T9kku4hwY1BRwbG5
8+UlZVMiaxi4+glFjR9smSJcddoJDOPXYxgqzoyLP8tqWLxqvnyJ51Hzb98sIA6L4UZcHjo+kttm
CHmOutzrQ+Vmmg1tRHUVoyVboQmZQxvZn3UIu8iZKiE3BO/FIWGBfUBnBbrvP9guCjag3NnzGINv
It+PQXChXg9XXxK6Y0lbJjYsthWfKiu4tdBpcA0Zoyy93JZK4wUp9wxMRdSsjD7JzVIsqNCjzFte
/0LRMEZQUivrOBYDFmtzmRa3EV/HsLJlrd0La1BVaClvdI4MJx0PuXb/G6QgD+HhzhP97ey82Trk
UkaiL5NKFd090KX/PWdp8v1jmGOuEkBSXzYLhYvLENrhNqkeksmGU/+ociOh+znzMHmps0NFK+Os
nF6TJfuCQBFbtbxqTNQSBw83YzgDHA7FG1I7AYtvb0yDVn5NfXk1x7yBHR8brqBcqha4lzZxsX2i
K86ze8X9ID5AWdTUIEWmCwP/LS90itKds4ca7cjXYxEQ0brBEFtxyojARilc4/M1oqEV2tGLnKxp
GipxtUVSVVg8d9LVyYIoYCJ0WBoVlX06P5IvJxL35ThxzKRHbE9Oj2l1Lo6PFJzb0gsL345Qss8L
lFH0KuZCAaj+M7sIQjYsBg0SOEczVeWbdtShSTsHIYrrPKWRFqXoXEmNtDpjQ5PoR3j1dyhy98uz
gw/Qen13ydhlDpgjNrenWz/52oLE9l4+jj46TR6uLXFNKj63EHGSnyDbhJnGM7j0vljMnHc3mBGZ
zitMzf9V27XsS8tAn4NGSti/NkJX5X4NE56gvKNligxlY//eLeOfzQBndpDZBUsl8p3MtPjGXdMZ
66wPKU47rKQzwiBQknuJym/xjblBgVdtLSyAFKcd7eTQLyIa58wnLPQa6wR0Z5F/TaQPcUyeP23Y
ehbJKKVNoFOJ/KDufXHGwMsPPUxrS0kpHckFhmGf9zd27IF5zlLNvdl7sjRJYaS3rxDnQOxf75LP
2rq3vWFEO5sZrxkylE8VKNtmoAN8A6VkWAWopeWtGRCDyAUfppNSSqrtzfL1zXzqhqNhY5Ujb8+P
5xjHaoZEEXo7wVS8Vgs9u/MXTaLZSIY9OrU3eRAXF9uaQB3zETJD8gFbt9WrHbnxI4ZEW1ZjOfvp
zrbISrIJhZ0bljD5fIU2kI0caaiQ5j4eL2R9yC49RbiULvooKcAzJtSemJOAqf1pAwsruvlqvEi9
L9lknNh6oD5qynjuJbwPfuFaP7it5nYr71E+0/reVzkQqk3hftBv1W//YM7jS59xKPjE+fEtx0eb
ybZx5eBdYmrsQei6QvrTM1nqpJV30CrAWOHtoxIxzC+s641+cDw8or6GCHP/q56TMMp26Bh+MkeD
T+HJlPVgl9Kfc8Db+s8YtBh+oLnt1TCASOLw2Wwu2YdogD6j6msFP8RaFgbjFrWmvdS1SK6oWjHe
lWy58dSzxasIrJrm0uoRrlRzf0I6mmXOwuiFxVxy36wSvgynmOXumM498sd91GZ/Nv0mYDxXCMmt
wgpyhNsznOPyBe9gNUINd2rsjeTih0LN3NrOQkaWx08ZiBRKWa0pDnoPn9geUog0crRHt2YfFBDS
iseCkL8uicaatc+Ojg9Pg6VvKsAzKzZc5HUnWAEBz0RfQVTc/euQ0gVFGdjv9RDQaZXkP5gznYUC
AuoJ+z/SjT0YY3Wf+kV9Vkp5BmLJe2Sdh4fMhbeNveL6p3it2lUgVxA+GTrqPnM5r7y0besj2UWf
J7osTGvfA1E5ZXvhfvr7NTpB9bOcTlUFlBehD9jkhEnditMb6A0o58pmsU5qQxaiENzLMe5yG4Sf
TNRHV+i4hmm38638k1QW7VldYMjbl7YqGXtudIvjVUBEdwM808UBv84qW9Es23DxMjkIWY0GsVv0
mUhWm2wHha5ZJHj/BmexoVD+R8hQdR/mIUSW12T4I713aYiTt0w3yhXRXynSjR3SQP7+kFvsFumX
39666WmnA+8RZzhMXwFpOk0wteYBYKCG4+gUZRAzIvQ6Jsv52Z0RBYQcIxYIDMEJZwTujE1VlFwa
gxGgfQYsOJ4C/0Bbk8+QdvGLb+3NjOHI5Nt1zfeA2tnSLOSEBDLo9OBU5ncS6CNZgSqlCu7Sllgv
EYVUkgZ+R2Y9SuVlBM6EPZAzl7isNfDDFhgxhLdpztFDefH1v+b41wKENLnYYaDdUt5rU8Dl27DY
VH8mmJ54yWpPL0V73HcqpRLHu69cCAN6sVndPCid6KLdsyZrR5Avr7sc2h1+xBiyix9WfPRnnAIh
bieKyTv243+aeBgiQ8UxCiYgDyt0DEiGBjDqb1wwNDWZE0k/VTZUxRNB0KwSXJZDfZl2siFaqodH
K+JwpBG70aoeTObbAnaAA6b8MEqGgF5GgK3wPF+t6yPlxCARKMC5INiK5Ra2bqrsO9HHV6eDPZPi
rjo3w01Kq9tI6Ys+OyLJg3H76mc3DpTXI//rfofhT4pVeJs6+4YMZ5guo7zpDvnobT1Nblky8JvJ
XB2Srm3OYVPh6n8JaB5j3nCk3tLk82WqXR7d/V3pQiWqhRJejfFUHlmzxue8a7Kd7yD/qw0eorvp
L1OWjiobahA4TK71w/A809l4VJmQ8EvnL73YyYofbXr+mKXnViSkni8Fg7cSKUsmeSGXcD2uu6Jr
H3LRcLQD2A6KRe2dsZtxbzQu+1OmN+FbedNmPUFS1VdkRB2gj4VbN1It8qdLD9zm81+l7apTl32K
3iuNVdw4dwqL+PNTVoE8CYZhqm1fZRvv5gBczQfDY01QrC+kYG7aPQZ6Rz22bgZE1dwTON9zGwVW
ZeKoMpy4o9feY42KL1vgwhHh+F4ypyElygY6Ma33g7tiEFK22CPLD8/7TBUy/dRTWH1vYOSu6J6i
8M4lfg50z1O+ySY322rG1EUfnfbY+V0F1RImCJ/fX4f+2Boy/CfZ+7s7pFENC2abBKY1a3Gcosr0
lqP3KGxr4zxM6hgh0byw8P+K23T1L6csfuV0vxaAqHIlyj9YhfInTPT+uO8PjAzyC2mvt3PvWiCo
7J/7DDtpObwO/VNB2Gm+jPrNFbI2uqO0YkNgVAPYubr3vv/Y6/LqmCuCeUv8Fvg5/auhMT/g0D82
KOcWbYOoodxP5jQO3dy9YfBeQGKalVmHOSCg+0CTAo7FJXM30Y0ysMVJbwuKjhHH5muOXPqr0K3P
xN3w8vA7b+OTlUym1kK3BcUsGwYXbDpvsnaVZpz38WGHzTEp7VIkQTm/ocAbaL9CowqwmBABa7f4
+eS64Bw7d82vb+7bKiLKtgWDWsySfqGgo61oQMpsmfLCyw0doHXpqXB+mWzzLITMAsHNdmEAp+rR
IFJfBMhDbxid1mWSrtyNtFwn2WrM2uf/8AKrGVbDHJu1DWmysmySO6r5OBrEUtyyik7BTBmX4p/5
eFLru4gQITx+ql5ipi8AQpqyUP1+A8fbymCH7QT5KHbRDwrgosCNWj6QuzODtqmjdnvIErT2VDU9
RC8lEld3tUc/GcDHZ6XaMXictZrmavVWGOiChS0B8y9vGGAlyTK6dWQ5jiSa5wdNE+HyHPabdxif
ihxXsSPrxYVHyB0fwgE+JRGyAk5ViXJQES/XC+1nJohMsReAkyUXctl8ebyHsu4GtdavHQfCkOXX
wPyGM9OqKV+cb2TX+L3C60e/WqTS+/l7lzoviQYpVGL/lsjCAo1eEfyccUJNugL3EhkhQXZ2jxqo
mUN8mDLY4jjMdEMk0FRS8cmWHSQpejIWUB5Jwfn8iElZiyziZ527KySg0Oz4pTz8pgLf6vAv+5mr
3Wm5iE2FouN2+gtGQxlokg/6cJBaM1KmVDFyqRQxr4fsb5yhO3FeZdGiQXznEvImFSAiDYVCL6ug
vonoSnVXgmwTDPPtRCgWlKOtkzs+fhDCki4B2idHnoOZm3Ysb3UNQDWocL+ad38ZIxCtktLO75Hf
uiSdCbOpjTJEHZLfeN0g3G0Z2OX9ix4NeF9yeJCqrHVXk1ycT7oDk+oQxHNKnRLRcgZhhytD1pUf
g3cb1b5TIydJYyKqith2Cx+0hoZTjJd8z5GpRh15Cs6xyyn+I9AWy8Znd1LxTNRIaIA3gvkCvzrg
QKwSsL5KQv0HY59FOgIVRJNx2INC8/s3Aqv7jbiXDq1PFO8sZybkwFjv7DMAgLtw58uTmZ6vQLp6
QhFHJ/GZMCxi1FBdIqO9lutxmIUfLGpDXvA1GSp6Ydtajmnjk35FezAo4jfsaNIFY+0O9ogbYpmh
Crmx7PpMKYwbtwC5FdaikeVOY45Czk/gLm7eKVUeJ7SZffq/roiR2tSCxxJrxFURA1B/dP+Rz+6a
IYU/SE+3+zBPQYNhq7rEvktnrItYGnohElMadk6wOnHMyNjdYvTOmUE6GOwCqcGpayGpq1gRkDmY
RfcCjEKBMw4uJW5w7OlBAwLqejVP3H9Xcp/uMV449qK4FHAa4twbo5ea27z3VjN2X7ZBzAYQR6Jv
bkHZzZr8uNIRoy9TexVKrbe1+Fgc8f4t9ABgzgcG1YBg7SG/AHi6OCWAjtvQhbP80LAkf2EYIGLY
mjpv1CYAYWHErAkamfhWojJ9IFjfEVmfu4uXzuSUsx3mzhiR9Hx5IS4IppYCXvN/m+XISWLH8Fd3
RmOGHHYn4VHoCbViBwmg+Et8L51ClHV0sZj8O6oJvq+LU7EpYzubGPWZB+Barxw5S6UZxMC6ejcd
eUxRJJc+iwfypay/G63msPaMoKJkdKHGVzWFGUNk+cid7ZQHqI48wjrc51ILC89ArQCOIGRVjgmX
nKR9SPN+qHfw13cY9B4Qd6wqmsB1347vEbaAe8E3UbHB8pZbPEEG/nBBLDH4QRXFe2pt//aBSCrp
QnN+pSZMGeP2pynumoaPcqHqdGJFhQSqqHZ82/TsXPM9s4HPXrTywCNeHr3gxaWIrwIXNuSQ+Oy6
JX9ZnSGlOuuB0x5iqbKxvDlx7lgypaAsn+RBmcJJPopoSD5Yh6bmIcJ/0itDlcDdewpt5nPUqu94
e4J9Ro3Q1jY5c2ECTXrEZy0zJYGMxTj6lgcRjNFTf5bxzigYpR0FMEOgWt0PL0xno6idCBOqqnqn
a46AClfBHFxURPEXm9qBbepBBmnZr5kduX2OflldTVaGCqe7YU5wix/EH2chnHfzzzP80eJtlzS2
tKaj5bqmRPkuHuLmghXjRzPugNtJbigfDzyfLWpUvFaN/meBl1iHpVBGTKReQCdVeAm7zpul8UZ6
oNtk0AY1Op9uwKcyJerRrgdpzE5CiIhhcMjN+nycFulhYMRaseGu+AZKkV0+ypc/i/TIlLMA+ExL
cZEcwAICeKHMxCGrZ+kolSdJ7s4dKs5NiYZ19Y+Sbzz/q3amJAYddjitzvKcWUN+FIgxlAS1CyTb
iZn9dLT39MxzioZAv+PFFLYd/ljhNPgFnJE3gBls1tkfoGJrUcrD1KBUtd7YvHI98FmxMnuGI9El
Qa8MVsvqM2g8GqFhM/nkX7PD2JBUhuv/Co9rMQGokFfVRzhVZAiJkIEAYkbhR6ycnHQj5Lbvw5Jx
OPem+6MK4nz7BUUhrru+qWDudFH8xfYk9+mYTq7qzYgWBfKCn0Y37vnKx+vae4exIOeAMNMwWfCP
XsCzA2T4gZTd1f1z8g1ooNmo0Ab5yJp/G+7+tE77L8mjS2EGxGYzYeX2gftkcZWTDLfZNYPjktXc
eUJBfi+9yKJrZedTkv8e7GTRv7FtAMcVu7HQ/4rVer6cvqBljGG+JUTmH1P97xq5V61yNDR+0cYK
Y7K9MQPt1G9XpM3ZSmTQtjT4qRTZvd3eiu7Uin+EQBSlnibq+mJzvkYgaNmP+9tOg+5Vw9Kmv7pG
fy3Hhf8NH2BQ7FWJTOOZ9PSGgN9cDYYYDDVrvAgooG9/znHfmkWZyyjmOWSQeINsvAUhqbOoB+VB
RklZWDqpBK/KoCiWpClqw26xIFJkwOuqk4Jg+WhItNjhnDdSdQWUkFyJALtfZAI5awiiGCOcaADj
o+G1bOpk2Q2o5imez2GMXr7M0mtAPp2lesWry+2D0K2rZWQMoWf6eppVZJyPApT2kIcZVs5CHfRY
f2f1m6e/VBGQCK71m4Yh9CLAaKnLL9NJgwun/6T6JkLaQre0osN0Hh+cwb19YhdE6Z1//d49tAFg
Bm5wnyNokD0UgMFtn57cD52CT8wli4BYda9JASuss811jquvpsmfcx7ARr6r1eW9knz8DFwG3yMw
UdzMDSSqfrq70UBBfRzyd/nxsdJJj8sAYZawsUEfh+NpR5yDJieRolVckBKELNja49PEf0VFOYho
B5KwtwgeQbIU1Tc0PWIh9WiEaJtBIb9Wp1dzS0dqJ8w+84iKJHB6Apcr++p4Sky5ahO9it+C/TUn
HF2HSwHxIoC8+dRdGho/7F0sdl1/JrpqICQR3NUYMHuYD8WXMpO+S7+L8TPbUMCsbeoR2oYE5+dI
YmUI4TTKdfr3U0C9wt6NL+Xc3wNUoSaGdCz75D368CPbq9UoxoVfdwRl2F2J4ccZN+c8sU/OPt36
PpCGmLdAnOoMQfwbvsNC7zyypdpHTFuQFTm+t7ix67L6NUDqLTo7Ug/YYn5g5hSak//6R6wSK48Y
G0OpTAGxRi4jIJRApMyRN5JcyALCmeWgs+icGbOOZGGbhdCDheDqCo7iv7Q0fJwVBuzyaxBGPaUg
NMLhn9tBIYiSrLmKoYnK4i0uIAdyi5IEqpIRIYCBzjzLZ6tJ5JDeNbgx77mxwbtCpSKkSqYVsVWz
O1S5dI2IIHocEctdyHdKHJKKk4tTaTMMBj2JDUABkEQYrhIZwYt92jm6esT1xOgTXGaKI1JtUEZ+
SwQO6qmKa2/SHB4QA+tXtC78YUANewHCvJSCd959TMUxH1/6FKxsxGTQ/plpOdfovtWtpKRvW+MP
hyRrpp7E3mz93lQHjQ51tFyXDegCas6TpcoePoNueIJdiJ5n8x+3w0OOE7Ot2Hla5I/4W5OJVM3k
Lq92DOnU/Nd4h02kTOQ71kfzvuj+SeaD1ukd1wOj86qw9BZBFev5+Mp77Ng6vVilzNecxondC5sN
PQ50CkAYwloTZmDQRXB07MmLhHQ/gnPBmErG5CWdQwsZxavH1cqSwhcewhchLmxYmbS0jVEMqoGQ
WH/VNhMUC7bbqRK5rMWwSXPgnL4yQ6VudVrSOXITc75EFErY4RpRosvJhpRj86RzatbYZiwWRW9S
hZ2hWarxiFrs+unf9//dbA713qQ8woFaygYMbmr1ge8y8r+LqWOFulUFM3/EmPpAh+4I6bUqnUeu
8W4pw036psRVBHhmfcsKYHZeNqFqBc7Xb0XLf9NukeBSnxCruS1ArQl2XKDhVsmaksGWVaxbH8Tv
dadmv/VHbbycKfkGuXjnCGO9bBG064cykWJeQ23WgoNVj83nvxbqBVk4YrmA+M+01j5j0jMBloN1
QFA3UgNwKRQaixkXDTNvHBg5OJuQjNXt2bToa32mbDQDepGMCwD/e0qXE1yQvYNbQIqforJQ4Cfm
H48OuWpSTijGv8vO/WCKnaw7+UigZAqm/8FKbIdQ7pfDUvavpBI5pIhooggLqX1jUqvw8IsdqOQG
2Wul0QaqpK5dft7Q8lw7pUYnfkM1MyohpaRAsEzsbFxSi8oLq1AZPfZYF4dm941lXgfR7hHCUnRC
tz8urrQt17RaNrTEa6+EBC+c/5lB0QW+RHNlYArjWkPveUsgqQjVz3AFgJcM51hkuiyIuf8xJd5n
V15UwMrvKtqJ9COMBBRp3KriEhJFvOrRfAIrzOcDuu44rfSZAMEZZho+ww8Cdym7SAL7DvWqcZFv
fngbye7d3etGHeCDKC2oZ2YIpG1JAZrjxkSBDyhG+ROTHcUkC8Vm48NHDGH6fx0B7hKF8wVVe+pX
R80r/j5clo44Nxn0OMCctnYh3q48qRChjhNmgof2yV6UASAbjwWnuesxLXmiJw/8ddfLO2TzChHL
oAyJTB4+iN0qakrAHtDMaQybarZCkgb8HOhiPLnUeR2/lPWV+vBnsSkg2DMhXYvbAIaYddUa8x5Y
PL/9C4y/rKNNIQ2ZDod/ThPkhuqKFG8XinYy6ys3V6PaDVJaXT0K718OAJbIG6MELN2v4MBx0h8E
OTvu3FZeP4lID8pGx+/ikJt0MFR7zBV36W7SEumTFW4XttMKOUHQyhQ5gFaKR+9IzJXLO+o16KrN
qZOP8kaShiL22w13oGXDHb/3e1ZSvij1H7M9VpQ4K7sgqnvnwEtc0kdnOvk47WM6RiPCHoG1KcdY
HLGx4aeY00yZlNkOCY1KHlp3R2zHzOlV82P9zQWfrM+cVZe1oUQhxAubMpMoO1lOpBiUp4rMB99H
VDYkcyN4WmmWyXuP3iAy2vTZ59XavfzVjaICxY18hIEeWfaN0W6On7LlFaGlPn6TfqvJnVdSZOwn
Q+2a5ERDbJanB8A7PzJZYiFgkIddwiBDyIQbrYrEhMSzeXLU/DFDQjXrbZMTKkYaTzdvc1gQMEh5
FWh1sWMwKwYuBFeE8szP4Tp/52m7o0LjObEOipuhY1B52+3LCu8Jd7/taS2K/JOD5zrOEAeD1Br0
eiAKeg6KcASxuhZwUe4xTgnCLMdLEaGH6m5UOEAD7LdhZx797+Y5WpuZFMdYkiepqoXos0T+kv09
suwgWflf7db/kvHTvFFJWFox0p1oXBTseYXxaaRqMB27PEoZqSIUmvuGEyKwx+9/wf3+WINTrl5/
iGqjLGIstQqHedFgcoa/Gm6BBJJAL2Ta45PRaeFQQqM+BqbWs2fGN8JNZXpj66N7Ebh3CBMS19b9
Qiw9EOqh7EwXgknCUxE1SGSCSnG6kepYgft7kSki5I3vdZv6RL+i3mc5cT5goJMMkx5bP0M1aC9E
HYJVmXWQDDF2n+H7AsltraTYh55hs7TCujjSbKxEGF8Pq4FL1R7RNWIXM3dzA3xybqSc88L+FsAa
nui5azghjpaIN6a3nl2DLuGiWcJzh5mcKXzQiovIk+SGiQp99l09nK74NL8o9dpqby5yeOZr+nX+
SaYoV+rUMFhQeAHYKG7z/HJ2l0gTP3DveOaRTjARyDhpbQJ4w1gz6tgcLk2WVSNNYxobOsYl0F/n
NuiQNtvn+E+0AYZhNoQ0xNrqHpoMCMdb3qBqePV/pa/c1P7RZbX3OvDT+Kuc7ksU0F9ZVj+h2nNQ
I24AVwkGem1LWCvJSw4qRWolInp1+KFzvzEpJ5QAGP5n4e3T/06wiMWy8ywA6S3yAzCZU+SrpIM3
PZm44RhV+FmIBhS+R5vgrMhlB7CYd7gMJEEeLGPVSmO7m8lST+7+GSAQWl5uTQOwEApyggMZP0LI
c1Sm0ksMGQ9F5b4aXa9wMngri1vSxVHRce3c3hAYvvm63PfkoTxvLicgi9q3WmlTQWdONUUjuE5z
1jcUCqUxQgYcprW8dfNo3dfZE5l3YZGdYrVkTU7otZhyh//q/Wps4WjbhxypTCKAXLNPwyj8Ud/D
5Yw2MvUMIIElB83FlGPRiGbpIaKX4yHHB5fBHM82X7sKuDbizOigaytNPq3q5Gimv6Rtgdk6HMQ8
40XTAzJlgF3+71S6a6YRjxbr2WDTj2Rg6xbFROufJ37Zqvbx1GL9yZAxvFogg+kjfGSIeJ8Jcsy7
0zNyM5Su2fObCMbf7sCo52L2CZLqUyWzR8Rk2RGr4/1D2VAQC5s6aTwuMdp/wcq0bQF5bviTdzu9
r86bBY7euBp9O48Rz5rFpzmR5aOMwIquamSWh9UKpUZFr0V9tYjWPKldDsHWD+325nJecg/Tf/xH
82rYVkkwfmb7tTUy7+355YzQdRm2YVR+bXML8gxh/yJ5D09fCQwUK4jk7BaX+2/gcB0N/5fh1hiP
V/wktabQGdHGvyboWmMnmslbtCJU5tm0W8EfiVmRh8cDcwNeNHZsTLnRh1rp3G2rjboX1uNY4RWj
QOptuWLiXetlTO4Q6o7vbImiEpS8a6PpRRNyvUnuYn4rod8/eh/11AdKl8qfXKTLKr19JZqe+7/a
n4VSX4et6dp6k3397qGmEfYGdxE8/Y38szWJ1N4hiQvFawMS4/L8A28PahmF2BBvc8EnGxlKsMH6
rwOQO27BkKNBCzt65gMufGOkjAi4FfdAtrQbvJmxRX+PJ9xgGpEMFMowYAqUMA/s65lknz0FS++L
gDkzdRk9uR5SNngadmYaefk6vPGKaygulhro064622rGGxY0GKtPveox1is5WTWFp9Xa2z4YVdZy
99zGG1MMCNuUvW9H9zqmwvSCj/4mfxzyNmzELxlSr0ltCs7xqgiDFr8b3uWOCHETaYQmmqWkOJpd
5XnX2mzLE9KHxB9I/rWOMmvM5nFJAdin4vuShe3jBoCUqgYZE8G4hc7e2NiC06MUL/BnDDDn5fPy
cduVXvH4ZSCckk5Pm/eEO3KpaUr9lY3d9Gf6HbipLJD5xNGFpJQcjriBV8euHjw2e9ftHMeNVZ/Z
omIIPGMss7FxwJWy+oU/1Ta2G0Qn7ZcUpWEzBRK9DRcEGOCBiVdjgexRC5vx91lnsFaXaz841umi
kKwwct5Fm3OkjpW9kvcVRb8mRR+sbtP/BUM7J3NzpuAlk9VCc4DIi958ZdcGaQwy+oek+8yjf45S
Vg9mUId9gm2Fpj+d0DhcEJmZeXfBFOf7PNsGsxYl9Q3Kh78yV3AiD0Jt7uhrpk6soIj3M0XLBO6n
Sz/9FaZZ/9g3fPgIfauAl04LMV/Dejlr15uVy7e1/KZo7aZURYfoNZmohN+VESMRYLgQPI/Vwkmk
jn6C/Anc4iG8enOiLNQf/H8w5bTVs7/R2N37QkUTUy0WDEETir1WB5gPS4W9IgU3JDYB+ohojzfZ
B0NderYAboNyAIPRSnzMndl3mW8hzOLzWa9aR8MsSdE4kCaVMqzcCJ10zKusfUaWRjIcuE6cReVh
nW+V33uoDpis9x9VR41vmibRZRwRFogu3w9+2C+y/hgSKTeW3/X0TaA0nsPvFlyCjADpPRFUXEWq
yqljcWMrFkHWQ/9Cs50+gv20qsJxTbqStDJmGoXxl1ff90iX9ZD9t7UQrMFKCZYoNl0A/qdZ+/rH
9dtd7VSh4Wyfgql/3gDg4LdiQaPup+tiL5iLMa4avyaIMkLVYpvnbeijanwxJ2cA7cLGCaRTYV+I
rxcry3oTzcD2CT9paM8X5HBl3df1xtYIr95DChym7zwwyOYZheSsyi5iCtFZ2HndOy8aV8UWBNHv
GE5YOgIIbAlB+xGXftTkEfLCPmtILhGNzzudwrgW/iitXPV/SrvPeloJeqH2wgUje1Vi1DtgC375
FG1mWB9FgDB8lVfG/A9KF8m+hnUuw3lsh7XE6tK4MfygqLphkJ9ocGV63+UORjE5j3tb8Eqmai8r
eGyCUcankP0kesAYftcypPeCgmOdT7MqTtNxBPnDMX8zGV9sHmHx24/6jxhknT0KAA9+hzFP5VRH
I9wHCPGWXaW0ale3KwoE6nD5t+1sghEoyezp+H2MZga0a0PTeH0992w88PqRiHXOHuFkvXKqfW0R
0MWj3bp2Wnnk7BM4KNi/2NuwZUOF8wIj0KzEgwZJ6YQ4sG17CdbhZpN24OLrNbcWFDX/GBa15byO
o+1jPLauGnkfoqcxv+bfrYofjwanSCraOi5yQQiRD3KO1ltO1Y6J6AzG2n6Li2AJV2ZeJYCV2Q2I
jCuVJdgoTmCsFJ9x75z8gjtm4+ikQ/W93PKVbdumDDJe4PEV7fFI49Xd5EoqULQAIjJKRnjyeQjU
MYxT2pnucjeyQqR8R9b11j8EPxvoRzPO2ZEtyLY7hDINqhKZTmrkl52uFFB6JvOs/dbsr9lz068G
frAqEVoC2yNEwunKkpQniy4ITkPjy3RvJcfKV7pFwsjMfCfRYaSUODfpQ9cVtUPDfXZQGRnyP+fm
tfYpCcs6GwZ3E0hyPB07us0pvpneM1G/DXled/vNR7dcxRgiNQF7PCYuQXUCZUd5I6QFRyPzVwhM
/ZBCxv+fsjTS2+dmWIzWayO7msRnkLsE1DFDXMmiid99UdcQXpGDR+FawLBZ0ftHuOo7zHR32Ig9
cBI56lHbn5lOSVSapEzGxTAK/BPYLCI573W49MlqHOGSUGkwebx0IaqJmkF7NZ1qncD6M99mcZqG
2wSWutJ63v9Vmf6MQaFZi0IRwF19ZLL74EHFldBCQEQ/pH8nkt1f+DT6Vnnr04lxSJuhMF/lwe1j
mcZWjEdGamgsPyKZTpoPOmBJlEb7/DJ7MMEVSddyRBa46zNpFnhhAKW8V0tbA9JdJa9+Yzxc6p2Y
V353Zpw97Ao0I/QYUx3TOd7VdUihH0Dz5mterIEXQWZt8NL2M+JWs2qiXv3l625kiZknUaKz69K5
nABZSo+QzLcUkpWrcAznPoS7WN4lDp8K6GRWf8Zo0ZIdEg5Tpcb9xKHED6caA5gm+0kxrb0y/3Ji
SZGAmS+Ttnc/OaapXGm8hkxEZaYMMrJzcSEfDTSSNcDdoNFTo14wm82trG8W/SNEr7w3UliwR6++
wmjMGhHCY/GLRYxpv5+aOmzdckkRaetvFK6MCB88gpE3gIa+lqjcKJ+hlj4LrK4Lo07FQ9e7tRZb
W2/Gh2HjdfX68eJgKYpaGCnzniQYkIEAR5p9W9v8Brd4Rn5UG9vv3Y9YyifaktJR/FEODEs7w2iY
f/ggLuYJKeJ7Jf6MgzMc9eQeLkrCtGxecw/Gl3Uxjab65ycPVrwq4BGYjfuCvhTvmSdyCcrduLWp
DZRDkQZHEBYGR6yJ1O5i34oxuoUW3AIgpaBLBECaGE1B6n+N6qvRX3kWRRi6Q0gapQ58SOyUdBQx
4UJNs1HW+wGrWiBGaahbXgzXHQSylJQsJTHVBikS4j360++/QJded7MuRFU5AnLxQfxiT7aLcFke
MCyHGNPLyVeAr7F6LRJHgILQarNQuRIyoH47KhyrllcuCmqgOgadYcmUqBVDYktXAZYb8Voai6VP
/XWaUaXgdeT5V6DgqrPtYcB29DHlbWjhNCar18rDbPxxH6NmAu12aAXwV97r4AFVZ+lZxP/YglXH
ctqRNh2PDDw5WEW5sqPQAo4ZTfLBUCxU2inN8cvlU0h4GyM2x4M9o6LnanQ2ipdbXKstQdc1rWvn
Kf5ib8ONHje5BS2f10wDsi+ile1DYf1/t849yXVVC18hs18FEe3XtBOgwVK35A6qtjvxjzG+bXIc
5h3L9PF/cQMv3lxPsJwxrF8Q1Jp+6LYmHiddOt26QzSPR5ZOZ7a4DMWLkmpzi5ubJ+GJOad1RvkG
fvAqPrGsKRYcxsU2krgaHsR7hh/fkt5xWSTYsqEBCkr8jRzBXUkjGKdJkCJvHUQIWdasmj4SkwrJ
xg1nUSwA4CinuI+jiLmcBSSG030lfhffPNiDmSsJpq4PbPbKVJsQKDBxw/o4YN3aEJCemfiBEUvA
VjFqCgCBCZ/HJUKZdXtuLkjicU3SbUsIh/nMHE0oe+sWzcoWxEGcQg/VGVpnFewsrqyu8lBt9ah+
dIvWn38nKGrUDuBrzoLlYDV1noXKfpXbckzH0xWmMniFX/uMSEeg/RjNJuUhjA35CSVa/+W52nRE
42Diub5inWKiX7sKy7WLk7lt0ZsnC42XS0IRiiiVv2dl8lbsx8wp78mjv4c9AdlXYt3C8uqfmO0P
cx3C3G74bRHcD3MKkKSpe5/pukokwudj7r5UV7R+7eNWrUttrBJr0txkdiEgoWRjA4N7QSJ985W3
GeCgg6BR9Ug21Sou42Q4yDrvlMPSkrvpruLQtvhFk6wOkD90LEizgGZm3k0K1m6l5Y0EfoGYkrh6
4LoliN5/gocV+lSSQ9y/+G7c0U0sKiQDrNKxve5Auml7vX9kwq+iQMkptL2CMnKqHCsQHAQv4Gcp
f15AsCdwYhTQTyYifHNzLC0w5nuqng2J8qIHjpaFtCHEgGLXcf2392VYwCZHlcnvo5zCZMlQGNdf
ibQgM+HlVzg0BT238rgRXPcmSyQErqi6dchXZtjKbSmo8k/uMU33FCJHLy/U1ovxQAj5y26ePV4Y
U8SmDj8LSyMjvQt61QQ3Co9F9RJvcxse5nm2Chr3VFHUSZgiw+HvjXSufqw8vBeyzd3cVO/I0hwd
FKMWvSjq48eeP7qzC+AJ3IqBva1Pt7mWRmmyzdn00kKTQhl8nYWchRsYATQYtp0tvWrryXozrKd0
xwifqyuo4AAIwuckjUZigSdq3Cu5SpT1TK3bSb1SmCQQobjrK/pvsucZoa1FfDvYez798XA9FgbO
ABrslVyKfUWq9m/cApqGGJhindoZGwBqkb1ZelvO1CLzvAAEwaR74Y3OWNSWCDn4hbEJ2n0XwNU+
SdfSHVwjIL6OZBaKG9cJ//DtwhmWu0tU8ON//Iyl7QsbudVQyp4nOc6ReazhC4hPWfCEL0C3xnry
HwcKYP5N+O/Ha19u8NaZyCoJkRyOe67f74OxdZIdPGtNMpw2GxrW+NCq6aXemiEnR79KFUt6ZlhJ
tO5K9Cb+wIn+gcQtqt8ShNlykV6kBx6Yt/TWOS3+395PF+XCqVLpplhIkoYFxPlzxkgc2Q3ZKpix
D48CJJfZ4ow5p3KAv9X9EwM4FxIBxXPcAZ4tkjyuPnn58UvuN5B/5FVCTufE6jxTM5mfTjoeB2FR
Entc3VN3vQdT/BoeskIGs5Omvj42HJi6xxKKY0GA6jQgqj+wara/kqYSC7LDvEV5+kawleGVJioC
V4urJibij9mJJ/ezKpJWVGAufDm//Vu+ZyDtaxNPE6SsB4zR2zF4CdWVxkGUDzMh5mA80s14l7aS
jsmCio33HLhnUOJrq7OKtpCGk0awzvTzk4g96HGXT+X0ce0qa8EQwDoLL39O5isZH0ANKAh1ZDee
J3B/lF/Y4EYXn5ScSY9hbpWGmMJV/Klkti9dWn9XsJXDztf4nHv+BRPrqLNXr5c2sHjNrCzLF5lT
LkXdxAgQ/YAHuMk965TiwEdkopv7uEx1+LmhBqxkGFna8lrvpH00mg4GmbxVHO8Wi+SlLCaK+NBL
Qj/Ijty30bKsxMM11WoK0tF45+QHrhKuyOsqKnkQMqtm3RYTj/82oEFfkkWjvoc0E0vDwGzxLG3v
ki1IuKkvmLVP2e8iwkP0n3/pCg7Lq//4T2CiwzppG4IB7+7/CvORjha96rdwEw1H44s6V4PPERHB
YBRt7/nzQTLBJhVrX1RGsPmfiRx7dBdh+HYcuC9Rl1A8piuI0eXVj+OkO1bK8zoGPrndOw+dPpNL
Jxkz8m4XK4wNQQaQEYdxKv1SfLOnok8YAbI/bCdGyQtvKtPSn85DYwEW9oGda60k0Var78+dwdJo
+aQBTy2MS5/CMIrh7g6bB3R/haZgNm3GSKJx1Ze+LoPqyp2G5l62hExp6JVsx/BI9DTWXfMuOt6/
8cEBIxYt7wiCGF6FP366HO0Oobb1NeNx5JxsiGI1eq/cEnCl2WPj5NStDpAYtS8NlkYEKhkCMg4c
jz+W0ws6u29J4yX9z4dMTxytJxqnRZzkscW3nWvWvEQZYZ0cBBSOkELIxfv6LGcOkdWI4QBGKw5a
6ZC1B3txS17Ojt1zcd1ks6CvW0x8mc281IWndMsoWWoHbwsyi+PReS6mnS+MaiHMNxe5msD/L8ls
Zcm+3pswWxUOyYl69gA/xcgG1FSL3uV0iFoyOwxB6hZ11+gH3UBMYhfSwT0qKMMOYHVi40ERqng5
GFDGYy+XoB92ZYw896cxHx3gMRxxMOlgx2IgB/U89ppVgrug76gBpU50Z2ccz1Zhb8x5/HDBGHRy
KGiQGmXDSW14jPfpwIJ88jw45sdRUrTvMjAOUUx0rxzSKM7jPJjSPAWUynQG4otwe2tgQnuLTA9a
zoBSb8Ld2aRsT+jevKkzlF4LLjx4qWPFwoivwDmgCvVLajRlKtHc89+SnRHMqlQLyVvbA6rG+YeZ
W6dHa5Vc7KEHVSni+GFq3zxV9/AGIlSwlNHp7fLcnFE4Ws0qbEYn7gCHGoBnK+DZFxb4xlRsAmba
Rzmzd8GOVcLrBIbWv1NpOjCechvBxhYjfHsxPbnwfEAcF+gV9jKIj0McmICRSzcyb4xPt3hN8mLZ
1pEgXlti8auWS95bcPovw4yx/l09/UcvMhCE7KPQh+k1Z8THol4CpPFM20tX9QNgD8I5hy3ZZUOX
+XOn96KbhJ4l/rNt6aLJs5OS0dH+WlM4Y1xUE/IuqSg1r8ZJrCBAXQq/EmQtlBeU8EM5va3LNL4w
cbNYoDZ9GYFwYzTUmKyE7KAYoxGeHzoimJJS9o5hUiLbEQJDBZNDS2IXiTNl6FNVPZ+PrGwatk0s
2t2O6GGG1nlvaVCN4qWaLbC5CrduS6psoMpMTx+LPRKOwZivf7jjLu61M72QwH9OazK2xgNEco73
wirWAf4Nknq1Zl9rb4gaGLByXenS4ewsjF7nfkU1ZVmXfWTL0O6XnA6Th0x9gXgVin291dIPZ7af
+3RUFUpheysHm9I7LNwrUzacuCotjRSptVZgsnA8QszdSzhELsbdDQ3PQQSY5ikAWALNKh5QuoxL
daSJfL4H21kFN/3AQ7xd/+yk2a3WqDKf2WMs9fb8I+eoFR2X8gcnhLR5jLND5GVvAeFxJ1EFrkxZ
3fWEOpPbpBXPvwgpJu2rUOk09r+EexMIr+bp8NHVDNXhlqygqPHUqRT0KXJGWvWQ3OxpbIfkvSLG
qvpE20z9c6NZy0MgBtIQi2LVXG7lwU75FP8NwOV1fXqRPj0JTBrg7YP77mfBP7yxekT7h5+OVEsl
2QhfXxQ6BSiKD6BXfFeOscGJz/HKgWklypqWVFcqbFqFFU21r2WoQyitY7vNGlJDfDVww5J9H1mD
ZsBgGndd4+XfXVSVJTP0WEtq91U0L+QavRDE7SbontH+KHQvkGUGAtYo2QM3sdoWhx+UnOG9hkRp
Y7MIL6iMuEU6eSSYuQhgY5tGW5Ox6WejfpTudTIrftE8IXsCAh4e//8cGK+iJHVhXAQg47H21WRH
zB+zvGztOAwYdD0W9aHzleUBNem1gjdicb+pn01UNh7SHJPzpJZxztW4klp9cRxZwSQejUYw/q18
AQay50DpUzqHWOatVJGHpRPi9Y1Iuj6C6V1kC8QeCkckvG8Q5QxKxYBD+PsmmZCK8Gr4GN0VI2yX
oG66tA0KjFdRCWbv9oURnlBuz1tnRRasKVMC/+pl6AwZxiw66WOB8DL1G32iv9oLP2qBrVkxikr+
g6+Lwrq8WoMJVo2d1gcl7bJJ78whIJ3xBEjBCx5e/+fxiCxduDGzsgRe95saBLtehXHXKasBt5wn
fCwmFnVc1g4pcyxflGHoJ7o4gt6hw8aO2fdS+HO6hxZH8AAPgyJdJ4wogKTUtW+QNm3bSjF/buQj
XId2mqaSGdqjfyg0R8KBP4ojtYm8AwRfJ1wt0O8jEal9P267i0trmKjE7MQsuzl51csSOPfp9TTX
zTyaDGHf67y6BgGJiIyL3bctWnRXI7+0tWdiz0m4TJsDCSZH6FFMa0zhwrKTkTbFPDR2FxI7jz9P
LWhkQtddvEQn+v/vjMi6zsKptgS4bWUUYnSLREwvxQJ/jofdqMD60WGVQJS5kviCC+NfsaoYmzn6
9vAscGkkC/FjkdaYC1AuORPSO6vzcbu8tqb/D9ISS/kpbFqY+rKfPvmVIRF96TQGWo/lCKhGTzZH
6opK8II1IfRCEZTFqK3SVVSAD6ln5yM1TU7dXR8rWFrAkhBjgAJLdNHmx5HwPZ0g1src80dGCjee
Bn5NiET2xlTCLzJLkev6nBOQAZ0MgxtLsk+Isd0hjhtb1Fo4ZuQffYuNSeNi7Dw5xOVZdLp4E8ZZ
0NuaQ5zW5bmq9fNYpKkI/HOtjD2TOP0QPqkMOJzxa9S6QAl2LzIQaaehCsFX9s+au5PqTwSSPG5V
pw7JuLB98TKYWQfINNI95Rnu3TeHvV+jB/gEOYtcfm6Dcsv2sBqOZ4/2C+8JCr5/z0OMg0g6Uh2V
2qu6UPtKp0UPI6n85Y0dnhCHeNxdirMP+mAhpujrFaNARG2d2ZQPjMJ3kmizuYcmmNLj0TmhCtSJ
vaRrf7HyDf51zFnoVElcnzswx6rXyXdb1GOTP+KeMMjOZwoGlfnAkAeMuoRMe8ysxwtRAcT9lHwF
q71N1Lk9q2XcGom7nNsDiPJm/C4A78cECOKL8B2TS5+ArKoNhLpMPa0bxhIft+loFdgiXDke9FEU
H1IA5gR+Mq4EpZ7Oqm2h/82/9gDTQ9GNlE7CxTQUJZww4p2d4t80zEjoyxSvXQMqFz4AX7IRoq8f
lSRWANQsJuIV60avtXipSLyGuTcpHDX/dtQhdmk3st3jkbP/UlcSdO+dCbirDFeS8kpIfdt4r5v4
dtvXyoA21iZJKcUO/HzWOvTera/m+DKyQPQynWx/nwlXSgtIluZwRxVf0FpbXKE/u694bFmdYaYJ
WP2k4DUs0B+EpucHv9G59xoLGicPr/DFFXK/vD1BcGZbLbA2AuPW5Mw40RhrWn2ylCW3sQyupBpd
z70sD1g++CrD62AvYdXjVo7fBB0jp7il7g3qtV+vmtmX+0Mhhsbjo27/qsYDo2F+s3rR1yJbT2Xy
+pDQr1xqCXiPrV4TzJjHnyi33+JDYN/wNA+qa67aLuCvVVb4i4PBY1cWVPJA2VwneLRI68j/ldsa
vYGQ6mDB15ad9wxFCqAQqmyqrV1npsDgB9IvyEtlZVtPhv/QqCyjkRzG3KwMH0TQM1cOaOKZKNOS
1sPrE3viqiLZQu8KDz/gSTiBs5SLR1r1sE7MArCZJol4m3sjm4GUKChHVGFBJwAHktnIMqZbqvTg
RDV8QKt6X3D+AWjPqu20kEIxo9tYY8ugi0rGCkZOxil4x4fU7pNNjlWCJC7wNXWuY9YVMA5WL3Ar
zAhwmJXgOX/zVrANmUIP2LVaheMzNHLgzYgHugz8nPBo2PTD1A81hrKUedFQRKiFrVLbYLRx637D
IwL6puxhrdp6JHsOECM2GTT21s87bvNi99b++Ub1/hafE6CqNVjA9GrDw4Wesjd2Qp5LVh5xVuO5
3aXkd/eghY9FpU22sMXxQKVBCk5mu//gZ94lmIQq3ZxL1Vl6frHPP2CkbL/1OT4LKxNPP1LJEll5
BGRi46reuOWy6RioYnnlkVVfsHpJfYdQhpsdJwoP6TcfcvyGpvB7qsvsxJJ1Vm1DQcajnKSI3Tx2
MtnykJ7DhtWmo/5lzoush/lQtIyLaqIt/byEPVF+gyVfgbY7yWudBgPtFiBl6Hv5pR48bbU/fIi3
oWy84EKOAumcFY326+8S5Qx5JUpOMVyClE+bUF3oWcCHjmkFMfo6SnuFLJPlMXDpnAgu5QT5Jwcn
5IAgccPgma7iJiwb94iwnow99PCkp7N2/rYdG+4LwIWdeeROzgH+ojAwyXEE7h7GbX9CrtkbIHPP
h3ItiTV8msK3f4p6AqBFXxauzQlAkyTggB+Ml1UV0iJDwr+uPRXFB0/tduy60k2jH/jewFHn1QvQ
bO0vB6UPoZ2RJaZBTw5CoPr0ktErxUGe7yFSZZWrQo2vLx5bkmi7mDxn7dKbrBjvI94OI+AsFPum
qZhbscomdjvwedKWp+y6fY2Qxx78Yd1K8DQPzmwiRMB2sBPXVcsyvKkZ2+yW71JTBH0RXvq7z4IK
iXvmDpJ1S68jrPiBZWDof0IfnNUh4xkQ5q74+43ky0LoFFrsAft9oHBSe0tvsNq8xyST/JLejnBl
WOMpxUyBg1KWDsuCA9X5BInEBev86rqHY/vM4RfDmaLb43Gn/Xq7kCDK2dNgQrPzDn9eM0pjuBCP
8veGuU8QBQ4oFOOd0EYUaYaVfG8lNIS7qZl4H+uOo7ULANkeWCugYOwR9tGfwHOfUADAmkn3Zat3
rdaf9F2L0wnz+vK8qlhaWRo5Hc8KLPEpUDL0kQ96WzDg66DJdF9Hsp02usTagxLC2kRpelgElzp7
GWyb/WHkwGwd2hRQp2IlSRSd3/8b2W4G1C62yZp68UhYXhjcQdG+DTqsjYuKWAarvek9PxBklaU5
st9aNmYmxg1oqUD9bRt6fWtMj8nt3/OBFQBrquto1lFzZylBdZ+4rV68PzpDz7SOqdT1IAA+IBBt
BtLTsw7cMkXakZ3nubthDYNyMnn1Ma03qyAZPi+j/XOl+Z2Uar9vKrhGK6z7nv2njD58vwPqGku3
UpqgHpmaLf81A/G71zQNkHzGOoh26niFwgxfirnJuWjoP9LmPxJwCmCT0CzAnsPXhtjrixfEV21y
mQmb1on5HqWG2/V0m9C/HhYAebxgdsS0Pw9E+BhYk49bJ/JTCuRH8mtXeV9+vA7Kz0j7iD6sWFaS
bTDCNDi7TdKju42NMMBRdrzqurJRx67jfVe9mA8zn1ZN266Foa0AdPgsEvD9/x63F2bV9R4L3Nas
DjkO+hTQrlxOJgxT8F8FwYfAGCti03XPHn4/X4QdF1DOtUk1AR9jLhLf4ea2jE9CDt4CyhpaN/KO
4tlKpTdDgr735Z86JW90jGnb1Mr9bbMkDNUcZj5FUfDre3Xo343J83WwkhP27lzKkHdyIoHgoVkS
91s2raDYDaY18ysrDs47D6FrAukqDnYl5hDouRWz4WGjfx0/VjAgVQ6xz2pzuM63aeMzzDkgZ03H
vvbbxzkLpq1oXIQH0PzQxf0GpM6AcqCzdVP9Ue0vbA8Pl9v1+M2p2a1VTQPVPetnCF9IDh6HPyWi
+vRFFjLO8MmJbln2q7AmkxPppSK6BHgdxU0nHaMUbw6dfDRD04fNh+Y+LQjUO1I5dAo5hIFuV0v4
gadNo3ORGBGO1Gg9k9/hlEQ7fX4qGn/kof7Dc544aFb4pwX1tPEAT+26qvEq/wjsAIH/ID89Pi9B
pITtk0cG+1W349ANW243bMd2e9uewNSNuKXfFfEXvUv7RYiqIVtj4Y3LPBSPKXKAESqlXdhMJYiq
dq2cRsnUzKnu3obeSEe3usj8w1aGKWetHqFJdkDkeOvagDgw3GBEVUS+wBhLiBSl18F/rczeLwDu
wLvXevZTUrnt+i4IuKMVeyw/I75n9N3W+dstqK0Ww8LOdfCELjOiKvK6lcZK+36COLwAXikTtgIL
dx9+h35Zgfcii55fnToV8tzqb4pLoIvnKR8Ycx6R2+YaHzM3BTZgqwdEZ/1xFmsuFeuuna8UxXUL
RNSTAELTaGbbm4HC0JUpyF7AFGArQiEugp8FqDbQe9ARxz0KEL3mz5pkqA/njvF4GBN2kZBnLBc9
8v7QQwbAjmDM5Q2sxltq8DUoPCefDl745zvgneN5Bxr9tXlhuQCBX7l0tJSXOeeTbyx06EuhiXoS
qbAdi6HEjGqgWKNYtvz4sBQJgwW3QKIhF+XntM66ouaAlu+YVXYpSlJaGQebfBkcaTzpE3iLRsDD
xH1DEr6yyrw8bpbhF5HgOg+kU6SlITHH1s7thzoyFMq0Si5vuMs5qFpNdE1jeKLS8Q/mbO+2iUn4
pen14lIKDHl/I7ShvvJ6PPFxBQKDPG10R78mwUMYvcIyD/66qj0cOQ8flpRFRfNUj3tZ3xMQSqiu
//K6f6FbWGfo6ARwTRy9CllE0iZdV/m0ckKSzzzqiTIrsYRnWCBdMKtFSlxiM7nsTwvAxvPkSFmE
TGGfAqOYDas8dgFeR6NWMzczS/NeQ2CzYhiTy9EHA6D+1BSK8U7wGGZp8ybXDLJQs15YBW0yf2uh
rX8KFv35LAa3y/eqXpHDpG7WLDR6qJN4e5zrzekK1Bs4HF16EGNv5Y3p/RgeZpZeu4q70cHWsWC0
WUmTCv+SAO68jV+BlPxWOkL3lj4r7HremyTAaGUUuEWqkN1Ci7gIe52WQkpJLiBQt/fjBIEYY8RO
H8BYCUcrJvmlNh0lxBWpIg3XYfaEidSsm87VilKo7nNvfZdPO9dfMMUru/IWXrYzJD1blVqfJ6yE
IF78MmJrjw4RPByl0wyuZRMeLCAb+OB5nOUkLtY9/dxhjLFQXmt5NSipp7hYuW6wLXUfN50viyct
JkmQB1ck2ZmarTrnoebbAhA2zNDDYiOPTF4MdByBAO9C2c1dxdIPgMktShke/OtXn/5B+D3EZ5bj
eRjd1bI7yne3yehAip8E7qKATvqpaVMyb50GIHMEZmCNR/54pnJyHFixjhZudcnXTtpYRZu9TO1J
arifF3CuFNbNHeSS1sbTUbB+vZX2AJNFn0xPgG3vNnk4D72/P8cM3VcRKKeRC2kOCxjBxe3uap7X
4Bi+M0UwO8WrfazfT67vVsdRqlZ9fpsXlTArTPczckylP30goixvZlEzjrJ6bvn/Z457S/+pncV9
/hGMygTODHfMnE/42XviS5DWDA218Wr2SbEHvTQxwN7fwLrbEFHXkhtqotIO9yzyru/wg2Le8vEV
WP1/HR1kynjGS8hgz8pEBp1gS9ZUIsXosl5xGzZxAquB+BSpxbzLLDK9HRlgMiTlALw9rVaKLkY3
0SrASGIAVxuqvlCYkGatexx38bAOP7RTJ3SIrgjkQy6ccPOmI4EHCndKK4gyYJ5HBuFhQl0fX+lA
rxIizxSZpRs4s/RPj3/mLPuCWF98JghdJ+Am2BAVcnV+PMic8BMV8ih3slwlfCLmP2+Ktv8eohim
oG6SSou1rL8yCeef7yGuHy9q0bWiozV572n+qmnk8Qu3c4i0f36C5HtBbYQY5IZvwWmT9d2EX8MV
DkoJHQmoCdRkSmbnKpIrV7x8A/nTURMJ52Q3J7EpNlayA5JLqwfgkn9721vItZxwmHlT0d/ejntr
voc8HUPmFsuHfdtL68vJUgMNOzcNLdaPvSipG49osTS5gpieUk+3102LeysRMO+U84R4Z0tlO6Jm
BOa6TCRpGmpd1bXODxC/5BnSOxOWWj913SAzsr/ie0Gr9zSXOXeZ8g+rzMCwHXLPOVEatoCg79Kc
lpHJ6rEFAtOaPgnC/g0ihm/WgTIPSM2QuuVcDstznrYulTO4U+fS7BcJi2+Vg89deTTqvh1dm53+
wFY5bxNUJLNt1IuNu0eydYwCVz0xmP+eqIMy14HGkPK5FkASgq89pIXoJ6svCfmrXmD9AtIbxG2j
ula1yc1iu+HV1HwWmwNsQbDk1N1KLSsxLeZlbKGp18ZjL7l8s0A0qbGIQyPnpvRMHGSKQMMk5nxg
go0vD2Cg6GRkYJQlgXpDzUN4n1l/176aTAGrYloMiDQSiI5ADJObQYHFxmnbhe3QyMj8saFw74tG
PiFKjeZU4hLQIjQ55BzxN2xV3CtsFINoSzWppyeeTLeYqEImCMrjcYKWd5rq3KnazvFtPzlVq488
qhtcsk9cwsdeKt6Ad0El5QSiiTZznQ5iG0+ZJ2TgDMsRclOYUdKH5z8WJjKQQZhshSzpIIaEcagb
ArvSLMn7AY9qUW1VY+meTvnDBrlnriUCpLtXNq5ILJz3PD8Zy9UeOYDp34Gbssa8iekD9v8kwdUn
KUgceiF9b0GmBClKRbSlQjfS6nhqxubl+MItpnyIGmYKF6VSw7iHyoAmawHnpnx2PxDnjt4EQ2VB
oTjrxKWy1KWJhUoK/ZUv7jBJ/bY+A3H2ScSDFZrwaocY/1KRR21zX+DgnGq7Qql4UDTQiu7sdDnI
aMQEK+CbziZBJ33HenTcW1dmbuLqrM9dhYaMouVruyRK0DVc2Hv4pKmu9YirLwv6N4RkwXp536Wl
j6NP1rK3PTV0sjqj3QSjJ8bmg4rtMGtDkSYKYvUDVVS/hEJbo5Gberr8BAPkmPYVp/V1zxcy4y/G
3Nm3sz4FG5pC9/1hmJ3ihuxgUDucwbZRWtW2zWGUneTFr7Gn11gqqAOP4vAAciUrj+31IuQrNT9n
qIoPz4vhMGVEbI4DRUBg4iw5KueE3TWxASr0gs1eka/qJlSlNUQBmlVjrGWI76RNMHYFezBM+DmG
nWk3MiS8SqXlAv3U0ZT+I4YLJUo2aoMz8z9WlXQWam6sZ78GZuXhAj3kioCWKbKpNwIqzhmB00M2
9AaOiqRQiKgws1U+q732VyUJKnPchCTF9Z28XiDhnXS6bupM0FNJqmVrUwwg0z1vTHOyd5FLav61
uSIRSVLgszIcFaF0TmcFtKAAdvjoBowPP8vFFRGnSWO5xEeB0ysrJSAGKhaKpkEIq5EyaKlnN9gd
MLSQ1hwe4sPnfzhljFuzsoy5u2BTJYXmFCfU+pklY+cZG37XEl6TgiFVRRHr+CXnLbFdZXtlJcOs
bmpx6MzUH9aoMeGZ2KEvQ8NyN0ptzxNpOk2wCrOUYaIUXnBhUbvIa1SHghLtxZRbC6dR8I3Tyojt
JHUgStSnRfaBpJhvYRQk9dnkxk31J4/ODSEFcfim/w6jGM+B+6+dGwOzgV1UdZy7vIAxS1Geg7yi
oxeGCwBWs2nPR1sauuWhgQrDTVTGTLCQRO+DW61oudqhAUaApQ7Ziw0hXWF2sz6T+cmLfpwAXuAk
EkqUiNMp0NRdByMZf1jtSEdiP/pLzvfgQkzRS2zu8ei3D1zGtHc+LtjZc/R1zEIQaIXo8rXG+bSr
146D5eVEjVZDFtgQ+x9V1GFXTYqSPDn3nJIuatZDwPM854jg9ioEh0giO5lyDVrWzd9dIqKzPmKn
QBqTCLPuIqy2A/SOhXWDvXR4z+M9Usz0Yf+McqtcFSBfxTyTyZvUCa+jwGCyM2Nm29gx73wCvfGJ
ezmKVkrRmINhhyUs+rLpddjC8T7WsVxEufvVFi+drKRsHyrRqO4V2j/Dyq3VVcz+wBZj5k41Cl1J
oPh62Ubzj1vX/KAeBiUDr/8INc6DAM5AzvzYM3Qx3kt4uqXbIJ1qPRkPh1U3p1/YUMAo/RHBYgS0
GsTLFsvXViF185tQAgfwndqBj2DofWHjhRYGk1wtrhWpFoj9DZzpfgxP4xJ7KNQaeYEu4J81/qsr
s4bb0eD0sDPthFD6FdrXKYzoFKcwRCS1NNwvSN3xk+OOHfQ6nt4aiwVcPIItHCr6wvWsK3tu86S3
KdCzKCj9npq6iJXmtQhKty7Tz1G6NhzhYYHc0EVYxiQXvmd7iNKOhe3tmFkoHd7EhXvySPim44yB
hBHkIezU/yC5IVaYj21VBZzkrLWsfHHLMyjxPKoy7e8iSx8KWS0sJPhxdSIB3beINLChxZ07dJZC
ejmmSkNjncNRASGXoAc7T7d6WPz7bZdQd4nBhN+dT/p0zCbTS/35S75zD7fbeKepZ9hSOyu5+MUV
3Ay6Hg+jLhRVqllv5MkbOFwutrBPwQ8WSB6PMxrxmQHRLgbGd2a21Q84NynhmWm7b8grS2qY/waf
881nuHyeVJHBbd5OFUgG8ql0Y3DCSPDV9UumYRzA/tq0F5EAEauDX4QMrISj9xi+q4MXJ/hm3cFi
ab8g8HVW5SXnax5ntfrf70u/jkNPCB8zlC5jr6dlvZA9UnYiNA5ChzJr1Mu2zKdPOplF/BxK4Qbj
uDh9Pn0MCiscCsdKBS1g/ROlLNk2EcT3gtbo6VX2L1gF0qNKRcvYKqvgOUZiVqA2oiDo5AFXhm5z
u+1hCMW/Oq/3S5WWHaOxxtdy0gLR3UsQBVHpaJyS0xL78d4uYJxeOx2y3N+levJDjWtyxTm8aLEa
VoEAMYtT+xRlhI2B3JZRiPqfRJ7HIxrnnDloiY7xH5M9ljxGj0FbRmqE+ZoxY8GfToTfB5dnSASd
Kfh4rRCnlDKFdK6t6T8z4GyNlB3gNOEaiZz7RmIPqaz4JU8jzYAKF3JBwx++CkhAmIJPbUAuGq6y
IuFhkTygFZ9+bDLVf8i4JXgREAvAP9nb9AQSTbdXQdzi23z0LSFZKSRewDWVhuNJkkr0H0V3SY6t
fPeoXQuGHRAjucaxFkkg+CJrAMMZHC7Ey56IP2ZrJhuAOv9JEO00NXyFbXUoa9b0/PvK6pCbm/9H
d39MYOZsvotBqQ9KvkbPewYC39TFDmk0kgGtlMOktC+xE/QG5Lng3T3BqStOBszqWjPIdke32ddW
LwI8s44Arm3Ji3c90LAQa4Cx7H39iH0zTG61lxWm7RmOU4hY45pvAqJMb665k1yyEy2WW30P54JJ
G7gUYcnLCshpx7obyy6Q6LybLqL37l38VxX2Hrb2/0CyIY+AOHwrZx1H5uxSEBerxo/SC+0KL8j+
BfxQS1zXcFSzEU/jfSbJTHnmUSbuzIWwsYXwuzcBEG51c3/vhgMLW9RQAOEPrNCHu7QqtH0wH1Zn
UmrR7sYxxscvGcbj6DpHWog/BWmwiT2eh9AfyW8wNKbhjEJmRWumntSKDwOwUdVzQKSxgx8+jTe2
bl/3PKgw2hRbiNGwM2qtDvivi3ihQMwqNee387aU1PXVP9dvQMWOtCAwqdMiHRITdURHjOlLXzMS
v4Nrd6S0WusKNyboxxrYFH52+AS1c5kAn6hLHpY56jgOiWuv9dxfOnsPUJ2GUCyi3VJzoHfmLu0v
zAzTvVPl8b8kY4DRlGN8no6nzx+jXwxV9yO93/1FjiuTN9m0fHkPoQwDHyYNQxjfWEB91F47dtH3
Uqi5F0RNhp7GrTRlarNY2sOGCfTXDfJn6xNDvdLr9PS3woK+zCntT2YnKndiahSO5VGIBGg7Tx7O
j6QWeYXQ3u3mG/5ho/ZoF9cODmfv2y1AdmEXTaadw6ntgevoqPm4lS0gv8bw/iYQgSYyRihvEI4h
JAsL1jPaEXfEJ/kQq4IzMIW+CdZQDX448RuZol2mjlNm+jkoG7OmDj8i6J7IoqSlA953OcIPUHZz
S4wXB+Utn2b1KIVLATmd84JRD30DUJcvu5rvOD1UYJAkg83MGxoOYZqu8D+AAqk4P9OUPUWKI11L
PtfmLxHasCo+JZ42gJ4QeoTPf+DgwsuhyCEQJBVHyXCIYOZbqnJ8FNTj3ETO+hYjF66sfS1wqtxI
2A1FNz1ZPnFRDcY9jliJGmgqqVr3PnCMmiv3EHK0cKPhregT/wM6Ro8boAP6MN6xfPy1syLkF3sy
odDuAFl/oawHJntLEK/rZW+pS3hmcwgsS/JRb967tprDztC+f+p3hUV4M05wJMOfEmj26xLXOSCW
90UxZq+vqIcfJA+RKfI+9sSvHCGcPvPiI3xPgCHLlaedhdbn3xS9qbkQLwRR/AqB5e+f9jQOpT6C
SgA6s20lfCkfjvtUG1ue9GgSpgKBCjswQaLxrqPgdpkRGChPI2Hw/fHf8IH2fg7vz2CYqhIhQzHJ
yYl4YxOgOIMmkMAaR48rUTOq6FxEDA2m4O0T+OTdMX2EnfAzfYCL7hLEJLaUoUPTSywFwjsyNSPA
X1FXdP8nMoCsAYMmQ1Tcfmq+tlxLMXzLieT4ByUc2/25x1kAh87HQQUHcFbnsN1YSWXjnDvyh8/B
gEX0B4l8K/F4rZUjYVfj0WKJkSDm9cOaqzvvfsNR7dp+6mrTYK2oNU3AsutjJFQ9TG8KYp+uP0wz
kwiIvRRHCfRiEc77nNnp1eooKdscFL+iF+W9CPn08E5YfdpIe9n+NGI9SbQqB1xvCyxz5gwbxKNs
ZTcqtvwfbZM5KzFzfSm1UvHyxknrZZg05dvSdhE4jLumS3DEJUq7m07vmyh7HI/iNDmZTI5J92/F
LKZg/okEPps0dGHC0KqadGRorW6CXsKh9Me7L/7eiYr55boMq6ysoK24eWjCLSfpj8g5Y2IDW+IJ
PgwMOI1HoRdMbB75zOtuQQD9qr/ig2F8/za5l9r+sPdmGCtO/aD8GAZocuxLifEoAux7TmlQ/eH+
IMWlNOd8F0o2G0o4/ok6cL7AhHBb9RhMhaB+bRMaRu39BPHgsq+G482AMrUOjatOmT780xTAB2H+
N0BXs6zB63d+I6ax/T3pyxibdEzrkeVjKt7OWIac/9cpW0xu1XbVcp4aGe0AlDh/kfX4wQUzhsGZ
XDJEvbfLLjtZ89vuFrGSpEcQ01O1G7wePUMZsRnbMd3YaF2VUbiJAiX6Y+a5HJcUEntzDdOyvJRW
fhqMjql4v3jk1kGD0NaTDrHygj2xOY0cnIJOT56cAmS/Y05KTgIq3VtQD2tk08BivrJR/yVRHcX/
YrYu30flTTsf5cSe0QWLqfhXK1BkoUhMyoH5wCGVB+2YVGhtDcq+4LcSOu7zY7H7T+5+Gjfv4Jw5
kuU6A4FBEJbAWHa/S5pOkdL5Jjqnc7AgzmuBktAUvRrbXj6LoSd4GR85Qv3q1gOQwkK2hegKof9Q
3SYHk9pWhv/iXOaxj+n96FKxjxUkMgPcshIVfM5tlhhIl6N1jeUNhkHPrDFj1YNru3iFwVp5qxKN
AmbM+zvLJqEihRWiE1oxtK1+xobgE8ROGGSAwJKkUJKLViqWD018m/t5bJyrNDoKp4zWrt3l44Y2
f4Oh4LzW7IlSLc4pLC4Ar7EKZtb8tnlsG4Ry3YL2lh5b24k5shtX5cxHW31jkWPILMOBA7opEwui
WeyEBN6JnWzYyI9PDP7O0mnHKjJgNgfi+ERiI3TT0iJwKJoh6AniIrD4Ae9RyGA1+p2w0D7vgX3R
/ra/GjPUHD6zHoVR1hsoWLTD/Ps/XytdqtT93/QmdsIPiyqQQFyjEur9LaqA1q63DAPe/8Z8UO+z
/pbvzsKtszcPqNCfoItreMLkHWVo255WpEmBDmPAksfUKw5GeHapU9vFijauj1dNHAilTWrPGw6X
1xF4gAPlwXvohnvUKCdL2plmgG83lcOeVx2RLeg2pjLPE1+P7agaxZxGtr2K9NCI375i+vfUrNGf
cZhRB+TlEFgFpvd9/QMnjJgTPOirzy9mkNa9mZk4gxXXEQ7puu2zFZdXyQeoALhiwX57yVTKpqeY
FBHQDhv6MdaxN7R1RnCg8T6BFJWYJzxGHXFwHERGKqW2XDaqdW5r1XbdynMst1DXKszPXT7Ba85O
3lVjQhWQy8hsyD/fQULLdfN7kLbXzhu+eMgLzw2dZsBKJtNmn2Pkngr3zCMqWabXJ4s5bO4SX/WP
YwEKoMpz6zY4mfrrjWMEBrcUP2o1UICYyinTbJ0cZl7KDfMP0W3jMvvYu9p8od5z65BPcVEHozDf
pqUw282HR7iqUqTGccveTDg21roFjk5TRL3awnPqQQ4+m0iD+yEb6/kxUWbH5e2XZJD94vTbc/Q4
cMk92z94vDQT7ItS/Kg6iNTv9wPxk0vouExrNbxvD4DvKaZB4yTBArLVFSI9VAAfJ3cc1H/cEAaf
rvzxuedw0crKFwPjUNgjQpQUooTkRXo9Bj29sfPXHSusRRR+nyzWWRs+Fn7k4VoqOaYT8lEyM9dv
340atmitiNP9hrN6sWBc6WG4be43+Fzl8tr9btgH8ZaiRCOUMAxhLb6nhIumE5LNwYZiSq8yRAsS
dgirGdLv7DTAb/ahjvp8SDcwrSlJidFz2t08Z/uFYi+nrDu4B7KB3vP9g1/gUIhhtHeOmf80qeJH
tlR60LxXfmKiXRH+4SswKVwG5Sf5JxZgHX52O/zzpjh7tvzqHM61g/GL8ryF8Jyh72ud8o1kg/Wv
LXwz/5vuR7A2zqpV1kD56JVaqAb4BQmPwbpUgjk/lM3MX7nW3Op5QIDdAB5755MxQv3ZS6KrKCJY
f+akp61Hv3vp6wMUKOe+17fO/G09t4smgwXiLOiJneq3ZGkWErRvbLBO1kVlxzKOUALiLRcdGVOy
qok4yrNZDPWEAPHNW+HMo3W1+UU6GnMBzbdHwk3NkLCySBw7hpnN7Z8Jezyp2+mxdSDkVKT+EapU
OynxiDbu9cqoVJNOtEfrUwooj5M9mxlilnqXt62pyYPRJxrd15bXPoFY1AtHC+X0JD0lnj+FIup9
1b2fI6RrQtGCUIA6ArW/KHUscWuNP+kYrl14POEhvyOvLbyNJ6PVC6cSt/fglEVrTnQLH6UVc6Za
7BSSzhBl2EMSWcfOYMvLi84c5srjdo2bwdAmG+NbKQhuvlNRH99lS1QTIN86Ttu4OBm9+N7Ctwfe
bePL5XlyLvZTBoWjkFP7qE2f0Ygs4unPL38kaVMMw/YUUoO5wVXWwjbt0C1jk23/vBvX3Af48JGb
dnYy3o/uFBbczAdVNyQokNIv0wwkU25QI8yE4wNSXPqk1l2VfDPVaEQ43CrWl1FOVj2jfPd1qBuu
OOC/GUqA1+cVK000FR8QoE5zsITQXhXndJ+y5PXFhxn/yEY+RXoKxOEgO0ZnPTlAwz4VTl2U6nGV
FmyzXSbQNO5p7ZxJUGxuL3DoPerBlsf1KDuQaskul1NW335G9Y2B5UpWEiuvolWZSeVqlqYo6KlI
jP4kWlP+KHDl3mW/VBMZyYFIQH3CxbsaYrxo+jJyVOOCTncATRj5u33xocZMZ4fgfb65QKivaWaL
nKhSX3oGFONzGItZl7ci8TsDZdAstkxpoFrBldHK0gaplmYOYDWGmuFqxpoR9l8MAEYv4MSWeVgr
vXEi4IuDL6Hpv39HQgPJ9A9Nv0ByTYzfkM+6n8Y6uvKj5GpeizWcxUgj4QApAyWKjIKqFiSehN0U
qoORtyl9GX5rkQXjB7JQTKtkMHwH/JK3jGHJrt2qw18/Fc9+tHwd0GEmZc+ZDn8V4hka/TPGgrLl
6CPMOG2CVIvRTE0BnmNVunPvftfRDpH5zuqmiLDrce7OVtKT+KVYOkKJAWWRmH5dsTixC8n3vsnr
UX1eF/PrEXlLUDOGMyaeLCzmBW2bDiTubGq3H7cTXrMJi7MUA9NKbrjkN3LirFoBGN48Uahot/Ws
zkFl67Nk62i3qqS9qzypBS2S//Lx/ae04YRxCF76dZq4gl0Y9/e7+dclMRpco+3XLYW9l1aQMXRa
qjdY77MFxFLKYYIgBiv7XrCmjrWZ8R8bWy5JKKvKRjDQSVP1neN/t0fJaNftb43uoAkGLvUrbSgm
zrbEndgyVc5SArlO7Jzrm0ohNJyGLvHRObR0ou1FsYvi3mSsPCVaiMxtL9JvbjmLffcL2Ekyz+U1
M8PGGFNBUCbAOJo1piOZxG4c2SuJBUYtKXnQL8WpS7JXp6NPs1zqbKpyug3yr8DJ7HXCvvFjv/yj
oTYDBq6Zuz4puUd4szIPbfuE+TmzX9R+i6qydJpMx4gVUho2Pofr0joVC7ncmo7G8Sne3CcHo8RS
7MUTbs80hFLzZCTGq4DX8Cql1U7kuPDdmzboShLaV7zcH1TQRIQJnQWHLfd0teP6sLvjna3KqEF1
9+tWmXa5dpgLyQRyyUd7/XvMxQl8TmbTJ48bZO85AeCcodDCOqBd7MAscAU5UzeAbQZerUmregej
6e4iNuYHIfqfF5qGEDagcZTVQCjRif442ZQGk3+hoGAfzlZIko8LmAvHew1G6g/RLzhvp2UN8gA+
RcTnhjDYp9UxEXe/b1IK6aFmHbcf50e7sBnFnyVeNVggUwBImBixeylTIIVmfILzg2iyrcpe9SgB
P2Tw38PqYTvADhhcwGXIhRRUvl8wZ40OudwKj0vuUa7IhdWNI/CEAjQE6VWOrGXzpn8fwBnVUYEk
Mqp8neM2y9wcuLtsM4yNyXbn3zIDShFoYiRDQF07XxDgzUyqrKK/Pwr819dLpye/msoh3ihkHlPh
7dCNneu9Wk1DGCa34AesTRMAKw6AWpZm+3zB6rD/jzPI/40pHGBw06Z0xEMHCnRQ4L22ELlOk+5G
14znNqYyGYRFtORG0GCPo64gaFNqu/gef8BwDQS42YN9p3mMb3Dr6OQzhQvLNCVF2qZSIK5TtAUP
Mb/Z4v1KxpKX9Nznlj/1XxY23JN8WkASZWmBFryeUfao7lUswkMFXhP9/5hMJV3AAz8ubDgxXAjX
2K6fQEUQ3JB8ln1cwLpI0HB2PrMdq24XHchUVkEKRkqkVB4HDXi5Ajv3fJtclMNYQatiR2b6boZj
fvVNeWHzZ0tQY/62Vr0/C2JnDrI82W/vNElimQ7swGQgvrNIJOSu70sH0EcF5bceTgfwZ4nHXoFY
WoII/Q6g+o8X4tImF3PMUc75q0O2pLovxGwyklk3t4UGdvbCxpabeCOXAzO0+0mALm0pJpqlRTm1
FrZXHfp01ulvv2wxk02OBQjB8JJVILM1iifk5RaAtnvlu00LGl3kvHDC2Ax4ertO6r6m/1uInjyK
MBQzMy778S1iklwa+WXiWf3UsO5t0mOHJK8qrl381xqZuJFVFevkdcbXPTgEiIk/h+GRuayFMQNn
5JjXkKpKM/8EEC20iMwE6XoqqOxVlohO4DctKiTg84CGDTLcY11cVzzX/fw380gfJXE+ZrLm1B4i
W8UUOic03u+id6LCiWvh2WLWnII9/tSF/1Q9A/I+qrZr6jLrgOtOY+R7UKagZglA/uI4S3jqvMIV
hDKa4jjQG/HHz4XjUyVhVZaHWON9dc+J16riDG+uQQR0hOSeij1qp6cafqxshuei84NOGvitkSvU
mUBSvLMw275scaX9sEGiUc3n/ruAEV5YJPbMH33j0ejjDdYR5N0vrjM40ccCYjE2/IaTf6S7QnsH
YIU56ebJsFbH3ZC1Z22TbWZHoWNM66GdtJ1w3cjsPsjPNv3Tc7k0V2RV5ym0YiVLKRbCMLd9XlzV
KtNt1G9Sps9VN8LekywHyJ15KUoRf+oy/dvjHkaLQHm34TGrgJQHMpcxUbHY9YHtskL0bIwKTX1U
f63kzniH7IHdAQ15LYh/KFTqSMHHOekmt1WPB+TFLLl/D3nWv+q3jAd4W6Hy/tDHiZDhz8EAoUvP
JmkGyrSvuU65AgZ7J/WMVZmUG6wtSEFgAXa9l9NQahQT/bzUbJKr9lZRRX7MMQSj2PmhdRPlK3xf
X9JP0T0QEAOqmJyco1s3h4HxtL5g5QFGxYMm8t3sFkZaje4D0NNut0URRVDAdsQ7PlzJqT9sscJn
sc6EEC4jEdNjO20MQT6unETDGbs7B5So7AFQPLqEkze143TOSfkk+eGzoeokFLQLFGpK3WWuPI+p
3GRxaMM+AXLTt4B9n73L70rgB3qnVuB2QUritJCAVGHai3mAvrH/nZrHqW/qofUfifF4z6qbWlLA
JJDTfZnSGoZ6UIGh6+7wZXO3NKH6RWM9+Prp6SVZ6TWGc8d8gjxuieYklojmTWj/WtxuddgO+cSd
yacyPfN8GaWRIV1h6ppFH1X1dID+scs4C4HOF4WzEJL4Fa2bRI2DJehZXRd1qAhpU3lMPfBIDywF
aEFufmfEN5GvnSOp97KPNXjIlNBoLH3gZZ6ekYrg3pZjCXSSn6i71g3CTzVDUu6/rZZSWt/R0ALR
ddyKTWwUVhR0lvAoLJlB4PKEZwXi6wrBxkD1CijWYU69iFbRw+ls8NjvRgYa48e99ncyQ0c9qjhC
IotXShTHW9UZgd+u5DfYkKUGSy4td0XByGAC1jxn08v52U/mWQHwi2kNedfyDoN5FNCXB8B0vhsY
TK072XIAX1kZElj+Q9WtdU9VTN5FKyZVknKZW5ntVqOvVHaSqf4Tw+GAHz+nm+Thfa0hwzfnCdu7
NJb0NrbPVCKVZgO/IkaFjLTw7f//z/r5UhdH/6wPxwLt+Xq+HxBnHdkDxKPhJvVp62cdKTWNYGSg
vYVZXUpuN9zyrtQkGHRawOzAMJojL9qiFDk+ZX51QIw7JcgTZwikBmFbIf4I5fABYUUyS0a5YbyO
pXIpMhHclnza6tMZeej7AdnIyvyt0zhcUE9tau4hHr2rFr10FNHXuc4elyb3bcXwxmiTfl0nBYlK
zwd5uemP197GreCxxWzQGBvsnbnWMmJrNBH+RJCqx/XCMY4M6fl07aoMtY0HfrLD4EDCJFf+QnB1
0Noqa7XwWRRDmWJzO2/2cnplBA6EzmtCOVSBBVu6Dun+5+Ki+dTu63r23XKtL6C1k4o5KUCB7xE2
loWraA7HemIY6MnDmEoZRPaxz2pXrLWG53FPVkeTokK9QgQxJ09bpplWtRdePyTRaG/znx6nKqlP
0N9RiuFUxvg7BP9BjoRgbpX4Wj+wdtye9BQUrvji3uAyap37sZSmzUYweoTTd7BhRpd693dC85nj
O1oeepBP1p8gQCSvW2ratd66GkoO0Kkc4XReBjKoTaO3pfKxlPapzXDKBVQytMQo6mt/PjJOsr0M
a7HKWW64E0HVAZ/z0BkOrmHnjZoeiF7b9TC9NbG6NAboP67iOkRHfmKV8jv/gV6O2kd7p/pQ+yzz
tC0ZCYio1ELnnejJqQBvqRk7aDnO8KgthGkKRQHW20aXnhsNRTL7honoJ4NVdSSXrIqE2FGeEsIG
Yeqrdg4/9cZlE7SjKmMstmI53iZH0n4YOQRTFIr6IDeFKBI6qwIwXf0QdvKR/pynIb6rqPKXDOWl
8B9WfGySA4FvPGoBVEf0GK2gjtZUmSuPw/SnJ88EOgC+zhVFZgX7anDPA4KA4Ecfmvc31EX/dMH+
9wR27t6EK/P6al8n/WwTqM4ac4Eh43l0U9X4roQgz1OG/tQ4SazNizvrVm8bm4eGrnhMWZEC6T9Y
J4SzrCU9mS8HAub9EXRp2YZtQcq5Cud1aTEQtJS8zfqm3Stvq3jDJ6I0KRjLX9TogAPxReIVNnLK
yKEj383dkNTB3CVDXJJxku5dQn3DW19bK7GxeexlEqRMN4HPE7qWhfNwxuY2KVKZ3anzAgBpmlag
omuJlKwAIXCo/mfRKnV1aL2LX+/YE2tJVPING/s0r8iUtVIT/VL/ath3ABBIbluasikq7FLv877z
rMch2QXh8F6PERMBcgWbLuVSEiZLTxHkqO/Utq20kmd/hI0F0e+mG/m4uwXHhudUvmZpN+eyUib1
EuWOfJganq2GXR8mfXEwiLkjVNG8pBXUzBuavGJviy30GoVc3lWgLcACJX6SK9FwL7hb58bGLZ/2
gzFqrPh6OR2wl1Gdf3rJpEU3Jx7BKv8wwi8V8MOIvWvutOhzvJF13nZGjkDwTApQyK0yZ3fxpZqd
gvhCT8DyQ22a+Q0uZSH/rnuwFt+atvOYa/lZRkBq4q0CJIl4bQQONctZfoOGmUHXOYYCf9kh+UGA
/FXvXbJG9pmczwnzRj6Pfd7cNpEfHDVGXsJERnuZnptlPAS64l7mpBgIrMiiGxbbAeqJVj2Ugg/d
psS6jOVEFn9tGlhj7yHAwHYJI+C4bXfmYzXjMTw6NEw1F3a7duB5pT6poGTBQNxlnXJFokvC8xtr
0duVMTWKaKBOR8BsBIcE8/WSAZKDlKEIN12zbdpjtzqf19I6qIDVOJgLw5K0Iqwt5rgFVbizYV2P
+a6jizdPLhq0sJpd9eU6inEMJRPrZL/1PdWgM1yh/OL+H200Iiw6jlKJxlA2YTBsMDl1QYmd5vLZ
V/bomcHtCIOG22VfKR07seG8qrTEdMlggheTeCluUUn6StZ84rrZVbcV514X9DaqgqB9gdkdfqmj
qxXA2CPVG9JCpVJT5xCbg17/AyqV/vOMNeEp+pJ/Kv8RMnqsuFDKi33fb2J3KEr+qGWUoYsTjLvt
YrBpNSxaqxp/V/SZ+Gw38uyDaHLllR2cMH25UwHuyuR9Wpp52CHL3yuAxbVziJtd4pgWdJVOEH0g
yWkh/5R48qTDFhcpESFiHPN4KLaC9T1GWIabRB6BhBBiSuzC1V4JnB3O36o8SPhaQgx17iWbivfW
V24rS5NxSDSbRFwld3RcOEAhq8SWtxBiwCsb0rskK5QHtR2JsNbPRj3U4eQDh+5nkfASIEDgIW7q
bfkF9360X7XZUg/ArAJ5Z47nlxLQOvn6lkgLYuBsutOlTl90PMMH9TxGLD0TUZANZSNUPe/kK2gw
8M0mFS4muAM+2T+KpAULlza2pHw3u9CEtiHxx7WQdiaDkIcnAKaF+3qaJkgaNkiVyHOfJfbnqmpe
orq/UdnpTN4sA0x1Rkv8xL5wW96emtXukX9/C4IUOMpnz92blpNMxIofkkscBxuUjLuG/wyjbIur
IBKA/5G7ItSH0JkIB3IBlWlOr4Iuxs96HDuUcZHnU2a9I4d9dii8z0tkkI/rSa76gzxLr6aQcYCm
Y6+C0NbUjSFFZrQvJqEuKF8Igfvp94vtZB7DCmwKoTQyehtIQS1uPpQGHj3uVlFy98wvGrkC/uE3
DoTrkIgYRqciFWjzKAum3cGNZhFZOKta6Aq79FsC9bOCbG7TkrKUWq4Y04RhggeBE7AwBbCa7r1C
j8F8c95axm0HC36amL0HOs5Jbum35B7529dA7EUU5hGHOJ9P4s+1QvqKWV2SM6+BUpF8FrANr9O0
aj/Ged75T5Owq4AydNF9BgVg5hMraM0vX5WBKfT5swBlyVlYbq7H88klIpjnNDCeT4Mgg8Sj/7hB
a7v05Y34uISQ54/ibutMNXtKdvebyoilMfK1/4/IKlR8OHYmm0L/yXPSj6kyshBXwpNXI1ZDF8mR
BF8AhblKgvi309GY/PcT21KI52GSGgDr4jP33wf0iCb8JJrpBVq3zUM1KSGraMxvwmWr12KzlGul
xwv/M1RAEX96O3WvRRRJoQw8BZzk753Q75zZBfnP2ycsZKnUxZLOIdxO/aZcRewkQV76U0XqefxH
eowOQt8qu9AOb5uYWOlX+TE5ceMCLCMd1JcUwqtWtovjLBDowDV1vUH/52Wo0oDMzzkt5ThQM+wQ
m0/OYNCV/f1OF7+zhN/6h9fV8uRYcUAcZj4mvrCy7q4jdNmPy7AxYVx1gvkKcB1fEK1DMyxOJUH0
0zShT4IBEQ55sxTICc05PqQsoJa2LVxUnW7gvy0ls1LutGGMDpb4Y9gQlCTJJ2WPo/DM9EZAvgsu
L/sh4gZN6pfAZHiO3WgOTc2nAxOfXtLyf0clT8N/xVWMKaJyZonBEPdc9J4L9joTxyLI0BhiwX1h
PZG4vVaS6EFJcIV6ctupa/a3XRamyPBbZ7NuqglIDtMgVNAtbyNgUyrPKBeRRqAWmdLatY8Wr+w4
617n1Qb3MAIPpL5M+XgDN9PG5PuB1gZRN2vI96OxZUrndcua3/XMzMqumBNbzb4/S1WJtzaQRoue
l4K8rIt5TBXY/JOIbbEDEa066dEE0memXCUEKpk5YCSJ09aI/HsJNUhpb6MO4WIuN9Lt26QULzU1
PDWhFt7UXiSiQLI8eXOoBPbSLNFDkTuseEtqBXQUTQN6xHOaoFcLzsEOdDiMv2HHRFfZ+puz8KZs
v/b7N8v1+a07FIxkPctr+t4RJnUOlBuUWAnrvAdOM8ayQsmGL4zB4NT/Ayo5/9+ky1qlW8nYxZ6K
dYKXl2Aeo5qt/2DVRB1RDjgMrKN8DGBeXDc2traqYam/OLQKmCUhMtdq/khVQgXermVVbCN7pU7m
GvvlS5mQEBRH5pHC8dZng9DhXkqkMZtcXXsFPwfKA1CMEIj4jA4NsoqEBddFsyy5zAMP3sfL8ekU
y3Zj//c4T7N1zge4IJ4zhO9ut9NDjIuScAviJaC4ymMzQuDvhrmXt1fSVkdPn6utoJx7c8BvkvXX
lSNJmOwSxv1xeZkezZ2+3SfYl3vDFTSEvfiW3F+CdJtHIUDrYFRjyrQKzM0qVUr7C9uqJ4yKP7sl
Fc7z7fmSGT6fX6sFBq0JBIdqEGloHNmxVJceY3C0xcx3O89SOSY/WCeawCd1XaieoLrJEWX1uXHM
OznnFd6YVyi2KGgQzkLUjNmy67wEGo0lRYMddHcNPGDCgWQChqUDjTCl247SLAYeCJ9oGVeAGnab
IV2o3kDGnGqcrCY2Xe7GcWAVGDO8HxbW6XjnJ7aagocO2fRBYhEMErggBntvTLDdDYo0BHDpM4i8
KQOy0SAdEGZt5ftuKhHH3XfHDD9MzFR3P6S8h6aTQvev3EkwcHarrMBpUfj8eGpcS8MyezlL9gB3
DLfi84PAMoAjAUXkBrACEaWaDmXshnCtHjl/o77OV4Cw61My98s1NVLMtiJt12DltaDJevL9nZWK
aOwB50UC/OjSjsaSiqzxLBiVJm9QVYG2AcZzubnpQr+0zKoypmTpXJuXc+JzhhvXrcfaEfncAHfK
qfxct54fjODqf9ztfp+l1GBoX9T90MRe7dBaOFPucfoq6N2GlcGOAMhU1YFSf34tUCfM+7AbpnZr
2f0szUEKIwpGrIJtagO//zSrTeFX4n2/JeShOtCRvhykxa55s/zB+t2ivTDqPmOY3kWWIZXjRrs7
5BdfxDS84nauy2skDLWnWeOJ4sFmLOVCpUMTCwm/YoivXXAtZuM1rQt1iGLC0ShTPTDzp6xbMM3P
pJdiwRcifnmqJzerltpvYuJ3g6Q2TVYQiA790RJUDb5DGF++9tAvnD2t9PIU6lkwGgS28fYBRM6S
iFnubx1q7YThUc0CWKlKFXcSh6iMp77TQWg8tQlt1KYq/6NKBBtoIFfKMSdUZb3y4yq1LJtZanqe
qMX31a/n/DtQo6oyjs5dJdKzezvpG2pwcNR63b2lxjnJ/QtNjqKZjhNmCPtdk1CngS7OLeged4QK
nZFPhuyfUutURXfFR+xZVbj24dr1y9F6MhJnnBU8MBFpyvHNHt9JmkHk8/r6+eYk4pki+si5bUMF
nsRuTPOSlsAKZdJUHjMiLUh0wTmgxAaJvRi2+ft/RaEDAvOlQ1kdd4oS8/mXxxBVWy2u1YgO9Qxh
wYpXh0yEbWM3KC9fu/9GBI3e/12UBY2RPxfiCDrrcG9BWnDuKCNMV3+9dcFV8TGu0gLyd6NKpWRW
eS1zkUfdgaALK/By2gCBPrWEOq8hvNoCajWfoULALl5wkccfk4xJVMEditpESEBylYoYVyFlxQIy
x9SVn8b7kJEw/F7F2zF8YVAsycZ5Z9BIiSyqJBPVXdqnuL704cM6mP07Lp+6a8r1mMv7HIESujUM
ITZ3rf2tPrdSM4rU2lQ4xqJ9uJ0wlb230iRVexmyZjX+Hek4n7xPzgKw4asy+GRyXN/jyJPRaq5U
6c+B4GV+8nWu1RpsZat2ip8mMNUf/AygnzzhFABFTvGowbA22eBIGq0DrPU5NltFUAy350QvhHth
/IuBQtv4rIww07NdxwKySFXToPApto/ciE5NkfZvNfZmz1B1wwEE3JQ15T6e3qHT2naTnBrKnHZ2
5Qs9cyX+b76sDzRsgqfpo9ZKz7+R+LH2DoHLdvuJU6IkpioRr9P6OiLQnJ5LJtzv7d9JoJNsDZib
jNH7DS0lv1reu98waz+CIKuM747ySLjGtPvqPrdt1xLOPWNyDDn11sRXjaflj+5/+2aF5pfGfnXK
QAY52MpXA4aq9Vvu+BESCBhfDUdiPz4E/LZHjn6zsdPT0UC/pOfA/CQHogVtQjKrOryMQ9Yah/Bz
b6ZSAiwEIXRdhbJOPLn9MJIas2QfkPsJ6dD56XaQ/mg2pNEgH1voDrbXfom7hhV4T+IMM5QCaaNc
R4rEpzYi4ka4E2CyElK3nYSaU+PjdFC7CtNNumByxWaD5eUr7wy+pfM2Z9oTCychJGSQn4Jd0tF2
4nvWrnl+wLWzeLMZODFfhB4rb0TPC5Z+1nRa7XvB0kVuBhvKWP923D/scOsI8fgkveOCjmO6DL00
+IpjP5QMvyzFbF/ezYTnCjt6mmdkn6JrTD00icnXUnHbO0ypV6jRunixamwK7PISNCRifUAarqY9
uasu0b7qnZP1ObrfnybhopxAz4IzKYlsxD9yxulNRdkJXrAzEJMwz0ifKYzLe0Eh/QNLof/wqdtL
Z6NJ8ddXtFO7PKo+bMdHKR7G/sMFHN6ffNmhi1g4FBzySR1haqUhnU8Q5fWArQoBaG5d47ambwXm
qd9uLjhV5wbg4syiSjEiov52ERC9KqytAUOcH9PhHchHC6DbciX+vdh0hzdzkTw96l+TUQWjBG4J
66MCNFKkwE0OVYrjedZ80l/mkTnmBkuztsrZZ9CcMjoQCVxEdYNHD6CWD7uJTylZ9TwUI/OX2pXz
z5LnhMj7E9oa7oaPfeYDyuDnkBnQMaDyfKfj0VKGn5C7ul+IY1GrfEsX9U79UhzHVOVtiYE3w922
0dXSeSzFqPE0XlzKvon9oDpffVucUIxTdIft2ZhjIivClYEpxz08AC4+DyHE6Fhx3qzKAKEwXPHA
kJigTCClERWWucDFnrlr7hewN1Dkl8+R0Eot7oI11PzgReIHUtmwgi26Dd/3/ikNAhJpavoKE4bs
idOw6cT0j646uHSz78Nq7+08jQdeyByWGzpW8btjHM6Ln0hJmeb0Mes3sP71Gxb2q73dmMAqE2fp
tli8uJEvk8T9sy1stYGiGSeAZcLJl37eBLjsnpw/RG7ezPnGaXse9UBz77TAL4BQYIvG9uOwKRy4
Gq0pdUZFxJ0j+qnf7cjWcRStpJ9ffxQZsoFgtTRTtVDYq+xAQ9pyYI4HmNUA1vJIzethS8DFKLxI
PvpMEB/YIgWy8ml5kL0FKqbifcTBCPTfLr3Rd/jWMdxJrPnEcvsaZlSKuargtdvQf5Sr1eES6G85
anWnBdDeog5bEZ3zQg6TwCB75lX+WBQ+H8HS/fDWWp0ybSk6uuKaRPJVdZbJ0TnkU4iWL9HE5KTn
7YwV06d2kuce/WGDcomG8Y2Jd3q143toutuYBHY2jYjk7F73LtHGN+x019YFhWo/RWKiyss1KA0E
B6EW5KH69aQYZciJnwLYpRbflkHSBr+2dt4lLe4WKec4AdKsG/BpUcpajWyzEijRFzEysid9d6Ng
0bJiCNEFKpJ7q5LnUSNb1D4fV4kRavIKc16+4ELjYIl+cscDU60bwSP0HbvxBqWL9b6SWnM4PLHA
jYfHLFQBt+NgdWl+ZqG4zLpq8bkOzIu9kcgeqBUOVYiFrWkfcZI33TakkmEYrJqn+D2B7oD5Dg/r
h3h21MpvykvrAFiUiPXozUOMp3LKwjrI64cIB0jkSXgDrqyOZlejLTHo6Je/dTQxNSA759dx+FpU
WW+tcPGNaW3WB47oh7GAD27q0Difk73xPWVG6o3+7ePBuyHVaywGkefTaME9+MUm61GONd0DKwuV
xhJpCuiMtcJeH9kU726goIccr2N1xmwANqtHfAOjJbix8EKBYOq4OqvX1Zy8RVw0Db1Q6Ojyqhch
MsVgL2jjc61Y9oAe/XtHTjSMd4O+MDFwrirGaHpm37ewsYKsEazZrG0/TNZGDp9C1lbt6KUdUIu8
tX7Qroeg3osdR2MCSkOt9OWbJjadnBrLrAv4u7JatGDiSQRljUi3fq6th0ei+xPD62MbmTaAMP4W
LcFuhpHhglLshbWGz/YxbSpwHlXBKYt3L3/1HSnhnpiAO6tCzvk+5HwbgpKANaKsSyNu/OzTLQBd
sGMA5JiDaxxD8a/EcJOhkDdsaKaQdqMl+fS7pjbN600QyeKj7to19jdVR/bNvooWqNwe60sDetXG
AesxD9sE601qmponmqU0tPxXqU8Ctzcz3uxtnjw7KzK5ngGUZ+k8uQoZxpw/BQ6YwO1jmcwEkQEK
J0h6W2C+ub469ky2PxEAyUlDaBR5PJEAJ4uN8WU6Cs1LZ3BmEh2oFhBk/lFP/1Hk8a8bfjJttaJr
DFojAOsaAUelZ/121DM1UwMvB70KPFaa+W6t7ZgQUPzp1R3a+xqfXMXplK5AUUYHAKyHLXF0sRyT
4kQyrDerzEDtvG1aWxwR7qQVybL/Xy3RPzJco7z13el7zzw2u9NOPhwJkdIb8NAB9j4XzQ5deXHV
+5ggazmA7ZBarsuxX8qBA3qPwtz0rcKyPTbYhooWuSqKJRthf2tq54ka0SDHw9GHvCUkjhVuYb3L
cQYoMiBsD6v3E79wwjzTesLXnY6aMjvkIjIGtu2Alz1I0IOfBgXo/OWrhg8R8VDcsH6LQDA+ri8R
m1OV+PpMFCn2c9Al09M9rCj6guxjJTxcaGw5GZU/DCMGUo3b8C2gpZ58bwY5+GoY+fvE3VKlkQrr
3LMSECF6lmsxNT5iKSiqZj/4a/4H2VIZqNgR3p1i41CnZP7Q7Rf9IWLwpmyRrD+d/6GQbZdO745k
FTPSr9Dwkktk20g3ahWCfusMXVPH1o1ED9aaKswhEg1Q+HHQYrSCDtidWRc+i4ELErFu4Mtq2E7u
akQ+UvtN1V+eSrh+qk7VnQ7AYvnMdc+YK40ZmLCko6xUtQ9N2A95BEOlH1iO7YOywMHAU6an275a
YKHi0cBVxzF1R0988a46tlq4NYNg3UxTePa/8ZZuRbDHxKbigL+akcCwwVlh/PGo1qll5hvoloQr
w+RZX5o5HQi0bMLgiqUuRA0uHwKHGGh60dJq4piozWq8iyBDcniVWoC6T23a5lmZ317P6cMKuNuY
xPDCooEG9jE0COPKxpAimuOqAbDoyLWIoxVPR5btgaEuVXmCeA4vKyjamwxhadMKj3N3v9+o6dDs
sUfvAzZ/a9MUKXB93SRonL5tzrOMZ10ols+Qrgx8YYuVEmIyYUDfGca/LrjuSIQZnaKnzMrojFj9
AvVv8NFm6vATd6XW6Bl1QT6k/EM9qg1SHsh8cvizpqYDFR12rM58LBIh3Q4lflcH6sMQk+SkLh3f
1+zdJcuynp0I393wO/SlxPrP9uXtyZfP4sIEwDAyHz+KOc2IuH2pC2AkoQjX5opml8kG5TxIAk9C
wb/ayHyHqKK4XluhR4VGW963UzBiDtjPIiPJcgLUL+54e+BKxIVnfyOnDfL9tgK9YAyDY2Hyq1C4
oqUn2xqV4Mm5g0TpwBvQ+jFhNvUKenBJGjHdATZzODrsvnLgV5NcXGRqT/BBxnnaMDCkShIx0IId
FobfkzUwN0+goza94DJF1bYzI6zRXSgpjWFpxDVUe7vZ2oHJoRgtre3s5sJe7gWiV01jszdzViws
5TgNhsDlQl/Gwf6jogwIjrQnvwCRCpHR4TiTYbLJAiNCtLC7zgB5suw7pROoT9dpK31cje+8icip
kEsyTDFCZN7OYUsDHQvEsvIePcmoZiayXDnzWEnW7zmzCohUmwd+a5ZIxxrPDrDmjSGV4VTnWb3/
8L0zVtdkkIiJT/qjUe7po/PWiW7enxW8jTztIgO26j+G7UygOEAXxtDdh7mWYFL/GeCSes11VtpE
5alxLT+KEaXCPk6253eDWrfXX0CoceyKLa0kvidqphCrJlqUH087ypHkHxLh7vvUkoAZpay1wvbs
rwy6aB+7OIQJt11yQJ/xl4DkQosxOo3c+DXJ7N0jkxHR5XwOzd+R70Wb9Gi3z+R9IrL4BkkInvDp
ZKK41OSq6iCR7nfj16LjIMlauQz4ZzhpiOmGKCLDdS4WzQ+EJIySmAZEFElnzPd2spn6QCLR4F+/
DTGJ2igl/OSfmQwWGKIm+cBp58kAZMOi8ukjmwwumvax1VrgFKVNatXLFABHgZjS74KcYdmY+20S
LPakc4/THSXPsP5JU3lGmMPrmQiLSvud9IGhrOM+tcAV+Pxm3LdpczuhQ6i+O8N/K7lDmuW/u06Z
61mts9u0ej5Kgf3i/NHyse/d5tbA8QxnilJslTypJ9QGnjNgZN1ybc5DHx18PnrYacQAhcJrCq8x
AuGFjBXoT34tcqJEQwNEfnsgZ7SygQwuxpJxKSI2lJy1nmbp9mihv1uOFh6uzTengHTYFd1DbXtP
vYpGr8uMG9UNIqL0Oa9iHQgmgkpTNKqk9Nz84dnE0dmnVeHpouE9LuXjhfmR6RPmzY/eIYSVG5co
uQIeuslcrUs8WaD3kAVqkF+3F5kCQWCUW7RovzOq4XVwL2apxI0SXFP6kdeP9cbNnoPEfe1VjMOq
9IyiYWMlhPkR37gy4S7NCtzeELCT0OGp4AFdv3/5+cGQ5OmrPjU9pLPxC+eYheUXyw5x6rtsCIWi
cMz+AgqRncy9mjD7H2A9PEJ3oiQ3MGvWh2D+nas473uwFFBv7zNDHtxyX/5QPgos2bOf7RLcMvnU
HgZyTagb5qVLcp6GjLWtrYJYX121E6udtwUXRAlYjUtodMkpTAT/pFuFFjGCR8i69bqO7vIRB1gF
ah6lZ35Xi4C5D6PVQMHjM5Du0bg8IK4sXdZ75EjbvxtaTgrzZHKope41S4YzTYnfTv0S5ieMyoCG
xPUDxGdyRvokj6DgE2Ffc73OSDrrmElwHidWz+ziPwjiVtz0kyMHO58UCD+FhfGuZY+34s2Cs/Gj
skJ9aE1s1YvVkJ5OkROV7cuUnma4Pbi1K74vFh6zl3mq5DiM5zhaxjoWPWEuW1PpaWiAduwFdjzV
eVVQBfLZR59fhxf0QnSbHDswZjJ8cptQAReaLkWhLfZoct59Fr+es9KkSJPGASVEp4etnYDBlL0u
UxgTxUhd1hyiBgzGmMp7TpLdIafHcZlG1UEfIgDhxxYFHJiXL58mcBmXssEJHfdX5nHmLH3gPnXe
l2bgGZSz1Ge/z3Zgf8mI8qKWVLoXhWmrzfkYa/lWviQnbrASrDDFnUBxGQfXzWvQTLqfmUsh2RMO
b0W4tegxWMbk0Z6AxL6jWIhTtcHGAnQmfvO7ClBc4kLKOdQoaIuphC19wLGl3K2d3s8wysJfuHbZ
H4BweMl7uuYbX6TK+8qAU72fYblJ9GMPBYON4xmB8WyBfDba5IT4G7QGHs07mU6CwNzuNfSfCzax
xCzRot0fvLHvIYpLzd/19Wq6pxbSlgj85X4ClNJpUcGPddPD47zH7JPZbclX0dMFCPecFUH7kRsn
naDjFs7gGHmMCU4LmxSjUniWopmUxxWu8N+v1EIdZez9Ku52nEA+2YTROqost94QDhIXno/zw8Dt
FVCHTHjeY9lKwLCxYXjPV84DaxjGZACsXRrBgS4Q0Ja8oH3XPy876gJBTgIcE979QayFcN8XqKw7
MF3n35i5qVDSB8GzP7qTbJpR2v0JkcdXWl9xh9Q9jA8UUCjtdLfE4kYWf/2xGSnQfhjegMJ0JauX
3RpPgwc0jnyZjEGX1JjnAdCNDrvoFzVL5C5xY/stle2ATI23BHcnZLv1gBelssycwlQcKgiGQq+8
hxOcnDIgbIl2GuX/0iPprrgP9TIACv0/cqcIJwjjOc/dn8bZoLtERC/i4IPjQO/I7kMAvy9WhR4V
zGQ6htrbjN9/BzjT6MDBEPmtgXwb4Tccu0yQL37tBOP7OVCJsNJHc//0u2IRGAHgMlERNgrMzDrf
ZBzyZzKbEM7OLQxf8ToBymBtYydsBVbax5imXAyVRzBrU3vuE314b/FFza1oo6r1I6Hb90cx4in0
m6yaQZ9c4g8HqroXh5496CaICEqfAx9HeMIgIBC/6HhClRxRQ5WaKjtRAZPnWXXkPm3Ykh8Y3SEd
BYJ0OJ6q/KWjZugG6PlgKwgLhXmoiP2O8u3p9OyRwdCjhwREMt7la5B9oe3m0HucZshE/HPJVLYt
52zdOLEaVLwUc+NzrCfaU3epFzJcEX8GtNsR2mqCdL7Arv5YrVqfM1+qwI0bdoO/0M9a3MsMnTti
IbSrMgqRWhg7Hi59Q257anb5RfT/dLsAv9wjJ3MzQgB172RNLKvIVw+XZu09R44vPRfCLf5B4lzE
WL8EnfugyoxhW58hPpssGyRb+6IYjmR8tnmhMBzuBCwM95+7E3UJBFgW4n9uHiF8qoAQwN3zu4ap
Flq6HRJLAQNpiyNfY4bV9Yagktl9uvBpw9g0WcG4vszfgZ7z1vHRk/nLBchn/BfEttJLsED0ZzAo
ZvhUn0oLN50mprBFss64zYcFwaA7xCigN9nhSz8BjdRU/pjs1d/b0KkcJ+jpVbGQ82UXpstLcpHG
Thv5ZfaEQ/dOqt8HUoUmrdZPQ6eE15GxOXoz0hOs9r54CiGSZ4Uvn5ijuf+3FJZtHf0sAcOW6miP
v7FwqxRRTZ7iAJbD978YBGBegUrNxEhE6n3v2mvrVBQfhQyTpYuUiERAL5Sli+vnXybrCb9ZVy9h
NilFw0NYRT10002tnBt8jsm+MQ61kKx5r+67fBZzfx357KI7NepIUpe0R8r6St30hCcGIaSSHpsA
ukc07GBxewM06rPLUr3FL9fCHIRBHwJF1nY18VzrJhreJfQJImuK22vImHT+Twz7qLd/qENbCDon
jg0lVi6JhyN1E+vwRHwhyUIsTDYxkFnr3gZq/+8sbo4XMe4LgpXCoEc4F+fn6/Bv/J1t82xVVSoH
/Ak4OvwNOK+0ekGvJdf+E9gVyqO0WRlZTIeC54YlBruEvCdaoZaN5TWOqtOskJ+O8qrPzQXcupuC
Dh+tI4LKooEtVTbU0vzdhhCciVzSSMnsdyMBIZwGf10Bj7ANcMyjk/YzWf2QTfUENuBQLu8kCcX4
I1F09+PL6HB7WpgHxkeqeGbXcV7kB2qTT/ONK0C8wUG0HRBRmqW3AQiM64gHii8guuc4M0eZLGsA
heWsTcq/cE6qVvL3bT+HxsEHqK/Y2Oo6OwAFrTndtpO+QBnk/M0b3gM4m81S3v2S7OV2GvCLcTLz
ocmzgIFJMfs7gzXkDBPceM6O0+bA+EKTlpEkwfjPkiw+v983fS23DERw5iD5xEHPOQ1Pkix54YZY
vwboPR8UbUwkXjkTq5XGmS0hvKAkwPJzmPA70Y3zQjmsWICZbhpB/s6fI8WUYw9vVe46o63yI/WG
ffEJFns5GfKSSn1Anmw5orFzsol9QXojTDPqUV/Rw25TY73y5XR1GyRxRuWtAdln/j+omCmEgJ7f
MvmMXdD3XpKCQRd6GJI5KRlpGjkZ0KBxhE2GE9qWnt/r3LIVpmJIwRbwKNrTvHKzsGu3/hfSZrLh
TQ/nFmEVs4okOifojZLoMNUn1c9fBumTCY4ZedfkBHGtALglUXm4fglLqbWWxfPj7Ad/4FxVdrNd
4rgZ6nf1rSGlksqkEy+MyYZZHuE8QIchF22kOI5g5ilXmJLx1/a2OsGTwq5/MrzSBs0/xugp3niJ
dvDMpOdOWAA4puOdIEVLBlekmG6IAApkTFiFZq7KtyKBXyxunviwAUySDMVl7AVkwcLuZnr3GIcz
3hsC4HP/Rd7Kjo0wXF7/5CemePrNXlIEjixHT+xFleSLI2FpQ4LyP0COXGdhD2Um64giO1IIHAn8
Hh+AC5Vj0kocH5twExt861gzsaC1tPAZ2KoN+pP5bGAkAzncOyZwZVBdNAacubxZaNDjTjU8VNkJ
JWZ4/Q/73FhvW2N84lZP02DV73QLvMEqxI+AyoC0MxrxiqC4Gc2UOR9ydxOwh3wOrYE7wuv2BahZ
uqX+JYpIcUwWht3WpQs2PedO0LdnzMWiOBF1+7yPn1nemskOb3yV9aCS5f0ihFWhDnBiUDq/b0vw
bHbjlCuiXIn+AR0YTcy8/SwWYIIn22XZT4g1BiC6Z67K3Soq5q+GIEsNxuNkP4UO4pIHhOo1zk5g
PudvrCzqt5Xojqwba+j39YkRPWxEsQk2xMKgyplg27/osj6C+/dWajrB1sal4Qc+A78hRJSiRYWx
NIeZWrNnpsyBHebonC+G21zeZXjguFDGnJerxyAYE+dygDH3KEQCbd7pXrDVMGLjbliqXl9Ch9c/
ww7e2E+Pxi2xEED4eUQ2IunLORtfwF1+vJkkiwnHpWhQS+Bc1i+uprosYVNMAOMK21XKuQnWxERQ
0ztBAnnWLpfrVDgESa3vjt0o7WEDLmpoYRHnaQIqxKOb9w5Q9DWCKdBYgo4mTJzrJxlDTAhSSd8R
lXMCPHYJnQj8Zd6PIUwtceSGKUK7jS2jHAE7nLZPAaoGqjaKWXyScjTZBqu5KH9hjHGdp7kN2oaW
eT+fbfmLfCShffgocXgAGalHcEcX4IRAUkfudb3vL9Ox6myADVfwxMFrP7q3/y86tpZPpfN1G3wt
tFCNKg4MXSiRz33oUaPqPT5mSXV9pERnsBkchzcsQmDS4O87P8qZ+MMzG0K03Gih5WQQDea6zJ7f
rt7HE3ubFTgjFHLECYh/sItrV/uKWLa/jZZ5EazVlpuQdQyq810Ph4mz3qKYPfL2g+sjfwg5A7rf
KVYaDCr8gyIw3l1wn/p/g89Nnfm1Wkb/JzLqVGcbz99dbsXc3R9H4ICuC7YT31fb5c0lwwOWUTUd
8OHqEnruAt9h8mWNkxbMEJFI+IS/6uWHdge/5LE+h5BqN1/JoMHwBYcL6bF2vTJKfx5Yd3okvYiS
Y/0tt64rjnXlAYyTTrhz58WxA8caqCKAjgYR+LN9xPijDuSsanEy8nKbuLgRmCjRy3dWgRsybp7I
tX3da1Vw65O4qAwsPbYsea6SlHpyJqQ1xCRd45a28TU9H3sDQoKgrAT5E+XgmJ4Jf0bDCLD9qoyf
u4FqC0OZYBXjHX0Fx6bK1udEqQSS2e38sTQYFwocKOXgIbWyNNPM/8q9kcd7XgXLhNnlg0otOVt4
JdXuKub5bvq/YXO8zNM+UqJG2/4VEDBR7hiLGOEp8xFuT+rIvTtAjJVxAhqreb/6tjObeypmhU9s
dls7vmL/XWIxPTMaxPpisET83T7A8vl8bvnx+RSFIaupyYzwIFzxnDGWO5HnQH3fTeLNTosKGrjv
yH+R3h2Gx0k8JSENtXnBBztwPse6aqRdVBgszGCc49OanwTRFG78ErWSeftTcLo3164bz4FhSWJz
Ov1tS1zyV6gFeZHg9/lBVzv8rNN5t+W03Sk1tBLP4ajbldbfNAzRBThmXSOP3tAlg8Ua7tl1qLey
8YiZJy7lvsYNlu0qrTqYmnnzNXeI610R3caGEpXnUEF2PKpAJ4hemwXII3VyFnOGzFPV0oWLf3OT
AHfgclKKUeZtpNxaGsThQqIxriPBHMkdyD88rBpm9YD/24qIU3zDiom6cC4FZteXixgj19/FRgvH
WXCz/9OOShZH/ZCIz2aX1zhfx87PiRbRwUBJ/vn/K50iLgoFk2bQfgbwMDmuWzym35Y+kIhdMDNA
onXn33a/0oETDR20fb1kVer2lNNPhpnHhECteRZW1w+5PsqrvEVXvo7vR/zqqvHgL5kAK3qrTDYh
jMduqtiW3errMVx7jpVQ5gSKQPWkDv1r3aWPZaWRGvWIWBep0hcb7QlTK+xkUZBPGwDJ5/Mu5m3V
OIgf9XzTgKVCJuxxVCVh1LN4OmwIxz5KIju3Cwb2zFgKNEMaJMrHJJhzAWlPMRFc1g94m0D/eS0g
pVC4hxp6y4MHvQSmj7E5H9SK8bxtGrSEQqkB3g4pn3qJ01gjim1W4tZI2a5ChHRtaajwdjr66MG9
nLJVAphgs+cacwUptdh238dm0LaUv0to9lwxXPgj2dO89R4fRj/l5fj93JwpYgRqiV6KLVYuMLR6
tLXQimVBaWtowsKhoONYhwSxeSbUkR9DrdQSajxgmVEZpn7Pr5ZQSBbfJtsuNu9zP2K0O907OJns
R59HMfjYC/q5gaZ9t4OdRgu8drW0kBuQpL7DFmLsM5nmBVG7ZqcdnZ3wryherTPd4CsqtXw/jQN/
sOsGQawn9ClXi2wNal1OPNaXCCsFNvuXm/+5Sg/N7CtEQOkiuKVBesVdFtmZj2bcoUjygFZTt+8O
BMtEqd31uxzp2/COAouU/mDbchUVewDBzcmMAUkET7bh0nmqrdrm49kDpQ8Le7o27F5dNXHzsI7Z
fOuymAaAmz3VDiVGpxr72/fwyZpxRrtlBxv38WO1z35hqHB2x9H9wYKbLmk66MuWBIae4aDkYxBG
aGKpGDT03vn3LU5fxrNNM2wGQAIOe/movxZjvDNkqPkJUm49r5t44iUzd4fH95/S4MNg7y4IxrXQ
5IzWR1c3bqfHeBi6jWkoSH+R6pV/9KRpgz4W8YI3svoSplCfpANVDZcbH8P+x5iJmTIOF/fDol8h
Gcz6Vy1pB8ZxKnNzMUtdY/zlsF2D0Qkvu4z6MqfU+9eea8BToUJiQWe0YzosR6gdqju/8Pzdv055
oxFWUfLuQawVYlt6jTb+4NHKXrs3Up3Ab2mCRisVuzfZcfvuLvSnwoO0bQygx1MA1Frj1yx2oCGb
vItNjIWzN7dqqIFhmLyau56YFGhvO3oAwoR4zcmBI+Jq/+bbhcESkXVhYiYbZ56ZG+BeNzQ8ZRB2
jwA7gTqZ5S2pkmycljCIRVrghMDWDVqa3qrzstKy7nwrYPSLIRvxAqtvbrC4r7M/r9X3i2L+gsgF
k6Y5r+GzPVr8SbYLLqr+z/MM+GFStqSkEiTjifmpjEUEjHCQjFPF282IZvs7ESKzm4UHBrcN8xz7
WPrNT6AYJb+WYY0T4LJkRi62irNmMnD0XdFPVlmO/Oj7B0d7J643/Zubnxis4E4M07Li0yMdXuVk
ND2pnZUGCHCT4Qsyj2s984KtsWEDjqY592tE0i51TF0mwJKL0LR2ayd4ORkuiteFFvAF2TuZ39c6
+RJxiMEe0miNEcdGQoEdaq05+IIPkjeEg846LEAibDdlG+BXAu9VPWpNdxDvDHKpSma/yZgCY7cM
59pgMEfZkbos2y8WpjkROzCSA+6gEQb+Y+BU+g00YV8Qgr87PAf7cRNvuE2Rx3QmHKiE/fP7IWle
IXyaR3xE0IhpVfhw6YrbaUjVAZCfXX9vw413wG8Q/fP27P00aCxbr597csjX23RMA9iu9pBb5/KA
7+9ahUXB/2nDNngCjQLrjHKC6+MomKLE72K7Gq1/am0Z9HxNoHehMszNyw/wN/n/YfiRZNvZwxYZ
Drd1XMRNDtE+L6deq7l2ngdeNPP7hDZ0U8paLn8KSZ7Vf8jRFbpZUajywYKXM2wNZyUrn0qGWfci
1/8kFUIwZSQLCT1qH5gII1r5apXxq99LY94E+k4j6Ie8raIJBWrHq6gQiWGRbIVrayQ/foRY5/aZ
TqnDHtRkKhmxN9LP/2FatX8ySLITz/9u/hBHebUS8r9fsKh7jS9WfC7uaHkbzFGeTgvh9FpVl97t
+yy/wCw29LMh+j1Kb6xTNVabC4r5SXSYrKbCQFAwI4H2VapPGEmrkZgcgj/zEhuUhqfg504V19G3
96rBOFCt3KwHfvomgwiVGe6ca3RYDt+w44oyOQnV7eNEdQ4Wwy8SnWyqVbPfzJnzJVD6HLNXcHqH
/HknyO+JI89ezFrJzwD8i8xA+7cVHsiwNpM6QTJK/1aaYenppb1p5cFIDRMAkCZEPXJv+ux9UEEz
Ld0yjBmpxOXJhLgWCHvgM2kH/s7FkT0AzhrV5Bw90pyJUep9jpqYvhZiM4t/LbaEFZwD32uA3YOb
0el8cPclNYx4r3AtatkxUNt1shbwOZjiq7+rhe8+pD8unTcTwk5nT37bkcSokKR1UQnDqe/vAIe6
CbRjBnCfWNfYL8Jk0/kRART/EUWXAfL5/nHO6ZbYUuqPLeQfw4Kehz1dvyuUMaY9oWgPFgebsX06
MWAweYVbF9mbtX1eaHI5w1AeD5VFJCG7wwKlpGRHv0XgxS8ZS3cjAJaaiG/a0Hq021FpvT8EBHky
lLAo+AdayYqmEVvoAH/sJhHghlF8knPAKdj3mKDIY8M3ArtOlVNMQ2l85nulA+89d6W7XZxqtRVo
1z6jS1ibIocSaNlpiAnxYI9ae/9XT+uon/E86D+CYj3SmJbWWg4IvVL1+4OtiViPSnr3gmj0A7yB
/zjrir5TGw15rWjx9H9ScayJWpls3xWd7rVPqcW6E1qj+9NqmSXUmP9GqIPbOePReqvSY3MiLFgH
yVUw03lv6iCJ8h/oKddwSGHaoevyEvoLKLcRUXQ4lQW6fISRyzRPbkeB+RWtBfTLwmYpBqX2TcnH
vuB0OOiyPqEfwSLXNaOmiIMZP/ka7GbcLKw9LFe1QY22bOqQOvcg5OatDN/CiAm61fZ0Ws1/OvCx
dkSDYHA5Ys9LCOk/oURnosr+JFdxB7Xt5/d/MXFbUnVsfOhtfjuarY/WKeXlXqXWefDRxsPOQlSX
VGltNqU31QtTr4c/3QnNMeIJkNVY/XcBE011PlxOq23g+dmGgm+o2sUEqXoaRqCUuEaDFPYRdP64
roS4hAVvdQTxE/dAavNJ7bwjpTIzH33xlJ1SD2e4dvfSN12WXu4rUrbHGY9O8kVdfe+9WbIqb8Wp
E1BIHB5EkBP+BoNsIxyIScMmQACeWGxzXo24ou+eo8cGFBqb7cfWsuHCtc+Hc/b8qBlizjD2/6S5
NQnWjxICaMAiwsfVvrP4HnmPUP8kDqsfLdjS8O67m9eXco57Tvqdf+ixlW/rpvhF6lI5ij1OHnqk
D0T68T6yBFHX7tBrTTuVzd7xDnJ5i7i1GARhE+L120Vxc38CL/T//YY2rKaJGSTh8czZlKw+ll6D
4rF9k4DdJoFEVIasXf1+y7Aixalk8hJXOVaGmpJo40Qiw9Yo6ndK9IS+CItJb6CCzcIv/5ORwMoT
/1PoNmKkj1jV407wigAMIBWK0NeaRHj4SF63vtn9suStCJMk3oPyIlzvL44U+SSKk6EE6EexO6h/
mjPg/Gaip3F7IHVL+BB2wCGFr1PmjBgbDWggzqXhKN8SzHlRhkQB3XiEBZcLCJrMOA2rRS5H/898
oEN3TLCpr9DK4pTDAeHa322yBii5KdWwXlwpYxl9l9JraTBxqwfw7yoLJZSSLux0R+ozoL7blowy
IlEPSZcFaNkZfeBATdTe01TfkYMLsiVS9ir/LulHDShuT6RaRveOzPBYvAJp8EeE2EDn9Fmb5lsd
FSfub/fSxCX22PfRyTy41cPlDLbsvKvIlWA7VBkaHtywbGAyxB8aH5vTer4YTH7XPsm/7EvzNq81
8gB098CjM5W0wKpyLwzhNbZrL5bJ6j5/wgaa8hZUxabP4EbeGWZSmqcsHgXdfXz9R8JFwlC/qqeq
ry2GeYNdj8C5/wRMdr4/aN55ZNCjkxxcwyXUAvxwNE0E+0b740410Mw7au7t/jq9cVPlAADCpMGg
9fyEPxQavHVuJGmhAXqzhtojv05t1abOhFhj8x3X5K1WUf4L6ckTG0hpt7RHAbRJw4Fk3KEgvkvj
B0Oh5ZRxuuAoLPEZce2fXlXHb3bteSXHw7+MhHKXfuVTGuzt2gOoShjlEAgY5K7mF7+1x70/gCcN
albMY930tWHKjdrsfR2lHUm9SzegkxpYhVn2meEb7PppeKrkCTRoNfmmVf/d4fy+025w+0a0UY4O
vIOT/DWogISc1KU+Sf/aG3sNvV+dzWma2Sjw3Lu4tdo2G1vrkRnvpuuAz4VWZpsMOrMsPn29Ec4Z
eO6592bQoiak10eMz0bgL7aocEQaeQKgut8hHF49QiCL0vwKFPGPL8qs/yhhFZDf9ygRa7I3oi75
aKirvVJgBZPEzsxkv7NXF9ShRdauidNbUiznvhZixkH25AA3EqpP7Cn5UDgykiUxGKxAa4g1GMN1
4Zm1cEfOMIt72AX3GSUCt2l1oyay7SBaq8F6LdxCTjgOZciFzt/rWUEOSztW0tB+bIRHQ8gVvjKw
q6edzsW+HyaHG6osWs2f+USqIGPlyHJYqPizrWp/2FA8pH1tdjoNW+Vzjdb6Dqb9I5T7BvHxUJj0
qj5f2wFS/3LmoM5LtIQR4sbKrA2rQSx9z9X17FzZh6ac/891BbYyLIsFBbas6Hz+rI4vTwg52ypK
vclhWwTtHbIqDAB5f2IedGrqu9IJ6J2rrVzIRkLC7EzjiEGqnogoqmCH9k3oC2+bb0IySk0I+d/x
GqMEs310itFFmPZpGW0pYoBh+Xwl2rpLvbT2OmadHTpXWqogds3+sJLc2pG7w1ZUn3ilFfRhzUby
LPjsvEuGEZfPxmCGynebbmmc2ieH0BLZaNct22aPpx0YrN787KtWEJscSKtci7Md4OTaUk8ZbTIA
QkVYuZL1nODKr38n18y0dp5INGA/L2CUbo7eJxwAjU0bG8cVc4V78dHRA+J2qVhSIT993tXM6HJ5
RDk+uUEgDsUeGrNrgViNNO6Yh+e1k+YLhq7e3C8ZbJAGgpJ6V2RQgB8gLl7xylKeVpW/xa2tBGKy
27gTbgVPR5JkA5REYnbm/T7rOrvL6QcMi9UvIRq7Rw//YL6D6alJEwEzkQoElVwManauQpNbKuGS
C9q9oX5BrtFE8Ugm5cJp+7OexmGlNjsiU+doH+fT2CgA/PBWNbAQQc73k4XJmheKinuduXCgbHc9
XO8YfDQ1GneqUo25R+cpd5N/0R/2kyvH3uFnikwV/YKqgOyHNmitoMnCZreeCp8DYVoKHOjXUkIh
XWA+Ec/S3WFR3wOdbT8ith2aOxxc5YcOAjoTyPmnh8KqpzWvJNIqjPXlpyJ/awUeHTeKi394zFYd
cjJZPHq5ay8lMdmuO+2A2gzQ/5rxGWUZezVbuwpXe0xAA+LJJswnYEK/hls+y+yLZecyZfIJKyiI
zeeXzIVLhJGkrkbSnj1LUNvF+1VeZdN62Xe1FwMeS5zZpwOhigR8S8dsLT2oXZQWufhOjyGid0Rj
5hxbof0u/f+DcGJFk4/e5WCXwXUr2bhCYdy09GDVVFvEPAdL6G+yn7sUjdGrueqvmj8U0oGhOP2L
Mt2xg/Zyki1x/bzBPdSlJuwv7jzcZOOFnJTUw+RtLmy7O1FLIZZ4yILZrnBkck6aWTiq0k2LHBls
87PG5QWPIl1gK+qgUCcw/btpso2mqVHKpVYTNIUEbCcNJLKxAvxg3JMEhDLt4ro+s3Qa52nOZMRX
r22GMZW760396LWMzewkmuOdxa3JY+094ADVUfbnrUoxa8souDyhDXoukduRRVZ0adh6660QV4c2
MPk8M26nlKT4hOzIOIy3mPpZFMO84TQ7b+lVqPq9yd0CimGcxRo5BcLr/c53XsJclCTAAhfKcU4n
J5NRQNogwX1vFkX1+Zi9FRMHKhZj5MtIB88QkCqo9CeqYG4rn54nxLDD3v+6ZUVGJsIOMiA0ffpy
7FFVm9MqaSqNm6rLfiUkE3UGMjqRgRmxYGbhvCN3J22NoVuIHLJHRx0g0ICxRTtnRpKrJP501I+C
UGzGVhwof4a2gfwuj5aV3o9z+bE2ub2rzLYYzKdVptEixTT2I8k85cUGcXBcBUrireIdEafJjPB6
13in9ZkfYPP9VkzI07NsAjQ+uygXZvib94pE9LVGVhP/lCihuwAb3gypp88hZKs+EkJCqkUBO2uP
wHBq85uOH3ycYJNDebrNQtucYpEVESI3D8BSe8LqZ8zZjS38k6QEmu6X452vz5DvQzzg4qlXfIyz
64Az/mE2bkNjhrhgt3m7i0Lvpu+s+0gQPnjiEV69nvbB28bJo3BsWGwYeHfFfxGnRdEuGZRPB/Vg
qeZcPaLOPQId5r0mxIR1clPE0I8gpXwUDQXr5D5DidRSJnVcPw5SmnmzMqT4el5PiERU01QwKbgt
7Un4eagVMIlHFdd7eoVzrg3wwg7oW14lnAfMvtqofD0abMowgqDmKPMhkqesEn2ovG32BrFnq7gJ
MwVGke1zo8U9KPilnMpt0BPsBnAntf68DuXbPIR2VvxXcULXCfHyMA4a8wWqncYbrzIuf2jo/aMv
icNsQxS7oMtOH6kR6Dmf1FYXwBkr09D1lM17/7EerJo4+jpVBq0T7z48NO6LivW1W4OHxboO/ZOe
CHYwzRABSuoSg2YTfyViyvx9RXJRC/FFeJdL0eutB1DINNN5VYC6a8KqIhEwePes5oENvec8gCka
+RIt+3FdPcw4VOeirmmmwwxKfjX8uHkmteOWfohiWyDKMpNhFrw7maEF45xaYBsOzK6vdrzYcqWY
s5ORWhEoa/WFW4J4UFsR5NaVyt9yFb/ZggKjGbwieEqTk/2otksYk4Jw9qOz7NT5IC2QN7EJn21S
sZ96AbBItd/sSqAU4dM2aV9eMiN5Yv+afLZ1YdkocvzTdzoHVUqOkA1b14HmT0F9X8pRLr9QB1eh
EFOgYQrMTgfJ4+RSxu2eltHqKxfuTe971xo5KzErELSjP/gdCyAYnK3aiYwyczC2rX1hJcxAS7k5
jLGT6wXM7OQpjaeohStSSl7XlexeeyGLr1uR+KnfHaPfrcJlI2EavZXdgwFnfZAWIQNueUSBKAoH
j0tIU2kk+iZ6v7RcJY3YT6rBc+I+vu6E9vW4SQNeahIEitLHhBG/G+vouiwgsIBT0crXouPQrVZ3
uvQsqVyKzxiAyAzJXnyXaMdJosXhyYPDcCqCqU+dAIcGohUXOgbmLkKm2k/sDOUtvcvUJFQXQnbm
jtTEtG1QktXFdLnrQwTHHwkgG6zSF3OkUgzJgtYf7hUSIlMKzzYipBDmZqKUd2w7atl5DTAx0bhE
erImZfiBh78Hy2OuzOGCX04iNqbIskdaXtv8xdqboT7Gti6J2x+Ey6JgzI1oFZHu9N5VLz3EIUxW
7qrQXYkp4IFSZmrdU8y4zOEVhSBr3EjzyK8SR7KguKRwMOL7h4Nqz+K2c+AQgx7k5/fxRVr33M1V
qHE6VjHfMzua0MQl1tfAPfZu2iaCuJ+sWEacT0zmV/G+8u1IegA8ApZke2Q7eJyX8jhlmI0nktXj
T+FcwitF3w7wJ0yXAW0t4YN3PT63rHjVszeynqneNfCb+hvikFlND3b0DveXSlzn+W1pAuqKUsTl
t3Okb2/4zG2P7lOrUfbLPNQXKP8kihuN20joYsP4eKW9kq66M4GLyI1Xm4Ik5yQAm6VYqdoLPkgM
y1qYI4M/Y2MreV/Pl5OyJ3y/X/dRs66eWmqA/rUO3TFDdnR4JP8pJv3Sus3pgmkTdN92QoO2bnKy
B9EQqzKkVggXKHB1uOAL5deZv1VhDW37FIExEwj6ObemMoi2R5CRCLNF8aT7xGqijPs3haU6bSVU
aUpDFZo307hR4aW8/QwOGB/vwzVXpmd6IosXBBvozuDgn2MGZBLejh3CsRvJOURkS3jXMVXB2W+I
R7IisO1CIrTWbCTMariVKCH9Qk4fxdzBjp5DYoKlXpqP8rffZNY18jaeS0nOHAdglfvi2ytf/J78
YF2qxUpbfo2oeJDQ2BvQ8o2LkoZxkeOEj64AKxYLqbGrSsyW0fR7juO+koeyq4ZobqKIqyslQ/gj
8U20kxZUW19aRKFf8lwKYkAwgFU1LroGEQnvw2F7cNPbtjptf/9wmiNLFayaW02W7k5d8lHO2O40
b00xsT8AklCWzPpE3hnPEWY5mcQHncIYuh57k1l6ARLRLceG8A8akSKEZZWCTGhILAtkKG6DLzij
FSgVaHf+nf7I2GTdylH6uR5BEzmTRmwPxbbVP7pLLhVHG+cmCdggc2VWTYCauIqZvwct4wCuOT44
x/R6nJYgg9Fq7tAGweJIxglB9/xnokPK4KDf3F5opNXu4RtixB3NtIJm0h8zXI0EYguZfx+j3/8l
STwJSsv7Lg+YsmK2c4+v6X3c3vBivqiMcbTcBu6w3V29uCdkGaqji7ltcv6MJhU2EP51LaQjTfWt
Jisg//qKSQ3/xU1mOD0OxMftvaFdsieqvtVOvdMX5wiVcuZFcgIOQf7Qi8uid0TEnzf9lUhZoec8
4jLTP1GmQIJP2XiPiT22foxqtb6xUuPA6Sx3ZKvf9dz7SBXtyGbFY2h60qZrK5dmNyeC1AvRZwZd
TrZCofNzAplm+6xpnifmL5lo/8Y2TN+ldcUysC/a7nFY9nJAYl63RNAhgNzcZl3H3bBkCDA/Km0C
DoSveyuaFMha9+3XGj6cFY9V12LbFGySOZNRpX1+YpOrOUs7recRiAfPPkQ/zC6z/f9t7f+HRwvK
aFEzAt6XeVWHCgVYkBIMb3l3xmAoDjihuxXbMNZBzax1jh9OEyZ8VmpcRSjAL6rlkb1eKO7LQFqr
+LnCO3TrKzT2AZUAucESjmYVC2eBSEKkd5bxcdNtP1P1A8cApTvi1q+XxeQpftp7xPbkGb05+bdD
itdRsSHHkf82EblQUNRcbQQkaXVFF6QqGQG7xhe6WyQIYP1pBH/RwCO5A4XC6zW0Zf0Fx1J8I5AW
+s+cV99V/jBphff8V4QBTGtf4wGP5jns3X1m3HgIJf2AaFQDqb0jNOrjGemBk+wAbWv0nI1NizE6
Ce4MPerXTjU9unSgU8sZAMl8oV1zM9OHnZVK5FJsuvYCQngbmg1N4hKtv03QxkCRlBcc2nXPhx9Y
SAkrOnLksLGLvmt7TwhUV6MnwKvDB0dLSmLfxoHMtstg9yIpARQ+x++nUydgwVuTaZ4akBnga9cf
B8dUOARY0wl8LimkUIVuoBq4pPqlY+2hbA7emwJNljPBeeyZDZXo+X1qebf5qPvCnDfjlsPIxMRp
L1nTMirK9L56tIB5yGGp0auOMF0nKNJ0SYnDw8oy2Lwt0LOJn2DiWIIVPXAltx0MpEeIzlFP7WcK
thshBpFG6tWQ11uq1dUh9kO76n6VWkCmlND/xWIx1Ltf3TsOylIRJH6X816SBJuUcdQi9yYzQ7Dc
YVVWhf+SQdUXVmv7BmMwBY8Dp0CxkdDmskkbIs1uE6485nrDhseEQxGeLRzu3oPeCx25ikv3idnR
2BWt1Cq6wWyyeCmQDN+qJhnaWKOMMwRCnQ+ftx7QpH3JGHVCqLPouyXv19EGFSZCPXJEDydiN1+c
iL4hjqeF4xdKvi6QrZ74lfE8WLY9967pTRgZteKt/j4pIeX6m8W8O+6+GjbnkrDhZzs8uoP4bg2h
P0ASPvJGg5pzkUnLXKGsxKSPNN0KlFh82BADk9bBwdBZgCVQYQj3nXdXF3yq2FtxRbbOhYGqtIHz
gkn3WKNSS51RlPeHf8a1EAkAS1byWy6Dg+j3CYUYqRG1HsAKcN2TJWFxGCd7sKEVPOx6Yyw21IzX
Y5wxj2hNVG2SC4Hv/fe5P+Yl2zQsuX8ebR19h9L2FHaqJGaSDmEyZD0xRrngll2Y58edoUP0UgyZ
w0PMLh4mzjGBruWkTYT8TMugkLnOEo+wFZ1PphFf3RmA8UxoWzHLYMpf1TplD77Dz+X4HY9j7eve
QyctMlu9+GAQ/2hpfqtYRqv1yAuHIqwoWnCnXmG1i30ulESFdBijdizIbgqxxfHd9vXzI8wdg8zV
ilpHnE0aNdBHhcOqiW2QILoV6xmqDYBSTJOGTXRToctBpR5II0vtx0ofmVFtwm0stZWTWeI0yAd2
4HhZHisspN1Cs+G/Ij/zRI9AElKlOG1rNT5V+z0QiiM3L0xIyw0eiYur/CrFo8fC1MFNanb0ESPU
5m1A3xGSDqg50rm1It5e27iUZhzlDhehW/cCg8CQ3L2kclfUAAPca4I8eDlUUBPr4ROd7YS2mAe0
ORNkXXcyXvHNVHEHgIyb9C4x5i0WIpHPJH6Q9fuD9+zjOl0fNtJvwI2U8X2YhI7mbUrWBe3zLqzm
xn7KvkEZfm/7p2bjexlMeF5Ju0SitO9J9NvfSDXdPoKlXcXk6REvovVdnidKbVY/a1OHm6wLzxhU
aNhojlIwFAUlHOA+0xm2zePrP+IPZeH51Xg1OiLT2fFsDeZinRJXuNJFWvFhVeshwoAo8ZkT3bPe
WMUa/al6twFuqje263o5TUj1rVU19JQFDThKyj9nTbpgabJzHLIVGP9B5qGjBxmzrIBLlhaYHESR
B1qF9ZaFvWgyTJuYOanHupYSDjiIMNOpJLiGdh0Mlkn1pvFMPg+mz41VVRz1cw+fu4jNEni/U8dY
MS72o0y4TRGiOhUXH89kroOZQ7iqhQMKib8ZqyeJhiSRl8vfdsWgVT29pp1UrqG1ByFiK0TSxAfm
6rxaj3Xbo3J+p/EFLHBAJ6rBwGCmWJExoPxiKfYvt2MOTF9L0czVUKNfnCts+QNQi5Er9hpCFKUE
BMcNlN+RD/GAdSC934AZ3Z11PNYAsCaV7QvozK2T2V3xMiTDCE5Ro+Z7cpXdiHMm2usfzubjdwXR
L3tatI9bUZEb1R6Ocd71eJ0mmzLWhXw4dt6TK6D1g5ok0jIPJccRNUcPJI2VKi9VbGukE+uMXf8M
1wr2QmLkyDo6j7h7iIrvwHZ+VuNFrA1Z51XIXwXlTnIVFu4KbJnmONlZhIRhvZseYw42/d4eeO8/
URnLvGUKAjWUKAY8VX0MIwlhGWPKlka9+5NQ1mHzrha+nZl8P+Kifju2Alm/Nhas0700MZrImS0t
ueqVJusmy+Ipc09z/gjn3tHAiwIvVGoc2o4GDuHg1LfmF0matDhBziV8lydPTVfOp1B3i+mYuFEb
T6Sc9vJjMcsaugvBI7SLY39bC2l2sxaiT23jVQh7CFMlbTXliFdnQvj+8d+/gdMAeXLo4G3xufU1
5Sh1bTDobgv5CeWsH9g8cFW4gjq1zqKXXkyuN7p25nz+YjAmSKTeohGF3DRMQERqO/MDoqd/jjsV
6PET7+OQ7cNozzCz48MsVZvueMcdlpIqOwhxoOpiYC46ObTUyfC2b00TrJ9XDZsugCNZcMuYR0RH
sWGyVvxE7f+SgbuKyDoo2DB6ICPCR4f8xbMKbNlOwWfnsg3Vty/mwvWsDFii/9Bc6gv9bt/HMNVT
7YFT6sg2MeFCu0boK0W1dXfREpeUsv68Wobw641I81mz96NMq1SBA4Lo24LlsMZMy6DGmXrZEZAk
tKiRkYjwDuwIGpxyAuvK/08lfLPnfKn28NjgE02UhwrabaTSWKm/aXxpPSe/FVrBvkLG0mTByza2
xpIRCi0132zTvS98CN6giaBiWYsfa5xKJMAZmAKvgpKazJ8TpNqZ+ALxpgaydy7TsbXxSKs6Msfd
4IPThKWckcS+jwJhhg8Tx4zyHM+KUIzO3jwAZxvX0nNGCSrsVEA3uMhb2lo9xhPj6NdaDvsBKjyc
5EByMCgZOD1oLIOiNmMeePx2yyq0a4EcmQL6+2ZVVhj5I87M9qJozJffXfQkan3eLaDsVF2rfAIK
OXpSzJszVKSYKtaK2xfARw6Vjvn6bIsGWaSSP0tSaQ5aT6/aCwr+8l/dll2B2FhIaqmMKDuLOv4D
3sOBUjvUjCvo/0JO6r6B32L5TXb0L3IFLE6EsXCmTwZFte/ABYJtZey5YfHcG6wLXIE/0i1w9gEU
UQnrpN/RuW0nH6sTOgXOIlXip5qdLFzwIP++JD+Gopm1pqzbuxKXtQHV1/QxjccwW5W8eeWeIjwK
+Gm9cKUEP/QtaUdpp2FPRZX4uAzeSNF6jUPMZcQJFuavb3bnp3xortkE6Xo6zzctk18bAm7MDGkD
1UD3qqSJ7/pBpTu1SMo0wSstSUPHMCdJTG2dFqY/UqlbOKCOBQQh75ufuqzYw50zH+jUyCUrgQCT
+KVLaBoa6QZx3hHcu7wlHVG0/pvg8/WpvdDxAyPIgOGdPbWKZP2V4NrgusXIxLEdG7tBPb5o+PuA
+7OCv4xsvfjNRa+1WXcQx+gVGhihUnuQbQHpdnIS5mGdP0H2wR2ykO9cbhytl4cJLKEw+fHzZTTN
L5+cYeeGdwirX7LBdSBh0Z2+mf4lMilKo6QkZwhwJahYd/AHyNcM0bstOp56xC//snlGOYtaYQOr
vn8JnkEQUD161wfokBdubOvzU/G/6XgJ9vy8CpkGjtopP+FZms+IlbmOiuuRtEAxcSFcdGPbDNVl
46nQP+aSlEh1nD+pESjz4Zxlz8mfARzuZwekBz3k+/5qDCdKXTmfOD6YJsF7HxhZq46bug90Wby+
3w4B8FKvqYhMqqzW0Etj3cQcF11fcQ/RAzknNMu+vWH5j7EhbrzLpYJ7rV9FBUtD3tTh7AmYV0Hu
GHx26p9/VYNGxoIr/wXTi0j5buBwBz5q5urJTG1de21NBl7rPd8MnAT58380JRj4kSvjEEJQFPa2
A6HkjrRq8sMRbgMUCPEyU/J0vY0iTDyX/6May8TZwAfuswd88ji8B6OAPtp/fiZBK1jy8KuMQvDI
2pY7GVm0p+AVwqIVJD18/wpOtrOxsKs2nKIkckqAPhI/Or/5+Yyov6xouvGGHwcAV6if3pKLyf+B
hDge6qyT1jjQX0phiGZrUnxDuBGE0QLVNSHfTJgdQc1Mzt5+B4YrQGjbekqPw9EcEQzu6Wz78cRT
NCLzSY8ZxtCzaEoVV4nZVs4iIWI7Yqw50QvKzm3FWVe4Q9xRzG6kFMnTRtJA9GWfqVT5dHZFsPkz
ZnnIdrYyyeBX92+gc4OIMFUmhm12FKynY9xzmgs6VOpbr5VdfsMpy3KSLjFppEwuCa/gX691isxq
Fg1WnrMmWCPraffPPMmkFvn2itJmAb3a3e4HWUQgNA/+rrJRZVvc3e4vOskBp01TXQEObWpZxmZ2
vqYtR1O32Gu/AP5tYRPIcBum9rO4xzR98poYfb3Ne67OOoevTV3EyvKiQj+OUqbnoV02goR/G2k2
vfVgvNfRZAx9pP/Z575FgxizdXakbfS5/pBBYRM2TzXB2tXjTK+a4UZuxYzvOyy4RvO/EtUJanB6
XWfh2t0wQrZTUeuDVdXvJyDMZWAAM0VP9ZA7o4bTxxyouoAneF8FpQAY/bWpxAP4h83mfxjNzbdd
K13grd0gPDV0W5n6pvJSoSsLmQ69Uc2Exc8XUvUlGK4+yA5RwJdJeyqwXmM3PNPSckgGdgAAeSmq
HZNdyZqIOr3rZVDdmwa95ccS1gMHcir5X5RDU5qxVN6peszEWCkUoGIy7TcWaPcqobaxyAhmJLKR
VpHWbAs4YwV8WkDuH31pKMm+cglhpXJ7VM520uYWYax5p9P0kTzrPhZpDBEuw8muTPdtRsMQLXCc
wPLkYwukklw2jcNjpWZkY7mutPsC8Phfs2AIPEgr6Ggfn4JkLMpYGNl4zvjgiyQR4xCWXdEoTUER
mIyit1trZ9uAA8xm3Uo5WAT+kqOb6BsYoMbMsRVIs9KwMrRIo3bv6UTI+JNQCRMXgbylYBIPkvG5
s+KVLwWt1MnjOe2Rxw/C1LLA5ypqbS+p79W0tfx1bUhpX6QMuhSV389qn/QSm8vML+Gp/UwVCd78
LqEsreW/l1THbPT+bw7d/DDylJ09wrGlCwq4O12e2GS+Qk+Qx+z9zf9/BZawZamdvT1QSBnO7Pfc
iWDMXaoCq36JCeojeSAHduA4xRp9ClFJmEV5hQT0TeQIPbdlvlUijI5LgFTalFn6Q8dsrpJZmjXg
ZMg3RiRK/Rqk8Vs8asJLcfMqVmksroVMZ0gYEBlmIxQfRN9K4rj4od3aiXjRK7qn5CXBxPnRt2Gn
9pwgbu5ASqB1u5frw5rFsCu8cWMc83nQF0S+H2xxyYElABc1MIXcODmU9kYH3Obwva9cbeBenvBc
qcXp7iz534Vci4+cml9aKyqM4Q1e44TnpXOfhSCO0xqohabVbW7/EbPz4nXYrNvfnf00yLaLhHeN
Cwytrbfo/g8O23F/xaVk8az0aKSYobz9HgD77f4GeP7dgvAF0UYyyM2vraVPbXhqP8ZC5TtuasTc
qRa/bfQkWkQsbXnSpGUygS5BokeBfAtTVICgsEwJNhFMgq3U1uu11iPcWeO8d19E2KtkrwcWjhtQ
awXh20dGKwjehvBQTyPRsRB6zH4TZRAqqfGXDSzxxQinhhDbLkxdQ10TPskqVhMvf3+nOI1mEOqa
fwzPbIqCFCd50S9bEb3V4ImUdFsRyMRBo3yUB2FBYdG2nlIfN+E5n7ohhIPYUn1Ts08RoHEQlB3U
RszgDuvZfMmWX9Xe/FypbEpDOD3XgUn34stfXjtiWPb2eDOyYqycpcne+fay6j95BmyplRWcqflz
IxBVKzv4FwadC54bPWzoDfqQcAjbirdgWQ9wzpbUj/fDckVA0jC9fccuZNPBoovg3xT5aO2bfSG/
s38etSzPRhRgmtBWx4efBGN8Bi9fdWAwRpoU3Lea8wgwrBYCqWO0aVNN8dBhveqkdBnG912LWugD
1HfckHDxOzI3TRT4wjraN2OxjsDis55AYcBQlv0Vj1D8u/vTJY3/n8+cUMELv2Lpas0C0ZhDNcWu
sdzjOmrroL0evCvJHqjHBofyHw/f6t3tx21k7pbg8uxgsB5wFn77fiSD0FFItX1zxaGzL9few3+Y
fkcS5NVf2mf79hsbspdX064wjO0T49D17AJxtDzn1gnYU2ntNQMIJSAX8kGnjvONljkX8rUn4afN
AuKIamyXjrCACr2AR7u9AIJuOd+kzXUPFfmsiowYKpWaRvqlSfHvw2wkPbq2o6VfZINXMWY276nD
3IqNrJQR+GWCHagtK6kTH1vMR+aL8wPmMa6gruiREdoxDen3Fd4XzoBs0LsLcbGxFW0ESmK3F77z
HreKTyZIjgvuvLkVr/Ie88zA1d/t64PyrdXgTbAUV0hcuY4aXWRMcHBbnt3UiBxynViMW6HSFq72
auHNmAPkHo5FJ13vA4+jLhy9uUhyyPmD0kQDpzD7abS6ZkZbTQvKaffZ0fyJ1zztB1nOdtHN9X9o
gVLN9qbFlNrf0l5kf9Sgba4durmMNQ4nPx0YHMmyXMTy4n+Q7i5S9GxabjCVflrUUGk6f8rpOfpY
jUj6zswXkQF5n64CwRALUeJH52EGVbdXOuVdDRHMrzUKKnBQvGWHCYeAaZMbUh+iRhYGi/6ovaqi
3Hy4vApxSYqM1nGaExGFMrJXFJrA3oVnFAg7cNpgu3ZIhhZdkfrJyGMvAnpUbdlupDsJjw5A9Syv
nZUOgr1Xyh/xRc8M5gI8io/ZcisYPWf5lm+l9RDdbin6k9omR0XF1mZjA8Uo0yFo5a2UNIoQi1VD
6dKFCvldaJ2Ipiafw8mOA1CfrfvDSYA1lyXXqD6lZ5Vg+YJZBi8I6qGRfJnPf9WImdf70j0seFH2
kDoB7I5GDwwm4DTFl3FqnSoyZuzjlQRGIBVo3FcYckWKbVyt6jr0u9qB4z9sCZ8pRoaRmTY196km
BerTojEFePO7eGXmZjwfji9tNef4WiPobep/aX7bv7HPz17M2/DbMlpbHIAYRdEAsiMEH+3hpnDJ
GsWDpL/rKlNTPzXy4O6lKGPRi76EKf1eGJCr0+de5Wn6bbb0tJUJ9+IvUJr6jA4lTAivXONRAXbN
eHw4uQDr54UQtCUDupDmZo9Fp3OdzCEgfmk7D8mgQLQbCcy5eoXz8tZkR8eXwn10CM/sFtWGGssO
D7oeqtOZ6iWQB1aL8TqyMBf51AzeQtezJWzsSQ9lzjjWtW8eLgTVXPW3GaBouzwmtW5BGb+sKwRP
neZ3k0up9pwo67HgO0E2zTIu3njExcMbXj13fEy2yfZ/uEb3sqIrDGsX58gSypOsUpz0p4BeiWMz
eJOJZeyj9b2PFlr8hDwMpO1380Wlb3il2W/F4J6CtoRIkU2BIIZSracRb2VlL5CIb7JLz+/5gKN/
Nqzrbj9mFfj4wo8I2n6QZhjKE3J++mgCf5TYdCg3aznBfZ5KZIqGJKa4nON0C8qjaaBEouSD1YeK
HACIaz/qPV8H9EO9+5sHqpNtGt7yJmCegqT5kpnQ1QTdfq0fpwJ+qydEAzJDilkp/r3pC79kFroX
TEIOUdJxvFIT2599y1A8ZOXcbBvGdNokchB5AZUzsk29HT77xmhGAtVCbp7ZlUXoIs9uogyLVH1d
4s9fGjbM8N+Al0WnQ0ZbpejpzP/CgDuGJ0f5cJw0gGcqyyExEPfcPxqRs7l/WAfVDpBlidafShvV
nsEfpyhfaol9G6M1J5IHFUYDBHb5CI5Bd5RkwGoud2DpH1VivdG3faScF90IckoDdC1zESQzogzH
dhOzeseauxVPtOemrZL2q0xiJKKyh73q91SQI+0T/j57p/xwpUISoSe5YH5UIPZmYMjqyY8Nnump
sq4nug7S28mQ5QFlpw1pmLXLa/GJfRpAn+KDPskEx+NY4srL8Z7a82YoxFQEToZ7/CDpyEF5zut8
rUIERg0D9C1+K0+OxdsC0HRQjSU7owh7t0in1aLn5QjskUOJGo4KKAPQNLHytGryCrRsCOdyZ925
TXA/T3nmlxtHoAzWa1Le+O4Kt6geeBwAzMZ1Pdq7mBBzV4f7pMkyzHUC+3EYI1+jEcbzCKlmcblA
hv/QC87qbn2b2zReDH7tnmY8XJ/IpT7mSGiCvQYyEv3AGIFObAeZu+1yUPuoVy/MOp0zkz/N8u4W
0Vw9K/ehpYCies3AAVFyjNsFvEw+9Xq1tav+VERLxvufUCRYaHt19bZZdY+blt6ew9JxqXUSbeJe
NRfAdGX4dR17rnDklLH8KlAi1rAl5UlZPjO0gMxRoq3Cxtr0BlAB8EnUUqz1pIsa69b1W0OQOPC4
469aU2BJx71PPzELZWXtNdb0hpAIMH6upnqfr8/Lt6jBQmXfNIj0ccxv0q4Z0MfJxIqMc8hNnHFC
zFPaGy5aFj3uMgrBGKP8lzdHLcUNM/SC0kDoq/hVpeoA3BNdSEPGOkYgf2Sj6JWKRfYtocmyMddM
9xTMlcrRJepq/dpkmVoaOj3yM7/Q+kz+nWmtE5hhx6ZmV5yhzW+kCuPAZTYUtMinCpm4JCL5mZ/6
R/nxHq8LGMZ1Qxld4EtqH5rqmMCrc9LujOywQAj0MK2fn/UE9WiIkih9u+SjMjELQTDd2PAVLGpx
mHGZ84uKeqrnM5878i8VfWmwGQA99cBU7KD6utV3kuN3CMdD671pfb5pvAoSpl18aiEZCQiDA9xp
6ix2vvwBmZKYJr/YMjEZpubKveYAE51rsxv/f8FKmUIw6+kMPL9lCXMVvu9wLDNLDUNv9nBkC+Vl
T7mmcfnIMha3zaBAdTZSoAFqwOC8wdxvgJQke8+ieuQvXLZS524XsJijwMxISoI0BsN7poHcuzjR
fF7T7jtmE9TwuEWDZWEkPWuCbXyieMKrrSJWNIuOsp4ATIiyDWkFMU5c7eskz0hheh5M1sBkeP6I
/4S+PE6zm56u4vm6g57IOqh+s214kFuhgVTnwSQsj39iWZ1C1iJQbUNvss2L5Eu2fNLu5mQPdnCz
oW5S7Is3iKaRbnZyX2ymi37lL9kXXXcwnJs0F0VvXlAtEGAwnpwhM16lXUeQkQ3EBo7zmUsRX1Vw
v7/4tIZukn6/fGVeFEpCkQvsbQjiqGGN+6RUKXIL/TI3kDzxxj0g3CjLYZErX6/3VDyvNH4JZWTd
WidULj5H9Yalz/Sr8R0ZbYg9z0PWN3tsr8E1gcL43tXMUkcwq0Dv2zcOopXtGbtsBkYFH8wiooLb
484mVUjVNhN/D9KBzEmh1HfmHhBMZIp6HGS7Anc7LcJfAmTTFRsLWnIsFvzuc9kZqRiK3VvBi5H/
6Ipkzwe80ukKb1W+Yn+Up1Yx0LjVzmMghmDo9cvAq63RoFgFTrQWL1faLqZYQq/4gdG6NYzzA8H8
CZbssSc+uix6aNrYxrRHyHpcqJomCHQQrZSGciYhL0Y5hdf68uYUlcC9ReyYjOY+xj7/A9q1zVSZ
uS6J42a5QA8J6bmGdiGGXGIG/NdVY0g0CNTr6/AtckoA+kDJ9I6wWlbdvQ0JtUy5awzbgCelgfGX
pRz7LuIkc0NZeQvr6kw0WjZU+oJKvSL6k1n6Jzt7MR/7hip9j82BhLyJOR04pQbufJXGGRGuGleQ
ncOHg8xOgsALlpe/H5KAVYa7v85BZ8qv26suIZrXvoszXhverd1nebe98ntNOIRLppqx+0ZU3eTg
oeX+TIx/TVBAeTFWGE3zzcDosnhZMldWzLgA8pcsfVIpnNjhJLw6VFS4UBjqEQmrc2gMX1gzPPm2
KEv3bD9VeMPRqgL8BhSxTft1MqMYkZG1s7H8KGRfc2bgHJOlLR4WYvyuVLOWl4SNWEuPTvRVoLya
eEJ8dzhw67dOUo1LyBfwec1BzyofcM4mx9UEZuwBFSPPTUMfrarN4JDBwnc3aKayCuwnVYCypx8o
1w/Ia00dB6DTT/A94tXHbBHHYfWwdxAnMgBER5qsltx5W018/WAx1d3CQ7bH4KBjgIaP55nHgm3O
j0FAXEYoJWqVZ55+dNdpzXvvR/w7xISJ/IfPpx4uKcaUPVzC0OrA9Sf7304jHapMu0oJA1fcIw8d
hQpSQQv/frVrLrMhue4U6v/NLI7yruL8m+Yi9WfS4j+ls7ymvhXnjd+6xDxQUSfkzDIDwLe0/Ef6
RI9kzmcGbCVlA2ESNk5g1p/GIAxks3B4+Wwq2wDkOCZ6cGMutiBGl0vF6XXaBPgMTml4U8JeXw54
Ki7OkyWSXmBvydK7N0HREAlsZPul3etu0VzdvHzNjxeVRnVk5fyPE1ZNKsxe1yGmB09HfQiHeYRZ
VpNaVNFTzoL6Roix9K58rAyWcDci9JEFnRO788CA2m8uk8mNN0Mb8DGUBAGbWW7r/d92YV3o5d8c
GMHAL5mCsniBrAwms1WzBb2qc3U+trStf5BhisMvqwgM0Wz6UCjWwttZPnVz5aYbdHjf78ssUY1S
k6NFO+w4O47hQBqR2NZqT+nKGTpoeaFBjFf9eyUE/prYHYmXTh1fnYgq7+0sJ1Lt3JzNEQP8eMfC
PQA+mc3o2RE+Id+ig80Ylgom1wY86tYOOoOyhl+Dji/1L2dirG9dykGAoMEye2Y25GVCI6oNQzPq
UFTuPA4pSHEXAx19rQ/oOBJXjcWlfJ6aPWFFELToPj3kJkcPyv6pjC/QFlzk7kY3+2q7agJG4siv
rYDvM09oQDZkTeAi0fL7EvgWDak9VaC3m3zL6oHHh17vHkVaodki5RjmnAjaujJUiaMwSzn4aHnM
3EhPYZZoN01jmaZ8890qNHt8up9QXS7D0u2xHtiCGc6Ahud9AyUHil4FVLP7JkF8dUxM7keVYYx2
RdzHTAPH5k9p/l5VZ9M719kbNGP0szA/elZOGN0S4o3hYw6lm+H6vLZoNJMflZrmkC8nttFbP7KY
fXL93jXvxWC3LqZYBiLohNSs5XbD3XjMrVTwHIMNomNu3skGawHGTFzscx9RvpEnRGsh/FOpGwuN
fcsIFZHSHGbWlJ/4J3J700z/6HLVRbThSiCUcP8BjTO4ynSqoQ7KNiHVlrIeJJobC91H6HKMQ7/U
NGN0mYnmnkq1iiL+0l0/R4110d+VoeRHVU1jRJZ41EakucKCKyikUiO4AocCHml3fc+xTLToNHZC
309H37OIJgDBBiYVM+Ek1zftXov7Gd2SSDoLQ6tZSxqhWPR0EZeS5pXZ6FdNzpHq+bobki3VeUWU
e3QUbFKZKDZHdZwJxKMARKPnTmF7hkQIQbReKwJxgE8/FsPL8B9tPwYkQHcgcwuWVKRGuD0NRD5J
TKU6vmQCs8i7u9iLgc4e47XLLSWBa2CvH7jJeKqY5v4+3DQ/9S0cpyLFqt6cQXgTibABt/friazX
UhX4iCwO87a1J73wFwMnjSkREkNfAcorkUqxT51xIHt63xGvi95+GdnS49iixCLBnvZSynwgEz2C
WTbCNkRSq3yrBXFTg3WZbz8JT1meUHnnpXqBKMnQkRofYSt1Cp1SfFGZce6GniysSxu7O+E19fr0
t+Ozs78kqMKXtog+eNBb2Q2X03xxv9V+htf7lh4KVWrkr3uvKFTOYN9nZRUPZtLTNkWU34CIKT1Q
8Mk2z7e4dN3b6HcXW2BzEKyEObTYl7cyAOQL1OA7QLI/65onhUUvjCWiLjwuleSbX091DwQmKtCK
U9vFVQuzTtY5C0gwwC0K4jdGIe7ICrBs+gjf3l5RcWhZ+aZz/eXO32cP8j8kRyCNmA40+ETxoqOs
viY2B1Y2zLoJ0qgRG1gCEplx4Pt19rajX0Q7E/Z4FBjtuRQaekO3w0NDXmJCZSzWakYLh5rLx+Pm
uefh3XqsRNcuq8QsR+rLIqzx+l26bmIEnw6723DMP21XOs0Ndv5xVUE3JGrxEobrbdRi+LCZgQCF
q1AQDGWcR1DDSVb/gJGtS9jFk/lkbXEgKUmctzu6u3Ix3N13AuqO+i/ENcRovge3OjF4NLsI7aMg
d9tNZ9Bo6ERdRzP35kCaO1LXJnAASeri2g898BdVFsck5EgiOyyHHZPqULwQRA6aoPJQmvSIvIqV
/b6NarkK682BpKwxid89rwaQrQzUhETzCjtvSmr9PK9a/gqykA+0iYfWnge9GWHbR3fHuN/3LuYp
H1pE2KHXbfaR+bF66Uf7h8TB1sYjRYW0sxqBJMd3gcAV71V+sK5W/OKC1Btoc50OQLdEO3dkPZCB
eJz3tdve/N8kXr/J42Yrao/T52oNLqeJWaaVIdfHs/1k+Zt0d0yyPapKxuOX+2TZD13oE6Ft47FH
l/wz0vfmRCHYtqVxNp2DTFywmE6iva4khKMDuFSEeQAmDFPoXATkp3XA7Wv+DUVyD6qPTs0dQVI/
3NqvlX5XOl5TtZ8j3VOdknQDfTrKdnoDBwrg6AayBAB1EMWpx1iAZiUZhzPVORgHFlLQvxn6w1WQ
NgLjFMBGBNeAG7Ki/Jx1OZF/+1PdWrcOD9+OlODTJIL1fd/bzCSu2X7iMvElzpqRYvck9yapDLQc
0FwHyR4heXOdbVZPWsFb1ehXC1kyH52wqe81d10gPbcyjo6+oFSwVeyN+siAUiJkvBhTlmUp/rCi
Re5vifP5BnEcEaidUNiPwE359v8hlbJa71LQLPMRbTYBmaZrZUEE+oiL8h63oGyogqK/lLJ+V+j/
u1YoL1OvUnaH06REMMyfwL0sYuXPT1UXABEdT2CTl3d1RnIgjz4QSX9nEGTKJYd5QiO7xI4Rnp0b
/f9Pr2fRdfjCeONoive30PIV9pgvD+0v+5ORJJtKyJ0ItJdJbcgqx29lgHh7b7oTE7PoUnINMpBI
Tnj3Fu7J2Vr0wsfl41y/DNUV0ufn3j9F+mN8sinPP3qD1wJo6DPWIzo0Tr2Ql0tPoggIPRGlzG9C
qjR+VHyhcjfT8ReKWsXNiNBQ7NCyyaLUtxJpcY+ujlZu+zBog07kbqv46Nrlefoe7APAcQjB++8l
zlPfCnNbQHhkty8VU6j7ATw31AxfxGm5t8GKSQsMj433ES5z30znehFbeDsZdc4vIxn02r4Ut9oW
mEIcxBsyrfFRaELiI5Kccy5P3GuZF91F++icZ+pEvYzypf/YFSIUZROUICFrukmU1At2Ld7elacG
H0FVXVikqVT628lvWQpcUWoWlP8dHvg8uzYkXYUfmQB04StphucsdtlIskyi6cVYSxLo5W60woHK
05vyBx/YfNpe5IRjovE6qezkCWW+URY0NJGtbwzl9OTf8JbTyaWbtf2aj0/hyU1b5zh+2YJku4ZT
0s6MvdQWUkek7ddrq7dMMugxzAvjNd5DPfpgT+dMyYX/gEk0I6QZV+NMJvbkf7iWqQE+z0kMKFFN
NnzML95je4kcm5SPqhoKqNz3JcBuZNVDFcVdHPTGZNU+PE8WStT21kSDtSfntSj8N/4XeTSbK60o
mgC/MoGuQdRJLPvkeHBdXEGFb6tEQvZP0eBKJTXLsuxExBjABd7/l1p1QSY0IRJ6P0DNT4ZqEErn
pU1ppz0+V62MLU9Umd2Gf+w/mgJOGd7q6N8pw0iBf8rphuSYco5iEW09HYzsPTSArv8zdNb5vhMK
9Yh/BFevHp1dux7ml1v+atnTBj74PXqPMe6uUKPVxzk5vzetsFfUlZACa6phyXplCP5hqF+1Yv7R
L5YnGL7Oof9y2TZU9sSXy4yV45ORXepWSOQ8wh2OKkJK6FMlfP9a/SLux57AjdgTvplTjI9Q8F6f
ZGEf9uUx2IQVRgJHdEL4/dgsxPkWdcwZgfkZONnboXj1GR+SMDQScUxElMTSTWhop+14HpRDSnLQ
QBF3llZm6D7wzpYzHcmi2PiIH7jwspfQhQ6EV0xLgOrMeMr2YuKef7ly17nMKW/AFZG++FLX0CGg
iCdz79l15hnBCvtxuW2eNUSrGE1AeMudNCmNynx/gRdE/XrySQQp2zyAgyuF94WY7c2uRPCDYcfV
sIozuCSgs+5+LBJ4KX9uUSIjnyyN/uN4Ecz/5hhm/JWKhA0gSMNVkx/J5/5Dhaz+NmMUlOQdfDto
tL3/NPdc6U407WWGc68yUc+ztCGdxxvOvwkwjAuV/CSrOKGHSuZtxG/7c4OB/UYId/NA4bpKdcYv
ke/s0AYpdqFPO8CTBkRf8xbQhof1dvkPws/T92DM5BRHUThcP4K0KwiktpcgQ19Ysv3COS8UIeji
parBXVR6znuP9O8gRqAYfdaIJmrrvyr3SihEV/ZAJTCfZo1//BOyU/7NI5u5YZnkXQoR8wR7pZxc
+qpHlu1wLveeiASnKmuV4vyxgbrRNwpsf3H+W/e/dotf3BIaUf4ZRU0TVnQBn/alVwOqlAX8itT3
y2eLMPW4DmyrOxBrrn44wRKoPKLA0a37OZNucDCSMdleG/fGNONPlLB0Jkem30kRbBrETBdPRW8U
ywdTsLm2UMgGObVSRdr5bMlDTo02KY6vePjsN5H6wnSNXufC0I30ewEI1CdohPIqpGF98lG7slXE
ehWmG75/hYLT8GT/kyGvVFoUkWDscfQ/TlrfQu/JkpNwUahnNd21Vd8Cx+uj27vbwHGtKif31pna
+azluq7QqSb/1WzyL7RkXErSizJYFBav8J8/nHpsAO02LwWWzntPGmqSfDRKgP6OnrfGWf66Cn+O
/LBFiYeCUhtTEvwh5qayGGQqSeceGlyGpOhESM1Ere70LKWUUWzZ+Ju97PdnzilwE8bUbAIeN4PG
yeZLCoA/ur4QA/4eKAJqsC22EWh/XZh1G1b3QSXx7zVPMaJM0hr1TwW44rdCSf6x3hfGD57Nh1Tf
vS6G0jeHeJmm/cSsDW4yemlZ8zaT2kxJuq3jhptIdvkutlMcFYciT/As6++edjhEkJKhj7hawLre
zqb/hIRN13DzpLYAuG8v2ijk2rOeP0k/1/wXEgZPDzeYLkY7Rpb0D2QYUYrzxhCLj2EfHw/FRZx2
gyXotPqk9uTEIHQ7i5VMw0+0jtZh61xT+/AigFU84IONGiIXomQvNKd/Y/w5eqE5i8zl2qKMayXd
WjrvtHxaTD9WreJLGirgDCWZ6ROvC9YCaEBDbeODTPHjkadbJT3hej3BTL2h/CwAMLUpz2tFpsys
toF+hKo/7pM5EyB96LRJij6JDQx3hSyLspilktVKZPS39ptadNkclAfZts510pXhlfgBYnxZ7joP
nCU8hfW2VRVkKt39w0PtbmAP4pTvi3QhpeIzxW4cOnsbsEJlRWCyUsCCa8ySoZN86LSUPDwQJuBh
x3BU4TZq+N0aAqfadd0mvDtu53da9204q7BfAO1C0KnQFF/AVD77OmDQtb8P5FXK+7Sd1qWtFnlz
nYaGcdTft+y4sPfDgYahGFoE68kT50kHZrG90+0XA9FvhSa8k1m3xxsgwwxTo/qrB6n/wRBGiuVk
TAcqABbD253hX92J5FuNJ+BjZeDKbAtgqP9NHT3/23MbK5uYD4FDSyE4+c+5EMNsbYnD2ZIRUj3y
O+P87Y/+xShZO8gzwPzb5Hkxvat0mVf5VRBypSEmwfd9J59mJlsqHjZh8pPvZG6AYkVDTD3SbGU5
vrG1i12rAtDTGLfhWfv52Cg4pC+vmjDLh5xOJOUXUTJaHcvvjA3XCYO9NjqKfhz+a92BLm3ZDMAJ
Lvz0qlba46HeYBtxZd8N4CvQCbQGNh/kX7ZncziywlwY+veyWyQKPY7SYpPTIWAE/oJujrzqJjj4
02Wsr+N07bAqE1PGB1+jG9lcP8x7JfX5RIIh9JcePMxCtZS8+npa1iy88ys/tetzTDoah5q5/B5H
NkeXaIAmWviSLJacXlibEA9nRoO32i9MCeODbI3SNEZFT2YSNCRMIDx4fG5LhdXERW7XJ5Jt9f8G
EsG7gSgBezSzxnBI4GeOaSd2HCexSBV/g9ZNi+9hvolOK9ViDNcHN+VdhwxBz0QzlQ1ydTBL4Z6c
SB+QMkQR9Wrr64uVVH9To+I9AO4KcyVS5yhIMQlLvhy+ZjVS7z7M6vetOpdNFwyfRFmGYqVj5vQU
LDo6GhmdK2Wpa4iGa8wJ4LR7IV9LJx+HwgsgPUCs6udLhoBqQkPKUsTQp/WdQVrLfCRBL1RPun6t
P4rddWjlWCHULYKzaOESoAoUzkhdWUpTq2YpZlhKD+U0CUC81vUCbXuZepCMbJH6Uf7pVLJ3Ctx3
PRtHiUUqQed6Ya6Zxx7l3/w3vJdV/sDg/oWvTrq+Ko2zo1Fw/gdezfIpUQ2egATHoXGsFYtw0Pwz
UI2k74Zjt2HZJNi77OvU9T8y64Ecc/jCATGPUIyQSZM7HDiVpxLP+A47prHRRdBPOAaIkhorfwxn
ta37SOsEuXcgmop1hJ+YQSxOEooYj6sDHyuXCWiDlyYiBkAKnbvsxp3YwjGbWFVwYzz00F7k1Y49
Mf0fCdGE9RIg+DAXa/p38s+XXoZLI9WSOvWLub43snZ0DUNgS8VcFr/ht262AtSy6wR42lsd8IsO
Rf+/E5o4ihzk8msOMHUnr8SeEXg/tpx0t/OHevzfCDGwnVjgOf9l+lxVi6t03q6KpTcYHXpRDgsp
eHyi76XQvrrjxJaP2DlskDxtcP609tt1DBAmmydADvgyU3/nFKKihTPIeSJhryPorJ77QPF0DvEJ
clG65F6R5REh4wnhA284mC6hjhndBqCrpOItTLJBz4uJAvEQDVLEeGerKCvawQHln/i4nzRyfVp9
LF/rWGdfDSu0YVavHFSbr+iIqlf8ApLSx5B4+IQckOkNOTZolBOPRJP15aUPABaxq26+GcZRwLs9
5oguH0Y2qQMpV3sWcX/24qcNNIoA7/1b22VBvaySla0wXc7zNCLmpti0qzzHiNpQrGm22R2XsgLt
+kTe6oiYrjifbPsaJ83eKXklDAEbmLr0MzndrRu3mHWLiRtaYEptFj0Wy9DP61j02utkwsWsSVlJ
P6+KvMJKLHrdc1dR0dm87BEhBSeRXsCik/yTEBLaiDe1hCvp1AyRSRgXPcaxJGEONqrkinEa7HkL
UoVnYycCyo6uSThPptQcGbPTPA6EevZz/zLbpuiiFRUp4+25ucAGvXzFEVR70IKHkJjzAhLtWUOW
lN1nMK7FF5D/p2j7EbEqp7ElNy8CPlSIEwh7T+DbxGivKLutxrPN87NuwaR3Ya1JnfnumwmqRJMs
sYUQyj5VRr5bQah6kBtT7JxrJtqEqZ6Ah4LuemtFW8DwijRG176y5qxnV2BjDz/bk8Ofk8MdaJtV
uyeEV2YU33jXiDaycgx5oU4Tm7MFPJNEyu0LE0MdtmipGCnKMpd2c6SFLT5yoExLmrzhjXjCGpxp
s47Evxjpb/zIQ7mPCIKAk/HjfWEd92Cw0SoJgF6IsUHQ1yOisTmQC6nHIabx4HHVdDlYTbboyOje
YSWtyagxPEkq3+U7Gz1jwekR/MYH5DeY3PPJBNIKPkAHFbqPQyV69XqCXgzdMoBYGvRf5fOWOlbS
Gqz9m4PwAnIOjSjUjPVrSAYjmmwORmQXBZp8edDtCq1wZoOvixQdDXPy7TtukY23fvrfzYenhU1V
RO5Xbv/kF414fZMGrWuI1bp12t5aItjY2pUZV4dZh9wTafJSq0geBLAirLLsB4rQrRVyWgWTgKLJ
MkB+RjXyDCpfc2Jtpk8FMKvUPTAbmsAfdM2wcbo6jY8MppALIXwbm4CPgI4bjvhQozmn8LrcvazS
Y8j9rmgqbqz1M9RjazfBvPEqGovniqqdQDw0/A+VQmcNwgXnqMtZUycgYWGszHWMNVv//fetFTHp
VHPnx42GYO6DPpWC5CFl7Pl0WWrko+9Oibaa48BX/QOoNO2c64dfLsuPmyFOyRBwfxMMgnUt+FCc
G0KdV2kmT2ZRbUNcA+vMx9OfcqwbGoApKiejTXLPeYACr7GHS9DEVzuPhIGN9/HJQ+HYg+pt1359
saNiK31Xa21ovkCtceXH6BRMKBFxxnvbh/9HXJiq1Fs7K12qitidKXNJLRiSR/01OamafAyRP2iG
yYjnvNgariiQEjDW32dfmAx4FtWq8flXoT/S6ZZFjbliASQAgjVTF/N5d+jMINU3AN7nj2/1h6D/
QH57rjBwejtJXpkqTFsFDZW/d+8t+ug1dgJz4whlesNxJG1PqxZ7kSM3JpND4i9U1tkbEGDJ7fmy
RZzk2YOxlMyFhledLeA3+qRydBBv6cM1x0YmEWAzrVTMNuAsNDxrDAsWbwbxbe1vD5wISyrGNjEX
Hx0Dl/7TmelZCx2ekPHiQiUcgteY63X2/Mc4bt465tEWKy05ARql9L7E9XJgkgzxPjhoYbYKkTvC
fYAdfO9bW6kjJYXnyWvyQKLf3BzC7h46gNYioVYhGdqUiIlUcuT/AkUUAGI7s9FPYlzhaV8FSNs+
qdsps2zroDbuvYg8wtexKlr9BmAi7PgHZlXReHDxDmAsykjC1AE3Q625atvw6eDulUkb+I62hO75
sR04Cm3rmp1Mb1dltVDmnNiR6D5oG5Rkivw+N7m7AV5k1GTgfzeFW8e9FHjmdKQIP94T1nuwpUw6
596U0UbeaKqR8uqoC0gTo4Xbl46DvgRMPInM0CWzEXYPBGKmzQFCbOFUkqiqsv5mMSYXtDC+q619
WjhYxNDWr/MlvO0d23wlKxZj6V9TP+xeHZtmJIkUeMFAcAESJLQK2CKVbw4lj77wod0lm25FeD2H
TejmnBUwOIas5q44UJExO+YxW/KuGYtn8JxyRZ2aqbfGOiwuPoBtbKtMJchnTysyKBH3DOjQnolw
uPW1n2mzQv5Dqfj1AU5KREQGP5iTMXpe5LFn6rgwIWd7RRvG5n7WqoifRd8W19fUFCavFxN0w6yZ
GV45Gb5vSjvwswQawJXwKTxGrnd0wWFSdWDRLTu2yrEtmEMNsjghWgSbOqgXiBBd+4XCY5813kzZ
UM0yxGMUfpotjDjD6LBL8ppSBRQ7cf0sGR9hRSQFNWI5H7c203y91bxBz6Lp0SmGlnBb2LdUoYUv
yyr05QAN9RPyfnrOeHJj7hS6gVrPQvWziMT3ZppwEdLLKsdNh+pRpKcuRQmz2isgQyGJK1P+jLRb
1uIkgNLlFq6/hQxw+S+N5KqE66SVns6/ovUH10pudZI0lKPNx0z9GH7SydRnMOXdpKdcvsAe0Gvp
x/5hROdiHJDa1ikreLGhcbbub1NNWiQQdeGzwE17zeQBSpLNmBSxgsXJeeH5VpywVHsj0qGcLocJ
MOsjLWtgFpRbCwU8/3MHQ+P3TwWF7Hu7/EvytLr8rhaJUMC3VvlCzJONSd7uAGzmCqf4T/3ZzIsU
ediOCHhU/G93G/xBS1ZuCPZjYyriiCsxmInq+4pQGrw0e/eTqkr+DM/Tk0M+KneR91nqt51sVZqR
Ip/2UP/wzzSZxhkHT5GrM5h11vDUuFou8z/W1deIUvFuDt10itXAndo0wl1gnX8rjL+ZfQden56r
0v80Ih0iHKn0z7qX2rjzPAqkRZhykiPCYCnd1f8pfmkEfUwPHiwI9LV19bGVROVmjNCItvxGIfu7
aG64QiIjCtprqYZZkgwxuczjAH7XEKg//Vnlan4dFMgyhIEz6RJnlV6Yln+Os9u9Gk+oAU8QLiJs
FlHjvGDqY/6kAOUGYHJNTHyMRzzmsna8RTGFDgVtTjxvNj+Ct74ufyld6FX+ZlaMM4UGmeqPTjXH
Y3sGxCSFP3CI7CJRvTLHd0fa6iaWK1too/1ItxY4EpjPw4S7gKgUU0ZZdilhsMG6cmX9JLnraGH9
+W8pGdhj4TE24gyWjfUbfQSXzSPLaNoaMN55f7kGFAg2YKx1H4n0KVg2bbdigj62JeGubwXGicSV
dEiEWpMouy+IATISb7BYz2F+t/yxH9OsWjN/nSlYCLoTKY2ex3gxDgq6+HYr/IwQt+FFaN/i1F2q
o+yW080HW1uinnwO0x96wUXV5jYYc21lVPk1WtYJPo94zHkO4YuZV4677m71VRicor/gcJIIr9GV
PA2uVZvxYvaZvxbOkaesaZYneud4Gca+DnXjZbno7LTYAaQGr7Kp3f4JjrSnNGALW+52pKtEQPt3
7DLu1rQ4IQHvE1Cujfa3Km9Hb1tJdI9G6Gn3lLBuUCbBsDTgWLK5lXx80y8C79kFHp2uYpV1IfS+
IOvbS91wuJ/q7S0msnb2yffchyg6u5Lp5VDugZiKhOqgstLFQmZ744jfGEu0pai9wNdlTIj69rIp
ZMqaxYqTYddga0tmw6rDqG9FMxMDmihi44q4qJmneRQI43KxgbKTNlUC34oGe1aRV542XFxOLIPi
4i0hnioJjSlUaVC76BshLJ5b6uZRuNflk8q0h0kjvFYgldw8YwbVuX0rT+ajgX19QGsONpYL3MQy
dvcOQvQkwtzVrQoMkkPd0EbRLUv2lmN9cabuv6StRdfKqlGioVEKLup/Z4S4EQtQ/ufWFeKiOVK2
ybgWnTi7gVUWzHj8S75vvx4GME+LqIPKN8FbhTRYek0W5VsUwHeUIBBr+02QiIzvNYuUlsmjKHIh
pgNVWwN1AC+xxI5wudCwAqS1xSjGt3tHFSEES0n/jBYGTDnV73ULlNw4xgRfB905V4s0L3XA+YhD
jQqUcL3+BmfrZ4MqH8mArseL9KUmY7HeZ0qV2Eeq7tUOAT54jn16n/nvfWCf1qrAmdk0GAXRMoeq
7llkZGuylv5bb2WxMMNTXGIGvgNimy3YnRTdczmoTnV8xhG+xrgzZWtEYrUfA7EP61OjRaaPi6hK
BWmnvWR3nEfIEHw6kHvSsKEVkSktSTwiTscdOY6zASXoHoSMjjBrF8ROzt//bIezJrHsNOYa1muZ
lyCnIaTiz5+1YAc4oOiF7vsagbnrrnWz+7UClxzAST0sTt2fb4mUDZ3k0f4O2UXrnaLXO6G5PRh6
ghinLuomJq9FAeEjdhuRY54ClLMRsjaataQEEk1fUBlxZCLmtmL/mcJrFHMvvGndJ4/QqBk5UTvp
fH991zcn5ATicpNY5TntFy8OGHVghqlKaVW5Opc+4/iuI8bRpdXOtJd5t25ylgHW7I5PTaeAKK8I
SvfLV36X9dVDdwC56vtAbZZ9T+7Cn3iqesaq0jLVB7qF2uurNWYPicF3AM0deX5/bbduTUH61Es5
khDl/x84p0mAb7/CDLwUT2Qwl40MaxnLQBwyCzgA6/NEoY+aXhFP0o9iLrXB99jT0p2Bh5K+PeT0
q8cxRoRF58Y544MhapVKNi0SJ7ixvLmwS9SNmJO9lLXtDhBeO7kRMm//h4A+CiDnio0GfZFKQ5b2
yncBOj7yHQgFEONzfJUbpwlK/wbgU/RXxDFK3fF/UGFXURNF/8isSHajB8OFh4V4ceoyXcXW7ugk
EeKv1cn4DGbBkJKT0FxWSzQLNe6oJ7wgWok2hGZOrz8BcltBA7uOg9XqF6shvPl28yUGnjccz96A
79PDN2A2jgzJ4lpOaF7jV0r0U2TF0wnun7JnkQeINj6Cgs8QeKcnEsqeiUDJy3FnRhvGMDIf58dg
fjr1rELJ1SHJ2MAPNidM/u7mmdZms4AdrqDYocXDMTGXiOdp1Kx30px7wngk/sbDlANKjmBmS+f5
luJr4x4YaMQrFE0Cin+ZotWoA8UPirqT63mhAL4Ddk8FkwY2vihGk1EeU3noh9R0wvS5EuA69PC/
BztUsazj6Jd5KO0qNiFkabiwJ9Tq5NLzQS7whO91Tp8dgHBsQl7bv3NHsnjvXKywYV2yeQGyZWDs
B3MwrobdiBk4C1F85PcUQ6qmnfgHpRl/EBLgKWFpJTqEYxqOeyt58sCaTCavDxRdA1EJ2ZFHS3BB
pvbJvI+6s5acl0P7FfEicD3M6U39eal/sE2P84tI6xO7T08Dlq3780fn9RvfU0/arj5Hlg6lqgsU
lwUJEOquZ1yaCwCgwyKlYSqEIQGYXYDgwZMse1CJfPO8OEnnF43H+iNv4M9x6q0nKYPRFmKDQFLw
HGe6ytwZGilclheuWns5MJ5x5me62t3etbC4OBxa66D/4qoDH/20x3STel98eWCcrTQLBjaX1Pjy
eecGE/Uv/5ZNiT24US7kxTVfdMn3AALVT7JTs6LWJqFboZSWGCqWDdBdNacozW7iiY34Bnrk4Q4I
enmXI8CHWk9CvoqZL58SSC4W++bUOQoA93XIhcXVdS8CNV0j0zUzztUVR7suEI6gV0zATlrCZ2pl
TeyopFhS+jlbgzkJEEj5s0TGKaqW/9dbgjPMp6nnW7LgF9VA8ehA/AsVOMESM+8jFv0w1sZptWPl
ck7N/5V0TD6lbjy0MqaRhP1N7zBRRnOIGWjmhtzzLGY2TvN0zP4bcb1S5fNBxXbZ0zJ34Gnm8hjH
5aqhsGrMkvN/f0heUYOyqvJau/+QbDnXcOypppRJqCsGZJbO+a57gv0GXX9OPsVrTl4UisHsDJWZ
YGn76aY7OQAWQs64JbJ8NHRrSL/jC8eol0yvZ8UD5nSA6+tTF1oUYESuedIG9d2posO7L2ue5bZc
Z03ndTXgR2sUMyzrhXxdN6nkqdvBJvht+uW9qBHLkSe/LW8SOSjVeoBVnOTr8ww4wJfikKP8HszM
uwcWYbsdNZd2OHllDPbTCqoKenG5TNIr0hbTLYJ7LY5V9yIML4VcYxhutFwTnUvubTHR3B3lC7Bx
TnL+6eXUYSsMDJiGpI5QS/5HyH25dJgVO4huUy93bM5k8/g+IvrtVfKtnJW+n0sY+Ia4fgmzO4Oz
gEecc1IMHkI244ZtzuHrrIlYRqoy91DubV7506yo9obbx8lWt550EbK4emvfTJ/FMTli0wJYJnh6
/iDnv3pTPFfs/fHBUamXjMdJGFKVTMdBZ7GsCNL2K6OT8lsS5mLaPROUHsGb+kexntN2f+NPOqfk
6pxQABuWqGnq7lMfV3k09LLgKDupNB9ND6DQidRkm+w1jkEfhgfZxJOHjIdgsxwTfboBFiXGyzBH
7mQkP/M8fIWGL08/JSujKNKc+4b7l7ZU6UY4RfB+jMVLxCRmz6dD09C+AdyA9I7Bvwt+DO4l/sl6
eK+VbML/FvSPfXLbEysW30Ex+9LkyiWDxqPVgTdm/TdKNQswsbW1GA8ZMSLN1x5lz77UOOdDJcvz
3daCqjPzzD0ESwPqJQvizJDTHGyegWDOFq3UtXnyWOTSH4J9iNl0xTPCKZkmlygP0Oad6hXRJ6kI
JYQt9SsgCKMLZx+cY5RuScW/tf/0PZZE0eRdCEh+x3TRrXVArp0u15Nc5ukDFHpNFED5PkLVnfJa
Yz3U2mCrXfkMjebGId5FSs4N3LibJmQOrEoGcYq2Gd9SE3RoXNq+lqS6U9m3hCcuU6RjIB5WOvLK
WulBuQmEK5YyWj+m+rDYeQyfNYLiDKMFdH20g7LGO3bpyyn7TteW0EAlEde7b0igl0uSRDqtOqET
I07dhgnE+SvBN8Aiomn4Um28qw3uRmYMwdhSazPJBePsW4tCUX+IDTEv1YjlS5y8kKwv2lO/H+O7
W8Nr7DFiAO/y2BaNJcbl8JwGQfE4mKg2r//3k3FhHXXmE3OTdRShdhvZve0J/HlU7ZqRv6ktZMJb
+jIeYetCOltE6d7T3TJXmlmUfdQrUJQm59lKMkRak0xZyhgVxZVYlpxfJvZbuWsD5WScP1f7Sncu
BJMzmt8NSJedjjnwpeVdAXca1b2pWMBwMBKh+HW+Ksk8EA6PTkVCRJIDQ9fZIrvemvQmgS3SkQK/
xJXyC2cGVX9EB+XkPIZzl7UZD7Q31cxCHwrPwTkMAVaPWZ0a0/Xn8d/8/Tv5qUgtgWka1AKSdqUQ
7Jt3Jh4s7iagUf6JZP5KcEQRa2b4se+y3moJ+4ecXvMfWdkxEQrJzRRIA5yO6v3J9MrHWXBFNR0T
8CT875PRK8yFH17wJ87uKwl1sa4S7Q0J/jbp3LXkVqB7/xe7HKDZAZe4nsW0JbOETBH9z50l9zBZ
iTEAiWGa6YR5FcPIXykyRhEolaFobjm3OlzBy+W4GGwKTZ9+Wc7nxX9hPvso6X5ykVZp5SucJfOe
bbvqavc6Gt5OOxFxm73YHQjOiYshDxPj2iB5SvCl62v1+5duPNJL2QTIZ88gDEiP2kS9LtamHFMU
eIkvuVqQCaDkqMenxELC9eIvt68tsRiRiozTG2rw1VGslqSNxOnWo6W3AUHvWnI9cdg4xrNb5Yw2
lYkhEDamEBk7y/ON2Degrc6CGEQq/yYeBOdmrF27CC8Xjy/ZAIl4JuUS1nu0zxRSqANU3wpLGrOp
1jytEmUbrFSS35OGmQEdys6digibZtdQbMkVQSLgTIaQpCKCeVJVFbEkjAdr5kUXzIIXx4jMcekM
xZnXsxhx+3i6+GtaegpREjrKt1pz/hhsX2fjRQb+rPg0UL4MCIuzcAH7Fkwo0PK/SaMjYlO7GqJK
Qz3LyWZZYhgjvbJt8mYiyNbNUOx6jLgj25ZGGlq3nFdGDswm/OSFAUHt+g+GOt+Vybdn4yd3FWP1
kOz7d9SzIdiraZ1K8U/s1iqRoy0pWGCEUruRa/qyLnqZbMfy0jkYQKVFRD3CQNgNaCuSGJOCTfmi
U3D6EGFr+Jtc5iLoRoLPxucrg4w79me+nNECuoRWdcfBUaknTE457j3en+UDEmkBnemiAnGaJP+K
DH6lHOxWitYK6iYyd9RMGkQY2DVso9WRV7xmzNIMckigURUcS2UcW3Q5bBQn4YLrQiyudaImuTAW
dTv6v+jmGRnhlZ/SVaR0IDFluza05SUvCr/fDTvC0qkC4Zyfwi2pIeZWVKoexhPLri55ikF6eItM
pdFLZcSxJ/7rlaZQrNMJc3GvEwm+TWExyR4yXCrtNCku8VmoDPWD+PtLH74vbxmrgkgm56dvELz6
UaOpLMntcg3CjFeu8Fy/oRbQ+Ls3gVubIkfbNEuc84zYTj665xhRhDJF1SUZi3wvB6LQK2tRrwmg
Lrzz/UHl9XPoxVWAM+pHuBClHWAcT4B6bVpoB/cRPAgyid/0wAgSDFCRXRH2kPMMx3pADcmx7ICD
4pCL1ZcIt/yJUu2QcVEwgsGRgB1ns6isGvgpzGSsbBDW3JeynoSlCRsTcUdaaXQUsrNy410YpG71
yCXutvPRbXLIWKA/5XN8EI2vTNSbXyiKkbEoqVwIp93g3365ZNsrsx6o2oWO+A2rosYfi3QMw9V0
aJ3e90lAwZkl5toMjKVKkqCRpVLh9OxxualQTcYuuadu8T4pvQohijUz0SICEpI3HsiMFh1J4fm3
PGlZ81Rna6//JdyUpif8VFMM+83Fg/4cqdwvEojKX5SkHoZeHi1FRK8lVF3PxxzuLBk0npVQJ7R6
LHWnUJvkb3hHgLJI8PQEwMI9inIZKJFf8FgZjQpJthUbYMc1HbiiCkbvLx1qTh9RlwosQb0WV3ns
2rUGv05R1MiZAmBfmlyia4cPvEYdOmOnwbNPvpTR1TDBNyeePdiCnHHHA3TXMrS005jjLp8szwNm
F+ezas44HOG19aRrCYWBAud97V0a1f5eTJMSNjCvYTFXkImosIn0qmXigGihU6+URjpX+x6A3hlS
J33F3mgcXvDA2HSUV7l8/ZTXnl/Ln1wv4+4yBnd3TOFoxWZJ3L1VejG4kSAcglyaAa79Z+0ns/Gz
s7MXD210OcMfqIdkXD0aoo/3NhM9H0QxjYur3cLZMpQKJkT7J7oLz6SCHSfCRuKwGaUMIa93s8Ge
O1t0B66vs9ZRzGbBiUbIpYHkuUcSNStwGKbgxyJGwkWkjJYyM9JruZLfWqjx83FA/u0/wYA6GG7D
riy8UA02Cs5oEPsPgzEhl0wdV78BW1ndT+eW2XuTosGtsswBWp3v3UJK7yFPyX/FqYhH87PNximY
oBoe4OSmLX777HQR8ImP/PjTS3Y8n/yV4MnCHtiGlHWLm4wS6jh4FahhbkMas3d8KEPicbeZXDth
JsG9VjWm2ykatyHdhEWzZvwBJnsYgv//C5uFrLaCo93CsiAFiBEbYwxp6L/YCYWypS+GcAiQ5J7c
eKH5J96JCoZcvRBPyaf6VOkrBpD7TRvp6DzLSSbrGkfTnlu+02o7eA0lWAAydRFBVrLS5JEGzBDh
odp5DSb0DwnfMbMXjtMc//kFJQjO2DU9oARbCHnXlYcVolmY5Dp9waXq7YOQwDGo2d4cC7vSH7Yh
fkX8UgX5vD2zxMP8044/y6/kaPQKxJaDCXr0I8KLoY3yOkuCmqjEZSpq3DZiaut7aQaCMNmg6QfL
DwvO/uWxnavv+oJka6cgsYuag+MYiF0S0odSVqS7SB6ty0l0Ov4/qOa7UvOlDOkSsDaUmtjL6KpJ
LY/XF0kItZC/8WzOtnA1/FyWy6SKtbdiq0G/Jyjdv/Aum0Ey0XzDNbiai/HIB1SVdYXA8P7+gyry
buDwn0cmpn/0nqZAwu91ahiwZzCQHqsoYuEnIYvksrBGFF7PvE6BEWXyUzAf86XMyVvk5j9aeR93
RVTjNKpENs1fsGtZXT7NA54CtTWoT5VA/ul79t4d8B+YoEczhW7Fx7qK9mHd1Gf1QsAZdOIr+pYl
LhSOnNQfWC5+XRHHofJPnk2HWlLikAl+crwqRX00W/GEgcaAsHj0gsRCShgjt4fMfxps9fvNjSFL
l8IXmP2bzuHE/tBKFEAo/7M6IcSOdLpzU6s/guJpqz/3S4Jm6di2YwU24bGVOPPLecm67IGr6eIt
NyQYUJn/Br7Nck45DVqwRixHbYfFPE9wwDsOxKdnM7WmjtS8QVYzqmHJ9Mqrhmjpvr5CAdkriOFB
TjYSqwtTFdOVwme87glVcii0e8+Inx6y0bMyaIzqjDFlZnZu6/Ro/GcuUxbHuiVrd3wblxPHlX4Y
4CKopXGyaaTnmlR7BR9algQbVYZpJrgRAqwjidUOIyYVN2sH5x1iXDV+1z5j8sv5euzVYc2JsNHG
vL//GcIdM7IUNW/lIlnsSsR6ZjpkBMZvuy9YC1U++nxBeHKnxJ9tSDBpAHm6zOegRC1VxSd5sdoo
mS50ElfTu7cZScxh+voTcgPSbVaaLs15fTIg5ELOFiHKBFzsNl4sIJ30A8acNaoFh5kJ6SXzEpjv
3mk4siWTIfX831iNegMKsgebKM9zwSmzHw17s/GJnSzw+KvALag/XaDYmJlnv7O05UrjzuSNepoi
6tNmci7JnywHdezgH+LMWIfEhQBkEY51cqbcPGXi/1EHGHcQCoHJHzSB87aO/s6R5zPucPXhTvco
jCVJ4rYz5cfd1a/XCa8gzFafd6vSSxt8kO9cDKmFyrOrNHunyV3lJwNlgYZIMFXzA6q1HgSnUQ5y
NqX5WBwc6tmeo3fOXUMxx/WW7dpmZLSyM3DnveDKrS6Z4kfzOAs0/T4fnl/skdFs1WpbY8/uxSaN
udjPdqvDj0L7OTBEQ7tWhs4OsruA3prgvJQKjfLqtXsIVc45tRvRsooG5v6uwKLAJ5vAo+aDj74f
BuND+QvET76Ah5RdkwqEk8OPUg7fYxHKGputkgcgVoqHd3vwxWryx8yPpXGQSojqT+06HSAKJJNF
ZYI2ONtgT8o8PEDysH8fZ2MAfzQ8WyI9/57aAxuWiApr/ZDoDXomRX2IPXoJWvbT0OuNUknACmbU
OYUFKucdpccuemiZ0dMSuQzDGvF9Rq4aN3RktpqrdAqN4fPwH02XgjHaGL+1beTlrLayQk7LTOFe
qBwS00vmlknGE2mI9Ncbl9OzPzFh2xknLzHqy+mgQRelNNlkXqb5Zp73l0D6SRqwU7JmyIebFZVD
pcRDrEu9mCal4axopUWOj0qYsYNl0bOJ52kDih9h31XtexxDZzSWGnBzml8VwgWhNaip2dwAAzDn
65vz3e9sjth+9keNDN/dsl+WLesKjoVYWD3DNu7kK4KDeTjsn4/to7PpOxjzPuZ/NQxfapk6h86d
8sFVgkuFJfnbY1dyn4T6g0BFFH4kLVroqCPODWFoU+pH9pyuD2l5Kx8KcPn6xpxXNACsZC7yrNIx
DinxMYX9l2KaZQ7cwuYKQ5cAT0B1Snh01jLYttykr16DnXvLZoAts31PvCvSl7XgP0jD6mHvSTt2
4b95sYSPO6KgCJJfYwiMYt2HrAi1W8IjySKLBWdP1zu/HXupYMm/UqEaO7jnpXtoGoqVWhEdPPez
VZeEocPBJ9pwAxs0+twYca4bPSRoAEDzdb3fhNMGISCERBV3ET5nGVuJVDfk2QxUKRm2YKL4iu+7
H6G5NuKMYBmXAroi2as3ybD6XIIgul4mePN3rD+7k8fvMP/9jvZPmOgRfGayxUtv4pKJjcnQOUn0
WGDZYVWtMJj09lqDzDrjMdiVRTWxwOjmD9QjsZHFS4tF1vjZHgfzzMDHvzRZCF/KfhmCYUXS4fXN
UndYSu1pLpSzDcW/jm1kNgkpG/Bz3DX2O6U5wk4y83+waChtwhnNIodFe+sYjQLbAK+Cy0KyENbt
oxruLKZzyqS7INc+aOIIMPRPqmKa48xG48Y+Tcw5qLV+TDefUP12Hrxn5Pq3iiE/BX9YUYZGHMlA
oHtFW+jONNWRAQbH/W2ASPLvWYYMjIuVCbgtX8ns5+WtvLM3izyN//2j1BLNOz0VPcXfYDggD7oK
yrnoqAu5zt8wfbFoguDa+V20dvp6rKeudB/j2kV6HSPCQtQ4hhbS/Ud6kgrIEr9DTskKKzYzStoq
klQVpe31AIdJvDFhDNE/6T+PDb+1mnE+RciA6S8g6ftKKEQB3AWhLWXlSwig1xbpPhb4xWxb5EQf
uxQLaavZeGESg0KIMJHNKGmu+I8+shoPY5UA3Z1BnERAc3ErGMDyNP/NGnBOJL4BZ8j81EdR9ztN
faonKr0dmUIUjBBE1xbVYbpGdrHtuy1StRMa/yaBUC4PmDm94S0W8hMng4jc3XY5lPvp84v/zvUV
Toh7LIZPZvrP1N7vcRV76mXVbXPDDQJjIYIWqkZoQW5oKbDKHuMAQGGnzloBjeR2b89pccYQDCE/
e8OTlnIlwLtfTOI7BgRUKjwFWNY4DZm1BPD6+bnc0AfvJn892rJW4nF5bzJJjrc1mXJc0osWvc+C
I+X2B0QDIQLyCIoq5yxTDINd8NyIVCFxLtzEZtXSVTSkIp8wFVW4zMXSuOh/Wz8IAEBgpibQuKDk
PrjiX4nw520laaoCi74b4FMWUGTaj3xbEYDJIGCBjbC2EE1LfLYR8kUon2Bpo6/d5UKnkonDKFxX
NtM0wMKEgTiKuGdIFoj/fkZpSgKIN2JJxRjHt/imPJ8OA6en4KHHRn2DRBX7TkSruR5NYdowCL/u
Ro8zxPsZQcKHY8niKgjJM0ope0BGCeccQV3mZsYinDZ6d1WI8HeBdMPwKh2BkBrmV/fB25w1XBv5
Bg+lg7A46D5YNT5APHP39Jn+thmd3q6Mm+eNnoJuMLU0pzj6/ccuVis58IY4pPUxtft8bw33PyHX
0BqXVpMLXevxA8bPkOmNAv4RV024ZGJVg/by1/ukKuuz4dnhBVG8KfzkP7TZqQU91wroS9vKjn9F
gonj4/AUy15RXq3owJ7sqCRc2TkLpSWpnhB0orZOD4zEhfjDeHN0khdGlIjw42RymxQLPcjXjcLO
fqHwspI9S6UvYpElwqi9ycpzZhT6g0Dh0J92xa+7WKtpAelEmqbOTlaRnn1ZW98del+Rp5tRztoZ
WTObZlvsrAXDB1V5yU8/DAA4w/U7Y0+xrPZrGwGWSCA99yVYzwmayomSEZvUxlgitxwtBaz5Qn3V
PGeN8EE1AYsFXUlkad3E0Q60K+MpO1sOWiwrm+p7nbHZRXkDLo7rF686DINWZ2X4n/OCccBt113Z
awkkkd/+yChtppQcB+j1voMi9al5WwzZYjDKW8RqfGwUNrr04hc4Im+gLJZ2q05F9BA/cSaQjR+7
wA2Yc2xLowFa+uX1MLg8sOIExHDE0RJDgDdl93XCaNhhWdAd3k87VCpHfKHgeRSCLmZBJgDgZn4Z
yJyd60XT9k3338oz0JRcbNRIxM8sKDwMZSGB4T5ZpNpp42+QC816/xbScYervRZU/PCRKveFB4R3
a7D4wKkYCzuf4eO6yED8n92D7JVwsww1H+v7lKsgzbUiqOja2l8PvmUq4F7+DuLgOqLbL09yPVSv
zSTVdUlO9CIH5JLa9koOTEwV/TJNsZ+0neIn8oN38c5hCzo0hVGPYLAOP/shkZHUA9DG8RzsffPj
onXgF01jl1TWibJbSxYeIqQmm126//Ysyg7ySkLT19gzkbO27fepBsfL9OhSe+nNNeRMMe+LOXV9
3y0SW8mWxBto2/pTvH02QxuhIenRm8MjNN+66vfJv8BOE6X7Qq4RgaNHZ7/fYbAHbDO/iq4j+1E5
YrQiEKZMcuzvnEvYegkp6dfU1ac83znPjwUtqEJefA7IGxveJpAjT7ssFoZh7DGwOaiQNsTvMni8
+5R2iE5foxXstpqSDOxrKRgbx1tuQBk20CPb6FIt+8gW4fpS7AX+66sE3KCWWgWWFuFPIYHwVM1w
N7WsMKIrQ6pmsAqYAjkZ5wsaxvslo1A4HbAY3Nqw76Z+reIaz2wBbl1QZWJ0O/iDqPW2BrSax87k
gKuOXDM4eR/ecWbSnPsVEDoYrH3K3qWQgJDgraJWGn03loAxQNs7ef1i9RTzORATTEMxWP9J84Vy
eR1VuLAY7eGPUYajcDZIZV685tVx4isyn4VioylnNGoldEeeDYnzCUJclLiPs1dfeguldFg20rWd
NaibJlK10vF3IFi+DvBOO+89cjaF/O66O3qxWryW1+BkaTMBpAi4SVIEHRV5CwN6oN2tuQmyN+F2
ISzKDumPXasmuYCxH8P066bNJAaCIVxh9ZiTSrbPGdWzJOmQ76xMJ41YBxLXUhRDyGmPih8QFb+I
F1MjxcT7upv5OHV79cl6fIiOf8sTG5ARfnX0HKxylKVWLgVGIy+fsnQdyAI/rHzyKyth8k37kZw4
cgrVRlOWJGdSp2ZZ3dIGSLlzfguCAwVhpZijpsmJvPY7CyQ3NA6BGw2cC0KiY9IVePNz2/SfzlRZ
tga+a5FZqqCuOsWZS4FY2+LwgL13U7VZPL+pGH6vy7DpJ8yuKV51kfti8oPFLFgciiMbMSyrWFmF
0YObKEAnqvIjLvcX5cnOgC+PDZfR+kA7wARsd6SHJfNp3rG2DAX8ouSuMVqOOogE3eN8/J/ne6lJ
WaTgm6aieuUlYb+crA9vUf+IFIWHT3BzQKMD11BX/itp4PfvacOmm0gsJiQxnF2tN5Y0zxkNYL5N
H2SZu1MybnjeRcYRWIcgyuYWAh/HYzrNFYZTs7xlPECFObiqpTRw1F0yfFVXBYFwEHOmsU9dQaaF
04uW32uQWV82RGq6zFFgg3XUa8q1nwh3EzuyX7EMc8CSBJV8mDWZbCcbIOQgo4vBBatSQjVcJOzQ
oUsWRcQPh1jmVuNYwhSk0rJ3CS9nN7PgldV8LsZldhr79SjCgnBzA+AoMysoSMZ6tIbyohrjbB1t
Xaq8bRKA7c4DR6xZnBEBy2ZDswPxjFG7mn0eIaHhIdVtPZL9hwHJgO++jqP62ffhgjnlb4oZkeFs
SRyIN2oTd6c2RxjNnqAtSoq/lZUwfDknAeToFsuU1HBygCHyYUEn5/+VK1MNSQxgA/XSs/yUbL4g
QEKqnVd33KY4SW6nn4bNwhfAjAowXKOJhX5Aw2yJ+CQfLnTWeHQoqm+sqAvTLy1GNqGYX6YEyUQr
hIcdjU+7H/FtAdJcKcc6s4GAlKrHdTuyOQD+sgyEcNCBaTyQoFYS5XnWLKLyGAxtAFUCZunacWh+
GBiHakZBSE01R7KQvTmeOlkRn+7JXc9p5b/jxDVz6IVZ8GM4b3xHWJWrlylYhuygaRuMPBs81OMn
j8kqfMWei9L2qj6rhbfqONFCB830xcvvRh1wuiKQ1+MN81KULCub9WR44sxtE+pKa3O5V9ekD0gv
XSy0HCBM5Cl5vIblnwwrBMCzhShvJfzjblSzhr7Z1FSfz8/Xkv69nj/bhRpi7/BSNPCWUNIXAdRF
WcMVYIQVwuL05CW7KtZlHUP0Z9eKJ8GtHEQp+Dfq4aBwcLhGoz+rVVzX1ks2kBhJmDnqj31QeQsj
wex2IazjI+8DX9ebCip33i6KHcPOKCs6MU/YeiJ6w81d18ztZNo9XKxoY1qDwxg3C8tig7jNHUqw
JjaO0t5jcOA1R1dVUadlDcLjoidZSAo2C+OZjkniAQ+Yy2hiP6ZQJkCz/QSGnl6tiD8Jf5nD1xiP
03NqGlGffyV+6SuEn+s/VP+VS1zLBGHxkLiiwxloTksyl7LGqSKyu51mzHEqlpYiWP/6byKp9F+l
V/0cP/Mk7q85/a5PqiMosbpADR1p9s/UMlCb8ZpKGVYgirALs+WqjtVcEfEgrlu8LrN4+ax1ieHg
rR31xsWKzZG6CFWKP19HzbVVVFxaP9VSWrxLRr3yZpY44UHmoaYMFXgMenQ7e88ZE8T0qLg0prqw
w6L777ZPWvxtivZtEv/Zef+ZoEog6f1lRQe2RCDWlL7VfX/1Lh6sczRsDk4YPi/1dJLMzk2ovVn9
g96/gMvjP9+g0+kaRqXAAnHVZssaf4ALefkWyLF7mnHL0CVsYQXo3ljT/mMtyMBDeMNViNBOnN/6
MBJXa7Z+yFopnLwJ1zoZWFDhXkXVUjFV7Y1ANjYeJKQ9N3SUKP3n4/wFoORFtg8JAnE7wjuNqZxp
2gbgQXvGYgULzUm6ACu/Nf6QeZVpZY+0ON88/zl7ssj32Mpt0QnwU2reNCSlozZs25dQiH3gaJES
UyB28W2DzUpCQAgucDkkIbOQSdd0lvx/PDa8+hbwsY1TU3Rzh7W6rr/txBj9TGLlP0c4CkIbEeMk
/Z3R8bEAULiTnwEj2jH7MqgSo1PgHxZJCMHtNlqnxxwpnck+ZgBDGrCapEqrTmB9zzD8+4MJdVAi
zvDbV5qSqSPoOin61sWrU9nMuwPZcg9//Ycc+kGUvBjDuIbh3Ztw8txVr3dsRrbpAmqWVnSW+eaJ
n6PPm7UIPVI2ubybYgchRJsGT7LkcNNKz6AQxGUOlKUKIgBrGpg3R0/WeShmjGZbjMCQLOYgMEAN
xUwsyggx5Q6aU36/VOaCT52Uu2/6dNbvnydsBUWUAZmKEpFnB32ZhSHqsNSOrXTGbNzv+g1Rrr2Q
bFQWDZ2PUFxjNAWKXadWm1kzc90FK20in4a3cBjtPRA0y8Xo5fFGVE7ctYXRRjQ4wVcstIxqDgDJ
G69FuaDmJrXj4z2BEFIKTUZ1BkvVt9MqpJgnzT8oz5I4VJMYwK+R7vok+xR1/E6RIQH7qsCdTNgU
Ag5l1sswTVbkxtinnXIZgOLThE5qW42Yja/YWtbba3C3mglIsIqsZD3REmQxouk/6dfNzmWWKhhh
RdThmzF/sTf7CmX7w++zRVy3eI9DReEYrzPhpGrFr25klX6wRWX1qbt0g+vuBdZVqqcwZv0q3y/k
8JGqJPK0KRReeNq2xVgpdoqgJkAFzDaFny19CxZFPPV6y5F2oKNfb6ZunDIYzVkNM5ywT9texqgl
rHYWL1wYHRa3F6G4BvNbasCV9yFlSBBtHfW+fA4EG4VfoCFRgmPrHlVZOcTF+gR/KBsHtR+Io0M3
2bHvzNC+wbjfhHXw6634MHlGGpfo0+Vc2jy4u+MJ5dQsWxpTCbKQ/RmwNah1PZdunQ8OaM83dldC
7SsmaTq0JD9zF4IjTkyDXmFjrY13fIdGGklQPhCqeArLKxsPSIemQmphzdvK+8gYXx9IVACvoBlv
bIR3lVZRT0XFUmFlOsTfE8Cz+1PNFw/7IOf3NsNJH144znSblGcVtJnAOBjaQOK90AnzSP9UkCf+
zKt4OIX/WXp8SnH4wOTyqAb13BpRleu/dmit9uFCm6xuRpKmcll7tWKytaZS7wSfCLKnOMK7fUpE
aCV7y2KCB019ZROmFYL9a3HRCl46yO/Y9rtvd+2MeKMcyYae+CnBDoc/kxs1Sv7fff4sCp4HdgNC
ChjPDIcuPqqmA8Ys5PWphRqHvDggEC1A7+iWEYQ7nt6EixW3ufKV6QnF/IHMWqEeyJZvGFy5l3aE
pvT4moP5vodeUoMjU6SLc85dJUej7T3LwSsahjLyLiq6cF0We6jwBvbwqbm3gJH7Vd+q8vorw8jN
DHmKyThReN5uceqrD90ygEBDCRBfo+n0uTiJS+YhtKIAbt+uvCUYuCabA4rY+roLb6HG7H0S8gF/
XrX6j9/ox/kgOdDylCGJs8lutl4rjoY2dqpKUK/PzTSTO4Ms5R78V9DdXZ9HTqjdeotYqzXbXCnR
mLrVxigPRa/V6WflJ2BaCVrkyNYxmJnyUgCDOcZ2upsAa6wjDlQovvLjL0bu/+W3n1I0Fmm67CsW
bRoH8BrZEOEyiHbCIga1SF7wBJ4QFA6Jg5g4O8zv+RpL0LcicgUwrbXvlaK0lyxScCs2+5TAQZV+
2QoJuAQgf1Y/07AravSzg+3AFvfh1xGpql2BnHXmHKOyDjutCp7pt8g2OHrhjnFGPkdI0QUyQtPx
pPtTrt+1WjywQ+XDSTQCR0xU99GtepjZi6Th5Lxn/ei3fcEGrsd2u/O3fLVG6JHgikJEJe3vtyVy
v3DYrHe/6304XqS7xb2JngJU5GtfaS0xcA1rE9mdqE0yMFftmVj3GTID/gUi2gNw2ICt+YUyjxLy
pd3zQ4X/qfDPJtcdfJTmbV1NSVcDCcWskLxyKMcnWZKaEYINABpd86slrZ6gpuz7GYz/ghT0dsu2
L2hCYWXjL6zEn94v082IoGSTbYxFgbaOoBYbj7vPoAUaXYcrSq+tdwWr5gq7KJFdRkIqlW5wnxdb
tL1pRhDzsvrJ+CcbLraWsTWLot4FT4+twaN3kB1k/SIonqwYE6bvyx4I2dJPg5Bbdo7P+D/eZODW
/2mwISRF43WG8J8dlFQORWctI2sO2Iffpqd9lnAY0rlJn9SOXiiL4grEbvcEvcvrPM7yZ/ShZ/Pw
8XxFer79f8Dl5NpIUjiE25KYinA5ZRKqDgpitf6Esa0Cu3YKVJH7tjmgO5jn/YhdVG7Qc2ITkcHQ
svVb3cRIgGZiwpkqc81hW+dIzgu61rdMxTPW6BnfJX2KbeAdBORKMwfbI4JYKYleuInAiT+8R5H4
HKubHgPZ1mLuHC6POw3J+SxIGg/Jdngf1nyorl7NGQOwzo+YCWjeZ5vasM7vyz7ZfqIGkzG6Kpse
kAmhNAfZvaXEHWNoKwW/6OW8+2QLCg129Ht1A4U1MeMni2ONYtcEkD5VqYWyc3IJ7hArCVwfyLM7
PzqkWM+3z6hOYQ8uDuujHtdkIPfC+BeK/SXccU4IT3Iew4MZJbx0pyKWZ6W+w0SV/Zc/bQstS/cV
+onIdsMoIR8xUsXSkEAMx/9ZBkLk1pheQbsaKfbWZD6GXuzXraP/FzQJwo66drhD4nlJ9UXSgFPw
JkosNN/PlkxdNYdgFNE1rBATIjtqYKaYWhlpLiFCPprftPwlc6CUa2cdIiTbY6RWd2dHT0WBAp9J
fPtSgIpynFieqbl8EIym8ZCNMmnVCmHLMe39lD6rmehq9mO34Fsqjs4NHuN7AFFKcxOqCavGVQ32
UToJYdlcgsClkG8Heh2NFO8I4uoic4WKOl2TBFMUvlQ2Y6umxYGEOEI8JlelWyrfyvs41Zc3O08u
vmU9w9tg/PX5MSPGmfz/BiO05BjGxYWeRzj39NT82DnOP2fsM0Tae/MIKWlObh98MjowhgbOYQt8
qIBSKmqx3aGGkaVNQ3w0an2a0Enct/cZHxBRmLQ43/cZvF1D6tdN43/8SqQcbuNaSf8EZngU1Pl1
9bPCYyb+9E90wzUQPuQbq5t2Ic7uE15ulT6/L+O9XgpdHGSWOBJTwSGtt/uodu/EtP9FaB3bDPD+
rqxcJCpw1MW7Bu3kyMM04GQm+AZzpuCce0MWAuN8N1iJQjpSA8vccAuZd34NPyjXmfWjRcMXKg0K
1+KWXEywe6b7mdCcad5evjEMF8gkvksZfkrjIDFPmeqzsyhGPQ5Fj6tKZfuxVVHT59rM2Ucel74P
jcbbOjoxZA/s89D1eRKVYd/7s9gW/5gYTxN5M13a+FWFvVO8X8XpLVmdn5f0eA76d6aM+qny1nmM
inS0yaTzhraZ0d9UKSRD50+08qQsuRhmrjMRca7R9McXOYYKRRIiJHxe03W3tZEPy/6XwC66JYdp
nqizmQIIjloRIef2xvl5d+NwXqaVE86L/P84mpk/y/A3z6xq8naC1QL4tR1Vl4ImNxAP8Kqmd7Jt
YbEaQEKjKcvl3X5XYB4tdSsUxmBSmiHNhyAmmTjew9wDHi3MOFU2CgtGZBDChDwniH3JViQ7Srqx
tI/Jd4rmVeIWdXe4RnDlG0DfyGTf8/faMrcfGl/cK9orAwn+iq3joefDl+roVm1qXr62nEKlW24h
Mef4V4iOtdCgtCPDgqcXS647gwY4Bi4qBAR/v67XIBnQE8M+26ttK8FzAZ6bFAi0368KLu6t2n+T
iusW0ZmUeazu/jJ7Nq8oIDBLrRGDNJyR2ALnfsyRnsJ1mIdOziGeOoeSfAitK74Noda5adO2xBMP
oql5XZE1IELzk+UAi+8oNQZVu1ykpbwftdfokAvJC7tveZ8HBfsP4Z607Sr0wWS9s11RYqn+PQZz
SpO1R3JHM3oTZGkeDrzCCwJKbwfCdT4SxVd8tTPU8CEbfeffuUbZMofAUdTc/1gsgyuaCXlBwAIx
pXnQDt0PemsQ/O0GMtfIWSgxf48mBWGthKhFHa+T5D4z5ehxUm6rzwCUxLOT7JCvme0AEeKsh/wD
4eKqTOVUk2zE9NrwiGJ4dXUowxSfBKzCKCBw7tFhaG/YLEGqqdmd7+xErAFCH6nPDSAwltyegPYr
AK8OvJOb7TMz9HB6aMkKH0TIrydRkgZJRhPbdOt6MK3Jc746YhIjL6Gf8HuDS9KU3/zhDfdyT44q
Knq+uJWrJkui4ycOINvMmyDrETtZGVQ5v9zJRk766YCk9MnjacOGyutkqtdLI830i9xPnsu53O60
iyqAABJN0fe20Oyz2mOrBUnmsGS6e6WY77lYoNhIV8MvhBW+hM6+peoP+OvCmWY87luXHM9Eskym
v9w0ljmeLyNwzqkCe/QvfY4Z8JallnTYKGPfmKO3KVZcrHTKs2xbtuQLx4MCt2JSFES9/o4lKNuH
6E4yUzOAmNo0bCpzDjUa68QJo4oQTVafLM+ziR7JWTamgpii8pfKF9c9Rz3sRcoekgoIAZ1Qs3n+
il2z8thQ0K3Jmir4DzMznGjXKrXsNZaoPljVDtJIv9+0DBUo9fjFiXBdIqBc4acvtzwZ82qIGiL3
Hwl8UCtSym0Vf6SK+AGpxlihjinpDdCe/i3ewTQHisApXX1fuo09iCLHyhb/X5FT9VlrOR3z0JRG
5eB234BUdhpy+QJdSlDxCiRKmIPf/4JwVPKTtDHW7Z5qD6vecdfgpDyyFDB7VOesfzEC0PuCrFKp
q2FcyVWdmLm6pINhm0UyzrVLz1e+0akqftXEmPx38HrW1kbCVyvPEdSNYaNDzPSdPtkMxq5pUPkN
vLwT0uqi2jTwKPNqfjcgEUe6cCGuu1Y1D3Vy8R0W9cDCYUGd8HLadt62qAbrfrr0h3vBfurNxd0k
6yMhxEkILp6MYXRJ4oNr216xjPt/t3M0Wx3TcUNLj4JICUTf2cISc8B105U8SqpBFQR6zvGy5L7w
D9JRD7AD01Ef75QazLGrr6EjtY+5sbf/cNGC55WocLsGimtv2kh8QDhA/4bznS7FCswcs5aJNvNe
BYXFqduDp5NIfn6ZLcnE/4i8ExpPpa4hurOwjmaAvLJ9tkpTp9ygfWZDgPx4oOUuyohP6269Hfa4
AVv30FmMBfTTtnOAUlyrma/TchOY52TigsXRu747X+Bu/fNS3RzGKbumkV4gr324E8nBLz5pTbJy
D1PxqVsq1jnCWAHvXqpmON6xvoxS2/UM1U3axLzg9XwPmMYrkAVeOfWQtuU8Z3n09Uan4HWq7WHt
Z5XzDER3i07a5y4BhxLVDpXvQwZnk/p32Xg2z7rwoOdcxF72+LhxbGZ9ZbgBIsdadgn6Jxp+no1Y
SiIiU8Yi5fUsSkxD5WHEu53JDscXzeq/cKluH6/E10PcU5E1Tkz9tFWfUCkX55l5kk6MN4kIES40
8CizQeMf8zZ+KkwbiboNL65YRGAQVNujXr6lmczOL1TGS4YeoSr5da2Dc3VckAnNzQ4mhn2xp4xI
e2otr8DenoV9KUuA5zFgAkTJhH1a1qrz3yCQmHeUilVRvcJWQBM9q7DYVqcIbqaz9CtzlrNECCdL
1g1QUhe0dHj1caXQDIXKey367U4Cb7gFO6H/EWrWnkSlA4aE7fMtEf70MbeDytng3nfZWFAFm9wK
NNPs7HIypK22sWIvx3GaloCJZ7Jqu1M/mSIeV1HkspMLqJNGrPH/SUASOP5cl6otgY3ZX7/B71K4
/VKeLD2mJE7gd9YvPHwCiU2v0E7iHdkgkNVCfM3qK4Kw344++vX80tLB0oQE6C6gXM40wDxT1CUk
3lP0SbFFsE6UUbDHJEGyKyHnC2XKZd6mleRojmVNB+rkBkby+Ins1p6XOJhxzb8qUCJEXmiX7YSn
e6+txvK0WORODLVP8aPBXrcS3TYhhEe1wE1nE6U+VBpVjrFzBUb+YAeOGpxKzdUUFiGPfknp7BVX
S+lK8Uz7FvlOcRg7kiuChb275iN5i/wzt0egNkPl7mJmkHiWGY4wdUejicjtMxHqgV5qCYIhIROr
rHn4fX9iF3zyVigfxXLPLX7nT0DZ149psjPXriQBAjjCJtwGiO70kReDAuXAgltW78DlI1LUjC1X
4xkfutY5a+jWN+I+6Ba1JQpxwVa7OiaTPpbOKW7HbZ6OEHk0NYSWRXNM9PSACc2cvPQPy1XpSLnt
nCS9b6pSxGE1WRMm7l4rRlPjNJkkUgSTo3dHE4Epp4b1Pdlc1tnQP4Svk7X1VjVieyvziNCFl4Ed
eCL+K2AIuNG9ouhPZO2tsZ+DGEMx8yunXNswjaa9qvGUh+n4CTQ70kPhf5QxjyBI6loagJZmQUCu
Ng1bpXuEhYxz6Crqz1bYJg9rYXJAoYxtFJT0o5NIPmFo/p73lILUP7Z397V3DJ8TBrTQLLAKauqj
a0QgB7iQ/Jbr0tXiyTLGQPm5K47QiRkUECg4C8ofnzesnKwhlTLbe4qMcRawQZlgrNt1tYTsoRpp
/9w4VUkKOcn9G13kf1VUXFxnDasqtcldrSeNmEpuy/3YUkcflMq4TXBZ68XqmoREno+LtWyT3frQ
khGOgNxLek3XAPu0NfV0KygWgP+/RqcJ+5Ha46vW4gFoMXnDdVidINyfphXtPLjdinlOHZFfeLTZ
FiKzRxnxb9u+t2MZGzlaTTvzXE1UNJDeY3i7ttbFoTAnbYL30IqKiya3hVZiTN65G/u3QRXA23oG
7OGmMdMm3qQ4uiyk6fdiCzXgs017Ptgq0O2WkZG3zHhRIOopKFyAifxjqxtG8Wgt2at1b1nYAOTo
yceXcDuMxBPsKMTkNmUQ0e9OTZOcZVDaN09lHzG0ySZOnsTkzzRdazcZ6z6A0UTFpdlvTAlQRGXk
PXf930denXbRpY9xqovQg/Q6TX/B69nFVVUL27lHIWT+tBMlXM7JYO/kX1pFoWbOuA3uBWFOm66b
fV2o9V2AtAQ1vIOE4S61pkJax9Iqdocx9cmtvCTHwAubFV7NRPI0qO9D0FQClRioqGnmChqlzbTp
0k4eUo1BvMeIAW6BURaF3UQJhDluTrEsrV5UkZk8QHXlQAJJlX47V3jGwyI9pRoj6AW+YHk/g0Em
/rXYP0Ei2UPmnxVNKhdHl3skbre/JNRwcuDmc/26GweUTGQUfqb1Nm+aoG5D2B6MXvyYK5flqSUl
8QUzCVqcSHomWrDf/cDCW4nybipgHqu9NgTKmFUv8deL5wxThZojBk/QRoT83ftn3ngegRSzFFKj
cyP9bsUzjADF7D1B4v4rCfyH8VpZkymTofcRSqBWDVIbyOBOuDnIWE5T3FRjRYQStgoEO26SAPFh
8+drm2NBxvvATpQo5ycWITDkd4a4LIgXMjCfGd/pZ4lX9/VP8FLI3qOUOp1vEFpKEPanZy21K+FS
JX+2tQS7iQtlkugPjkBtql7kEK9PlbStGjjGjZitu+ospYf8XHNAUk+X9gE7sIqVEu+TgDMiqRqC
HfdTaQFLbbfSZ5g+6YjxdJqv3joCvIzZfnNAQcsp1sgkvlSgfSIZc7FlMkvHkzz74rGtUuEpnlV2
R6kJkv+ms0g42G3/zCOmqQmxE+W7QOn6jaFpgiQMiTqPpwiISNCz0zVk8E2LHYf7KsnphgHIleJS
qBW8/LSSKbaT9SsXgGtcX+q4aaDBwPzciZhawec+EqK+9niJxNSD0ChghBE6DrHPOrzjNChu5x7V
dDFwf9mkuZtNq7figqsgvLKLTmx815bOK183iEZ6yUGhXwvxpfG50JZIhM6YzukHBbkfZzqWEdNY
ioGaUqXRNlHYg5wO+Y1VM8wdbt+KygaYW3gBvWyNmSqyyk2K8tRpFgO3BIjgd+Gtb1ouYSCOfIA0
3MQz+jXqgV9xouaAAq8PqyNPRbTy75hldFOmV/JqJK20VC40u8vPgOmwiDMGzQSisE2yA4Ayntqb
XrYWr/KhOo/0jXJfc9cAhgeL6Y82SHaQCSaWxAtlwDSA8angHQZQ2fWFbjX6cRUubgisLyuyjGBz
ebstliAkZ1vaKGrHDaUraAwQ2Rhey6Kn9WIQMruAD37LEI/6AvsvrWiumFp60ocyr8diVRTTOkus
N1YkZ2pxWWX8jIaBV/v3cq0ZhyZlZ5B6+o3kQ/Mj9NKSTIej3RZPjnvHYn01lgzasGZQ716xpCf0
MJ8/WhKSuZZfZGslGYNZQLS4I1utf9eewhBcF2JT7Ezdl5eai9vYw+OOOCrkKuZkUyH4sTZOg94n
FrQGz3a3isOEvjJHZzYj/CM3t5fcT1tbefGen9aFZAT9Ap70yoTJ88Kg/dnXfoEo/mr1fNOFYNzX
4NFePpuj78dPbLwNFAwmv8rhqxTeGNsoeOH8CHuzxAp3fc/s39t6tMoGW7gsgqc3sMCVQ9DfFtEs
plljvuuR8rTLzqeiv1RCEbHKLkE4oJ0i4Q/XEMz+4NWlJ50R2ngeDuykFaKQ0SSH9zp5GgiA3juW
qEwM7Id9+nml+Xg9SgFwIrlPgmKT90gNOzvaXHg5+2YtK4wybogA+qyZMNwxualk2twEBxlaudal
04H2CSKSTzNLzD/q+1OP6etxPNI4EEnqgP6Ii84WxkZ4SAnoP90H7WkoX5V/SwVtiuSTRw6SFVSx
zvRiBdFROzVavi5b1hvtOdT4+tSBworEFB1Qm/t/l15EgJFdggedT+QsSRXZTwVPhav5G1MbnPAM
78PT0e/n/0+sdxQ1ZSJFPGXDqmLPa5fi0BwaJ4uQgyg/2KCas7Ihw/caox9RYqF7ZRUZNXdYLV+l
myBrZcFBvLI4ROd1qivOV+6rJ8pLcYeS6YCPCaUhX8XAqgq+AQ/vpwJ2NhnbKRo3tMfxJ/IrBrZc
No+hJ5WtSSdqgs3KwS/aDL20hHbp2ML6vgttA0z10klo0sxb5QCor7lbRV7aJylIDo4ElkKisDfK
6Q5ZNa/cbuYunt2hUVaiD5dufkZmd3F7RMEIrKKus6fBqIaUnZxHCfOHDW+/fvlSmtOfLyjI564+
nStXQZfk+GUbb+UjzUJrmAbqkgYWZyoGL+oFNiiZf5Kc9jsQdQPK46fZFtA1dNGLYUbJHaTn4lpe
CLlInD695XH0HM1j2PbSHVYN6Uw+lRd6I1R8cXkLYNjKhVtBGVzv5Z9JDlYbMFGHGI7mmMcanAbb
uol3zG1Oxrz0/5SNY5T1Wu5Ojr525RBaej4wjTJFsv7rZH2xzjooEWvdW8yJFl+8wzQVNpNkDoXm
WNtm+Z3+1fJmxT2/CfVICoO4r1sqxuBykMp/lhOIgzF9BV4B3Q167lHYG3ACfV4138n2LIHfMQRo
Uz6r9jpGLwa2VFebMEDSJ7nyLxbumw8ItscoSbUICc3C6hfyu7RNe/MwlpP9DXvsdilog/koBcW+
5/uzvoHkPBq+fS4PNpWlepci+SxwIJ6q9E18tLeiGgCxGv961FkyIkPLadwImjJfkUpndQNgP/fC
uVgrN66/Qt4j5sAKjBMhYk89v1i7GJm2RtuTKWyEYIeTWwauMv9Rj+rdaWlcBeb06Febh6teHna1
xevtt2hEFXgs+87ywhWz3X1ZnXOsFhPuygiUrfGQz7C4AhOeps1nq6Rs95ZuB9IcU7airDCkLlGP
xsX5GpXDX1L36xw3Y18/cT/87HkSREHV46Odky0Y7oVRZ+DmP9qoVH3byosQP058t1zsiGpOa+/y
nYpEWfwopE0Q2qo0zggdICjwZJmLPtV4La/X2n6jPJvEEUMnLaNi3hQep177mz9tjGJHrQTLA3NE
rhX9+/wXJrOFkFrAfD9WiEx67Eq36+TUQS4m8dEI3XLvRuZ9XdwZDSEckgOgDeRWj24MsWFhcd+6
6BCN9P14oRCb6B7i09XGED2zm2Cqieo5JGrAfr8Sfi6ncSyBH8pB7tVeY6iS+WprGTsuVlX+R3A8
BlgCFvyA272rXH340jM6tNjmY13Yi9ZSUG7ueBSzOdLK44L9lbon0yKwGcTml59hzHEmQMG0xlFC
Y0a3HvqAH1fQWgALvSRkCkfR2FAYOPuwr6G+gXJ87jYCQ4Ax/tXAz6WrYXG2+BSrtyaMdJCcWoJJ
Z/M5ghSDJmH6Z2eXXhklPCyIqiJcMTysnvMvyM6RTfUuOkyztiDJMHaad0AcRtPZ5cIlXdOGRNiC
LIo95z7WE6AQhEOEX/reqk5l758qrfYgNtVryX7R61Rzy5mvGW3uNnc76skCymaDcfTYcm/L+a3u
eMdvDq2P3k0NuHrbBWEHgrvihwz6tIYXKmRM08LkEA+67F/FoyLfUJlvn6+wEgRiR4eRYJxHDLiZ
O295FAu5kqDwrq7PDgFQp35WPXjpDI0r9M+ElzPUADMeCL9+uCy/W9Cr7EUNKsYrj3U/Xb8+kRRO
KgEg38PYFtkX4L5ul0EVnGiySd0Min0M7C1q+Uyw9Z6lbhxbZaqui/7zqUdBgcD1I7UkC/y3GgFh
WCfEzdyU2iwob6+qHuLgOqWuf2zirc9pmmkhh0HYdVngkcOIptimlvOih/Yt/gKEAOOpNaVD8qla
q/N0VB6y3gdeZTv4478riUT2YcMmN7wl9QnziF7Q/HNjQUJSu4mhwF84BCn1+OX/wVDK8zyp1Ci7
McxlcNShlyQnj6W5OgzQqIqwUxIM+ue9V4BT/EnegBIvIU5q7wLKIr4N4H59XL+xgoU9oUenmeeW
cU1irSb6j6w6UEcBUl1WK+5GZwMIt/ofM82u1u/ozhIFEB2U4efvDVo0H9eTujuaD3JhrXuy2hgV
lBzT/Gor7Ra+WYM7gPTOawoGNMB4ZomefIy20H4HhkmmO91LOXlzTLdyV3oSH7160o00U6wvGau5
O1xrmecYDS0MAimCCuGDYJVwN/A1xtVuXtKruhmucNDdrQNUpTdmsUQ6MvGi4bJ3hjyOetj3MGIa
SrkxsUeFbYFJKhmyHYLNsZsSiygnZ1mU/axS9CwqgXCluZim1U6T6lAIfPEat7z9I8sPv3wT46Xt
HXyhBYJWhfKYcBLomepwF4LW4fXJ7FGln1arBhrN0anE3cwC7C8x/+lwK8vFBJnoTStQ9agU2jhC
ZYJLTEsseIqJ+1cYkdEEHpfK3YW8Lz3qYIVd1smj5jfYKdNpcolWoplU1V+BDyKgQoKxRe2y/NtH
LFxsmWGQeHmuJw6vyIZ2NrER+eirD2muoC9VGt159ANQhZO5BewvCN8/AD9nyhgnA+hsHX3VZvzu
LBb2onif7ntLl03Z85ZMUbHgItPi8Skr8JT3nl6T1k7Yk6ML/uTGHK8Jtccxeh/F2W5M+EmedT/L
5MSaam2gUX0Nyleun0XG2xM4FNKRIx/YYJwEfhaqFlr5i10cDLUzrmYryNKASGbxXDeKVlxn4KIm
Rsw0Mya0wOCUxiviqNzIjtG7OcFA/I3Vzgptwiie6dcrRQ9sD786RWajBdjeBgOOsjTdc8LZ5LKu
U29aF5eqHDYBMEJ7FiuH5AGGojUr45Yuyo1Yi8c5URQV+mP8KsKi1cBXUay5iYiP6uU1zp0ETvhE
RMwKIakfC8G2peeHcygclqzwqtLAcQUqe8NU7CpKBnbqMNGMifCi9UaGtxKhpX5bm9BJ2Ct3aWId
yuC4xIliF1RUZ/JVnCHmfw+ZMCb4mgKOjW5XEwB2zDA+OXk6qEPTNVqjpMYY7wqQDifiUTpZL39u
jt27g52A94MepHQt4kNW/U6aVhhg4ljWdFFm9i7RJb6QPnnJfx44aWnwUtROGeFmd8yqx1FeLiXJ
qKP1JM8SczuovKZxsT0/2cJpKJNnQxSZA608E+i95OTYhYDXV9f6NyXOyiBFazwnt9X8EEy4mY7p
XuSMriLanv1ZZRIGOqV3hn8C7xQ0wd0J10kzhKXPNtCnR6QUTP6Ou6ojPc9tamoNohKVoJxejlHs
BEC/kFMMl2GrW6wMofGYTjT9b5KFxtEf1NBxVtHn5GMdUKxvo3Yozw8tcWc6GczZRwTsTCVx/99H
hc0/89EYkDTMUgHtWZLBLLzFWhAsgCNsyfovt79MOlLZoGcqrmaEer50XqU2HxxgRyWNUGG2I+tH
vMj89XjEjTPybkGbzWK2i3rcLa71ncPK4dfTHCKUrq1kuZZkWQMq611uPtiyTrUPYMPTrMLqo4YT
5sgHgn9bwApeFJsKdqGj8e6AskOfAQyYyZzl1IuS2R9HnHKPYNxQon+rXVq4U9rWMXIiYDPBeT6e
aOBTrdK0HXDejil85twZZqX7cx7DJjmGzs4kqd1rKmm0MV0VUffFsuilOkjkv2DaWXgHAcj8IBfu
NAFY31mx1pPW2ccFWrCo5QCs9a7jAisXnyCuLQhoO1S318uUmhThVUYyPpS/B5piyPjjqOUkawy+
XJm8DuaFKGzH+b86EUg4CUC7KVdM29laBlsqe2mHN56l6eDIBxnhcq/2YSC6pMmBzBmov30Fg04e
HqMugPYN6h+K8zmYu7jhuBo+VX4vntoXcuv9Isgbp3UIT80bfuI6GbVOHnYByr64kttq8xGkZAog
bh6rTSQbTDOPzUz8qK0PuFb8xuEM4o7YHUN2AJ2YW1ACawhTIy8z/LZl9YJ3lCakBPrHOvGdoe/h
vvJ2GhHFhQz0GXWP5TQFiSH0mwm8vO0MDyBx09T4i3enhPHg9/BW/k1OUmHSuJNaj7Gs2a6bqtTq
WclP+qDcnS3RJ/qRe1XewKjesVGvQhmyOhmA+yzgasLELkSqrvnOPqkMZKezv1aDAULZGwONFmJr
CyAmO9OTuwevRBUfwKxYiDlz66qpz/f/nxSG+Px8gkWa1BgF54R1fEWsD5z+KiM74L2pov3+Gco5
K0rBGwXSKL33oE0Ut6nnhH0MkJtJxCWBLV1Ca6h9bEgJIZWII4fHxxQMYtNOFoSF4YHd5vvtG8BB
mj4ghJ/gAf0UOccDVEkmuBUqvMZkUXIxawQErNTcElvrd1bveczxpfdhicZwejSLtKwv+jQCv1kT
+i6+v0mv576dJfVNdzzkklOtGykpvZJC9VYpkdONittFarQfNdELajZoM9t1ISKz2bqveOtdfk5g
m2EMEBAQRNkQfHFSAzFlwSVsJfadPWiX288N1TryPoN0ZXn4M12RCL8lY3Fr5GX7UJ59azi7GF+a
WdNkV8eFuz2C4343+78yc+0m9qRd7ahtpTBoU3FFDLR3T7NFtCn2Ne+JHJfhP6SH7R0qXwKhFhWT
xEbmEOSUfX46h+ezhwoQHeCemgJG+gl9xeR9zQFg2e7ZHvbW5wrcZL72IbErkIphyHZEqRJg/IGl
Q9YoHEfWEEO08TiMps/RuSHxUd/guNH+7qEynqbOphbcIpWfCSuU5nWEJYgBO6hOJt8aBBICgA11
libEO+Ws8MrOoQhX8y3jXwmEco050b/9h/bJObjtzDyZ+QoQXq3pJ1fbZ39YItalPvBLeCmA0dTc
vL6gUWCy3iYTj5z4VzBI1JA36KOtkgVIKw3HM65liHOBueT9FDwZTbgEPR2Xl6sbxXbivBZU0KgK
rLe/S+zoWWDee9hmHEE4pl+gyzg81/MXJgCsuJL17OAg8Z32eacdrRHfaXPevhtRBuBSjZ3oEoAt
wNSI+NPfkyF18dQZ3IQS5r1c6XPaJGR52h21qrWQfpDq8xyGZBQF4eAQg7s/OYcUh35sEL+ZH07U
RrdWiGMVNadQpTSDOYVt55k9e37XW3zuTzdpt/KL1VgkvG06OwK6NN0s13YIWJZJzZgJwwLWAZQ3
MaC3ovVdZZWyg6xN/7ddEi8YSoUzqBBhj7m5+o5zKZAZ56kUaobhvJ5pyAVKSStNkCwijflcDjRH
dIy9pG50bHLarTkTaqjbeAW96o6w38CsearxcD8K7Um2DaCKbmedozSeZBifVv2AnFvJJdZU+Xfg
Sa/h9qoqckZngS3yAZAGOytahRoGTcrrVRxKipdiSqA5ZA/OkmSl6edrm8OqaDypi0gaUWaubmyX
lxqPeAAdI2bl8EupyaguCVNY54Tu3Hgq74kwFC9C9EmaiwtT2hyWjBZLNNDjjubs4F0qaoypFN8k
2Lxx/JXjZye9MNA/p7T06ZC3k28oQpSznCQxOCS1R7eZanOz4bIJdsbonF09sdNTY6Tu2MK/qSEK
pAQD0X1qULwy7tyFUkzrxuGdoDllFri/e712VUF7Rg1itUgD/DU2/0RG7xd9c1I57v8f6O0X5IXd
impEQG50uH0fQ5ghHulms9ICxGINd372MJaDABuVi3RHVXwkM/MGkwh5IfShfnxP98yzq2Qw9YUW
iRx0DeixxvyDMSNAcoNL3hTfwrqMXfVlAun2hGF5fao8qFG4M9ykKwi3BIA6wUwjh8YCsBW/ExCm
GLuFwTxk0BGTwYcg2ADRQlomfOflqaPAxjFdiD71AiUmCHFXCcGygzlEYHeM7NpKJ1XUzq+pM+H/
BRUUFJqrLJhDFA/jYcofv5cu5kDn6IB+qi/GFEmLX/cnl7blD4/8CaL79VDFsEpGhYZXFbehlMp6
woHUtQu5xGa+9MUmn1XYUVHZxwFZKTu6Y1fsGn6ov/MkZrDyJ/q63EMMKzPe76/uqA9D767h7lI4
nKqL2aWkRWIFY/qfEOTxWlEipj9LOF6CsqjcSyx7p2s5Oh4xfP1AE74OvEZjuEhP/Pz05Kqbb190
bD4F9/ZDcEEBVfPuE6UE1I2L8TPX0pApCSt1HAUQasBPh55SFyQAjA8NJnF5RtzqtKidvLOh2Kcm
ov1qQlXjjeEpzSyU3EGvxS5OhgLOWbTxyKTzz9O9HHinGkLc6mvABgl0utbzzRFbSuP1ueRbM+iJ
YJOGQlDh2WHaRc3kO/WRGczdsl1J8Q+9tB3P0jqIUbJWSzzpHsDcc60uN9474znj7vGdaP+ZVCOg
FjebNfIJAKWCO69JDMxFBmkJ2NUS1G2SLG9c3h6USzsEpkCQCsulF1fhV/AOPiSL5nS02rsk5QZq
CPTi6xSu5Zc73c1nnICXBVa5iWYTAtaqLlzK020rpxGKxYOFUPbBjDU92QJp3pi9oYI/bTDDbiTk
wfsZoiInZhd7Qw/0El2NrMVHlYLYWolh68uEuBrLKkZxtb6SvPXt53tq5292hA/b5VIAX08xANhs
w0fkajF5Oar0eBD4wgFhdsXdzMpukfSef6lQHtYljWbJVqNMD3bm0bNN3G47TcQS0jM0nxdkXkst
Kc5Th5WGq4ur5nr7EgrwTIQixjXQBEsXK0/xk2iaHP1e7w4YeIFfhncnHUEW9LtjHFnOnVuFveNL
hy4snglBx0yyKbISr/n4LUkPrTjNstYyAt+4in3CcfOpkfkFX/egtlEzaePy9rQdpf3k8D+rySeJ
HHwcag6dC1ISdJ0UgCiXGCxJT3iZHZKXp73UO+IbyEY66kTCVWLO8SiA7EBXiFaIq8JG/+6gO9s8
AtFIRji1td/CyBezjsGZE7vG3MYZjToJptafhDFLoN6fcXSD/HJIygAlYs7wGliMEbjVvAxK2aQk
f6vxQQ+d0ovt6iFaDIA2f6/e+bmfjZM/dYxogq6vgE0nd5EXR0PgUjdW/c9XpzwZBkqlnChm/Smm
66VLCis80vYUrZHZQmJDI3hmN10Y1KzMfwsSQSbEzv3Yx4PIHUuDYD/qEvbLZpx6qY6o8htLpuHi
K8SnN53fiSYSyn//fOLeJiULFHd/KKN1B77DhmkuqnVcnwq/X+B66E3578J31FmEYuW4FaiH22Tj
1UN3gPvnVKFG7920k/VNcewUIHGEFYmTDbiadhuviSScLStbSfmQrzXlIBDTDKbo+5bUwojpA/Ps
15ucmsT7jKdoucOxW7U5ONi4N0KUmcLeoJXMqXPkaLT5+jsoSOpX/0LQHDvkxFkkz8/8N8mEPTMs
yGmey04K8SqIVZ8vPo7WZjSrb6/dcP0F1tgqXp/XqfZ/v5EZ2TA+b2msmB+rbbRkNj0m9V+/zrle
5Ggf222bhJgYBNlGSizUtfYek0y9uHdELI1Aa9cpfUczyRPtsdL6FsCIz8TAUzY0n+iXnBiKiPkT
Brc1Fg0RrWYhvC1xvP49a9dQr2Km350Dwu7uvz+Il/r18PJ5XP/GU2leDfAL68YgWBMCMYTWJ3Xb
sWuCW6zYEDg/4u/w1tu1t6nUGFyNdnNYw/jqNQ7bcRMKrRbsbPlIOa+Nu05vFyIBQsQh9FwpqS+1
7LBwNocUPARoWA+ZgZqK6KQp/EJAoq4k2Otd5pwDCG4hfKrSYys0ivVKT7EcAP3L6RxbOkFfvfbp
1lYtuOYHX57nMrTAanJLsjnNqXCsHtsJhEP/JAuRc6Qo/l6tKOw2Y4KSIh9pOapqyybFd28HgEm6
BANCgLtsD9KoXKJwVxifWIIZ2uAfSzufKWMLaiMXJGW+fRlzx3YaCHZP2bLtp5HZa0nQq/diSIPI
AlCqytToj9kyjq6YO7gMjnlQBeX/n2QtUusVJoz8R1cdGUFc32j1ds+UmRn2NSB83VeY89joCNmp
7QY3mcWaWkDYM9IaK1CBLz6iXXWbJgWuMfyi2iLC9nZ2LiPKkXtWjkcRvPZU5Lo69Jq1fnIGxcZr
ipRrhmihLVs6qFVo+KRmDwe3ZLnSsEdUh+7/w25s7nD7kkpDCbDE0+x8QMjQ57QzCcEsjZjqy8nm
VuVJhnZILdzF/V+NxLtp3KnA2Pir4rj5tqIn+lReONCu4ow0Qnvb07VaCyDWFH7acivgxfMzuibd
1dUAJolr1ggy2qhD77ywBHMwhAag2GLIYu40NFuIXTCJ4O2S+RnTUtPOutpmJ70HeG2ljbf16Pei
3pmJx/nYrZfT1SpFpMgMwYPe3+Mv3vAggxvwmXx+FijkjKfBW/Bi3xCaqXvuioq4et+aawqVspIg
PTC2agsPafiZjeGmHcNpMVitvVdeyQg+2PxcZo5OJq0Adtf0nwWlCfnGqjF5fepVH7OhXA0q/d2K
DpA9eoXLH9LM7sCIGlTsMhG4RcVhPaGHBBTUtOJNjzF5gESbaQwHsPf+bTFw70T+vbW6Fd4F4LrK
2o6b4MPyHHsbtbikQjYUn/tbI4uUI1lIjYt4LZW+0I3ELcO80ACya4OpG0N16m0FqIAo6H+Akmzb
zLhN38pTAdLk5QKp81pJKDjguf4L7m4HuAhmBIqugCz+lab5QE70/0MV7dx3JeTNqf/ozYM4BP4E
bFKG5a5s5qBaAAihNn8/R32SFyqw+98WDMPBjAjJ3J1XTfdE4QpB9n/24ZA27pPeeevVagUDqfsL
dmBf5oQrH+DmbQfZfb7o+j9VcaNwxJWFhglcyGvjsDNrwhn+YHFk1CHBziME6FQ191GN4IUkmy++
iJNAOhOd6QQZsnAu3y7e5LunaI0N6GriaV/tr+8Aehg+5q/TCY9BV0IpxdfqRgPquCeml30ctkTu
eEqfKIBv5p9Pk607zQQEvEOyqkkaafdCifL0LDdjXkacoU3ZouIDl6fSEH6SxrLKnmSX4iCDRcFa
p2PCvFIFFbaEm7QBBAX07H2czo/kxonmuOjTclm/KMt2jtFpw/Bs2QNBepaphjbpcVhxxJ93sgVW
rULRwDWMbOnEQX7qU2rvlqupUXWh7S9rKGJcwtbSOZpwA7P1nG91pJ6ipWeDQsJ0+mwNYqbH21DY
9aOX2Ad3jXnsC/AviPpxqfsL/jxjYOFeQuOj/sC+wQG/cs3h9YdsBLlFX0Q9Nge1T6fmPp/0uZEK
wD2TU1fuUR4zVQKil0xudJ6AdjMcSbHoS7ReACqjjRsniEEVo7iLe3Yt78yj6B+Ass+yj+flUtVK
g5RLB9KmM80zYqskF0RnmvpsPaxkQ8gssSpl9BOV473P3BmRybCmGv6AgF28MEoytVU/oY4yoKw3
SIMx+y+OaOd5UpjapLKMjYmWXP805ChBgCate1/6qQ31hycaa87YsK2z/2AK9rYV6NVRnKtwdpCG
3hwQKKljlANrTVgSYgXtv/uCqSbmr5Mil+JdObaxXmtAzagMMynuSrS/fkJ+tlBa3U3Eg2lpY+Z2
HSWOU4K8R/bfP8lgBL8CIImHCJPQarfn8Rj4nAvSlrcyOhxPBozT1Cv75q21kp/Yyd9bVJa0ClF2
oj5pBaaAt8wxQ0ynFHGD4KxsA0xe4RDV5Fo5JUSbJ8nB71Yl3s+RuYVpbwvH5pM1boTKSogiRXze
nCY9Vmuy1rIRBnAgi5bcaNGAwlXp25NrM9wxx17GyU/WSU8P9OQa82OzQZAleVN7qtk4Ad+CTbby
mP6IDcoOPY5P/YozweaNvsZ8VZSJGBvpo8dWrBhzjHFBhB9UkkHI/M9scKK0iD6EOV/kKpufG652
avbtsFlDJGiZzDxDXePKITAwpsAeIqTFpAHKF5uErXvoZMyNH2XMFuRAkAOcFm/wW2/UT6tN14Zv
qcPihfQjn02dYYZwQNlMbui1NnD9Fn424mAKCcXs2/9FjqZCz8O3t75sYfuIBhuE2mo/vRMd+kFg
GuWHwcAG9ZBcBJ+AMBj3uVeZ+MRuc0fLMgXsyJohQ7S8JCn9AGBxxqnnauQtP09bGw2Y+qe8W2CS
8D8V4LjZ3DC1xz2IGnCQZEzPd4RlJjoaEN/P9M7UD56ysQd0KxrPnWZARrfoGtBMFpMB/P5KWOOX
2FLYE2SlHTUPlCDRitgzJOz2k3k+7EIcgCEgomI0qdDjg5KxTCL8WawVxqNNqcwtDhsoJ6lhcZtQ
e717v+mekCCMR0I/Lo5QwGjJavihsES7pGPjopRle5J9TuTXHW+jOVqHnQCpgGO4zWIUjyFqimr3
CtSmyPmjThLyX68Dlit8cY4OBiFkBT9nCTEJ79IxfRlT8h3McoOp+jBUz9a/wF5NNrxcK17jbKY3
G+rZ2K83dgC5LUNoY82zGkFMxDDiIURsMvIM0PuZjuckDVUeELo1L/mG7Qy67aPovYv5WvxznyK+
l1CFddsCHdbzKL5RR/vGqoichWRevc30BcInnLS3i/RlUit2bciTNwZpbdDzUxQmxduftsjyu3N5
h3IABD43pOvsE8ejEBXGE37/plu5QF0hJf+ezhrF8E26u2vVDGMOEi9ER3oMXOYL43S9Csm+dHeP
Bd0WUDbRRntXfyIJunqp4M/EtC5Iw9OX6XiMhMgHSWTMeFANgVkvgxJRba+h6lyqwJXBUo0A4xU8
j2n5IsGmDRkTIJNMjtwfMB9e+EWFr2N7RNV/Md0s8si293qrCIKzJyNOp6io9E7K2FNsKQskItKt
sB4p6pI19PA5L82v34ObnSIejFm8kf1b8E1sv3VTe+vxhhpDEHoIq3ongeOFJ/CQhpLXe2oI8WAu
s9l5j6H3HBxZoEPJUIJgqCKRtQD/CNL91QsQLe9AGTObKdJVDG50AFpE99mbYIKT+JuZmMQNUgf0
wXKVxTNO2fZJ9wMpJTAaz6nVMtvQTXYYcJ0EkGPa9f4m++web3pwubC/LsYLMIrsaqnOe+iCwQag
y6oKIuGgGykrOsF2udfn9yGOEqk9fqg1OK/gIWu2sRTzsj3XuL7fc2aRPe1wLhN52tKMODic4fxU
RBKcEbQWXNJyWh7m9MvNMn8l0cvoXfuoKb6Mj1FKEhY7FOMMLz81fkd69rHGIfQHaMNtoQuxeiVG
DfFO7c9RJvGco1LndM4fG/paylPySjak+5UV8TrGvUX8NPMWidswQvrvsaazxPrwdtC8FrGIEIQG
4u1gLW5km2aYDb5WY2l2a4miLBN9hnY0WEX/B7+bKO1GHooyjHLlgHKvrqZmHmVN8ZZyZU4LHGaY
CdFhK8J2PjdtCy6prry4vt0zq1sSM60zlRL9O0sAYrce0SSQmXr+jEEbpOEJo6DWSxBIGu3S5RiD
FtE1nYRg+naGbp0+AP1ctKavQXS+iDYMyx4yeu7tLwJkmnQazp3xaG1ZD8w25Xt2/1ORVUDsk1Vd
wFRo6LqWuuzpy44Eb2/GKu3vGUQaOP0QUVKTC59C9Ixm8zP/Sf4yZnrxO39UXJ+Mlaytig0JlD8S
7j3ZivdtMkmOnyhpD6IrzoN40ZPe/RZuy/NxyxJSJQG3saNu5ZFQNpdfOK/kxGxU7MsnhFIuYlj6
+33KaAK7a33WXPVqTvL8oiwuHmkNUdIY8DMB4DcRXf10Js0bc3vKPSpepxCINL9P2t0PBd28yZt4
k1yTuYmSAeMd4PiVwsMLsNlJeBEqZy/FyBBh4FG5wL2z/U6bla6qXOus7eh+e9NpRCNtoA6czGOC
WYsv3a9YYsVQm+z9uycShbzVs/qg+x6u5PiFNg4fNmJTSb8/PDXwR1jKl8ZFES8PiSKI7zpI7IaP
6EhH6lvp3ywfrouTxfoUcUyqTlEjH7++ksXwnJ84TqT3P6fYS3cjUW8GPwfMR4avksCwbGKvWyP8
cI6hebHQoKptLvDnXHws4ESKbuOD35YeGy0yO26/fwwMuGwnYLKPxODvgBBxR4VW2sg8X+e9NNKl
cuPUODXwmjUdcES22SDXX8q8LAMS+W68yCDqn2vrUititqkScpnOhcjLZnBnOUSXQbBNr/UhGRlG
elHZRaqtCE4C1M8AQyJVljqZ9rhd0ThPkSThaWrqCM7IBNKx7PQJ0ApGv4ke+ROJZkIm/V9Q7Iyr
Hs9LbV1wg2a8F5NJhFpFVoLf1sOWWt2Rj9l+miR4C0y5IlVseDBo+ZJ+0/HQrzsU3QaoNip7pzLd
qChNmYPkE1D7M7d9q2gbTvYbNmFcrM2PhBprIZCPihJaSyu3OI3irswvDeKsfFP4t5SWnfeQRtI9
twxRLOUVdQFAW4fjC29DbdCkP8d1OEBiBxv6RpQVHCJPlr7jFEbfDzIB52eyWO5Kd7zU6kHWPnzx
GRnf0zaq/mqC2YHlRaFdiu9INCu4Nicwjo6wLOfvndzKo1JG2JAfSbahtKwAZ8Y8n12gtiwOiqr2
xzAmEtFwJW/bhAMDe64GJKyjcXTdV29bYRpXdC2NFqxOw2n3JwwqVDHdYGwcpZ2/r9WJRfspiPTm
iMHrL/ug9y7hF9V4xgzckMEIrmn4Ez2l8nl3Ou+2pxXfG5XbjaVz0Y0IJhebJePk4KrTxk88uYIO
SeGjBtWqfP8D5MOUk5m3mAobskynYmrhx92wGxm3+VH9EhL34UEQQbrCGSEXOkQ7aIJ+9TcjRHaK
9t5SCLoeoHGp1EPe9QgnMIun2og+AOjAV3iOZdiuXagTFttxCSDCE4sLhyngchcBrkdqWhMTYpW0
rKQp6MBuvcIqCuXO1iwh8V+xD94Dsa2oWSlwgQpS90HyIGvLbHXM4E07hJeVIli/ChlTvm/Z/mH9
UsWGoWtrpcUr/Us+eNOMFXu3CZHY3/PnSymiRn/b6vGNYgCOPg3CdBlkPF3Y6rDduBx7vYGJTAJE
cA+L/jPFDbTuEikoE172G7L8pWQEzn7Qg5Sh+rGNrsFGjNxwBIV1PSBDcY30vvyTctzdcBb5wKfM
QN8aHZshqE5a/JMwHz088rOHepfaFth25rZNaZAGxils3a3FfzKJ/NqiqPSsUPvPLmHlVojQwTz3
D5UCNOECuDYzbToaNaAb8C/bOWYiy+w2ppdn0Rucg35EExTU67uik2G1mEsZy3szFos/ORl+Fmev
/xPWrSQolkOVoyoEDBxLh7vO03gJb/DOrAYLBewES34wpSWP0ztfFb35BiGTuge/5UJZ9bIqos/3
sHRqWkMsxlWqE0in8chygOIL9hGxjgqZQ7sS3H0jG5Gj1AgG4ggi9B40YDXiqVJdRZF/pUk6CjKn
ltUwtA1KD5McrL8hKUzc93nv8hly+rVqv5ZoQSIs/l44TfQ287xtV1m9iJX6AOktuFEsAxKmB9n6
xP9AJ2+4T8nA1Af/RjDY1XOUJW4f8jqUuRKLCQBVrtMMsfxY+Lb8CvqokWq2AIpZT2gQKQIMV3PP
iDwqqQ3hKHx6KvZbrM2ZOvZp/Gw4Y+rwthF5GrgHjheRVF49yOd7GQ70eRXbWOfl8ZZj5NR/xFqX
COWkQArJ97qtB/6iCEgvhV9rhQsJvkbv/DBG0zPfiOBkxHoR7hUcT7yI82fM4qZ4V+rs1Fn2Wff7
0ADSjpmriiSUXQwWLM+nByxA58sAwZsfTLNaMqHaiv0wEffMjDHVOJ7aDWUFp+ueJL0jAwfqxqct
/xvrwM+nmF9rtYlp4EuvAJF7gTpACAKNZBgiDog8FjmKwoC9Qux9QwQaAGInmf1VvbLxY8qoCNa7
nONMgf6RCUxar253XIOw7tt0hVtjGDSzrRjz1ipFT6oONKTxtetTQ2h/fW3/Xgtm8/cFeabuJLKN
rCIpmwbFszf9wa16CPEbt0HReJJmwsY9J34bUbMS/z8aFv/7CVYeJgIXHcfjwerq+3ZrpQ36Cugt
SWSaUevIWP0HEtclLf4QvEvNZIbabHo1N5TyEgqHXwoM0M5b3XS5INf28GEglLhEkS2ba3Z1tuVn
C2sjgXhEcvkh59j4xx8B598KLcZq2IMAP8pEjPcUo2bajz/o0fjBzCOMnIjorhctzjqbv8Rf+NZn
B4CNuu/0IPGiIRKfGaZhaYdZ/aCTBLQMFSVkr9sdCLIkESSjSIetbxWCo2zUphz9/jTfozN9DmVw
C8mVD2+fTH1dzCaiuUEgSgqPBoJ/4mmZURfw/RY75PsTMNvjkQI51rPJxH7/uhPbZ1x8PSlwfjrQ
U20tfqaLXm9A5TeacbbLC3y88XDLRxY2SeWW13WoMDV+XhJb2rf+phLvWByFatYlopVkk5aTxZns
Sxq+LNFQbUX1XMO0hNOJOh0cwNsd333No+1haghB68fXBcr5oY2erEumeGgLjpcketyB+bgHxcKN
LWdQG4cZiTIQeJ/hVJF+7Gb5qcmrml5aQILWN5QzN0cEWgkB8F69q0Zc3HmCOpDCP2Y5n+NR8gXN
PtdOQ/c9AqGLShzGzP/a9BZnuaFHRZPzWdr9P55Yc2j1AubF1fUMZuydOPtZb3jnwUfDTrBojoi6
DO4C8eo4+CQxF4JhhP4sYT0nDFLQG/LNV7egt7Rj3czQntGsY5ZD5CA8bWrKCEZfwTaVEfQ96zIQ
4dusqBVGlkR+5xEYLgaFdCJ0AzAs1s4J/qmI3CpMj6dM/G20NHOsdE2S4p/YIUGqgjchprRzDOPV
5vVYARTmte28BsLTKDcHUep1BGqIbfuvtE7BBxKlMtIaqqn1Kf1Vnqda5HLTznJw9NcA6c+q4Nr7
BhzNM33onUqpQFE6H069W3kmpuau0wcVwqnRlPq3J3hagpiDZcZkKqx+h7XgDsT6em1es3J944GN
VvejZzU57fVrMBDWrlChQ15W4aR2AlDePXln00mA/f2WbLGxuBh9vdQ0XHSTlIxmVjgsri9HMA+y
mAKR5zSydGxVYf1iMytHO30v0pBwLJaUxgIv5vah3otHH9xPSMv9PoslHEbnnt5xTlzH71bWMZ8F
mc+dHZc8jwEZajr2/I0hPaytDoxe7n/JmUSSE8QM5wotbjiLfHNwTdfeTmhZkhiVuFLU/MUz6B2U
2cqlzCuuqQIJro6JgtEYldCFRSCQ2ecuNklDf0QYQljNxFaoxtdOcmVJ9ijLHGr1xDh6FHNsvSBc
tC+0CiMPdrk+GPBy+sjVOtWdHnrUMd9B9oHJ42IRILOmuadVCuQuXUtNZiCP2tXh0rqal31UOhGH
rrV48x33ZB0IcmEaPJSmFA7Wo2A48LWtC7w5pOWB03uRdVZe//YiaA2bQMTi3m2m7qUoo8FzMhK7
laDLvPx5+yDEke5yw25sFgD2T3Qm81SGmzWgbu/PxvchcEuPs/9c3jviOfEMy1PV13gq0MDRh2Tg
QEfFyj1tjcfctHtBm2IIBq0ocaytNHjeVun1UJW7JYe9swpOktOLaK46vDpanGQco5IDG730GOxQ
aZSk05d6N4/LL74VVtZdUQkU467pZYmFAgdEjt6a8kzDD+a85vf+DfZx8b6+/KLg2jThFjNikyfI
S+dyJRyaPJxw4qwcSWLmglye9Cf+Cr4bnCNHnM1xgH+HBJJ48S7kOrWAlQYP8zryFaalHqvI9Y0c
M5+PrxSrD16OmyDmIkb1NsLp2iFTc6+qo0IPXf1WmXSjG9Xu5zkP9MiJYOb8CGjHgfdRsk0UWpvD
/IIQQW8DP8PEomM2FkWvZmzwGFqccCh40iwtBJiM+Ik5x9XVPdFUcC4AShFHqgq7yfPkH/3ybzxa
4XFKE2j+kjZS4MNkc6S4ovRvA8IMWG9uNwUQmRSwmRArAsahOfKDrosBtOo9Gar/PPuCbjx4rj7M
XAW+UpbiP4P1dH0yop+8HZ9DQ/NLWmMoMWIjLGKbtf9igUnWDCnRVFS9yGtZeX+6AmDfY9zzpurc
x0MPl5ndp9uiDAjPPXyBt8y4qdbcw2ypt3yYhm1zKx8nSFKf0+ntTGDEfAXgLX1CIt1KqJGqjeCy
Z1bG1ZXIJFlYhU3O6HPSMEhIHiiZqW/6VrkKfpCnGCPEBzCiFzB/SB4JkXMQyBdrmgcKsanORfQN
dZ9OeWm+HTKu/1FiSlV2oSmUVgkJM3HvIuq1QXVeTzACKgI7aAqWtLlYMMqehW80ssEzU3idR1CL
avqkwL3vGqrMDyO63fr1xI8w8SXRtGNwogzuXurRjhd88gQr+I6PYr2tGWfSfn3ldHAfzxb74k2V
1og9H99MbkutdkA6qLBxzcC9jhK7YtzeZ4QNlFBV+ANhCuWdklJQT7Sc9U5dPnno3fqFg8HvkrG9
gnDt5K91o4rCJ1N0oGSnJm7UVvqp65AjvGS1E2ODLesZyOsP0/P7j7ZEa6eE77wqb9TQY6X+xQ77
Yeos/qP3HP8KLjsWIFeHk/UAz2hSjAxV6Ht3N8oY/2ayWmFNCP2hRMRQhZ5HRPxESUuyOQ4gLupQ
12v0SmA51zGufTJbHw+O3DwrEt/6mxHwS0EshG4uBPZWNieD7fO03tAirkyAt+s1D+Cu49qUxaZ/
ApZrx3RW3FrbFNBokmwGojY0w3RHbTSoQoE0IGFcaZim53eOQosDm+mgtapxs58w0qbBtcp6h6q6
3QFTm/+ic70a8yGqc8miuuUP00gJVEUmaJtKPEAPY7b9WyBlxNrgFNDQXi5nvno/pM1MsYqmVLE2
FPI+YtH4cLfjdS4W9k/2a1jpace4Bik0/dJgODuwGuQsY+CHvyxVCqg3Ih8qNiLp1YVYEVdbN/Ce
NcgHXsAjQ5A8+1xIxiZgMmovUUPGxImOLV+qOG3LQral6i95ew7ogvsT1TZ/fKJR0I4IBNVhuRYV
OQT4hAcVokeHirn/azwpCkH8eQMqZe7dawfCEcp5NvtdiqySc4C9NdhqBhnQBQPA42ltuRdenRGG
MOimtasX8zs+02jriD67+YkEKuSxOVs0VAkccQtVBlNPcGsihTLY9zWOJxnZOcRuB8U3mVvbMwtw
HNYtx0ZNo8z4+MCkBAT90iWL6L596Nu95G+9ugO93CRxwVMJ4fHghA8GvR/OOuv+nrNpr0qds5DQ
AoVJSGZe7WeALzRqmZkdI5Q/GH0RGqBXsHKiBxd9OPV3lGVBO9QZUAr4EVBJQkvNwU1qLNTYbpzv
1xn00EcrbJrukoPQq/D6uInktPT+iefUfjL7oGZUHgpMbs3mJspM/I8Fgp5ElTnFnfSBXhdUciIX
cEzavEX3bzH0IRPpyQq+OyfyPVDoka6TjLovDnhGq5+iPiPIWGtcXiO5LlLA62oggniC7qzi7jmO
CdDZgKI38nm4AE0GHu8T2AS/rGZCYO7nBcC7vFB3XTSpU348/QLSGp+MAE/pzSWrH4a1UBUDj6Rr
TM8/u4757bfdCxhk0I57sE4QdhuaOhbgId1irpP0YCjPEey6uRV3JXlg40S32fC0qoMbSvcipRaE
th3RWVBwHZv47BI/TbNBtFhf+Dz/znc88B2jrwa+lhPmkO3HaTLucp2ROa2GIQ3kdhIDYqWY8afZ
os6JDYte7OiGM3bZL2nIeuB1sOwSirBgrk3k10OCoJ7YjBVZOEEy+kx1pdF3wVTUAed72YvzO+P1
vAtpJsi1rdxQyRb6eyBxDoeSZXsy4SyT0weFslZh55GDbMZdQgWZaUM+kRjuLxEvcN8lGXbRFFwF
ROaJ7kUnOcybsqCkqxSkk+xcgzqj5Nf+dTGiiC1a1X4l7rTWFTb1GdyQ8N+y02C5ujOVAJZ5Rucg
mEcOjA1MC3nzn9ilcrBkxgAxO5k4k6extAMGOIwkhTPqOgs+c/bIpQpFi8H1VHfmyKPmHUprBoMv
eR0YeqFNo4HnR4bfIRsq4O6Mu9coUvVxjDgeVK6KLo0urtMRcQpRyt1VsBdhQWs6126UHEdcTcEO
hzuKONMTowDBxtARRfsDZ2Hq7AiyWvh1DR2f3ZltzxtEyHKr773ruQolNIR5xenKFl+KFHcLb3bw
qCAyCrOcubmkwlR1Ueh/Sama9OdTC0YMOTpMRsQR7uZ5rjHjkXq+VOTCMnyre3dq6txeC+kgF05q
6/2LFmcCAfWuY/f0r6WAvjOXvDki/exMaHsE2+6/3/vU+t/aHRRn8GWsIkRMLmvR82nawY8nhfaQ
EQsiIfIkKiZlK2GHPBK5WHgG42P0UFvVCzED4rulmd+U4Y8BfscaKgEjOlDi5lopJ84z2ZrhKKNr
3p+GAZ2pFt7m/zdcEoDGGsu0VWN9DdejSlwXeaVAMYbDNJgHq818J3/AfDoGUzoo0zuj58EIIzf/
gPdsrCGPd1IHtTnDk1UOLmS/CLT/NgA5xpxZBYlfizf6kNYteHzYA41CTFvqauLTMQPK0EsUqzr6
M0VAZYMPA1kgrZNCi/NCwt/FM4r3I/0KyKMna6luIxs4H46huG6zUJ8slReXbX7rjNRasN6R5wMW
jIIw1yxB1pEYv2OG9iKeAzK8JgjrrNMTUtf6KVr7T7d0A5j3K7qkSIGqAeGEB1fBFXv9JelF9q+r
JhvjNv2nKWDjMan5g6CX4W7m3/yc4x6tgKiQJYzQ/TyT581xx44hIfTVz4aplnpN0qs9W9eZx6mO
7hph7DgHEXceW6uyitd7HOyDgC4FvfZMHwNh+WNWmrPHkLu6yVyMz41UMK/4pjeSTdvxI0jzRmA+
gSvn+E8mq4cPFaBE0v8jrnm3sRQsejs3xNEHUipCvCOtHNWrQVoxsuBzVWPUEn3DKnLBeJ7WRFjs
QMjEZQvxk0TkFa3kpjAZMl0znZ5qxXosIPx5XnFkHZ3Q9ei50Gg33tqexgmfktATfPLbnbHI4Bn6
D0q3jLiHVcbEz/3hElKv0VWFTxqF0F+ZhPyQaQkXvmgMhuVbVPuJO9WwGdEmbFETTJ1MltWvbIGO
CBy8FK5/stHj+Up7DX2qyjYh/YixN/63KMrnku2qPop1mfoX0C9aUBgZYMaN1HHTQ4mGVvjM8iCh
fGC5TiG0vsCjqjjwFrBP2zvuP5vZoC1ryZv2oZDATS0qrwds612AB22XEsRe9/obz06vADj3YQwT
dY4xLN4h9YnHNVsvR6aFffKtiS9ryqtqs76tCkxHZqrn14UqbkrizSUpxBiK4pUpRYdJtDewjcxE
TSCvo93IsdEhbc/StywMa/4nRAYK08UoYeLylmZcMCbOrzMCvbjGZKcEWSOqaLe+06Njv3Zv+y5Y
ehzfEhNwUXB4+JuJylFqAZLTIOanCBy1XZwz4aMkIwkm+/1FdnHbF/QCrRRdqoDDPDKXr1UZmhUa
2q+klfw5VhBwQWunrG+gBs55CP3uQxw3SJiMLsUcmkslZ/FcWc9DLPCvjCLwyYMDYj2YspVzJuoK
F5HxAGYgYOgCWgC7AI7VcFP+0V3BEUuBPF21UsdAewV/BFno9enJycJVtOAsPRcWx7klDZLEdiF6
VqUIQhdJdviUxQk3FFdPjRxZYvG85qwQrbCJmM07OQbK0/aPu8yq85B+Xy/n89E2hrv96a2JwWm1
eHLBDfmZjB44NSloi7Gpr++LxpX7Z06W2GtgGgYA5tll0R+Sc0CYI946LZ/4B83l31SwXNocK0St
FdbKySSa9X3q/44HzXl+Fe9BRuCO2dG3C5fu9QYG/NKULvGCVS7ZN7GHgypCdkNy7WFYj/PRe/PB
+Fo5S2xVjH1UvRspzCm0+ZmbyCvpE6NVcrUIPDiatUUlM/If+/jnvnBimGFoyQvK/MGHN2vWRtOK
ikUpoMcgWoThYVv3BFv7VXvqMGZlrvcWYphORYxcf52Qo6YTable6F5cIy5T52tuVAa4NlKj7M0g
M36JPqMY5ef5pO84W6HPGCj3Y1HQMcY326msTAhtReRTHZMDe1dTBswLhl6K2/Ivfvivj4fYG7/P
iY/vkrbsFT/CEPyW+qjUWKLux7mYn2m1Y2keTxj1l4ojcFdUY3DT5o572SdLB70hJQcLeg2Mnkzf
PMbvrQ/I20axkcrWDFQGr/U8UseuV0hrM+eJCypN8dQ2KuGAsv1PVf9ueHXmp7N81XjsoxkATvQR
iv14XkYL23LW0kgrMbOseMAatd9JjT6NGiz/8rPA7V8GNEbnGnsl7vVJ/MT7tB0cetnKg1/OT3+S
5J5AHBJPqsnB8ljK0dbTH3xN9lKAnU7148mljDwHPXlJlDjsRUfadFeGN/pn9U0vQzVNJh8L7aZE
sDPmYh3tlH1xSNtcS+nZs6NYKHicHsOujbG3zCfl7qYH36ecMqZEXCQUVL/BS8ySx9I6SPhW8cVx
EMnBZ1FdGTchVpL/0TEstpceREw62aLI17anOvjiSQ0X6iE9ZJqnePaBdIqd3GJvE2dAN85YvW1s
DbMFyFCMuizbOf6lB7GvphO69birZChO7a5+ftsKJ/aJXKVQPSrmcLqcCBsONv59yDyLzvGCq78L
ch/2nbozZcu3xtVb+lrvbJaWSv0LTZs7SFCSbVV5ck4Ph5xaUsMq/jiVi6khgxL5YpyHYKQDf98Q
CVwgs8m5hNCrbTnjdqdxNDu6F4B1kPTPiRjsP+vMF85xnbDdDdqQk3J9t/8uxe72iyBH6QnLqmGb
3Sd1kWCmYTHSUfjMWMgbmySERtP8W+XmatQwoIKtgNGF6Dy8hQSozE7KAnR8Cp/vCbSn7NJWMXc6
diKhgkpI6Z5f8MrX1xhbnbLHiiBHI+l+kYUPQV0W/T3z4ES7Iu1TaagBONP3QxT6TlKA3EjUUUJQ
put0eY62ZnBjtfiPubXgEDw48rjAAnwJqpRAs1L7ZUzKBfPB3yX205aIlJO8MFR450pyAu01aJYJ
+lJ59I9i1xzdwo97X17rCZYjXceopq7HfLo2nF8kwcAD4wn9oSXjYMTHDr7if9my8NkULZ/5GiwJ
yunGs0mYrHMYOKr4rG3h2jXgHgT6UQOW82FbDC51WYWfdOa0ZmcH4WRB6uSXeLbZ8taCoqsgShSL
rIf2gQ37zqL92NVNCcQs1ahqypnIskSvMDitII/UH14EGwovemvus2ws29juV36ttB/iJ9MnE6/V
DLm0wU24AnyEQvhu/lgwelw0+csXChxFhT/O75hArmOZkjN7EY5rSigu8Fp2vSp8B2u2M9Q1TLPR
R+ZB313i99JySV2usFc2UNCSkNQZEyLy7CtJtmn+g+maQ9C960/0e83+ieJQ5fXB4smrL+m+Mb5M
mZPc52H0IP7C4XSn5itDLL4fB6l/GzgnUrIeqPsD4Dwt5yv/rCxPFNWvRViCM24cWUrWHaESEoqn
7XWksyHNS9OgeQBiiz9BPU5t89qIQ+ZdKIp7+STmbKYdf9r1FU/hLLIbsL4iJwIRCinMvhQ8BPet
prHJB5yrTbxCtWmmqHAHshuxxVjX5tI6TnMoG8epEg4qX8DuB9xw7CoPefcNU8RUjnmLf79oqq5c
0hhZDVTpEPPk5vp7i/dr7LcRMR6AICuakP2imP4Bd+4muFgBXzaja+ZV+i4JMcx0ytW3AuRx283y
zSl7eYIujEEqEqWVLcH+6XWGtdpDxhuyBTNB2WjONfES49oJFnJvRI9MWRdCCsJmeqcJ0KMv7GPP
NkdA8k7QvOoHFFP0dg6Ca2OUidGtKBsyKaqSncjnJ2T0rYCYqFM0CS2ma5qqFTp7CterJb6YIYjp
5jCAG9dHKCGULKLsqwUZFxnnnmCKCMtbUFU+3fYfWeeCQYYaNgAm8SOie5NBJzY15/nnP6rWY4Nq
vM2Z9pgjqokUjXEa8QUFzzRPei9h18YmT6JptCpBcZsbpBoEbw5j91FytXUgnRZ36Ypnc9RdxRpm
7puz7Ua75sw59yvo/ciI8ETs+BvfDAWIvYfr4QDWcOySPs+MS0aRWiwPUh1jc8dOBH92B1jLmJ47
uHqcMe7g/LRgQzlpCRMCDwgzAVCxt8E/VllkNt1AUJwhZnSL19mi9+N4dzY0SgnI8cRHueJpOCTf
tOpNWQKXp4HDDu0DXdn4nHkGTR4uBTuJ7tDOOaESwBsMGRlEw6R0R/+KW9F1teM5Yu+NxhCEvCeo
jkZVjrfs4GMHd/piB9bdg1HJoV9sEnof+dpHt4sN5IQDsXJTdxsYFaUafSAALnlflx6iSfNM/bhz
I78d+rLqqg3Y3q7g7JRbqIzwQvdhIaLCcZfuXHj8tAismQfsjIq6Buh+ozInU/Ghg7A8REn49k5G
oDKMt3RqgoIPJN4K51u5tp50wUt0uDPIvhTZxApmKqRKqpiVAnS7xPy9oqxER9iDoDmZIyNLQH0A
ITfR6utQPGKyoY0v8bnAduUK2GngLs+NlD3+982RHJNM+strPjiKO0/00tFfbAAcqos2ybY9Tehe
6nSg1wHl6Ke1XWieSoz3B5LY/KVQb/AiAZG4U1Wu79kYBJsByFZr+tTqMDVhglcbRSJwArvtkckT
bpsovuVwkUKyl/zi0sdXIwpE1tQ07PqtxBLP8pbbB/U/P7LXVjO8vMhojRVZUZ4tXx9bXtvKqc0A
PpYHN/Vbh6bgJV2bHCIzGJOQggjbRbLDPvAsDBXzWbPkHZx84Ayf0mM1RohlUF3b92YfbYFNE9ur
5GsMxm+9Ipid4XYNHuaunVAE/yNSOV6w4nhfIfbYF2hZIR9cpz6s4oGaV5TASXTkiUQhBd6AuivD
v9aA8HmhpH/lH+h99cXsXxRHEyaYSW875U6I2bTW7AZ7OKMn3g+qcUuoMwssotuNyQCWgFulqsKe
1ML0/OwOjekPQSy28rKCAPc+HnRuyWk3UE3+n7YKuTvdVNUkMsw0jiECtHUWZx4/Rz2Svv0xMCUk
ITbokUlZXkB8ZimsdrUFvavYObv31EJphBeg1Tr50mL/+MJV0xspbP0Bzb/U6wzTuKhXO73+KdQV
bDmr5YpzCXrbNj2OkDDtqBwVUOHxeivH4M9xMX8FlkKHjO95b9uJX+iCLlRUXZ9qpw3+WZDuRSNj
EvpJZPEYMwuiXZplLNWUBcULS4zMaFsLBJJpdBYkjabD8rPBeQj0QmJBAOMwhOjrCE+m7TKzQ/LN
NSHILhFW+MPUNj/Z3oUr6Q6Xm+Vx/z17LsjyxRA8wy5k5QKKUYr5tEVFrwPsFJ5TsEqnEOlHecrb
ptYLwPZztiwZehHoxgx4+bqeOCBUaSKTfinN+zvt9yiAMYLEhXyOmPZzI2jtUAS09ZOhy7WkXUs7
DvM1Q96N2ETzJ4r2OLN0J++kKlIFshHRZNLIWFTu73XkKE6lg4Xc5ghu0oOHy8J467JIFg0DiVTl
9aRdrztNRpAvCDRjQ07qNCXJdEZERLCPJj95IZEBBRJewY76lpEc4wSxb4nhvVT7dNJCflIcF5Y/
6pWR1okUfS/vvCaLsT5EsBIQszb54zHBv+IYdoqCba/DMvb/s28lEHa8UhS2y2GjV7Q4VnCodttu
4+Vs7WdUhp7ZYArPot/UCFdK713hlpe3E/Lerc7qOLPCK7AUQg+LotkeRHbb/GAxdDneGXaDz9PE
DQFUDOVOdk+yzQU/O4MkONOGjCTUv8KMx6PDE3gsJZJKvoSjQw6uDNJuhJjmw2HgVB9UsQtAayvp
7rDKmuDspKp7NsjgpXOYz5Z2osnwnkVQNPFcgBjKmw2ovhIv3Qrd74p9BZpjRlG2DHTA3dlUXGZc
t4WXIleHsQs/EGN1axAVApixIRbJxUXHKZnvtMaPI1fr+bC868pahnDqZMULI7ZbGkZDVIY9rk0B
5iMFs5hmbxaxZyPWCjoyo3ILOkdgzpxTXf3gcxqQ6v53Eik4adoylIu/WHGUCCtzWwdqW8h/6GqA
TX2L8rED41aXlY+/oFQGaXfp1XIWQgmMfeWBGP/pS7t7b4C8fK1rWrbO/UPE2W+MpughOCmWEySX
8LFFRrb1XRjXXns6c75QmdpOSYQEM4RTaSyJblF6Zf9pRyEHFzlWg89+/ibQBgromkkIDNO7irHh
RuF6Kr5Ihozoj7PGdbc33tjxfkKHufUn73VDI2xXb+6wP9IFaIMfcAQRGYNf6WOpL656uQUW23Mq
Nwt9qTE9MoIPZOFdgPKiufDkz0UieDFwUL8Lmcg5HDMpuTDlst+L1HlkdSnqwP8j0H3I6sJJykpD
Fq+2hMG+afrAvBB8iPj96FNQGOo+9IGJzKV85xTkeT9M62sgktJSSABHTsOHDOxrSXMQ8egjc1lC
uH+gSMXDTuILCkRebZfMeLlgxxPaR3QmD8P5a0jhLN7E27r+33RVMA970TwS/8POGuzi5sHzhXfD
yp489APRqTAotvN7RzYmLwGmpCC/DA+AzsyrNo2yg9GQiMcuMp7v7p1SK8BLath1rkVeXj8KcYqz
wCYuAfSmh31S3YGL5EZhKyJZkeawF/jkOe35YcS6yvech3BSHUSu7yXFWWBT/Dj6UNZPt189/UsE
AE82PxtYEH6KIoaiDUSTMXzRrsSBle9tRYkFeTDWMcDbmZkqisgvkxMyjmAfr8gNS0RVigRko29M
fbmu003nVj+hiK75/CwjP5/Z4mFXtXtlViK0YPo/lCa8PAATaOR8HD34XzlBhQDuyS4mFt5x7K88
HDPtzvl6ggUmHEubE3wrMAh93Qj8b0Z4IftUG4BYEcsiUOrCmJ692Atlu26n7KVlzhzwyJHigsVz
pPelBfYZfjZom1F0hk6N7KHEeD7nl9rvdYZmgqVLmFXOTPiBd8UrxPIO+lwCP9U5yoK2g4WkjBu3
aXOs2xfwP5QpQD1M2jFwYFD6ybSV6smeRhvEzUUcSiGrN6ua+wt/i81+U2MJMicXFW8BQSQ+onMu
7SMJLGO6mgg49XtpNYUqBN1izbvBmykjlSONBddSFwE4/Qh3wu8Uc60NnChmNaUd6WgLQPjOrOYN
/RKLpYXwyQxvr0llHe8VqUTCfJc//oDMn1lAjA6pjwl2KcQhQpIt8cdP0bAN9iz37xMzSz4NyjLW
m4XPCy4u3lhIU6mdGhHZAJUQAeh0quw44RmsGfazVKcSBhbCWvQujpyGRhldxswcm6ZzyXB7VhyE
HuS9GjG2fe3ZOt97QQRgCcs155Z02fmRP5VXHkXPFnUd2OzQfai0SshUiPWX+haCNZnS9meC6HdO
Dh2wjVkhLqUXr7eWf6o+STPXGMDdObb75qwJfVTqajqxyzXZsR3hX/ONoNoNyJ7jG07iKvwvhXLl
sieAqRoxiQ7f4ETl6zUI6tb5yMEBHnRj9FI0MnKUKq7Ar0UzGDoKj++7pAz0QGhOL0Vyl/B56AbJ
n/wlWWqa1VOrUxzc5SM+eBnnt9El1/Qob/3rYTbcpp4nPuGae6DRSBti7Glj1byhmlduMO3BKviS
YVKLX20xY7dUaaC1Az8l0pSpQ+pzv2RbM85vPD9R02OxuwBlF2IyGPOmQgPGVA9HtLj00K130iLa
eYYsjubUCCBOqrczaCX6mMZ6CqW8sVqKOD6t3DgQ+eRBcSC5/rPXEmtyQfG0oTBzPSlUqY8Hn50d
DGKo7RF8vf0dLa4QooNktx6lcaSOzdXY6PkhbA6X58ZLTf3Z2i/uQvTY9GGsaOexryADVv+/ITKT
Xa3fr74eqGOUH5d9zNL+ZCWi8keIdfMtRK6T+SCw2YAF0s/CemeoViJc28W16Qnl7BtzpW0w5TyI
4EPq3OX+CfFmFzQ7mmoTD6pv7CFHyAZH3tG0Ulzrz8LjpPb2Idv1nH1Zh/r7fHit2Omd+0u0TwgX
4MES50/FcaPcY5WrETGuy9U092GVspZxRJMtpFy+5n+Afbs/F9lniYyFQRbZW3ozoZsyD+beFASB
suC8DOsn9/S4Qu6YF1TOhGN02ye7kEy+2r8dNEQfpoAcMfOetflwr1x6oBzUdzGYR5+fIBjuq5Wf
BDMdvNTVEjnmILhJSHn11G0oLahRmoXfflxIb+ulK0WACuo4VGku6jyzALssMDKiuLtsvGAFKJhF
C9VOvXMdcPygXjmM+TpbtztvG8KBq2IgmrpKYq6hcfKLTTERHmoaH3JGFJBeZNbgcz3TNxivuB+u
FdRhvu2+rHx7VVVjbRcMGgBae+nABuMIHNDKyNvf7K4H6eLF5w7o6HczHiy2EDgKEfKqDNHuJN3J
ye7i+KYrkNrvayVIOX7KHw36kRjh5cCKu2qRV3G5fB2HZj39aKC3ncLXf8Okn3ZK4Wix5SSI5qYU
7xJK4P9FBoK0m2fYK4Vlt3LQ3VlCBZKefny3dS3RYEEbTtHuRCbpFQ/i0l8TEm5qJhOVrJ93e+gk
h8K9wEEXk3IS5AojxprUpa5da7NAkzGpU8CMlns2wE9Af7NcLK8EPmSLFn88kgWoV0Kz+Jzfblsb
m9/OleIL1EXPJPB/eid0tguBRD9yXxaNFfwTQyPxCFOs6/UD92tQS+QgR+/wrX9iKwGQnKuJVSvA
pZNxQKq3DuqowiJA0fkHlFVY5ghQLgF6ToVyuRPTSWw/3YpJ3NIF773agIqwu+yrHLAyOxJ4kQD3
PwkWpYH6ipIWKdz0FaVhbVSxC+3DQvZLuEpwpfTxoZYo2v0NUMl9wZmuVrKbVb/jE0ytehslvieF
u8Ci+Lm9WUu6G9gAPMSTW+IHgVRyz0bz1d4AbIvq/51viycO3ybqdInyMa/H/9ZV03VmiBTs0Yl9
2zL7t6IXqWfuoH0L6MFp2vKf+2wT4fJ5fN5FO/o757pEF3lbsR+Q5S3IGgDo+ACH0/9Rk79BTmzo
KPDL8tCh6xcb8R5/fYVNLgG+zgK1Ea6KDmNP194XjQZfYxynRjn/kX+OGpcrp+tT4qvDBc2C+JHb
U5EitZylDpS6O2vnz0TxTTnSIhYzgTFs/evn0u+8o9uyrgvDbIFEABviIQ1fUIMkxpf0CwErYU+p
VX59gaPlEWBYZzq6z66w1a6Qu6ppGlL9ncg8Jo1rgG5O3iHLOgGkei+lzaMEjuRgB0vueKqZshEP
n2Fa7mcpCc1/t364+xgNm5K8GQpaQX0TDYUdIZnrMmuu66wkmhGzuGwcvnB7Ec3oeISJpF4yQ/aG
B5qJVCOt18lhy4otrGjVzqvRBKIOYDJ+0/WH7ttHn/0xjdwFZePI13rA3TKmJBxfKD2gtZuXWZhJ
uHOwnfC/V90bh8YFqbqs8xUr+eqssLxSOGMRJMs5QO0wdOOUuqpTMy5JwgE4EK1RkW4Ecq4rAzKI
kW04tDT62lfZTj6JfoAPcLRTrWWyZQONjMkYyT5xTiNwUTeiZqYEH1eX/MzNiVuP2qppHO92zKb6
Bk7AbhkrJVewf5LtfsUVLkM7S5X4G5hEpVu+Mdsn07VcCZYGrMqzvsvnP6UU9uWH88qL93W7kNmU
FBVYGrLj/vtrSj0L4zP17jltWEPME5CbqsJrFfGGqPnjay5UcmOJukEjPMmhAHgTKv8K1zdxufkN
KuUrpzmjE/Kl7SPvgAMkOyWb0wVPKavaPagvMYIrhJmwwh9kLwNXuRBunvlVClTAYVOf8miaiH7M
hzchHA39rcixi4Ut7uMSW1ovZ60quiiixhSDA8Phgu6QnQJeq3lpi3Qr/tY7O/QRxpGTffPRYnDN
oz0+zDTY/bwlynZ+J9CwA65h6R6XadPLLNPEOQuTjlt5nvH8peO9sjlkSIfQcFKVPHk+yTVv6fkw
U3ArjO9nuqOXcXZSIsATsfBNjoN+pgFGqlnmeE6Y8YpB5NLpmEXrGE6fzM/0yUCocWfmJx8KPAzJ
GsKV3xSHdBJ1vlFy5LUXPi9SIh9F0sOYh45ALbU+ec3ybF4IMtRMW0qXiya1MKgwbjAlkQ0mleje
7GAJweaUs4jL1SFqQ+brPAHPPtRXQwIYLgk+vnbaMatUe2W+TQH8RTZPR1hNt6ymx5XRdqe31mv1
3nkneKRFjn5b+73jYXkJ60iOY1zzgZJQJovd+EHMbzM+zbdhG5fe8Att/NhaXDt7LebiYkl0xZ+2
2JTpJdin/DsgDU6K7AOMtNnH5qm9XI+rAdeqJN1LxWVoHF8JcMhuFJ+/8wmXsI67yMt5ygxAgMK8
wC8Zt8xS8XWeqy8XnDY8J4Xx/20BQDc2Jm3bs5D2lITgBq4SPlFVAYp1rxGZSAXoO5TTzMLue/C5
Qngv1g6zRj8ul6Rir7ydj9qVmHLL1eb29bT0Qn2O186tLS8CvyJr/CX0AeC6xnkwZpXBzgTTkBG6
kDDJo5ppwTvjXcY0mtt16MZqrPIQKNNFN5zk/11W/nKvOp1L+LYK4byevulxKojg/nNEHp4YE953
qkP6xBSxbuswXYYDSLaemaYkk6eqoew7246izVcUjj+7e1AKfWaOxeP0ysYCvmZfJGR09GcxhWZ0
PqvMbJji7OrRpqDSpCTwepwA+uzv5CQDMgpISjIa7JyeYplQ1YAiwGpOD9/KdGNPCIhS+HFdtx+m
sNFu+wASnd8BShPprVKdmO2u6S0pGD9xGAeVJsjL/WS/moFVSnBq8tpmBuHYKNcBaiCg7CxEoUd/
tHzbJgaUaIPWRzyfchdaX42vgDx4tAZ+PiiQOvii7ctFPClawYIeWkitvjGTU0pi+ttxwGrjtvs6
1B4jdtI/NvNS014RS97mb9t7iJQzXKAO1EI6Rt3Wxn1thFPiDSIx0leIVrXUSNHL/gl3qwInh0GV
5X/4mv4eZcuXCeCmQDBxDvJfrAwYeNURRbYRMcjiQB2bCZxYrKldBji+7BtsE22Vtd11pNmvrYCA
TnBaamVpIS1RG7mXUEI8SlEK3A9848yKX1KR2akcx9Z5jGvEKT4O3wgvkaQVWwlmwiBa+Et417y5
8Wi2jXpvRknGxm2sNoLMbvvmVSQgRxavpBp1NmFB+P5+xTW8hLiw7QsMmS3gZhLIJjqIo5kzKR8h
3IUiyxpr/puVZkrHj8qsmdxlsUhBnXQ6WmLSf+SMSxVVnYkkVS0jI0X7+k1fFcE4x5rdFHciGHSm
gC9JJtlF7mNfcEAloTh7bWzwQrvt7Yxx0W2dQdfzq3Ls5XvNwWoJgPbD/qqYXJesjahywirUkLhQ
fHhARW5Obw84XrHVMmefeSVB6HbQflcV45mgFZN96UipwHJNH5AK6JxZkTs8kD+XJYkEJLbLgw6D
Q0+5H84IqnXAVeeVTLeb509Bwn+jPytzb7BclkARxZzraggSVlLxudxoZzaJ8acgBCGqSO2ijF6D
VnqM/rZ28Yj6tcx8t+skSYDKfmfsQ0Es1jAMmGqUo1x3uV/2brPqQkWHV6g64vl/lpanIzBObB9T
r9jGigKiLfz3whlhwqmCoyfoUAEg1DWhe2q0FrU2sun0LldGPSlk/IcA1xBMXetTeRfYczeexaAx
0d/oQbtzDl30N5lEMORWyOZSpKOLBPZO5QXkGH9cgiRf+m7duN3mcL89LU91Wz5dnrjdRywKfltF
npYFRUKZcHIk51iKQiDOnWEM/YufH+t0M5G6OkESw2tzgC+SPaDhjdnopcX3Uqz+jE7xlaxwh6x+
/Xf0XoEc/aB0e/tzPRK7uov3Cv3R6MdrIhNpro55/EdNPzScwnWjzByqi5KwhGXEzdMS61eSRKge
xcRM+8hz2f+LWkdN8bFJdtESjUT1Utlv3dlK2Rd6aDwRE8ZYktYIRIfNCCPQWbpAYILVRIWRr+NL
2wcBxpE2cw5s8eYsNT9NZ10VB3MsrG9K0wCNW1UsvrnT3VCI3a4y6yNkXBF2DIgXslgkFeITHIGN
rYdylYOne9gzrhFzhs57Jht0En2z1BuJ9DfKNudsFmwZcqDp/thgrcYQcnM9rU9PQSfVowSB8Xcj
EgN6ab+xLDiyjeXwWxpCii1jTaoQBQk/UF1TOS+vueepoEEFbu93p6iMKO3dKyI8XehYQPEliFka
QJocMj7yEk5Y5zqcDsbEivLTp9Ek8g7oBelHc+uII6lFZnLGHipuxQaoxqJfBQmhp9KN8/HVmC7a
R4JgAloroL+IKINrUv+a0C97jJ3rq4Vw+Z1ISKRtqpbsXafXPsxBVz0mH/QK+mpX16+4vc4f8S0Y
e32JVyzNftA7RZZl8x7ya2bsJrdUVpAzhjGrhlpVT0u7PgXSG2x+DTJSwUiIgQqXq8HCCyK3YRGh
C7SHQu9wXRNfPNmhC2BKAV5i9Sf0n4WCcXI66v+1aIzUEzq4S7lJYh+vNuP/PorfoKBawiphco+U
gywPkJGOoPIzgu/QdSmfXEODXS+QTQ4tPA5jGyaJNIXU6GSgEJ+sm0i7jfZAH7+Hw9Ar8hYA7+iQ
PtNfUXayMMukT8insZeSAlJmn+tXpzWV9rlp4x/kWYPlkm4nbPGLfWVYPPAmXAMOn/stjTxcqFbB
G7azLyOTTDjOjSb9cPfx3H15A4XnOn59Tl7THyGc7nbLoW7XAVk5IpMcKnYMiVGebM2TwQhhbb1h
DJbLpm6yt6N3CDWau0Wpt1+tFf8LQqwdrBVk/NuJLAust7xUuDbAb7ZQuuKErGpOrPmFFtMn7WkL
dgbjYCJXlpdPVXba4KZ12cY3qsi7pi7g9y+Vx93gJK/4lW/d0x9Jtr9Vc2BtwbJ0s/+Hq6wfzfop
kzNRye7ZF/dIugvMWLz4wB9OzX2haq8VTZj+UCUWBeQCEla8tfyt4ND1bnJ8ls9b2P1UgZE58OO1
m7C0qz6m8WEMOka6N8KhH9AwjYUxfglmGKCxQh4jnNM7/+EtjB507D7wZnFXSsKHPQfdzjtPiViH
5HpJx7NJ3HIe6vFt+dk497jK6uVvn71RL5Qck8Z4IzTgZenpTN5XENfFEeJGM2FA27OQP/qZSuH0
yDKzN7hu9QmBQWOPlteon/FvzK9ToxJFB3E2iUaFAJFt6IuabqZONeIIlAwYU4GpczbnG1/Afkmn
wPSnlTkfj/EUGHw/Fs5rFjBBaQJPrXHXQsMzL9ypKc/+WkzMRhKE5zuAmzM00Dot4xAgQRL8EPK1
+4CjshyTG8R6wMI3iYzR+GuXY5YfQEszzbuaJiiYiOS7AUTzLu90ucTMbV2Dd96QvghQ68ipFYhQ
qOKoWuJ61vLi6nq2taHzSDNQI7dD5Tgw+8QCa1OXWpEJU8hrxkzC3fYl+MEm7ser2q67a464YDR2
+rVZB5hQIuy4d1fKOM1/uoK278doSVzzKHHJHJYc85AxRyBzIC6rDyTh05OntL0TOT++l/rMDP81
uyzLWfdxawh6R55PfmYwCXQ+ARkfeJlkmLCFXplWvODzdW6bUukGGP04JTTJuf/h9NEfGT3JlWe3
PBdzG+jgnoHABs/iNPPwvYWI2m2eSU+Thhc7dLSJOph52TXMWlNyD33mwBA1DUqOT2Ntpf6Gq1rx
gMiNeui/hzga33IObprIJau9fxvihqvmC0y113DD9lnNLs2qKsP0KYJjJhS/oVM4GlgwCSOQCqoY
PshXtW/jLsS5TguBENr0lu6zcjn8yt5H23J+CWarXyJoeBkLLXbuMYvTC80KqrR2PryZZxA0hg7E
LiYD8R5kKfJVVJ+a94KJePCf527zNNcBn1yUz+RC8prq+Wi53zc6bCyf1QJQfR9sE0e5GUBpuM5+
N7FMz9hHkBpWzPeXeGyXHf/OxXCuKV+wIx6Np2wqzg5msWPmHYRpC2SgwfortOp84lNKCIxj8uQr
+bJioN96fU7e+eeD+qeajI3biB05ct7Aivmfby+PEvgpRq5BRtaZSknX+P0dNThtgcth5iHwwRsE
929B45QWeYrORbAhQVZQKsQCyjGQuTmud98/KG8haiXEx01q+wHOC1am1Yc0oyhWX5po8DN0nKwI
FOiOy0U50BnBygbs380Uc+tHTin7xQve6GWPxoWdDKB6SAMhXHXMK/j5wz5E9PsDOle+ntHeMeBJ
NCsJtjF3dK+iFPCi2LJmDiN1jwzrKbolOFPNy5CC/q8K3Fho9wHxG28EplJO6t3V94Szu0sQNEd0
OeBC6bzuk/9KAyLpi9NwrBfkffxjgKPHEGfkX5U5pmKLJ0ylCYEZah0txmjbISLnQKEDRCMqwsZR
L4wER0bCVJ2T5uASAQFj3nHKVb24WlKAvIoww9izfj0XqcTu+sXRhqxbP8qYT2XaYeNwET8cDXRx
Yyvyn7CM08AUe6ioj29j35ObGLYOrDCEDezIiaGpMFtaRGRmcdr3O83G3oO/eCKui//ZRCBgm8Zo
8uyfDnfSemfbK4Guajv/tsHqmoP4Hv4J7HARwLycz49zHQJxYn6NZ7HLysKI7x3hQiHElCqSgWja
8bMVLDNKWry1qc2Vuume12BIXr5X35k9Vco+NJ2X8eBDvz/A7FX/+D2qUjtBq9c0WHzBuEhOW+IN
V4nubBOFFOaXRxkBzbNV4y1puvMzo13aPJ8Ozqq928cm5ZHMyjxmbSy5A73vGAg+4oJmahD4Cqsl
xs/la6GGySez031G4GELNKX3ac8ZtuwaC3Xoog4lxm/vLyUCmUDpfODQ9T4P69Gegg+Aiim7ULhf
DZmd6I7SYwzu1laoCnmf59UzfxJOvw+SpqGQK6odrZ1vRQzdAkOgCnXbbuwjXWHQjbEcrkWqyRCF
Fhk5/OssnG8WGq1jSBiP2GJKJ1ZV9ug+S5WgZTAmYi448biJCtogNltYUQWHFyJmNWrlCll5y4kl
c9tv4sYjY09myNj3gt5w2bzcvBtsfrhqf4v2SX0QOr6eamDY7aOcbrJ75NEqbPf7voe/YfJbOm0j
rMlYhaB2x9OZ3tKgXJr67f/2B5Z2quH7g8Pma5haGyLKos4lCbDSntuNyISxLRfFvtvSMz/9+7GL
3Lre5kyQJN4ryIgXwa5Lwm5rgCmvtnJVUipNb8PiBeQqmJcB+VGhm1OGwkqkdBlf/w/1Sjy2CS08
dZAekuwfxwQb+6NkL75y722IUJC6viObBh11eS3pVgtapMmyFGhWnD9sqcvWZqFTCozj67AUnU1i
tX28qcWVYkvBABPPeQytJi7u4IZNeI+mm/8QoWYyYkHx9h0eEKPbzaUvq+0TuCUtbZVYDqJKDWiM
f1aVYNKuDXsCSDk7LekkBvtRdAYaL3sQZkrnhFIwf0YYvybVmvlKOlGeWs2EgtxXTVkBxF7WLqgZ
10heiwLdKz0fj03oDad3+EK5xyTaPqcXHb/ClNg9ZZloLmM7zaK6Dk1p6NECblPnTYl6wCe2+Pex
RgrtrPKjSoiITpg9wQUQ7Ve/dUqm9jYCBAPv8Zoi5AoJNxX2FFbIBldWucDPOlOgbDSWx68aFboM
fvlP+AcOGOybKXh4Hg06+EQiiyLqpmcQfzMZcxu4UH6CXKdVlK2T+o0VuDSI1ozvXZM4SCdzcb5L
kS9uDf8Ub4LSU6AvfbhDwufr2anRY6fz2x/CHqFOgxMmw0PtWj7GQJ9oOgm/KmZ37bUdOLffjNZ5
CalycHspPacioy0jAOTq91Uzgi7l+vS0B4SVuellPkCwkFArjmVtQPir3Bx/HFaOdN1V+ME1/d1r
g+P5YEFF0IWrU45RA3Rtp96s/9oFWRYJ1Sln4oq3wvDtVHx5rZqxMn8neagX0qogNd2S+O9jYR1N
l4cN+O5v5ceQscrZF6uoZGjKU765cb32k6PKjqI83c3kHc2TGGyCqiE+2muB+kuQ+GCHSAJE9/PL
zbM7k27nxmnEaw9m08hu0e8yGUKf4TO+o4NyKKvLR4b/ZpCfacZ/jxChUNzfztpLmcUsQ9ffm737
/G9jUTwvTLT4vmupi6hh2+YKknil9XvKfODibGTh5xDWsFdtU73kDeOawoccb7cH3P64Iz3wGrB7
7xap20fZnMAcVJLZD2R5Bjx2MVl88Lm3XZ3V9DoBReWS3oerDXSrubsonrJVGZyUEtTaP99I7/pS
lhfwQ+Gu2RWUmSc0N3S63rmoU8P9kzAyAI5aV8+T0BgOeVqdxGpzV27bUNYguWaOPXRvllSvZEq+
AdmUklz3v1a3455GIJeYNEwTgbmyiym7TcF+VFMqJMwqpXqhVF8XcpP0qDUoF1o1I2MA10DPJ9Oa
TEAp35dssKOK41UXyywYXN0YWZ6ZVMVAl3QLIsm9vrad2f28m/Cip3HUR1B6i48GkOkgaV7/v7sy
zbtW068LC2+L7LTwe/dN/hdO3KVV+D0HPk1d+HgKsqmYwDbRJVvPb+j4IKbg8fzWYRl6GjpWk6AX
8rI0+SPDGkpDt6R67juJ3Twj74yHfnXKe4/AG42uSjEDTo5ZtKAmvJPW8Qe64RjhZHsy29dCSEH+
/fMvXV1E9wQ+WDrdcYNAF4Ph4ttE+jGSQ6skLX39gKLVkX8h9R6I4QsEiRneB/D8RZ0IzCGXo3Q3
wT0xteJqv/s5XvzIG1qlscPUs/8gB2DGl+zKFJfot7FEOVZSap/P+d95P7knTZCO3LY510mNR4+c
q/V/Wb023jH7aVIZzj29J9K+Mp2TypwWoiXxJmbCygmAC5ev8KfBbUGM251nUrecGQ7z4sXjr9R1
gFeQgN1pxCnGF/GKI/zxUHcsDDq9mkXrmzOnCQ7cvSFz0WHG465DJbAufHj4vh2PZ9BqcP8wvUTQ
BCOPq/dfGm6BiN9ZUWQkNTlD92FuwDHtzy+CJHaMIJYAZMwRZ+CJ4ziCuLA3yyOxrZ+v3Rb15mMm
NWvhzl8JlUGMGw/sqSTeBwQ5IvhnQ06+9rZablBnieV/U6BTBBpsVMVLdOS9r6juN3t766+xN784
V43eK5zZ+WRT5vwE2aF9XPTtMQByAGVe6rmnNJMPwuuQyvVXPJ+ucZ9vnS3bWK9+QWd78K2L7KOz
RIPBYsUKyw7kesvtsOJdKK6mZGsxKLIYU5UVVkSJ/DbzP1rcLc50ZxD/9qDncpiX+WmlJhx/dzaj
4Z3IgKO4YHX7gefN0H06oPn3Mq2en9bu+t0NIwwepk5JkhO5eR8FMOfqnI6YlisxBrKBOapqjNyI
mAuQt05vQtS6obMYCy5x7O0f5efvN8rK4RZKJAUG10ory7H26aEEDdGafxL4uqvI07v3TNfRyyKI
X8mGXBrTq1UKS9EURC9+zZG4OKDXsM5vgntuw22bKdIT4KB+kOy8Wn5TupLWMc0S+RORMcGc7wuP
mm2kJy8UbFb7SiB8FUCCKorz1xhUnS7pux7ZYBwi4S22JL+1qFLorH3JJBRE0dY/OEw4HmTwv/zC
lZt/qo/9FvnUu0TSTZ2/S5GiKkwYQmIUTdFBnjXcCaAwNAQUXR408KjU3oNKa0KdDWdieoPBvttg
e+zBRiN0GjiqvTS8I/dA6Nwnuf+Un2p9/+ylD11q7g4/oAOJZbvJsyDWt8dU+Ish6pmQTvqFVRGV
M8gR8D+AQx50Q2RvdivSGLpnOrReBunUKFp7jIh+0qIwH4CnC70DIkzmgToRqd5IuXbu3s4SlSS5
2es1KgudU8dhX1cIEj7+xYlYVCYA+/ZWDGSls9CARnmuNegOEtt0cOZZXmLCXFaftpqIdz7+54jA
jhwx6hROYSIv5jDFBF4MPIap+t7PgqHU+/i1lWYmHLJR0CK39sHdrvHO6lh0xbDHgmmuyji2nQBB
gi6SAKyJ4VuQIDYv7uQUMrH+4QHGfjCMCrph+dHxDewtP/4S/PUMCm4CiQzGOFn/fuflllfEJ2PE
vxOcQbFdLLfcdLDCA2R3DCLqEGpj6KhYs2ETNjiu2qvJ48m2uZHBsVo2EuqbTuJPd+PsVS8GJ5Dr
kjwMu2tShEzpjLhczs2EEQ5yJ/AtKnl6RMps9qaTuT+z3xLf1nyFbDSni+0Ymp8Rs4TxGx8+UloA
CVV2DyxMNAiFJFYF2ql+0H/WCUuLbwqkHzHCogw0Z3E47fI5vvs8fcAyGul8oUA77ip58eHKU0Qk
hdXVGzV73fSPEFpUD8qK/7d+YYPtKByPujVSSH2X8HyXCQLo5PBrxAvCoZDC7k/hSanGbV3AJYtn
tepk5iDwlbI57sm9Uv+zfQeANFgmB0rFEnUS7NjR/J0ZO2jx9tvemvgRcRCIzuWkA3dBIsbdW+AX
guD2gwu4e9fDHajBSVsVscMgIGXQlmw0LguO7hNDMsKCZ6j993CaCUp6MvRoghAPc1bHnMRIjpjS
toATLdgzD0RFiNYn77BmYSigpRyUqmU9VHW5ULN+jT3wktKd9Zi64ItRSIFqzEb4hrdPdBcZcVmX
wQwWVthuwh5gs/x6I+1safsWWmWTZQBaG/M5kqTIc6Ekn1uoBNh9b8bRLSbpJAHinueHKrLyzzDA
YyLc+0TY2I9YdIl5mL29aO2jNys79YEC8htrr06eREttZJ0eksmCMoYQGepSxqUt2EmSSgAWfyVB
oaQiM7lw7rztDLscXD5Id2eZI/NB+pHVZx6oNEaynoPk5I/EVRbwXqse51xvJSWDLhrei3eM6m1i
33Q75Ps+yDYnamxumqWFmYX12sDfQN/dfCX41ApAeqhQ9zMpmUOEHAzNr8Zan0jFwsqHAyxKdg2N
67/1MVM+lfCLuyYOyYK24B/DuOMwJMWAE87m4EuczZ6oxPSaur/iAEG6rb73d792Pyz26at6rQXk
5q+oqhuuj3GKYnNo+CXpHBgJ0R3wJMOBYgfwMtH2nMwiXr+iNy11FV+ScZwr4ea18XVl8oexO4yZ
EER/WrQYrQJzuXhwb+ffnkhCkDk4evwp0MQei1SRtISLQfhfxtWQzlrJjecIsoJ3DLPscCnpfGQ0
0YrHCT+waWLiIEWlx8JbSOrm2IyLtD6DOcMwpLkPWgd0v5YzmXf9QMI4kvf8T4vz73TCRodSKSfq
s9My6R8mkQvok+pegdZjMADlnzp/64/r9aiIexLDDtogn96jY7mwDLN0RsUuTSzcirVCUjvHydbt
qTBZRjr+0VAuFjdVGfrAQv37cuI6bhy34g8xgxK4W7exaVe+Ra8B+DM1roQM02apQZ9fopSKomqz
jgLLzH/WVNLPyhsen18/j/4JIPHdltGBUjfVo7aUYNFLI/yO6xx06V+Uf195En2gwMA5cR59JeMX
DBx8JfXDiA37HTndTQk1Bmjt5EhOPP2qmSyl69WKJv7zPg4vY7zeZB3oEHgvZeU0Rtd5OnpXNUw1
IkBd+2eW0rDLlnG2rP9HI4Q51h1EgobZRIDLSMT7LWuWO7NVfD307OM/I0kFmBQkG0KBZX8Gkzu8
uh8s+zluW6rxXd1O6+CjyH3CsRLoKZ9Bsm8nN8UW5IOpkBtUcLYwjKQ1mRPbnP7NAM9ABumzrprH
Pn2FUyoHp1lR0qWHDZxdSRUaTr8yyamZFgLmZJJVQ84THPOlWsW59jmC2lk9w8WMWlRmECNDJGMj
aOq1FyfY0wfAOJYhaTPShwpKr0QD0C4EK5jw2Iwuofcuori2hFk/nLPwgW/19WPFf9zACLbb5cZ0
cUG8JrU9Xx2xpN6sfM1tppD/ZU97n8xgdGKx05jG90n0mE7jAA5tNnLxl1Ufmy5ZidsaFT4kuSaX
k9HdIbm6pInQ6FXuGKKIoT5xWsA1GwGD6PJiTFPGLJKEE+60rle5jrQPkaiv5n1Gpl2IXscIwjAJ
KmVx9azx9RnRSb3N5BzoVM5Se8jS9seNKNzn84P6FbqJG2QehTOl9em2aKG56rEuxA6tDhHdkYN7
97c91/LxRXUIK3k9Xp433jtD7FBTl+TL/+V+ACKCMr/Xn6WA3n67LnxApK/MDcmQleiHbXXtLzeK
0yjEfdvWPKEA020zZvKbuKiF3aHsofmqZ6v/6irBOpLa28j0xhkoL7KAKyCmkU+jK7/6+D+f6VTg
LsG1p91TtVgvBhh+DH/rzitz65PlMbBD2UPkD/Y7T0DF3JvyDPXDho1dO7WiDODJ7f//wYJHgzjl
2Csl/jGZ0cSo8usRVoC6pIJIJkESXizLUElproFOON8n1nh9tWoK0OeoH002viLwBQGzWk1/AOj9
KuPYStDh27jpAgQV1uAHr15JqjhYGTcpEhGFIh8DULEPOHK5NRTBUKyi4ohGzqJWDBrET5uXcE0f
QZJWvWgGJaKGJhRzrEJL8W9ou1aEod1WEt0qCBnIAmj+LmvA3SIOlfQ/oEjoYCV2HpORQ0zLR7e0
Cbzr7Jgmdi3wrzI9o7aZpBHbTrii+84RmFR87pUfTSQps8aLp2KOj31L8wcVjKi6oErI1WRo7YUj
d50AIjxVjqz15e5CEwbaL9w9JRBkzCI1FEQxBxHd86b3D8KZ6l2zpmAhOnHzh6BESxpriXs45g0p
4zCwILDVB11BN7jD0TsSvZwpwVVVuYGqYNvf4czR1aJeWFWW1VLXBWT2orDbXuymjxuo6ATneOxi
EkZaIpQGRnuJcls+HykYMkoObWOGIMnDk9vCmLSTqQEVlSErB0CqsFLOetlDHP0hNO747YZ1Po6X
QOsgQG9JK7MdSoIDRztiUXxqE5nlryIjhBiP9/JbDNheNcIsM+d04RMplzR/5Y8dzlIVLe9WEmRp
2L3nqLc8doiGAk24ZwcHVwPGkUN35LL+qBYJnCkzjWV5yQ0cL0xwTT2ftnj4NLv/qmxPkFKtcOl1
xLtbsSPEBdgU1sZ4aUUlcWM4uUgt4fYlI1F/rmEcsMjpbdS/F2tnH7x8ETbeWHee7xLOBLaeTyMN
XDgLdj4/1j/uF9Ud7Wdoiwj+AMkyYYHV9UDm4G+FX3yzviSAaYMnnm2AnNFJG0yrkXhhveD2J14R
olBXNzTvCdYvRQgUK06Tk/p5EdAw1cEyKVmVeF4mhVLgJs6Ect5YIesqLfUt3VYvHB4tFNa7PHpc
NY8Xe8vHV8I+I/EHOhAuJVrInyXKJTlOX0kZykixaimU/GBhSYkjvDnMZp/XdlleUsbyUL0861+D
CjhenNgTJPfTePfH5v5l9PUFekraObEAfjDkoekJKl0VngKOlfEU9SC/wgW4/esTVlEwKYUMY1FN
ULLl+iM0pPQq4vYUS+iCjMRwEZEUs4zDOCqtnQ9+CMvwSdky0LQYCMrYOkdZ6SyJHFzPd9f2B69W
oAo2ckNB/4a3oUdW6tVavS2uXUm2JUHQliKhBwwaOByChhB61n6rP1ZpbbJqiccxbE8BaIhm4gX8
2eq55rw+p1ZRLDy7nN0Gr5k271nQnVUS3A+SO3soI+zTNGuKkzyE89qbumK9YzwB+dy7j2Qei59y
Q0h/jWglCoAJmg6tS42ukgCpdCpDSq1vbAcmR+gPWnS3nYSvv9tiGEs0f/Tz0YSUgtspVoJjjqh1
qxrkutMLfaAgf/HRWs2KKizmrJz3DT5c1+L7KGKqXH2xMqli8Y2cf2gnzhBB3zdbEXSEbJ7Vk6YR
wXYUP27oD6+LPoylM/+9B4jQ9XMeTM5SnFgoIgm9WFoKDDm8th25fG07/nT6iKXSAYT33M4vGKSh
ASDeBR7lTU4GIhiURU1uAUBMS6tdZxiB3928bOHQKEfRwBstrma0TCMrvaYLv5yf6l6vpe/VUwSZ
Pd9ShYXlnjbvKqHszR3Tq8lpdLyUN5dTAJ1Q9LAnfMW+3l0sDvYwfIb12f2OvHwmhFJ+DwKdvL0p
iU41v6sJOaEsR6zh1x6nnFgG6WLeVGb5U8lrDGwAyd2hO5D0Op+Ua5yV142m/0C6qF5NzRwxzj4E
P4uAmX75xniBc/zI4vSnvjphBERITJZ5hfpUHsmVQLTUM8k0lqCV8Udv2HwnDzmjLcTx/7hBRHJu
WeWUkbpK6TUtWTJL4Z2a67lMmBxBizXoDUt/vKD6q8BnYK1brkP/Z0Xiapkc9pXhTvoND6SY9d6z
JB//I7+RoNdr2rHx/8l06r7VR15L4mWNdmd6+uGxc6aEZkEUryTaGxn4q43TZQ3IW9ZyjtEs4CYw
nFxvSfdxKx8iEZAgGEY2uCSPdUTXs5UUPpmFRfBZaM0pUzIsqs9yd+MKXP1AHwW8ounytLzvb/nD
98DQcbuZloVO994ux+TktFq3gblt8UB+CVPhw2iOsyQncVVXrGxfm6wDISqBVVAxQZrrV/NgQ/xi
bGWJ0WETlPvLH+sSP15re2RwO0z6n2FYks34P8ZFLVKeJ2UDOZ9DbNB5j7GxxWeaeGdXcxvLQ9YW
z8b8r00iC2P5k+KesBAYocbYBin3usMxFkFKItg06FI5Ivg4S2GM5QZXxO/teAuQ0VF8MCtWZu9l
dVZM5ZoKVl38pLkCWmxwdJzqzBSNciHqeCfrYBwRx81GxviX/Wf0EIefzN7qnwxEacrZ6yu/ckMT
0v/Wr1y2NpUgLGZagMk0aNqvw2AePiaXhT1hAscq2gX88bxA8s4+6xOl9bAroXRxHR09BGxoh5Wu
wywAO1cTnTZN2nipwshwt1eFQL06kVnq2m1NJqVhR9VGPWfVvNvZCa+v9qCILSFtofHRTvLRd9vR
fcN1TaVRu0uNSOxYD701jcoPnU7s8NPkA+uEWwK6yxYg+OMuRmB0B6TEaUdpK6jOlb+EyFXSoYyJ
stsKPk6RiTm0IAKmTRvtiQ+xpn6wQ1yFjBhCkIgZp7zuBoxisepLMKahdh0x1gC7ToLLsUT7J3I2
92AlgcjaxRbG78sWmy47tW8/tAinyhqq7J/7juO8zCPnQG3nedOW6jaH7y5jjugBlm6k18QHp8mU
atxYoEflmZrdsb200Pl3/4j0kQre2ZWJUAxNUXRwUdrcdY+dTZ15rBLa0ra/jU/EPfX/QV61uNVw
U4kNgir+12z6/ajFrI7YjXJwh5y7JeZqMnwNipiRqpM52yRerm1ispBRRBPe7ToB09BO/dFQ05fB
bgfL51nVyfa6NT5tY5xCqAyz0jkeD9NooVx9X8DbMubdx5EynDI99t0sJ69zDqRpvquDe8ICGw0m
EO2rlP2wTaqJuVr+C8cKcODvrPdDOMDYnU6H1kXfxS4lJ4j7idXxyaLv9bVTKAWZa2A5QB/d3dAh
6ysbG7aCzqHRi/vJ+mAYaoT8vJMoeBxO2SZqZV2OiTtnSFyR6iAPoYEJ/5+B1/SqMAQPX1j7l5cN
XBZ+1/p5br8JatmItQ9/nUqhoF3jxFYQuL8hDAMsFuKNEcQLaKsoQx5OCmpSTQaTHGjt1u+gBOqX
8QLd7kzaKy4mAB8iOsodwUHmT4qgsQjpO+vtdplDfhTSCmdl0TltqINTl/zkn2DyaZqYNMXHKjfS
s5v+b8hGO17YPYNZ3CqAnEuixY0dEkOtDGwFyZyvpkC9UL/a/5r/3vgWCUJpQhRIhPNa5h9wUrx9
PyjMHAfqiWOmHRv2Re6VOUeJsfOiw8jM1xCJu2i7hSoPbvWC4sD3vCBBKzSjMkvyrTyP0r+s195D
F7AMljJSxd7XPdz+Q0IqABAXusq9J8sktHszf7WJHqysNFMptpggD6FzIS0NM6+5socOFBuNsUjw
DKrgtl/TOnCY1uFZQ50Nvfh5Jy3siISA8H4xaezy7sDmrfczTb9vssE/dosMVGaVdiuzD2z1RI3o
XKxozl+euPtx658Yj3ngX42Ja0WPsAERDkmLYglS93qgg4Xb6EZlH1gFs379Tlv5OxZ845Fy8HK5
PxNwakbT42rot7S1W5WgXIf8YrTVu5aSk7cwuhPgsqkes0bFhDPzshHXr8JmKJE24AvFp0kOhofs
Nwz9u95Pt0LU/v5pWv35NqJB7orHGStHguxOzNVwNbVc4q5H9hvjXqNmVFWwNcGABT4huEFxkSHO
S8zGg/aq0o0JstHLSXBykdP7O95E5Kzlcwgku7oBRzcBLUb1OqKWQeHC+pMMa1URgbTTAo1pZZm0
TMKYENU7YleXr+/0HmhSeE1lozcYnCa5iiqc2CK2b+R6Gw0NH+4tDAZEfyPCGhZmFZ6rxO6bAu0j
DNLzaCR5C8bCCFbr5qFlB3fXl5cUV/8pTvMmB/90lbaTH/2SbbXIFi4eRZ18PTJTYCM+k39p3FwY
ARvQDgCinDRrRg6FJzZowN9CA4dq4qD3YBja46QTaU/p1TH4+MsdgEPl4aF2eSqJy4aJD3lx4VnP
+OOKYrT/H+Tip34/1AsD4J5ZJFpHrxxnOzkqsF3LZN7gZKhUwlwxFEWyUCDLnccOxrr2EkAvBpKy
Yj6EjMfoFK4aMZLgjonRI7LNmwS7NNfK0icHTedzyU8ONpY/igufUwIYYxnel22DkObim0HTUUWe
1O0SDLSYnjc9jO5tURCnax2qm6hXBYZxmpv+ppqY9Ghbaiw0kIIEhYU7ZVnrYMB2MYw8EXaBprTJ
H/vAiZjjbv2MGQljmHjmBUaaASO6wwGOr4CS2VwX6fXYiIvFiCzoPlkWiYOG5pZAeuu7K11f/hAH
Ks5Mkv/wgu7ssqGHiXiXI807E6yfoXaRp9TwaQ5ADs4qmxn+YZvmMKj5rUeDphgQL8m4sC7Gk815
msmxZez0AjkswmzsHLCtQzS6hMgNyk99yUxTZtU5tWfUZofZzcRkVVBSnFUgwkPH5BJ51WMU4ppl
dwCRFS8suZ8uKKRaYAlh4mHMz8pCNwMQjKwf9MGO330Hzq1TijZQvvgrDByFmkgMc3zSG+4G31NU
3xgL2wYaJM/PQQaI6wC35TT6cZ4DXZ8baG9TUTz4I3awfzPenrHdo3uvi8Nd5tHNU11mQftw3tD9
Fn9FqEZP/x41ZSObn1t1YhqO+CkxsDdshrka/UtdeXYKQraNtsrweqGZmQ7V1CryeS4uMgbF5HsN
9xCVZy8YpAUJbmG39nZozvwgQRORaehBScQzKHTlqessc5qTnxjfQnqIEP8aYt9GQbJnnBNS9ltd
LzfbuoWAgG6rMpp21wu/WdMeweKgBhwocBKpI3wZuWjuLZUnPAd4oTbpEpGorzK0uWMHCXPdPXJj
Mh8yOKO+KN1mWXLgBQMXgGQPHtscYXeU0vXhFGshIFyO59x6QhELP8u0DwEiiTlcr4rm9On3IpM3
5pxxdu+D/wxwfdXLKIOhDrlqPcEt1eGVNf3VoXLn9O8Gu62IG+LtOkZTt3ylpIE6pKVmV5YGaZmf
ANez4d0feoRfPClm0zy4zhLdGVmUOuPaewj+NPN6qmWbvKefx9eF3AImx7Kg3oDH+katE5ZRaaHQ
020Q6kl6GxLJWQHyp9FJqNp9jXy6M0RTgYKGBP8wv8Eoy16s94v5u1+A7FiQY1JlOSeCyum388gC
s+gsuE2OmEJxUp8BVw3+6eGEwZ5cLSEu0KH1DmF8Q22n5DSoKVbx65NcogEEAZLENfPQ5bV5E/t6
nXWpIHnmB9X4tguWe2dLAVaidlnj939ebuuUeMuAzsAkOAZTqiQ2hBgFwlJilq+ac2hIjcIZEo+r
pY84O/4Sd2wfvPAT9kS5kVH3ktFhhOtgx+GD983K3wcRwAziZbvbP3bgopwo0L7gQGrUF3SM6OEz
vdqH16zg4UCRZpyvbuf8uPlsDwV2Vdg8sahAwydjI2fIZcLUJvVzH9m00O3uXUErVNM9CCTtr91P
HioQpaPgJMBl0VSLANGlmIp56i1pWSYNYCIyYMvm2EU738ZiRbLOu8mZTxP4LI9Lsir7nkPhBYvq
mWpNS4bfKxe31znmUTcjPI8sAqRRMilhw6273UgwZbxdqruUNf3ZQP1jpfOcQ2RAzGiXkguaEIyx
STOJmCBOlg0jVPEWGUWeYCkHbeTz8mTQtpX30RNv5USlQmrP+lnCFimmJ4N8dhRmWAMOYrwd+A29
EPtCSj8AaAToN2cWhgZiFh77kFWpKvh7Ig3mBk+gEn/D9BnRksUS/sTXgHQfi7wYbVPiE5TVPD4L
KbGNnyA0fj9OkYT5rAdmVd1xCz7uCLPz3TRyvPV2l4V2V40WirbxB7NCvQZCX4W+6bssNW7SGTJI
paagaUJWx6KBaKJppQkLVK6kRJGQk6QC+bf66DsnWXBh+ek0c06MVQTaud0uIfTmDHHPwWUMZQtU
Fi9d/bw22lh/GpLQH2Mu9W+OgyRsCfgO8ad96Zs6CnVu0FsjOR26AjldY4brz+X8JIB34PNdgi64
JJlD1oE8/GHJKF5ypDQuJmb2Cyhez3ZD+3L7GR7Q4foSOBtUUxHY4SamkEIb0AKbtYplk3P7G6EQ
y/EqhnFG3rxQ9i6LZv9k/q7PFKLN53ov00k0dqSPQfngVjBgxEeIk/U1cJ6aKmn/x+13bE3DKjni
5Rd0xUBZ22LL0OwVfWmfOiLf5R2bWTHabSyREglzaIOI4he+AzhColbXrIWBwgLRipHTMzCvdsHL
vhFnIhOsVsHlHWXQL0q3oMX6lYIiIbypC3BYRf6LTtsAQx6n3JrlJDze38gtk4CS1dDb52KPuLvf
BZ/djxPUZMDU4i35EFHnHdhsuW13aqwZXsyiT6cxmZEMTWLs/9To6CYBw+qQp+cu92XBbO07LWnt
luCqTR+Vnz27axzBpcdyC874fn5FaYY8trtd+BOS8Hg9QpmkTbQKcAlZ3Dt9olZ+olBzgnRXQC3Z
myL2sy0+/0x3K7ehk5f/5y27E3Hc/8xrwgQs+2cQEU9PkD9ZF2VRextg05sw/0VfwMLTWFtSb7sF
MnWKaSwROz4pfLA/ccztME1a5BAO9XdZ5urGj4vkGmE2mGP0XVKKWnvFwpxSBP1MJt2AImo5YfLf
GB19jWbGGmIYw2a5dOKFDwvzrE5En+RSq4nEZvcdoDF5d0H8kyXjIliu9041xvcJSNoWIL4OCuTN
Ki8xDG4laPegWPVplwncKpkKk3aCH8qjI12gNML93ToSfbZ32PTV3JmsCazbbYGHJLf52aJtyPEj
qJ7lf9OZbaKE4Sef/2xvNUDfNekGKP/4bQ6egSmlvE+eIMyyASQIhERfkvxSfzT+t4ermxfGO5EI
6Rs/QT7SzjXg8I0OiFwiWrfosc4o8EyXxanrb4qTBxCHyiXhd8d4TLaVSeV6Bl5rFI/req8zGs3Z
IBCnxeqUilTHAD3Hjqz4E5hW/d+Qx3jPlmu2CqQUqAaKMaecBGyg0f/7kmHSKSNhkAybNtqkO1ol
9TQO3EJt0bFesRz7oUsZqHcReqBvlSK2DPGzF1mJ2HN5QQ+tAb4Ub86RjQspqELEmxzGIn0eiY1t
v0RnefTIQ+/ge3wfm3a2qtg3VHYj3x8XB6NoaOOsIn/WXgwWXGa1latisV7Tx0I5wr1o/PzmQp7Z
5ujc9pSW4mVtyuOeNqg+9WItFihDg5Qp2RGgR/6IvZGnAwK0ruXOkllCKKaq0JlF7ZfXJuO/WolD
wAmiyMwO+oloVX6KQqruu9fs3cR9XOXrLKVZIsWLn7Xd460Dvj6n42RXfVPIjtDe5rux1SYtcCQh
ITmlW3DYKKTaSOVnBFT7UhVPq5tti4cNEU2y/DUa8zzfyxAC5ugveUZm6CjxMlgaxXbTiiOc+3mY
qR8mTiEUQLnikXiPmnQGwbkc9/24Ua11cZs8W8eSUQVckPcrMy2BBLv/DBrKMW+/oCRuKxMEp/Ye
Ny42pWKrMdRfBGSWLHE/9TlEw6KUuqZmYoPPZgLXnGAvZv45dzJmRjJla4MaqZj0a0aCfYvhNv6M
YPB52KtfuWYV+RELSoMbLPRKyolIJxgEGAvcnq9pn+G7AhjzELeuf/0neJ4FBE7u8qJWIxOeyoEH
iQnlkzXd7jC1BdipsXHcdcoa3JL5gbxfZDhLNaar0RAAv4KXhyZdZxg81NLE+9DBcLi9hUDwqha2
b1djLqbebtgCVLiFAfu4ewf+QSXMQFXEu39Xehjhp33wbN7p9M8zsrBrNGY63XLopLvFqSJmELQj
BDAkTXyCTSreky02ww94p4deZTe99afGFN20BV1tLm9Ct/kMkQTM+k4ckdgUMLYbAmI1+O0ErRXD
euKMRfu+aUinzs2SO9KdOA0h+NmpQHlS/fdpwLKJ/0bX46IEb5izoNOKqNXxXahYT9ypN+AwDuF5
jihJKbUpBq7PrlnEJSTzyyctf9aBMC8+dJnjPAYADcAuH8hRRnBejMlEuPWbd4R3GYu/ADyANZcM
D1DvEB89dB0DzmUWc4stsYtxojRHrbK47ckXvYOYiGUq5ON7Rdi+7lFtNJYrTzO1+0lWM9ZjuXVD
DgZjsw5wZ2gkPnwL486IqzhPV2p5OAT2AOhEzoWdF3g0z/HBV7McuGtodf0wor46WwOqMgiLN98F
zw25IvtSRc+cWkwUjjZ6ymOZhAciP9F6+AZboQqtw8K9U3vHBczGEc8NhUHXjhY7o3ASWRAn0eZZ
Wyr4Hcjs6WspDa5Hwq7JfcttX9wXdSHT63HjRDfffwjMl3pDBuaxeLErfhCeeN5ttTwgqi5g78OC
McAtpk0n9nifxtJw7pHsEy7dTWi3gIFYvOCqqmJHShornYyTlgNX/dMSirWXNlXo5sw7Nbr5ygJ5
V/2l9zHUMWO3FGVjQmjP/HaPT7wJGPpXJHFl3cRS/yJa+7w9eNQN4tdayKek9xiSvHnvoVzRiqB0
61H0XDJQFCDleKgOqYFGfWYwSQGpp8c/9qnx2S81npwZoyT6vu5Fkte5Qma2RIfO113kxGaRlzU+
CqbKodWmsppqfTqQFpYI29H43aqgxfq5FoyxbiJN5qLSvArT+tSKIvBk7Ilo3cakVrsxqYaWo40V
WMWJiJn4kTtZL34ZDXBcWPeVBsmvvc7EsyWCcm0xpCl2GSFYcmYnvXb7FbgTFb/QBi2uxU8mE0px
KOo4lym9Xy17ew6VqmlycNcsBMSOrykfasPH4IM2MmDLzzG1H114ZTVPylmedmm6Zc/5Fzo6DYQK
tShoT53MyvzYq5EnPHXU7diqo0HZzjmMkC4VIWdkUWzVf0bAvU84wRmRrXnpaWfbVCaghCqzS7Hn
L9ZVqI1fjFZFU0vnU4hz9zk5tAzW3YsSYCJv9dQv7Qvak2TjgIgHyoNb1PKFjDX8e+l89jfl0EhC
HAXehofzzpAam6JO5vvqCfbC+v3omRu/fE7Em3F0EDnRgvUxyWj8DEh6i3QGoacUII5S+Ppe2MWy
iF7CTlUADm6SBZ4my2Kgpp7pt8zxo2X5Jduqp7w9P7n3ZTK42VWH6OC/cJq+cfZPhXypl2sLPWx8
7aypUtP2g4m3zOrDVP2Gco0z/1cCtzdRZDn6SvNOCdYRO/pUh939tyrVKcCbMT0tQSQZv2YEuAwz
awUNv7bNJEpj8LWfYnjfOqW751r466Vqj2paeZr/xR7DpFrSqvB8SrqeqDL/tGLFu+PofGtxUj1K
Om73RllZmqblFRenRtZALt/1RrjQdRik0KR/PxjmNU+6kpu72QI/v+2l11MqNgjEwZdrfidTw65W
Mym0URJAs7VRwFkFI17zS4pN1KNYTqRj7zZC0NSLtIOgSK4vitlm/U/JvZata/6VQb6yDyEJ/gbw
MMjy9ZkAeLrQ2MtlqSIrj8gSIRUdj+6BNEUuMGwgU2ATqRLvsbFtNXQlCc+T4lVIwcJis8W+DK5V
jopSEF5jcYXLYbs/XQp8XeWh5e8piNuhEcP/lhSOA7pTsEqxVBVpibZ1tvxaOQDpUq+eDtBUhT9A
iLatmWAMfkz/OmnKJKPrKhOpvu268SVzbbY3arpj6fCIfqV8zAir/Ux9MhF0A8pjtwVGEIszUbhp
YtmqfTs0DvnkaXgCEipB05whI+eZ7euKMDuJ4By3TBP8PYGmmNt4H3KLR627zRAdE1bWzdLX2PNZ
3GpDt7dequ0i80ZpTBhmGa0uGa8C+6gKNEVqU0KE5YsMddK9mhpM/eDcz0gWJSpLY0v7BkQQryqx
t0kW2/8GUp7MxDRhYnSAei79hW7l21cOepsx1zsp99y0T1JEhfz0iJw4QnhprN73a3m0FBDqq4Az
jtEd2cyYDHeMSBzovd48TsetDgQjvPImBKrD4VnGM8eTVZFyHtYmIBt9fhvykbgVMLNmQvvbtzZw
G0aoPZ92EQMQu3vau2tNIg5FuSBUgQnMVHP73NpxImXYcE14bh739+kxnPIqhk+U+APZZw8l0gW6
CXZk/gsdjyc/bOC786NLjRTp8NAcXY2tur3PTWQtCkKBIiH9suYjnjQZFMTWWAJU0y/NQlZPOvOF
KdhxNhgArgIJkVSHb98/US+oTD06otSi5i0rlfAPscdvNSZ1PFCPXQST5vESo9NSan3m+hK/+oRB
drdwV7BR5NZjsrYPslqcncHeiF7kvlSoewxGmj+NID8fB+wdS5a8QrARUyZ2EKfooX+wzigdDMBG
uGHN8+wBrXb7uFRC6yfh0Hir97x2AfnQLEuCaODGctCX6i8jxYJIrIYZByoWfkSD8/h5F8nbDW4I
B9nEFE+HxO1FI1ysQUvkPaksO314KPdOIw4coStqrpyCLkroSbCjjAbbjgqXTEyN45TBC3Y+fbyO
8+w3jPJ8TWYJ0TwwoEvOb7+xpKXO1tKxkrqf8nWncCEJZDCIa2io3exJvVxTWI5qmIj7PrqndEcD
HczRkIBCayejKurKJPEnNEolg0MTGJ3zV6xu27brSzBx7nJT0XuK8c5G5wmn48SwxaUwv0oszTab
uOypACIme1KabmGQeCi+eyRsl2PlZqoYQ0LnW8JQj6urEa8ziRvRSJoAsayH/V9kij41ZB/RpZHd
ePbxCyHdPYyizOKgq70RpQ0749amLc5ETRsxujYvxqLvQUWfvJsSxhIXUbtvW51sCO3sLKVXRF/d
6X4dHOsusvITcyS4z5C9LoUIuiy97uwjNSa5F1hEX8XNPgJWB/uVJNgZiBXKHNd1ED+FXF1E5fU3
jwhaV+Yb8yWYefV6EjKNqpKF7dLk1Xob8KceqPleBKOc6QXMSLRwsEFwupGuTm4J4kQITJtfAntP
v/59TvLqiypxGUKDipBd+/V5gFzCSYahmWYh4ttpDNJ8vcC5OXNbO9brZ0W6RhdY5Q3d1JtJSOGu
X6+6EKRKWnWdCyEnv1IEj/k4S/T4f35J2czIBdRYI1+5RB2PCE/ZsKGmc0hZhii1Sz9BRpa/chrC
0ERyyXcAqGkWjVTTQVZp+hS1PnRWkQaDanRyfQ3xfGzkfr5yd2oWYd4CWKnl0Lg6NVDRlLjen3fo
zacOnWJ9xyVZo+afNNQYgYa/yheBWGCERcEQ7kYT4ZW7tOhiDGbhn6zYcnfZsGlk9FAq8mW3fF9+
KlsSTlaJ8+coIv3lC7U135qxMX8CDNpQHmH/iOEsVm3xdNWDhyPy1/oo9u/A14tAc51W8+HhBqSI
P2dBHkOnMUJkAHbHiEtk52TgVgQiJer/poaDeij+F3nM/c6I1fq40CVGVY7I/2/vJ2Rvka/XWwAV
UL2G58DeX1lC8TMGwES/ZWsrtcTsS9p1vFix9kKxDm8eh02EQ0aQm4MvaKL5Pplv8cilnq+vx9q3
9fVvlKslT0WbOmjwQaTXj5fnhYjiyd/xOZ5daRp4qmpaOqQLF/rnKUoZv1zlbQmNPVkg4yetC9yo
z9MytUFXXoTfWjLSgyeGmGMkBSzs8WLLBFYa0YcgnNyRBVpsjmxDAdD7Z4XCkSBGf6VFqwDxq9uM
gyIazcayO2Ckv5ZKhfaSaRgc+tePRWmB/t5S1KC5SEV1oJnX9UKIOAvSs7G08bnnp3Q3Sfc74ohe
UcfSHiQaevvqqVwnIvhxhFf6Z7FTgka8ivCex29hvLGEIoILSKMpFfF+MfkaQILyG860OS4BJ5Yc
rUioVG8cb6pI3IUp49dBinnvrZmMTAb3Kwp65EjPGxSCAt8tlY+WNHdknyZXYo+kWkTm+EMDZzTX
y8S7ZzrcJn+0cgj7PMzTE9Q6hdeE6JqV7aGVErEWCv3M6QONc8OrsfBQHLJX/bdBxUvrFSXvLIft
F+LGh0fqJrEp6sjqn459OHcmeMBseTZ59GbSVw8DBSTsjAqQAphhw/hqlnFhtx1p2ZryVy+3vJ02
0tGSpWf3j2JVYxnnhXO0/sXOau34CgrxMhWpsXZoctht8eYVfKY34TQBTc9z0TzX0ipLA0SL7wzE
naJUNCDJI8qb7md5ItbPYtq2bMZaeb6kHlwwhq01G+ZL3z/YFRjlU1OrhH+ZoUgzFyPMTDBVhdW3
blxNOLzqBqpvSckXafDjIXmApyMdroNe4iO0QYKUwGzVWU1C8tNqP6d9TFPzJDajtKB1NpxcBwCr
fnR5wdGAeO5pHIwMz5BpUvOo4HgNlmcuVgkLng/MybWsr7PgBRXIq0gyFez0czUWPZr7l4XtMIGV
AJRrtlavTjqTz44LW6A0OEzHXakXT0BCYhhZbD755f/gawJL1sT08UfQlDcULT+T4qdL+JKtVm9t
dV+IzZ9xTQTtj1UYEEcRDHk5RD0rRz/eYCl+G8M+ff2RtAop4DrLYFFvSomqBpxUPS5SgYEzMxwU
3QnWJZsbCd8WkXPeWZVIVuLBsY6l1/HcQZ9t2nfzzTkJoUSlBy0ax08HyiQ1WgIn4JdDJVw0zekN
vKFlxGSb6VOaEx0KYvDUO1e9LNvwejCYT30V0vBVnxtpPq9OaVVN3Uox7pwFCf1ef/Ht55ARKh5v
qZPdGlr+eJ1gRqjoAwBr3hSiUrjKZy/tDI++8f9FEKBlzR77myPw0ZvUCG7WCuMR/aCTzz8RcKc3
bVrPrfD9tMytX2FvsZwSztbuDvyuBAn7xRyhlyk+D3N7GcvaeuzpKctzFZBIEsQua49EQChFOn5J
miGKkNgJMgjqe54lEztzHPnG+XliPGOvo7nmTPvPTyNmyfa1515D4FrHtDnYaHVMMTlFkjOOEiYe
rL4f7sS/REDOw87YWpxmpCsEDYy2+Yglc4LZXNNeyOSTl9peazhwue+Osd1uwhkLydM7tWjMo6uV
tDb/nq9JlWEbO8r/Ua6u1fIo6cJNtJzkcrs6ixUAkUuqOq9A3deBXJ4HjwZ6/6Ofc81FQn6EcqQ1
Q/6vK2oRxg9bcu1sPe+hyl7oDJv64nlEsRHq7m4tcJpKb4J1H/VuW06rAg56vucbpwoYVaBG1IYS
zQO8h5NflDVOjvJ/EuUpOv48pkClCNPTLutKmPPz06glJ2p6nZEYuNSrofDFbbK7UIPlXHaPKQsF
D4GBtsEfc3ftRAMxYQ7/1yDQR+dAQvnJ8pPk8f0RPlXz/aEDzigJOZ74+bPYyjez/L7oK/k3y+wQ
b2cV/MLXeZhxgfiJuhrpEFPYbwINUyB0CumGRTgNZcjb+m0hO8GxJCZ4QmeFwiSSBwKCmXKdd4kv
XMWThfWTfuzHJ2jWu2uisvfjz6xrc3TzkdPq5OvTaMKxp7A+Q94atw9ASW932yvPu8zqIoR9l4xn
5UjQXliw5bbp/Agfs6R4JAoRvL35QCJDA8s9Edqem3aJxG2tRRy8mGwcspyffBUI9vNbMmJ8BhLV
92mvdIdfCBpbTONAQM4bv0jk1M9BBU/rfhDI6C4LAyr8g5DwbET/tU0rcHv0Axhg0cwK5cY43RJk
F52QDIYeIVMHNN5u6f15a/k1+MLgqCP4OxwFGoSmSvcXClqcsR2q6925g5Dpp9Msmw8uJiidmttV
h1/4nqxBfDeReDg/f/CgAoCbIjFphTls6YJOTmZuQmLiKTDwVASMrK4zQolZ3NYLGT6BpZRsfX9j
LJJSzSVaaVGLj+ANr4t6IjSDXYYS7gxwxn5NniXL+IApHq9qro+HUEXFYYH/86GB9WvFL/eVXJUS
PoEFUjBYp+cVMinUwqHxPfp61DPI9j2dlhsaaR+qdCqXG0RPqywlRSg7wkZpqQBTaIcCzkI8L654
sI9cFmAFXAjrM2v9BDBDzjKX0tEuI2TXvZCrXbw7hicEx/q9+jQN7jyVzU6iQ6hSRdDfCXinFicq
uS4Jmxxl++S7da52nU38SzvS1tqrtv177qKefSo4MF39ny9YWBvaq2ljjgnaZh1slMnNjIWgF3B/
xRLgv9gjKF/diV+zCSs4zSzuCd1tOMcyFtjx5A1Kv9DafAB6KEDPsCXgJ4Ssm2UNOepEwn/Y3AI1
Q8E25roEdaJscfhdb3SvR1hTizkiPZ5HvrUbptwY0eCjmLghV7ASqrf5zIFxOc+RRz1dHWB6SwC2
wOplHFkFVyWcII+T1lx3yQBgPyC+3NjscLvylX194TzoPTeuLJkzRR7hhjzrS6qRaZrKmpatZ6B6
A8T95T9tuKUWN2XAi0ELM9iRaRU+76jDaJFmj9yQQoLL5CgUkFIAhtqMK1yBrHbIcFhUpduakK6G
r3oZlH30WW3JUzBdCwKCmNE7lLWbFgBcBvnFiXF8gxuZQSIIJlBKfBBmsR1+M3skUvkvSD9MLnUC
s+Lr15FZnRdezubKiHJYtx6j5hem+bfY3k+6dnaelZbKRirmz7Ho7wu3wkKYd9kMBKIC2H2d+3r6
DOl1EhWPk6h1kaRhUgzTkvu6+IgNAvDmU9YbNArbuIBqNt1o07UwVPM2xcDG5d777n/fiVYU6EX0
FVHxawpVwoVqwr8ORNBE4nIqdieDKJqKSKNsdTCSbbmCpom0QA/ia+Zw7A7mCLhD0+LUqxqnX1Vd
nivVGAm19s0/CIZoL6IXrOupzlNPCeF9yDJ2Q/N3f4HjJUdoSQ8LEUCi5SUk/oHc/bFL7kZ/5icW
y3gMFUIFf94qfRQcrTNn62cnb/EJp5vn2/ARP2IdqB5AWIJIvJhdD0moDpJKlV917Lrfd76d1eHA
a2exyzFIQxSBiD+i3gHLwE1ZOYYx64x4QbZw/jb68zIE94jwY1uUkru157GyVeOefHjg5ERDixZf
VAoYAG4RYpwIhM+t0+6pXi86RYEPTV8T3GT5DLKHmvrScejOZ7rYYuD4VTrIYwyeR7itV0PSru4j
IG5BCaO7pgcYSP6R7LSEcRtD2BmeoSxm1eLFxz/JfPPyB8U25iDizrUqfRZhqFqeKOsUzA7KrJej
/95LwxUiL7wT/9krEQGVxLaZohYJGlmPIGWz++VGVm3FymubTO4RKeKsQrihonf3rgLH3MUYHlEH
vLO1wdxPpAArexUdDl3bSirb1F2gRbP9rH4t6FUhm8JJMRvKdpqH5BESEpxvD+VbZYodevxwWQJx
KhFbjTAMWu5uXgwoIoTMXNsd1jKcv6xXCrXDW1uQFb0+6BdbsFdHXgicjdjonU3v5DDvECMlWMzE
pfdncexgk9JulS2XVOuVW7OaKLyTvz6mqNr1Hk2+fdwY7PeZe2Qc+SJlvmEeEUzoz3HkpzIrbMBB
0Iz508eoSGpgvmrzepnvXvDETG6fRK6UfonLkGHMv6LAcLIRVUKT+KKubyKbsLG7E3u3ix1pAFAY
Ugm+5JTN4spek+P53LLxvXqv5RM0pH3j22iDvP3NklhSiueIT5hmBHiAwTAz5WJHBb/E709QGFcE
VKwHB1/UQVmT+09CWgpz9eEcig2i8OA5LpXRT5f5h8gXjeUW/mktkJ1hpXxeUG/lN8cdNKiFJGJZ
qjqQ/lHW1K/jOmyIYifmw9eHRe+mcN+X4h8d98lvfdQFHVyCC9MRCx0ikHQsImiv4WKXtdATRPG6
f7ZWFpvYNM2lv28CAkMTYfcZZ0hbWgxaRA8KKlrwVth6DkGRdQy1EPD7ThKaiY8NP+kh5sV4/dlD
zNNnVxNwyTtnW6wHWLV2aBXrPuEHbGTNTuIBo2cvU/mdo6JxLB+Ef0PJ/ssKGOnikLToN0sd6onh
fH9pCnf9QJksQ3hpz5xJ7K/sXB5AwaBNBQUZI5ObIBGJysuFcoUyM40SJq9x3Mscpx5Mp/WVdTdl
jPtOBt8VQOGt3DjtXKlH1oyRHRRi6WmbD03CA7+eN9BxVzqTF42H95fOE3dbw4vwZ9RBHcvcEyrP
48cAuYAm1dmg4FJXcbWexjIyoMNHhtjriFYs6aBrk7SDNdg9I+WUJrTdEdpJTIslkOqzJSXJJHk2
CgpyNoEiCpLeROK4ojXbZAIJ8Jw5Chn8oXLYPBuihJ8oOjyoQv/IG50oXcVV63PG9fz/8icdsXtH
r67UiiDtvCFTHllnoOfyN1kkUS2v0nl1Xk63WGOWEIp1wSY+FW82jhC7YFc2X2AUUbRrATcG6fS5
kWnDE1Mpwir9iTrpk3nFjNqfKdA2cwm/bWPGjx9+E2rMyZAAclvwjXHxziX1/OVilBsUbSbVeBMk
xKnP3UObSQKYJFJYCPnWqRcT4exJmRIHD2Lt0ChlvATPNA5dWhC6Hd+g98CnV+rMfy6DeU4K1x+J
V7LeBrdyUZINwqC08i1hgKl9YkyisS89WdTziurQg/gjsFhjN9h4LjRu4HByifMnmEVy59YRTjl6
EwWQmgdNdxkKzPPn7/g8yVKwxIFv0LzYf10tEplgiH8RP0qSfbWNfPwcUXyh6WJI4/RpKnYSVRE5
X8NQFM1KMxvpk3EQCGm+FS2mHYIvaVR5QOhOasw7TqjwpdSECwGoc3G8GORbCFQx1n7KL9R3HA1y
BwxtoGjcTZS/Y8yxMsvb+oPXB3MHgNqqWc2w5uvtG6r7DIh+tKrakIUVjwy2kgYN1PGjoxYXfEiL
SXVYoM0AnGDQFPtXZg9vxUKyWOF7HHUuxnok1uoBza9Eby1B/Jf3Nj9wkwQV6GscDmxB8x8VJZpg
Gh9CxYDIFG2N7vgXuPzt06y4kLnLqexWrKDaaJMeti4y72zJtsSZbu1AdOo3D3c1o9QzPfb6z128
j3CWi/L0N4RaA0u7OdfHpNexBe1mXhmZukBXiv52oOp0if8hA/MgSwdwVlqTo83eI8m1hf0PkERF
jbNM2UTf4TSsPNDexcnHRhhZ0HCTu81qJuN1hY3WD8AIAp1+HXgCxiHjxRCtVD1apAJ84lw7E/3u
U0i9KnlXU/ojLTTVAZhWHypc984pBn7f2CLoLZHwrrvaOvxDdYOZjmimJIvjJhJdOw/ds/enV5A9
bM+EvNi67AvcPM6dkhAC08PeEBKA1wG07PLhq8s7pbEtzIlWz06X3E2yzd2IGZdo/wjpN+BKjqYx
fy/yt5Me3ocaGA2jhkiqG2dTD05Vg0o7WoFKtCe+tb02qMfeRobwZxkosJ+kGjsASiqrl9+jwjH9
l1S94noZhjYYEqn6Fs5rQ6jNMQc38FvkmdnYyWo5DX0bcmPu7Lyx+u07dMOu+wLAR1ZItJx54fa9
J7NpFHyR6X3FLPQC3gT/oeLtlENUx30ujVL/g2buhJh52Te39Jr+uQW8sgyYdIPJsHfpsTgMlemB
KCbSWQNwSWT0TUCEdOwS4VyimRmvfAZYoeRRRzgLcfkeU4K4D3khw/Pzppd8GZ1W0wF+BVG5hMPV
pedoxdC8H9URZ0A2RCsKe/SXINOtoAxHTe3Bmv42nFrQgVxSP/H3OMOayvU0cLpx0WZcftTpyxpl
fC12OpmUxguYv7Lsj5Il2ytV5pngQpP8L119DLS4ZmIoepGC+Y2VxYJraWsdLrLu7r8DBkadC10C
zC73VcmDNJQh5IfrNvRdewWTOz/L+hNBj2OmeVM+qABrkkQ8OjB5JPAIYmSUI82jR5CqQPHCHgtM
10zxzJU5kcPZ73IhtrXgEoxHA92KxhLF31vvSbFTsA56cw1jghRzVg17oNtvujWXoWA7zdzJaFWx
KvKvbQvGYY4zxmwcn2/m/Ew1efbvEj1xeM279aVZxX/AzVTdOfMi9/yqvacx/9JB9zJA4Ik44grn
X1iR6dw4c119iBh9kfNqb7d42nyx8IzCbkFjNluwbKja9h2LGXot//qaU8qZ5aeig+G26lhjBiMe
LIVn/dyINIasFHbzUcu6vmUCNEWABFsvRQa2kUlwbLROMG7nUmoQJflV/S5P1WsUvNaTbVUsPJ8m
u4uUakFqKKqq+lk3aKdnmlJTATwaLBR/SzaDC7uvV9gybaNz0oQJgJd6Gowk0w1A2SrIUGlJFEXl
GAHu4f2q+NbEUhmm5JfbVravZjleoPBHzA7J+8NG4EWwvGyFJ1qF4U/Hm4IqvSLL3yjtv74orVXM
cC8B8L7C45TNm0AU/Tq+dCXVotQLLXa/DT3HU5fRphgcIVBZktlVhcZ8aJS9ZbSpOVa5F9jmJxoO
cHpE2zKiurxVJZmD6694X6XFYLj4aS72kuHFXJsi98xl+f3ePSxHKB+NFsoqCY9umjfs4qc8AHlT
xXuj/T0ZiWGOqRPsmgAZifcg97Q3suXazKvuBUfrWA2XiGjAkTei5r4ti4eZltozFM7riZ/WFowb
UJasCFkS6XlS31jcjN1Zeso076kkcjkBwwQxGcoz4ydKmvVeep/SK4NA5bf28wGxsxQ8xHHrPzxj
+Il+aMKX9oibJXFfsclYtJ+cYG5VO1WuELNv+RNeQg1eenUwYAqjepnER7FOUwMK4XTMaerHZf2j
TxanTzy2mNl8PsAzauqTbAyMeE0Bvoph1uzIdXYnUOAVPGnZHYaCtRRWKECsjiO6yMy3NBXYATx4
FtUhz/Y+C7iUzoFb0n+cwktzMS1G3AixDGQQz2+vfv7O/h7oMO5O4J2ZI8lR4MCA3JcgOuXvAzPf
Tc8+qMp1/kozd1pkHvPvwCVyUVCILP+tZlMOGQWf53eYEhvhzTDevnavw0YokMn7CrboIgxdGCyl
rR7NLCjIiyTIjIbdR1MyvqjA1EtHcyhP84xLR/DIj3s+/FoqmNYX8VplFCQ9tR6228OFfLWjk9gB
p7d3izSn7emZKu2aFaTyqadGR4JCTb3T+lZmiWp3w0Uk7e3q7lq2/hsgrp2xgtLgls8eQQp7xwio
8+H/wpcMfqbKbBt+tpzsuS9MVM1HRVMUDpRdUWol9z+R+KZ2yqx41pxSe4BuYWmCj6xF//e29MXP
FRiSw22MHSTrq3YnVsi2kZXij5c6/v6yJjERtzdYmhXmvrV1J5ET62a7Ye/J5iBZDSiUpj0+nKR8
JAmmzNV+g6XJjN5G6LcZSJlOtq4WRqs4wXRkPtO3Cah88oVd260pTu0izhTw6CyHUu2n3AX9i4vD
98uZWtuWDxbi0Ipa5bymym8SKgcgrDBGPRsIShwb39AmBaCikKBr7yInQrVrQu7ppk8KIsvPL26Z
MFgXo2r1RL9whvILAaDvYfdd0EJmYeA9NBfDq4wIki/TOWb8AFHlQXIDZfYRi61at8uso31uyMtM
clNIhy7ibJShj25hHvzxAizGp4qHdwcNxgRvCu8Io5eOiU4NEZSVB2XB+tvyMCJfpCcs5z2L17zl
EmPtApwlgqKg5WEo5wgpIQAjXcOSl4Xy7Fnr9ly1RqDrWWQGvDWs8j7t4Ds4b0efdfmJpW+raL0y
CcZp/pj5XARCBxBaP08K5nI41FKmBvx/7PbUZOEnpQf/HZsrxCHOUu8EHkf1leReqUQ+Jqsc4FVc
OCXK57wRFf8cPjYeeDNU0gu/leIdpnOJI16/vc/RqSusqV8bWyoFImVtQsRSV082/O7afoX0rXMG
pefkgx+a74W1TDEgH2eZ3hl3PPEziDhpii814UaOVHR+IwQoKpdbsoitHdxwT+oHzL6qdEKU6B0O
Xfj+YPTki4noicyhiBMJ2Wyw26w5JpGPfSSDTRLOx1Ut+fT0oLDWRUJQjiCVI/e45OOG6BPCedrM
tDl5pW9CNvvAWY1NqLnrDOOoL0xUktld1Qi4qTyjiFcJ421Bu/E7qprY6/tVlaOxVEAZ1E6S5FuY
o3ZGyupNkjQA3k41oyT8FD0/OoTFOtI9rGKYcTz01XUszF744Wtbu8jiX2Gh7pIlpxTydLZk+2+7
EXxewU//8nj7gTytrVNUWafGZCxFfKQTLR21Y9OBInlgcMuIqEiotV9D8kOVX9eddwYK6PWFSJUO
+XnIstcv7tDreOKY/0pmy0+vNohn6Ahj7L3zSOkvduBfxYwfq69tdE48AH8mbupYNxJJfFHhEvJG
Vnhxx7TZX5a6JNwMRn++gVvpPdEi0CmZVQulL3QW4hmeHgCIz+dVdvzYzoOa1ajnHdB1oo1SnTVR
Hd6OtXH3/Cjk4Co3NrcyeoQl5Q9jOVhCRQuFxhVfIjRXknwRtxPIb1Ug+QCcAqtYHXuaulSOjwnG
wRrowpLAM37LYA1fa5xfyAqQIMZg+lwe76HBFC5k7+TyZxAzXISZRRGteE9t6p+L84FNCegptowI
wd7wMvMN1s9iicSFq6W/K5/hhC2FPeQ03GKZCucXVAAXflsGPQPj72w1lxtw3QpnZyPjnCfnXIX5
OYYs0Md9bPtQAK3rYwSokBLmySaFmWKhYqJWM6i/VJaLUeZnL2kCdoKw/SoXOL8GCY/T5AZCqDAn
Jn1ztwlLP64Mb5ZNJIwM5ANRzTJrcZFb+t0n1UpSzUwFN9qpNXfJaYFud6J1OUrozmt7UfljKi/g
KTL8YM09bfwIYbJhcM2NGWF39MLLRJ6od1/NfCZkA7HFAcVbVShDeH5TawQxtg6iZ7VmPcXB2Jdc
YJoFKdsrQl7myuEB9ktk5Xk8+0GDq1muDevsd5jH4G2lU3mwYbvM7SkBkpOcNX7Di/RZAzWWWm3t
JmXatBpKyUlCT9oYKuvj8G1eO9kI69yxXfZwcjPFEbgAYjgTTXRs+i59DWwtGTmusNfj7f1DiGFG
1zH4yYEDM6fEn/IYEWbLGWGq0XM9VPIdrU1WjiyXyIhgXGzyy4UYwOHnli5I7W/RZI07U66zcjfW
IWu2o+l5z5kPGMJR88/eVtYm/JcGJa+X2Qv6sAOZpYj/YB8Ie0xbLDK/Y3LYGLaqj9rfrZadO32a
Vxr+k2S80xPup0zm6rj63casQHPy9bP8xcDWxBLa5GJHfvRfUQ+Ue+6MqI4B/nyRS8gOFm+8Hxd0
iTXUCCR2pwyGfXgX6j9zmgFHaZTs6zn0AQLY3f2iG5t2BlBQzZv18T9IWrFAOcDvU/qz8X0QEzLF
rqgaqI41XwfkygKJBa7riYTI4a3tTvPGTU8R7U0wos/XfD5dHOUCEO+drnMSBRC9JekEUOclamgq
Sq9g2MOTwi8LELmZNOQNW4K57QOsFN/LITA0r+HFb1u1E0gCVVt8wbEzjmntpntBd9aV3VSXg5gk
tc3eYJBmEGtSfXiF3zVrIBAkvgmOC0TYR4Ca9z6zX8QCTXD/jY/ksRYpXb2ndFQyG5lZIf6jgTwx
GTLTRO6tpYWiV1ALB/JWihLSgeCjqJeKZzcQWp/79TMNTr9oFnT1VNfRAZ5KeR1atsvARO6cdb5S
CdLX4wo9o/BfvpYCHUdah1a18sW9FWG4xiSld6lp4gmjcC3GGTB1HVLddgo4cDLViWhQtIeo6jyt
2TdiAQC7dUUrMT3jJ9d91pgRAih8eLOKgWirEC8Mjkx7adrXYfhFmMFbd9iuIFkCx6ux72YfnYGu
iTSOTaVrcfyyE4Pg045ua/1zBP2TZuNnYGq6+khUhIRE6zlfoqzyYtK15wFqS7CDoOfbEX0o8+bo
I+Bk+GJG/09LfGUEC1aozm89jlFcRnTa6nchJF+Y3ZP9vSJ9YsyHAxlaUjziwdDzZoyFDtrfrm9M
QqF7cTn451vfWSe6vd83GG9tq8b/Avj6VgSYkDPAc39McC/utguLkAMZnNQuDhw4MEnMrBPb/2zM
OKH+Ob8P1t9rzHekryWjggB44EAB+32oXVQVZ0d7mYdWaAsI0Ig+MORM82ztNYYiCsmDzsNgpgLq
hc9e++JasMhXSnUsdLhEXPKRV2Hpq0vYG484b9CdgyM3U4X1HYQQ8TT5KW/RO1505LRgX4NCpYMV
7CxE1DEmGOyO/3RFQK+t+tmLRYIbfpRJViLnn2BDHAspe2kBNNaWIP1bHC8+aHY7SQJqO8BBD0tq
rljRjlcFBvTk3sOfm/4SlC4mb+5tnudWVsEj/5W8lXHMVmaffBaYJmX0zlHgqrxn5WSHk2/Cza5k
fNaKn130PGnsaL7XvF8u82md0L0gxW6FHKgpWGESs6gYkkHdRT0UhjvNXNwC2EK2yOK91yfjGOTM
6gt+OtKqvHq2UMXSOLrZ3bch2RKLBsVjbwrfkQls5Nc9Jxwp/FmPJ/SqKGhy55EP11WEWWVqm2mQ
nm/QctpeHVgVT5SLzsHA5fsHsotYmw+e8CBEp+kXTn8HYNrsPc+ZdrdgyL9NLClIsz7udnJ27Ecj
V5C5e6mex079cWUzO+PRmV+7OTXtBI/BvAiUGaG8aHa92zv3hA1GRLjH9OWGWWLTTX1d1cqnuVdr
UeokW+MOE1cVr2GuunR1T9e7oIOKqwwwWgXUh/ez70j9U1+CcnuMxNVB0r+os691Vqud2ABjhWOC
LTPztHLHz0SBYvpJeK+6/vFDV0PxsyBPsquQbd465s8oXsLTpqAw/CElr429xc+FOxozqkzj8rp8
XWuta8ZnA24hhnyrZlnwYSxbOEJzOdOZTuvGHDXQhdG/UxqEWFR0q/Y9psXVpVWRJnq1nPirFdy3
YHcIgY0SDNyivo2FEP5D9pX7llfXnTvRJT8rFlJ5QVFZYwY6lnBq9QlYAnjPWfFVasup73P+vYZ2
wNDhhrjpACzMihkXGSd24V/9DMVzYR2dg3vMOzyFg5ML+AP2Z/UVfJIj9cT4qAMrROe0aUwu8fPd
Uy1Q0B4kxqGyGk96HzqjlRcCv4i623YemX4T1gBl5CSFMX7bEhqQ/dL95C0nA1FroPB8wfHqkuTh
ZZ2GMfRvuTMXB1Zt1VljsQcD7fjOcK51Hme29wIecg1wKngUKp8ugv3Dvs4dDXM0TTR2LDo/XEzD
I2Tfelk7mrMAmHZfF05NlBhAVnIqE8C8BCowzN0VZ1WEdUVPcdJ7mQjgeFraEAec7TS5/zMbT9Lo
tgjTZnhyevlWlXT2u0gNt12pvK4THCWr9qvLpFEeDYqNvdj8KyCXYb1OhlxfmIefuDKEIXiKi3Hq
FQnrKjmbCkhUrNRQESHbgdPCtuHfugATnCbajIi+V67fOSnvJ2beJzscvBLmCKJlIPjVko1vhQxE
/pfJyzV5Wfq+NqzifpJk1aq4cqkYdkwfo8p/t86hI4tnYjwydcOFjK9Uimv/iNmRH57qzT7y8prL
pOjRLcCQW2iPln0FptJySNK72brQNzr/ou7fy8MWy740JqzXQf8Duq0xV38BENO5p9iBxTIujbsm
Otjs+vPNtCdnOkH1P7UcTSNlQLyaKZWRCiP0dxvHkXfX7837kXFzWD/ds6ey2POiaCFBnMWmkOvB
6RjSgl2L9jtimgmgRMR9Je3XzKUfcQ+CWlIvo7qiKpUufmwOF7A69o7h24Iyz2/1TZdxNlftgB93
YYuHZEQyIyeNJli7OYV4pMO/CBQDF4Xx370segMdnWSsQsYuejyEwNsp0GJJmTzdicg/O1Hn7aO0
xmRXrt47JG2w5GfXUPGhletmJoaVDnkhC+0EWFL47nxEsx7wgsosw5J3RYvqou+S56R9CD/0nB+3
Jl4jNc3MONbTuV661B1FKwJOs/QoIN3FNXJXuK35/slaCOoK7KvAGwyZ/T4uodpVQ/OGjADMHS3s
3jP91X4Y74SCbL924i+l1o1mrPFjPNmh7WAG/iOraMHf+Xgc+23RVHbEh4CX3eTu/UuUDeOhDCCZ
PM8Cn5pKZTLPupcPXhCDFr495LdGRm8Z+oVUr7i0v0vovRQPpPmi5NAOWuSWOrPbSAUBNTQCPxEr
Z+9euDbOYggdN6cOvo5ehD0yi9iE75OuL68BSCqQo+rEY801pyeRMMJSk4HGhWM0BaO4aO+GQ+cl
tnkuEd1A1nkr0BqpOlC0wf1z4871poIsz6KI6d+1vwD7k9h5jZgOjW5n5Ml6gS0afnrrbC7ulJWl
+JAPEXoHndlmMJLooWzYjTQu+/2TOekPwNL6cMA0vpEmaOLrjyQi8umRqGL+tshADm/TD1vuE/zQ
7IjemDfHhE7lZKjz/4RsKcmgoLd1q2q9EmIxkO+nf142smHxEtkqqtyjOZ+gsL+CcRQ+AE2HKq41
SeQYjacT3jzTEfndgiJPHPRqWFTTALTF4d88o9Zh8sBpT/T9yhPGmsjoTPhlJWgxClgGzM/vzXIF
6G+uFsAPf/JwvCzGZqbQ544FQQ5xLtaZo3F0qvfTRY1CtlrathSqhBsSVy6m9QEbJa9hLpQPZeVM
RfhktUs1+heRqISbUhMuyjlxx/dy6Hsm0uGTMhWo1AUjoyWFCG4zESlLepH6U8KxpProxbX0LlN+
wLwvTqXe42YsmMgWIK55WM+2z4uwXaotCopn/8HazsyTF8x6ATUuJvbEfOmuYcjAMce9FjWjx6sT
QNjZAKtsaO2hlCSYE+SVV02kd75Xi7oMYs1OzVt57zlY3lahRKNGIJY4Hfu18sUWSYNrAfW5oM+K
j82YnMlBkYMAusXo5ZRaynVr4aika+nbam1v+6gakuLCG5GGUknHNCCTd8djuvLpEllkDbZEaROP
Wbx9hwzyAQBAmrPzxELr6BXR4XzvFJr5P3Upz+pfvz09QizFGEdNQM2NfzzTW/CqOkV8zj6gOlYQ
1L1L/aFsNUwIJCcfO35V7njn+iRqHZkPrm5PmWHG9iheDsOOaYQC4kq55eZfhjxAa0M+YS+OYoBC
A6V77QzoFBehsk4B0NitStD6ePIN7+nShuUww8bdFcu9rYxKoTkP3huIDI/pjNwEAWpKu+mOPDwF
RdaqcES54OuKAwuue+Xi+GE7UG9UDqO3dS8zF+SK0SWrWw5TZIPS6kY4ZLyLGtd981F9uPjJGhYq
so85Ao0zNA2hR6YSo+4ulnt1ph9/+6iha3LQwnX8oK+mi2b05lJe2+PmscemZ5e35bI5HR8OFLXJ
BjHiYTTsJjCX3IGCxRG3yAXpx7/NiZ5c5DqyVhFLDBu2Mv6Kl0x0TyUmsI66u+UBU3NSEMRmQSks
yRAnG4XTUtJuIwZgWWJZLH5OjaHXmLEkZew+PS87mKXk4zLamQP1uRVxMRtId9nFPjWFGMwdO26y
HXIAImbpSLohMTRiXzDpS2Wb2yHza3FQF2cfRM7udDNTVkdPz8TpvTRaRneO8glI73EyktwL+TLD
pGkyks+2SbneroIqVySBYnnoOHrCtZYV8flE5XPWM3sldfV8zoYcIzU/z20oeqP5Sqb7/PCDRlGz
lEBt5gwqMUn7OtzE1105SZbr+FeSynT2lFRycceC0WgnvEMfSn4UI/2DQJQF9G5wn4mD3e6oEvhd
uv7Zp8gknc0w0ZO4bGXed+uofkdU/mMD6anWbL61RLgmMgy5cVlhBPXr9U3oWReu26XLlUl5K3Tu
KV/VN1SYl4WKQ72RMrZ/jLO1xLpEF+Ca0zXhNA7idIF+XTXe1CtFJ15VX4AII0YE3Ad0l1rzOwKf
lc28zKzrhomObdddoqwrgHiJ4UzWtl4IXhk9sBquksIFu5k6vZm+ZaDzvNsfNfNIXIFu3b6beddq
5tJcbYMptGT+DafXuXNCVyGEkaA5YIMap5/IFnD2d8wmr7kBgRnd1OyFOu9MGtE7QNGUyJFtuvAR
Rkd+cK8A6SLv8RlI1JI+MJ3b93pEQIn7ZqMJrPUFOUP//lQ7YmQB394itNTT9tuwJ5eXpr56d5b+
CCnn+9gMFHonIgMEvPByMz7tZPYW7GS4evK3THKDt13FuPf6VzIO3BGZ5ZhOE6audNLqz0x+9UNp
FzDHTARRBO52VyD66NWhC+9GnihBQ2uvdVGHCurmcXrb5NnLBD2Ey9qyOQrsJRCQxUXa5vEVuE1M
p7K4btVyKRVQLj64UmdWO+9giZ3VjOpChXxK8yLFyTt+sSQDqKC3Dji3d2aO9U2xCbaGj5kO0nEz
UsUSsTL1hitlwPGgJbIOlC6TE4q43uFAwledolXhUSvadBXfxFamN6Tej1of8usmPOJMtSsG0+db
g2za5SuLjNe1l3wWtj/KMyMqzZp89GAAW/7JXplICHu/2qeQo9RyV0n5zY7vxXOjxa/IXFoaNcwu
ebT7226cfEDA1/U3ZY7008rMyq590y0yYoMjvPi7giOCkM0C5oiQ6akDyEypy2wQDgG5yHlU8lHC
htsXz0r5g4f46SWTGNZ/CMNE1Etf7GCT3zE1Ry0vlkwMXGao/gD0VIC70S+9cpNrzgPGOW/mXNcC
6g34uQexeKxnAPjhbwq++IOnXKPRr1f0bAn6WBphXXnCeIvuROhw7ThLdWTFhU4x5vqkUfZ8fC/U
WTd4zhZEfzXOw/cmBKCDzgGbcC9KkdqglWQhhUkwrvbbZ29aZvqBZ7vdv1vRrwUe5uqhqHte/TIt
C73uNyKX8rCkR4b2BOf5xhqoiGJQK1YT1xMyjESfYVYOcetiqYPA+RkUfa1RPh4oaqmPNscc/fkN
/5PJgtWEdf8glNyT2a+rdxSSLxMXN8tQvLBg9TwuFyxJQJqqvG1P/KDXDU7SGw8n+xpc3zc+1LOo
ld/X/IDNWnY/727hiO8XG0ecCcdkr1MugqLd8gxJkWMmSHUf5Iq/rPBzuBO2h6KbZH3COKaWr5si
kpLSCPQXA0tD1gL8+A/Twb48I7ga03NN8Rc7B8if9zDNFrLtebWx7Ovbdme0dsfNhNOXBwEbrhkm
oqA7j62gldoEdCqaVgrVZjILLK9jw4hpvZOJzHYXBdaXW+btayFdbU64tV7YKDSP3C+afENTVPoG
+cL59XYkpTQqn0XMTKPYkXBdQJhVOIm++uOcqYTWIRGa/vPaPEhhswmsWkdXa4HIjdo4MkLuSuyZ
M9G5ljLq+BxnpUWKbGkpWn1Mf5RFIwKBXvdRRhbWtjob7XYxE3KOhdFibSgNyYjDiR3KP7psol7c
gyB94hDKjhkp8xcL/6RfA5hQYA/ru7vy6HlBIDtZX7vVEGDCB0gayAUe32T1c9QqmcbAk4Ygt2Uu
PDzHE+LspH8wkUvyceHXINgIM60WJQ0Mt4ysIN3bwdnNP9DqzU0AmCUHspDyOHF8tUKQfpkMjX/N
bmhxrXvRKLUAjLlmP2az1EBqWvSkS8Gco9Bgat0KaUfLulCxV9a+U0+uK45Mvu9udeZqtQiI4/uf
IwuVOTWpscZeUfUWWYXYUkyiXIH7ojIjEGxidcC0TNXDgg08/XH42+Bn9Kf2WRnQnx7Q/sW4ezmt
wKMQr6rtU9F39p0sK+FcQl9qyIkW3UrWA59Qvb197eX2toYHGDolvsasjIlzi3AJzdlLf/s0M2fj
f9pi9BSkEqvb0ugkiG2BUOjdHsGCqVJiW3g8xs5eqmC9GjcHrOZa9oxxLfiYyjzZVCFQ/S4p81aC
KQ9o17HvSRCaPxJKEiIBZ2PltqLwzL82/pnKWv6hHwgGIA4hLpC35j+niKYty57musPC6FP93L1l
tNqP+XSTcgNAtLZQoH18AVBCqpIB6SGTXid7X7WTDVZEbZ7lbLKBJp3N64911iZp2z/rH+nTvZ8m
m/YbdR+h7fNJmbIWT2EIVhuxnrp70O+rq7UeGGNTM7AEWhFLrJfWW6RY13YY+5dvYAz5FW8pPJr0
y0NFokDpD5gDpOKvsI3CVu/E80M1xTZxvtW/RQ9Fgr7VLSl++P+HpxwhiNsL4irv4EsjpJ1Motdq
/jj07jhSlpOrrFU7j1u1I4pEYEPBGvLCuTbITBNzEskCpX3CjWCiGq905vi5Stfi7eKsZewDqtRP
axybHm2GiioeTZCEX/rJrO0Y9Mf/O2yXl80+Mrx0RPTkQBA8SzSabUg/MN5k4eZOPqa3h4mO4oI4
RoFGVhX9R+1d8u/XJrZgQtSzssLv2OpOrazYWxxkgs2nPYfEIDehgATOHhprUl5pOzU3nsmT64iy
PNprx+nnUj88DlAepuMGK0njHZV+psOEeQeSLRUEhuqUnP949sOd/g1rHrZ3SkkX1HdIxX1VyaeB
8L/sa5snMkzC0KIaaBsk0EZvwfCA7ksph4ZWn/oTMxa7bddxgL5jxWx9O+ucNQd3XIzeWy7CwSaU
PRyBVyaelb4TqH3GZ7GSql+ojnMDYdDHe6Q59Ia0HZui+m9Syt4zBiAV+En/X5W+BKT2nUqp0pk4
o8t1ZV1LCWtiDE+WJMKLLvBrz6fFsokgut/5u9AjNNqOHHrDs72wVyLByEU3FxYSbjDZdGxEo5SW
h5mFYR3rG1kA5ZWwuDvlmgdynO+OIlBoaqOVVC/65aGTdNAiB4gSM2Fx4AKUDbCn93Tck9b5n5D+
IcVBWq2yTYhNfnCTAMHlHzCbTOSfsmkvYIY9Fh+S5o3Imq86JZ45KvNe+AQ7u7w0idNJJbZXGDPT
oCU1wNa+93Cvs17IaVfjuFMsXyf1YO4KMfXTk8j/9N20l9zvBsjadGzm7f8x/p0WFfIf+Q8tBqNg
YBd5v4kZMB6fISxe+Z4hflpRd5XkLuzCtFt/9Q8S0zJSb4Lwp+ABNU9srC2esFXoAY9RMa2pgrPM
6enuQvGU0RE/s+j1/pihu8exj6z9D/KWm28LILaG6Ap5OaMMH8Ib0bf8vYvoCfKR2L+G1uUX/CCS
1ugrSoLlYwwcstTuWTQqclpEyRbSTEE2z/vZiDKOB+SSnhLbpvIXV/L7reDzTrOUR2y8ks46bdbI
zMdBoUSdlMM5A2g388cLhXGfE6lny6a9vjIhI60OObZm5R8Q7DspIigTrHOiUoZZ0qfmbtdT2eZh
jWozjMsKvU4m/vNmxDPYmyqBA0sr20ommWPjJHvKeuYzorohMTntNosxkLsk9wdfkhmGz9S5n/Nn
Guajxs50D8oBk4LaTM6J56KVjQX9PEFmaiaY/U9UX39N7ACKV5VuTvfqA9TOLgNYpnPhM+224QuJ
jp54wp+wSXuY5dUmmDIFI8UBXMICEYER2t+BXkPaICWKVllYVblFwRQaY8H1/Yjf9hKvlCqg39Tw
zj4F35BoZN13pntNR0TrYREQoFbN73p4AfrOQstj1Oput/Z5etBZ1797b3WRpepKLGd0WAPU++KZ
FOu/aNID3Aq3sRhTs0aAtlpIKiOTbIQp60hHVi1vFN5FdZIF7RQ+Kv5JYyEGLQuP6ItY2zSXnmN3
sMgx0E4MJS0/3UBRIoE8+olbZLuZjT3bItLoOKKy1tg/zCXgT0aeT6cr+6vEQAzmrRLKZVdPGBYZ
buhih7R0IxEB78cQtRrdGJLpM+Fa1r3LWAGWBzU8kG7bEX0pedVKYLbVSUsenHZZMGDy18kCfTNz
+zuOr9kEgD//wU/r2kDZf8oGdkjPe2UiCOhTz5bBcfiaoRwfuh9VtxdFmo/TpyoZjvdCe2lblIsQ
4Qx4hENlCSOsECHf3IlkevBApe+G2V6Hvh/M7LirmwzzjA8CUA6vgrlmTpOWadNCFvtvRmnh9wNh
lw+F2VZfhR0hb/wP2uujmeyzp9uzKVQ4oDAYjxq6poRa4X5ncj5j5bPBrefwTGDvpKDrdoZUlXil
r0tgHlZGFEePRkBQDawkn8PKCfrM7pM0nNWE8A4/Xrz18hnWx+x/dC/DkOXQAXQwLxqPnuZIyPhx
xt2L9GFmszuVB0NjdhwRbWY5qFg+jeoLYFbDqkxqWZ4ksWNEJR426MjYtqhOyqqXaLaEPcLd/iFI
Tq8YujvS5iLdRX8/WrCmkwECxT2z24rY0tEzDPux2a74kiIymO6YPyGhrhwomerMwssIdAjOHi33
/desvcVNNMtrfhUAX8VgJou9mOz0/KmlDmOryjnNGzbGtAhJ8plq5OXQQuHBLtvLKZimCSmjKWRi
5SyNebI66XGHL5lzkMSqboALIlSsPhm5zyADRik4XeIVmqsPTcarVfowrmUrUU9Tq6WHvJG0uKQ1
eudvgKqAsEGCoUHJg8gLn9/Lo2kwt8UF7WhH5KBN2aoQTB8dz8grBfoKN3peX8n6E5JzPsqslcsb
rTOdPLbenbzzUWa1Dj23Yw0TgFquk4GYP8B5OZcZLMds2UydmYrg3XS2So9kBVPDPZcu7awL7Xod
11L0yPYmL3/fPpWDmd+ByO0YQBoKodHVJQbPr6TwYQHFwAMvcfVq+ZHpKD5u6iVcSVyFj9PCOEVI
nID9Ac2U98xWtJYRSrS9lV0qOCuFh0Xq50sZWpHlZlL8S5pGj1fPHjZqRm+allIHMB41YqfDwfKm
ubPkijtBumNyeWCSp/zPgMBFbFlscw2WftVGpTH53saraFIc/MkwlkGCr9yffK1PHFqeLhEoHRfx
wILg87/+yTh+mmaKIx7EaixEwclmlsqCJP0At+VNBX6jHSYR1Oh6gKxznEZeN+3RdWnGZYC9BcDF
p9ng1BYTa6WPJQDlNXOiQry9hA6M8OZRSRq/oM4Q0r+5oXGH9VrN9Ip1uRks3GS/XXAi2UJX4CKm
j2iCTW3T9gMaeZW2P2vhjo0FTP22mVFYV/whq06/j/1KmhXR0JlFp4/G16YJOKHDL2awFCYr+8k3
PyUFD1Z+NKGzOFfjeTpN0rwBPR3CUUSR2NklQbMaVjaxtpkO26CeV4ekSl03hJJAtjC/LqkfPbO1
4y/KMyCwebR2sWeJxEKmn1c4Q0ZmW6ijyAGqkBYGOpYmO9N+hw5AGyrWEq3OZ+3v3yvslyIqlnL1
QNXNBz8swJQyVZiMrNJeKA6aU+q6as3EAnYUpD3CYz1w+QSfcdTEkJAaYow95spjsh3cHSserTfD
lDCz8dTpB/cce2x1x44Gni8Me2qxzvjpnx1OF6AUsZv1WFtNPNNfwlRCjnQAxFooaCx28TU68w4e
6FWv1h9htToyGNXJRfN+nVomp/1o2M6fjI8RQUk2bd7T7YtaMGtPD4Xyhhsn6z7bpcDM848rgV/n
G8jM388UUCnYRsIlFNrTRA3YqUA/4hyJTb3eUBhY/Ek3ghvpMjtMC61BmxMkmUWwnd2+cadmLizu
MB0/aCu32eD9rl7ZlHIIlTzZOTd3atdJAlWcpIpADPEtkjCdmXuLok17aAWEUFhicNxGoPGeH+TU
tVLpgURGL0IX0+Bf2IXPPUTU16PCodgiFBmjwFLbLWjYsAZLaYLyZZh23GY1lNRoftnyTq3gNvwB
VjVtMAQ6diL7H0jvIPttBI7qKSuk0Z0o/LKv4ItvkUr9XVKG7G/2zCHWGlwO8pdlYD79Oh/gcPGQ
YniuGOI3/5jmmQD/JWBK1c28/NMlmSzPRg6MgkLDzPA/TWfFfRzQZBX7Hv9eer8L7CtVRNdEacCX
3u+VepYXseuAuUobLmLlYPVl9ECPOqvtEUnfDCoLJ38GV6PknxAunTNNWUJc6dRyzctHKTGxX7p6
hxfygWbhoDSW78W3eV/z2bBGWDwkJC/rksV1BPdvK2e/mfsq9/2zKd2+BH22qmnTUuRDQaA12x0e
v39CgxYnrhtcZ9cOzyqzKXs8Q7l3cN20qoECujgnqNEfTw7A90c1m9aXbO8yQq/AQwII0u3RmrQS
jkCjewBIjoYLQM8DDuWS8VFs77sFkja4D3ZLqVhImXBOrVBKeWUPbijXD36df+Z1dvh+4xW3wmzH
79FT/L20LDubNnxPKuWk9qef4bw7wJQC61IUB4BlmBhlLBa7NVhD43ftVMicH8N6KJtKuogWcvIt
80h+n2D8wXEInqha+YXWj002Zfxln6tYXtZXru8slUtBepX/z7GqiMAQTfHNaWJ1rSt3L3En0kEd
2sFWpzwe/Cz8Hh2CuieDg6pf9otvQpXYzvxc6GRlUto3rByLcukRLhUq6JC07y3KUNWCMAKdAxsA
zkVrL9sTfjMcvzcamyKENKOE9yx/DVMZf6SaxB6XE0P9+n/D8vXIfszSK35RDu/6t5KSWlVfAHoB
kzFAzGU9M/UQQV8pd1iowfomLu5WfGDIMLA8XwO3UvTK8prLAsR5LZvi2IB4sDjTzylcG8L/n11v
EipT7Pg4uaRi4MbTwib+KK2bMeqMzE/m54lnFjmcSFh+5D8HypknCwLeimuzvZ28JGpEOO2HCCVh
/i7KATSd29jdxyUkQlcPQjbaJUoAUc0XC7xjWBTBDoZPlfQzBivVnpcJ/ODCxDvFaN/oQMAnXzVK
zt6PxSfUwpKVdJzsEKbG83NrN9ieuiagwVVU7SPmbMns+RgYsaEHEIA89eMwJUppiTSKwZu28v/Z
N9qRHjPJTl1YzbdwqQM74GYcUOTjPRAFe8Vki6B9TAsK20z6SKbo7TJMSwRbBqVEN+cuoFWFpQtc
GuKIRO6yddbbhdRB/7KSTN0hkEWhGngI7TIMEXOLg3rqTsEgQAN4A7mSO1fEkHVajt1br/8loJM0
EBlqAzYPgHGMtcIgNq8udaKp3o92oyUSyia1+MHNqWENGFmBsPnzc7bmCVKb4jIfl6Zn/z1RmdFT
U/fy/M2GnOPtKWw+/PaeAibimLWXu0e3Y+b+8y3c1FINwWNg2pgZ5wGNQDRnBTHPrFvVSRAWWYFN
+ifif9MNg+Pn724tRhVOCuIPzrWdJt5dFJwzaUKBh3S3F151yqL02VOa1IU1YAlFAG31me0iA0Qe
qVijABfcBdClGTZ9NuAEpl7yYA7MNJ1hJFU8vMbfA03UWoby+07Ddpc6lvYuz0G/U3URhzC8kIwk
ocB+9CcomGMsEX8IBxWm+xu2Er9h3hWqLSH+GZmEZ1tlL/DuhQZegtZDKNWwzv+3OY/Ctcw81u3D
3X6rIx800/dzUE9nDiHp6l2Vw8skpJWV29R1MMS32drE344JWh5j1hPrZGUgsXJULc0d0x61xNHD
ic4lTikCxeppCETw7/9Vt81HsOQl3y+iseghh41DGihyDVBuL6COt5Cn0D+At6WiQTA5ECn6c30F
tn+Om5BpvKFTK9P73HPKvxY3U1uJw24y8AUzT+OMb8BefzFYUTGK1NNnQ5p4mgmRkOmwpdr+eyJF
bymyQifDYZsQItDjGzX9j7Qdy9Y5T/nGwErcDNc0FbE2v82Fe0IyeSLpMDFX/KQDDJX+dxKXeM9o
bmoeoea8xrdVUPp4/Uc/S0nVcxe6NOMjzONRhsaRB3Aen2ieYI//b9W2t6+J5qSy/XzQ1k2+9mR3
E1O7xDtKTuQ0FD67qOP+6NgCI7QyJItcO4bSVlypYY8ZI/xzQTz/pN+bpeVixDq2S8KF04gUgLQ5
P5J8CH/XPQjflVBparFh2Syy022VTxrKKqj23IP/dZYA6KTdXF92e1et8RN0LiR8nGCJMrnA6pvk
4NW4hAef1DzYg/6QdCb3H+F1QTcXnDMDtaOoT6J05ieY7UFzjzqASEJ+ug2eB5hno4wJ89iLp6rf
isXte+8CVE0z89cVCkCRGWqGHOYGtJBTeZzLSfnxQuuW72aXytQPvPOYzqcxxIDPha7Id9fO1vRD
vlTOj9yCzGFMIthGUAsd72+ZOlNnFGpthzq9dfqhSwoBUXKlTxzkXOx1TC6lQddVVm/Qx5sAcgQI
NaJ7FwOWTRVYwHRCZI/CU1sFgB6x/+rvCvIKyVTiywVuUj41P3TdMqKxY2d96cZ5VbZHe7hIPOh8
EF2zThBzN0zPO0Qf1SUM6L28MEre16ayWwJrAxfZOuk3pV9FEdD5edE704VwRwGKEJcnDFcKkOW1
vdhJbdvG4YCnSNhcCHHhK2n+Gh/iMscRdI9yOvSBam8Mpdw6yxzoKUnt2/4aXUX7xuRhOt8pv2mR
q+C2lz26JjJsbUP+E7k4NSLFf5sXgd8Xo5MIl/+/PbWw3NUoRAxPYES4wlhBPovivAVrBFpxNy79
pvx3NU+jSfEmOqvvQf9jtxJJssdMB3s/ltu0vp9J16bWSmiJODdamulRUPO4Wl491huEcJ32QBuv
DuaYK8O4NmyVnhDbQueLpSHlo9bsulF5upnpEdCUji9Cp7d56Gzo9CiBhNzaio+ZZcUVwdovX85M
GydJ1dZC6SWp+EUvKgFud4Q36vdV/mBx/1HqtP9cNaBSLndhRUbO4qN6CQyw9Y5dq+gT3Nx6mwO9
jhKgSeGCDZUqv8wTBHMH+gY7x5o7M/aHaWwbNthsHYcS/lHpQkyjsFeu3d7nHbQC14W6Lat3xDsL
glPS34rndi4Nd0roArwB6WKhXER9Vqi8Wj0bcmm3kyOfHY6Dig/nj7I8sz4r6kq/KYSTuNgNQTU1
3lLKD4oPdZeCQ+j/pwtexarQGIzaa8eN4dn5/Z2doHPIYi2Co+lo8XdjA4F7i3sRwNfb3U6ZmtTQ
+gvx6O7Z2N8OPhMhj7b6QzWZNfRdtfoNpOBzqloF53zT99pKTu0W1/MAbrzQ7C9/nt22wHrGBeuY
si/ZKBjgUig0A2H8nentsCwuYVUVioObR/YQbn4p6nILtHsU2T5rTGCpLaMxOWLxD2FA9aaCCk0O
Z+EwTdPbjGdBxmK5UNZAC5gzIi4MpPgXPOvxQ4BtIdFZB6NZ/huGidfPVCyK9m4DGmMUjvXGady8
of4i+mW4HJKP9x87aMP0aIkTrrCJqsO4QZw2LWPFzUcDyxYwt4xNPy+1xQZM1sQwyiY5GYazOyn7
HDzsS/kqCpT7qlmcg5rUibINBrpmt56onc5Cvd8bH5EhDgN5dIUqn49f1rAih0cZT6kJgHTziWAo
lt7J4lutvpcHFZJmD2hwzWfpVTmySn8mGYeyTTgODLNMmvkEYp84yOWQJki96GvTgYe65UECl8Kp
EYUUeRXKFBCxdROI01YPDuflN3IAAh/ioYURb6nfvnHNZ7PgLaa4HtbcMtM19PIUpjGPrSRAZPUR
H0goTllxOw6jOBUZ7dMcEIjMIaozlFQtYBZrrobz/CEZU3PVspZjirzL+Rtk6VA4J3np2dXzdZTm
RczpQJBP4gCaQF1FqJo0e/XQ7oWa0tbesM4RRjwYf4/0EddEMKUrErBOE5a5xJbSQEw/uomqT8+D
rtHPqXzkVzSdYk7rryS8pQwxSjEBCUpOYVLlMO8X43Bb4GhqYgAfZknR02+wLE23KhYp3dKUYVyS
pR9JgCiGGufn86dX91u68/hcZYvHTg28p64oWYtropQIveTdywkCSBum4FUGrx79ujaIl87AqGhm
bnpdnzeiSFEfaVUGLcp8I8M6JiEbOZRUJL6r93A4YL4CQOxsU6GtoOnaVzBKi07oDt/ZoosQxQC7
zduPlrL5wfknAXiTJcxcOJZ4MMUk9cxDypdCWHzaKUuhz7hExbNrSvizK6/sjmX7dPOjui656LPQ
Ia3yVx8yPndEqPuUKJhcbquo+D7O8YX8iEjzoVEuCga59caN+Zqn4sxqNnDBT11Af4fOjLDIErp+
7R+BkIq5aVdxsdjDTb8bVmAzFBD89s/31V4Yc/OMkBi+Q6oFi3eSBStLJzjrY/1zN+I8Zd1//L5E
7wANcPEAaf/dKvCFKIj2IMSTDc3/BbZd+jkPqIFuROInzUlP7oTA7W6Omv26XIP9z7Cqz85DriUf
u9iciht5ff4uhc9TadkR6sJpmNaJz6G2AvU6TFj2VcE8b5ZEZWSfVAs7JfpUySaguJdXo0gjHNdG
UC0J2eWnmuWTM05AeilSt5kYTMTxtYPBT1srOTPFYierZano0YpLwVW7N0Ne584RGyHIa44M3d8G
phMwpYtoVlX79NKCUrpBakdOsUPX0ejT5I2T4236LC/Gt4+ypWYNNPIC3imC0+Eo3YzdFjWrJGFV
3dUndgXLy8Q8reYRD1GxZFFlxz6bvNHxnsQzST8IWByDkNDa0/3JnOPglGX89Q4rqtn1R9uYYzAT
7VQxxIpw8IQURlFHuqt+IoxtDOi0mqMKRpmqFgxbRUSLfFreqlDdQXdPjFhb6f28QqXZST7jGDb3
pbE4eF1YWrkfTJhO/VjHcmrA8tM7fIumRgZrwh9+oqAGuSTv4uXcaetNNs4XU21Me/vgns8KaN34
UjOgIxVP4SzN4NS87DCxoEDHU13B6QLwNSafVs0H+wWjElqaR1Drx6PUiA0Qmj6XrEUbdO0iuDb6
fgFqAzalP8b9HCzn6LDvXk4Tfuy5iufZOt6C76VSK7OoCtp1hAj3ge7yjPVLZSUySYNc3thCRRkB
xLeAixsXlnw3ovbayiCJ4baj8S8s2Exde6MjY6I6ZFIDInqRCg7KIXuST0LwEjgAv9ZsNUIw+PL5
tSmMck9zo6ByrdpejcS4KZWZNpN6kvoGJfqOIiy7bg407SyYBFQt9WmUqNhk+Yt3DjbFtYQakL3m
Ghh5HRo3GFFWZi3NTWB0tG3VVHEZZjqNYQWY5huVDKD+ohfrzlSYmXM0hq68PzWk0HcBm6tV2oIW
ER352aNSTtOHEh9lnikbEtNmd6RkcU0V+0bjd5JDUt7QhE4lgF0aauqmKU1CrTAH1PRWLutYOC9W
+kcdiWEAEUhHH+qnBiUr6FyvQhMzjIeNirLuOfW7uv75sALV/LG3Dwyz8VKyX7Zf9Osojj5dAb8c
wPOh9YVbHkjm2BndZmZDosYa937woew+ARULo/l5rvrfmS/WrlOlyzolD0tHlIas3+JBrZYxa4zV
dmR9BDUzbkfuLGUNBAJrsB8qDIsm7tXPAXir1BQqEMK7AGCndde4HWH0ydTjF0/Mdp5mk36Sp0v9
rqSHnWJXRt7cJrhbYTAc0H2BxTv5nEqGGhDBxPudcEdm9WcIhpznScmwFENkq422Yju1aDYApjPu
DwtZN6uR9kBdbYqSfhRu0+Qfxx2oFWpEo31mSZMFzTQmb61BEFG9E8PWN9joWaXLgvl31TAs0Ie1
6EedcMpuRvZDE1vatLwK6L16py/UkG+qgyLvm6UMMXMDPr+9/BG7U7vUslLVgAMZehUlNgCWwpad
mUXAsFgzLmj+UG5vx7JRJQ2buuyfO4ribDS7PHpAqXtggdiuPf6kSqNGda8xy05VluePwgSjjjl7
SOFZQ8LGOa5yi5oNJUoMBcE+WH5dNXZqEFvnSdwQHBs70DdDN13HqZLyJIoKUoIRkzMNX7jDEQn5
W32nApwetYHTZR0Rn9zwwVDXrao9iJprLgkbEXGvR0Pi0CGFE7MAptG+Y2kp3EFbwWDRXhSdTQxA
iGfLZb/c/g4nXqRl2nGbpv+V38M8c32VvsSOhv6AmvwMESjML+BCaZAQ8i2mLvVUYthJbpDcltp8
1DirKwRVCWDVx2aWn0bxtF4Ri7qgd4diOhebzD/n8h/7xKyVE3jX1zQE1HMyKOEEj2UDNk5blR2u
bfyCaQwCLT7uwiy2zkaADAySXCKsU+FhsJCgqF4f9Cq5izVwhEatIkz6c0IpURhiZtTYx1MZVrpo
IzJdsO8Hr9/graPKiyVoM9qVU49aj8WsUBz1n0CpN8PTGh5A8xQf2Wb7iCVu+YC63FtnTDcCS8FC
P2kxOjhuSrF7xAKb1bWXxe8k74r5YTkBcVwM40t1nwzK5wI90wwrTbZyBVHxDT1UGJj0tKnnnusj
gXmLBJp6DdgYHoIYOXzXls27XM8At8n8N38QFICkkyHG46vvnwreajU/aZN5C/pGPiqO0kFwNoVG
4OWymrB5JEaUL9cYjgJGTIZvg4C21XjLmZzMbuTyIqIMLt6ZDxRgpHFwUSdg5Vf2BhJN+qEaQj/H
J8e0vEfilpU+f4O34+Nkmr6XS54lPp7RgnB2tMpvCjGPvomgM7WE+U5uhPlUXjwCnAyzpnuASQRd
CQUGgAuS9/Ht4JcEqRXCGj0Z/F2HGGxH0xuxYfrK8ySoSlu9MOsazFLX2hUkstATFUyEg/x6iDVS
tIQEkjY2Xi5r1PK06TjvX0sioeSzHAhwQRQGZqY3cmw2h7Z54yzmgqn7cPqth0dmDeFGLczfdJr3
M7yV+kNqemntnRcA3O34FHPMMY9QSx87QimcrArds3oSCuV2Vrb59wpj4LVYVZpsdAPlHXUrvrtd
RuTIWrcHVvOmMiYj2yPGf9lXyO/DinIZU5yciw6jgSUakTf26+Cclcnoygsuvy+rmQV3ITuit3SD
Bj3576I8wawYVk4oDu/SXJ76pRjLVI2W8h+RGC84cKgEgTj3cUPOxNffmYDkuSCIBCuZaAoG3K+Z
gpFDQH158AvNL0V3sbZmjXl8T6DS7dM2CqHyElBPQ3Mp1oga5N78d2CChlriss35ZfQkxbav6TEo
tRZZ+GIXWllSC9cMiySwY3xc/T92QM4PLzvK/wfxfNuICoaDfSCxotW2rfu5nlmc+QbxjI5Y/z1Z
OIbLwAAGNkD84dZ4ZSl1c44RiFQvlFrDsWKuVDppG1Wv4Ejw5v5E+Uivioervr1nkJV4ZQWsGJbk
/oBg4G3UvZ10BOgyWuGfxRS7u93qhvmr3LUsPRGnISysu8q/D+hehQfJ+Z8nc344vcaGUsLEMVs6
wSTwW3R9E7eWmcyeqHjs+uzwRmnWb+vhwRyTO4kohR7zQ7DyHjt9EfFBhZCMOg7HGopr9/P4z/Ke
TngY9kusQhSH1eH3jA1p9X6uuXrYL8r2WTR7zcb5oK0OYZjZRmwPJE/0rWXusfFVt96QkAWgfIa9
rPKgfdTF8ORd+2bvoJ7mHoMFm45/RLEOfOYCHb/keR8uGXb11nfuspjb1QNMFfiroC+IOn8IX18l
D8JSmyVkVhrSVcNW2OPSLX8Y7vPKnXI3l9cWc5XsLfYHM5kb31wYwsYg8IigraRwahY4elh3k2r9
fKUKm+N5xoVB5qq2y0UnhET3EYUaou9NcZt9er6AEGJWzMnL11Apvs8jPvwoi7YMJLxX425yT/RG
H1h8CzJ27sgevB7VrsVfDVOPAcvrsLHBxJ0TBTIbqPl5551hv4ZQy3xQoSHv3D6vjE8+0HRxN3If
bE92PXGe95hsnGPkzymuNfucIEaOna3iLEy4aptgwOrdTSlfoGOHPw5e30rJpkRrhIWcpmCTGtgE
xw2q4rOrH3N5RY9BprQs2KsyTNI6YscsilJ0sBG2AQBAUY/yiV4XPQyo2R9ICAOiu/x207TMZAQ6
Py46+nMQ/OqdrowWbbFBSIqu1t1kZI4K8skHmTqXUtpKg4bLi93TMWehHEOREkoK1oody5Bzl7WO
k0/JVkFqLR0jzC7DDYWghFpLFDvfSToe0bdreKLvOcKQCTpzdMVR5d3fWl4QCPVg5lKQqvkJcwSF
os1ULvLwOfRP2k27T6m1gwUB6qenXDAC+iJLsRjlhqV9xlXdmVqqpYx0sTALbo/H75bL092ZAWaV
Zo3zpCs3T1UVVikxI4Wb1v/ipFTSW3i4AKapxB+cAtMLNMjfOOP0Ka0+Ks1wdObuvg7MNfrrOGQW
B3NR4VTB5Wh8zRr8YyX0R4bJ1I+a6wXMxEASL4NxJxUw2TtStt/BdztYpjRd5uOibJcxnpxZFJhP
rDSr2RSiSq/ssB++W/blPgZ6CtpCNH5FEIAa/TEorodw95KJ06JGqHQSs/TY85YxfgttdVZ/6fiS
cbQSPRDSfsdbTE08cPBZHfaObmX7K6T/BFFDUlOHUONy4FT7yYl/v+1mbXSjtfvKjhVu7KqJ1xNk
JFG6qZRMW+t2kCrcQwAWXNv1DgRS5bTa/hyb603mjzCXl2D+ExTNVW2TZ5pHBRWZb9HFoDkUxkZX
eZ6G5q/b2PERjJOk0XjLGQqLpXm4mn5Se1XOXfFSBHgkAKdWKsmDaT3dJc+Z/V3cX7DT2Xn0V3mo
UnAWDBEp3vOjKwflRPA5Wxl+CUKOqrQ9QiIdxAJEUlbNT0ghirX4t+AQaRydQrOyjqErcGjQRAbQ
7ukk0lpUfJwCijzZgd31DNl4HpdriZOBVEx6LmgYQ3jfBVd9Rd6+ro4P2FmjoS+Q+dgBmkNJFlKp
3UEZLeOI1594yl4VFmIExNMpFIcMZKBPA4TR2vVZrdaPSHRLrLU2QHk1B1mvPEiOqPlpOIIAib7N
dtJZcgoZUFwqpwwNTugRhd+I6Vjv5QR31FjZqmrK1/h241QM6pbbLAGg+PUrU0YkcwVT0mXrKgxy
LN+Z3fqjsETVH0j546edbth0KY5wOSJYKUdenD//6jyNcuofiUXt93Aa3Vs6LpfkE06l8KEh/frg
C9Meme0FG1j9qPLnHLgBcDBA4nvVigBIRal8JdRhAazrxhzejgNfd3UYbcWCaR6kqaF3x6/vvpWC
wWuyPCwDI2UbegrUtW0kZFQIG8RD0O2lyyFeIRghEXM6ju0XvChXgl73sjwtgNZBgIW+ZxKY69r2
sB6Z6xjI4Y9MGNL6764boHpRocP5qZuBDctkKd7vszIhWDQ6lrs6zeDsD2IkEcyKog0p5kt2QGmh
faQ2CrW7TmPWXLsMQfUggMUh9InouOzh6eDl8kE6nHIm+9y+DOt691WXRJNIfEkrWWwG6RRYjyMD
xYdS7wjavHxgPfytRVzUHEqdVSr/e/z/WSossM2QhclTo5uAZIPmir0XhnlziO3ZlVj64bluDA1A
kvNsT0rTjdV1M1OZLDlTUAI2RslY9HfHhG/Gmxt9Y8BYY7B2flnhJ7WYPfuE96ciNZWxMQg4iaZ/
Ywy3t9q/tON2yoOIcsqv4XPvqmjvIuEbwLA/0HnB7PhqDEu4mVlaro8A/Jj+zfBxD1zxt75S7CW1
jdaZ3F0itdupvvNLz8wn+RJcuAszQg0Z00PfU8eo9Wg+suWxFDZigQAsurw4yq+sRyo29v/UNe4n
uW7+enjWWidbrRyVJ2hiJtAhKsSnwjZUoe6CF0GVK/G3r6B3IpyIcGIIYHeOI9BBdHj70V6vs/TU
vIJKivdV+aJ8aVUjD+Yr8XwYIJU+u603XGTAxP2c3G75phbA+NdKTceGbXnYr79DCLRgbTn1v1v6
1pmLkWrF5CbLpPlMCTBgBzOfgyj3UTLicmrLg1dt4wMaGXy7+cIGvhIqSRwGGoksLftxSpaIXuT0
w2y0CIHHHXusGnTga7fxOXvB+atgKemv7hsNfYcdGveGw3F7E7HDQJkYl/XkmKEzw/I/s1v45Tne
HV4/2M/NOF7hZbU+oJVtAHW2AifF/T7IVXjWG5r2q+SmuIp5Xaf5/ZUBrnkpebbnQQ/uXh+7EJmp
AXJJxZG7q3YNHC7SdAlWzW1Dmr0P+vh5acN/wtk0+JHiyl8S9ds5kllryYVQ9nxmOxWlhmfv7Dlp
0Lksd5TZ0zo7KR2MgwvvolDyLRJmojEJDBqgyU/r12VlFP2wtP0MzEi9huCA7K3N+Jyv1N1KI0TB
gRrD8gJcn8FIwXX2tLig+qjHlMR+AlwKan7bSZlZW8HpFgHHEq7xIOrn4YYBTUaM+eBFxk6ROUSK
mPVxPymglVB3jMClkWdkaYlVZUKm78V8bAQ24rpomFOqMLvHzNZ2+9oHlA+I3A3UsFwzVdfl96az
USgY8dq6EgbazkgKQ7GhcUHZZ56NJCyxz5V/DIYnr+UWuJrXZsYN6MEkV9fWFiOWLN6UVTaSejx3
gHqEuPUecNVHgDlpQSE/kWZORdRXWSdp1oaN5dJ9Uy9b2KQFfa702MbtGJZLkPiM3GQwfQd5G/34
iPKpDN0HoSrmpvZpp5Kx3ZeLCd3uiUaHKhPq/+IDfu5zc7ct+RTzJ0EwebmStyyKQrFFU/4lh/EG
SB5tY0lP50csUZuXZLkG8EcGlp8ahtZUISglD9tyElYZjyhTCjoSyH0uaY/vsMOnwi1/TZ6Zm+Qq
dp5RfODMPmA50hf5WhczQWkN9Hlqy7CqUWpN5kOZV/Me6l+1GcDqP2K0PiPAh1M323NyPfiKdVfj
ugnyLaD7K/EgXjCXAZQ3g82BBwJZGxnMwG+yejpiPbG/k42Ts4w5mw2oWTvvDA6XHicC5xqJnxEp
7bHjJoSvdK8fT522nETLPqbu6GJIp2P23S8uIJixNclUglqwuMPyp86/OIgvVjCdr0tMB8CLUmAZ
FgKZu0basgZrnpwdGf2pKwAZqEfIGdTQqwY/IZq7FhmGTcfgKvL0uJqZ9ji/pMZp41LXPwPT+iJc
Ox4RH96v0OfjYOE8aWLmHBjAOIrDY5DP7xWmQIhuOOFbcM9ZxjJVuoC2l/hWIZyG2WCq7OcrlpbM
6DsN3E9loEfOSMWaHH+lDyJ6uyVM15bEvPaRCKivLcSQr9NFOL984YfQJ3bJ5rrJ96Csjy+gBxso
74vgWc/VBTQGq5LAQ7/m52nmN+Y2WaTjL9M+xa9gVJowfljZQS6ARfa4VqAPiZOX6fEYUQc8Qxbm
JowZzK74W3082Lapj307cLJx2XpGRJ6sW5SCl0Z/NGQP95yBLkUIBHYtiZA51gB9he4xnbHHJNzh
3RqsJjythLybP/IB3Zdd1ReTHPo+LHjpE6ndjilML2LheNQZ+zvWizNGMh4yQJvbqRIy/gWt11bH
u+VlohmKRZHlr7hdxje7vV2z1YaqgE4rsEwtnRHt3mY1+7E8HHVu2ENTih6mWjrWjr9fl2aTo0Wd
nTzluRlBBgQ9ETAOhIIxdFaqOgQRnGmEHR8dCwQc0Sjmv1AlDSMFdTTNyA71ent+iFBpMzYbDPF2
2PSQWMGSzmZdXxoSVxezm1DYzgKE+dQSztfaA5+NhAB4NDDHmhgK6zyG7mkzYRBZbu8eFP5e/SxH
VocktCU8vBrycpazU0KT/uuxoT31nYS8iPbiS7HA0H8IFLPq0LuGJPxw6cqsV8eptBUCZqJsTCz4
x6dXWw1XhYpBzM8vtD/Rb8gfm+q3R4vxLmr3YFkvtJvdsQkaYlTv1hl2WnabEuKz8cDl2hAtkebA
u/x/6pmxxYhnsh3Gwf5GLFpZF1LnArwQV5y9u86Hh31ujE6bl+OhuP4A/MSVeUxXDXBTaB8CwN7l
eP5N/dhq3zMaNP00zzT3cziCrur57xLz2/X8EMCbU2PrgZCpeplIz4d53+8hr7kwWBSbtMpmYcvn
OXMphw8aGbLTQk2wtTAZSTMHeq+blcQOf5PAlAXFQE6V5PWJNjFu7q1gWGM2HdOzn8FbriXpgGbJ
fJueCOWQpWQIMUiLMuNf1+AC2ZKSSjLOSuWVZU5Qr6Cj5AFslw4MZHBJz/SheD5Xqqh6zO6QHx/x
4Vk2ETaOU5wk2AMa58OuA13lgLHC8CzWeGXYANkeFu8n92yGTwYUsJut1Ogw+vN167cm0qF/aekH
7uq7EdqwUWl+6GhCu+cIZ1Wt2yZLTF9OJoRJJdKZL4b+8D9FA8gVbgNIAEqQVPz2/ZpmQGfz2e0h
dfnFBRHb0Fze5Oj85i66W5LJttZ0W0aUMM+ZMVOCDR4E+iE0AbbSIWZA1HvpBuTZCKX/oGHVzgY7
FxbybMqApQx74wtYZIEVvB1XmYMLbUGBR9IsmTzlz6SYjg2nF/+NT1OTXVRKNn+X3+z9+B8fVTFS
X1SoPH1vJBZ5eGsPRuQ6WWURkF/A3JecGZ4lRLfFYGVh53BHT+aeU2kcPy+jZY5YNXlVKsyRWyex
IucoKzBId/pv2sY8BhMpyuGPDMPFqwANXAr3DoLmSg1hDJuEDuu621DLJ7e2E9hXM5PEKvXp1uUH
kxnQ7c/zKQ+PakoAxmzfik5EdOLel+6CvSxI6E6bmKENXRBszH2ENvV/8I/7MkufoW17u2RYpAbN
had8maVefYqfdA2Q0AjOP/ZWcNLEqBDDgw6Oi3NCEhtNTYLAOvWTD1n0rNNptx+iu8M0bAM21JGL
jyGb1zRop5t1zNQx41EjoXE6D4uOUorG5lYP7CpUZybeJoW/rCDXFqVUNP6JqByzttMrm3jiKCbN
YMfgWHAtUhZCj1LHYCqDJbr0lQFhPpstdv+MnS9sUZLI2f409YLPE0CqOIZArC0GUekP9inrNkk2
mv45WDq6X1v8RGhOlsoAXBnGHx2PTigWRHv7XJC+tI59SGNolTlth3m67hlbBz0z2zgr7AAU560x
l5KM40a5zgwkeEzvD6q9k+59Y4CQShIS0A0eCzog+c5sqAoALXpewOrUntF5VMGscYxIzKFjBtXh
ygoE7z1ORtMS0TR89zjkaXUKUzrXkj1MZNvnf9/64Z04CAtMHAxneLYsV0zsa7ge/6chQnLrteGR
tMksQVxy+Zh/ZW9O3mTxbbHRkDtpaGruazCe5GWa6KtWTGUuLjoln2B3ZxtEjhdXnIR6duT9LO+Y
vW7B9WXH+D7aMCzl2+Xn1HOIZfGDHtc6T9GPLXeMW0KFsR3cJ21PN3piWyuzerJ1XRAnf/ytu51q
rHA8em7gFvtvwbctQdCG0B/uuQ44FC3R53tX0j2sMPsdCJWS5taQd/lkDMOOmT5lrTXBp0An8POk
95ZO5BTo1U97Me0zchTq9ZUJZMNaY9FfK0cBRXnbyJH4G7higE7aSnQN7X8eA1SKK85oKEszDY6c
oT45CnR/zGl/Y53+KK3Mww39hbaQ7bkIYcNInvqi4YkOWJIWYaKrrSTvWhc74lbfNdJcUBolWsft
O3YIcDjfPmvKqBEX6kCVafdhmNMznHZRfD+fczdXL3HvVTr6Jx1FbXbHCzqzdrVjJyHuORE8zYXN
RbdE26ttf06W/eeXcyEpZ78wsNCZTP1SnHzipqZpgVy+lioCtR92n1scVdPbpYpZynXuBg9jgRIV
2n9atCblLfS8T37P5rVWt0sN3UFteGV/ORcPCu35gsKsQByR+rCjrlQj/Pe8W5PnrEDXnbv2fFft
YUnFD3MtP1TI8PXt/54k0A+yUXogutKOZXHYlNnj+mb3+pxWgHoNWZ0ismKWWLfaMDNhB7I3kY8b
GJvH7WVqyzOmt+GVTx+cGTCNYo52F9i98jpiIj6Mb9gwRylbtW1dehqDM1eRAXbPAvjH6/ViGoRm
Y0OPUSyUN+cv5lVOdYj9HS3DR809n3GZyLc0uRPg4t4rKim7495BO9o+P+8cWDmMyCrLtDS142AB
2UVQYsUbI1EQ5FPPnDGGVKPHslLMfNM++SLGYUP/cxjTaNohLBTV2SNeUbqBgWd8kXLcVStKInwB
NUl33ycJ1BkbYPYVbKfQ6+1WYNhtA6i3OhXyMFwiI+MrdZCCCoF5vWzL1WH4kaJCCwfVFhyBJGVh
4+oyEhKCNZ3UekOgt1rqQfnVeVb9y09AEPJPaq0EQLCYwcpiGLhpI8FAF/6XGcxRqlNr28aG2XuI
mln4AAZQThk++GbHhEBZgZ0sRnfJX7dW6aHtcQWgrcTM7tGID4iAXBY33I8CKpDu5jYomRUiOX3n
a+G06YeUfVulzeBQeq4/WTNQIo904TDb0lboVR53ac2Fb6FaUHOUPj8sAv4/8YbaNpLFDA+BooVf
OS0MBr5ybtcKWQX/FE/YKrQQfpD9ClYu34wgTzUQ5FFnqeawPbNg3AyoYU/HnWdGOzQsXC76VVmC
mSgo8W2XFIGJ6hoUgau0ZJGe0LKxY5n1nJ93I0/zwDqhkGp3/JUQwBjEjN6fg2Xtmffhye4p5M/G
o62eSGum+kmHLspTQtdXg4FCBjTW2bjoBI63SVjVpjlQGt3LBj2i9pxSPzhnD/BzDLDhfHHeVSsn
LcwWY55Tb2KhjK8Do++GGmO4rbzQn1WR2AQ8zMXTDAA0hu05POXMqk52o8HemUGQoXmBXvH6NL+s
zB99wQjrPMNhkpkM2gCK8TE07vcjFrir/phCjkxc91iQOnY/oQuS7Tza6EQrX/oECCg35k3FEFQ9
4Y/WwHNVnP07qK001XEZVvjxAW4bEODdJKMhaNDaPTKw3gJxWwIt0z6tUrvBEokNng7PvxiU0mK3
EHs5/YfiyQQ74Pro7xOe6Ot464Gl2Xkn0f2sjja7SpgVwUKjeEsyQ6yLce0x4za9swwoyayo8/9N
MTpYGkH6EiICGE9qTQ+C1I4MpckavWusONpVGxSLFAi1ZQhb40nrwV4UpA+Gyy6XSOc11F4RSzDJ
2nzUredki6RGM3Ip5+rLw/dex4F7fxGaTiiP3hnTqhUFtqyExzI+xsu1/DlWv6xSRaTXPWRDIlkp
0o2WydEIB95b3j/phoxhZ7DrwX5mIlEsp/i6EtVak3u3pDxRxCCuArmb3/qknkvfws2d7+XdhW0b
GEjo6FSSQjpNWwt3Ct2qt45QVosxedKpT3kekhgtYHFlS3Fc/LESqToZsPDR3ZxgcVPIBSOh+wJU
nPL4V4DOi6qsgRgzM9Tzielj5rS46/KRZrdrPK/EDZtETNsSLBsFgDKRFjSXBqvu1c9zXUHcRu54
n81WBziHQJomA88WeF+x8VtpXs0hPq6JbkGv487kgoG3WguUtiy3gIAMzUvjfIljen4+EwxB/n22
ivcqGAsE4fruXwnFUmxnN1D8ZgKac5fggNEl2fyOE6sZqs33RCNXu9cAurAugCreEZUCFUq09SaG
/kc/9MaV6rMHCtZ10ES4d4wYxaoiOWJ74cVPdXY5Dj/JWmyCRrCLM2eDu/4TRijikxpsfL8w+aNN
QwpTXBEThInrRMAiDvcfJWFoNMBTcUBktO/rM73Kl5WGd+l7eRXneLI/bVxBuZ/txIsjhQIp+eFO
c1+Hbq9RpBh5hL6d+5/4Qly/TfAVApQaldVY4xCPAL8KxvehrSFzSJZOAI+C3Slf2B7vt6DuNsZZ
R/tnOYW84iNEYOxwyzd0EkXFDmAfiKNXyNvYi06SSvO7PqJHPdEulWO3osjALD4pdUROH7GlO3aq
Q5a1z5LeaRjm88pQR3bbp2DklVYTVK+tqTR549R7WdKWLYf2XJCRB51yTDXM7lT6DhSjDn+Pj2Yr
Uy47TixTdwoVAtOY0pcFaiCIJYHbZZfnhhEiZrpVqJ9RLYCmBv0H/ud4/BwbCrBhiVucpVq02uO+
oW/LcdjqNWsuqDEAc9aUpguA9xYBZOcX0cvOBEKMnoofMHg2ypGgmxS9BLtEdeocOpEiIU8RAJWN
OqWBPvwVVBhfSrBA4UaFBS16pcOCTn4bb+QphRqb7Pkqrl5r/kfrd2J2ioRs82uqK2yG9w67yU9u
YSXhzLfpE6iG+8cWdQ3WLQx0zY0ZbcA6ChaiCPmRUYa4S/uilC9CQJccHlu8fLNqA6+IZeZRAK/f
L4Kaf9tAV7S1JrMPrEE9Xlzc/dvr0ftpKP9nsx7Im9wTPnb5MUis29x58S9qk+RPGI5FS7Pf2OY0
bV6+PCchX1M5PXc005RhiipM9AoaOyH1t2O1+MUITWjKJquptMLEV10swMp4PueiNiCb0lQiv3o2
53uIE3R48QV6Bhxo5hGtVhXnF1S4obcMC+zlH1EmvKzKnuXh85ml+4PyMyNNfjf4C137Cra9BmZs
BqZ8RyvxzJ9wOydX8kVfRZ6otGrWYWLPekZx9/njvBaWzk2752fLS7xtimUk8XLckR1fBI9ziB/h
W3SAwISP7xqMOKFtYZrgKRKO2W+Sl3cMyreN8zUx/JJdi1QgUJU5V8sANHuFv9iRwSyh9nUHnl35
mUqEPf/xyQGy2Nq6SmPSDd/wYUx64R4ssDFLOPuJRtpPAwjpBKmJSshE0O5QtaaMiVP6k8GMEMuU
0KMkyBK5J7BMvJxDtM72c6OTMUCcikj8aeu6y5lw2uiPRtBpB3//+8gYYLIibqR7s3e3APi/+r8W
eOTmfE7bTw1qPvPLlXPk9sY3CRNOT027cy3xsCP3A3NysI4pcAbR+n7VAS4tkfBHuvZJaCsqwVvK
RBqEbZB+ac6Oc80+reBdTpp8JrhI4Q1ISUD+fBhygxxvaGOxQWF/H1gPz4nU8Xj7250kTdxF3VL4
qtmEwf0p6mz5E8oHRDOCh2PXT/Xd545VtwcN36Bv0f+N1OsFu+Lc9wDKDuQsUsV6f0dJlIf7Z7bG
oDAIWhJ9Xin9zI435Qd0zufQQ1Zgg/MFokCiV5tLL8RWjVBSr33jCueOTTaPRtnxmOUS+5kEjCyh
euDEvAUXRZnvxaDBJ2KfJLwMDBhgMS1w9CVPvtSF5A03a+Fq4g2Vrju/z0TrATvEg5speFs3vA/H
00WLpDxoyEGSEhtLomy50TxbyOvK/2I4ov82VCcV5tSouJ0ZVvoF39YmHLvSKKBx4oTt2indb/Nj
OOKKVnp9tDlOwe9mi1Apt5ya9OcCulYEVDH5zvVedOjbECm6C8Nsm5PmAuht0n39kJbqMgohbUr3
83BOpAIxxkMeYsF+5ImHxnY6it4ucEsxFspesD2EuxJn9wfSGhdcg6w1ni3DrKC4G86v2ZMKnJf4
TdZCretpSol/hKV78Y5oi6cdOypSyqUCglc+bXRBodf7+IPQxkUdjednK/y9hpiTkTh0U7jMqoOW
v2G/KDqVMJ/FXrC4XyRyqcw51jihfYgdiAVVL8RSEOdK4nTkb2DDj6wI9+OZN/aQBoNufCkXSzAE
6EZ9MqY+sJHDFdGdm8zn59V6M+mgGl6JXo7PQ95rRFoctmFBlZKU3vCVOuUtJgPyMi7y9UVrnY36
cqlvwE54yT2zahFM9xwCdOG87dYd/dVQAk0iyyDkUvEWbzDfzPD/VR0sgxCef5ThMYfv2a3I6pbK
F4/qEiFXreHKV3+GQqULtniTf6XVRAYH6n75GeN3MdSuJz3RRE67ckDjbGzWXjkTMdTWlTlx3Gg5
ZRYrroR9oGzfUZbgneikGzZuL7bIgEAzfnXcrdUVx9Ifohsix+pt671IZZR0IytD/c0trrDzj9kv
AEmTqo1BXNbvY5ssS9G0A/dWjlF/sWY5bfauRzpgeMeRjtRr4P+ITAs8cmtbuWBRwdn8KJtgCSNO
u3QyY1uAuBWJXWau6BdwMNz3nNptwY5v8ap9VLOvvDVEqgUppPglPzWewCanMDAQTwc++SvkMPzO
dP3ANMerqJxjn7dCXc7+dBq1ETIy1XdkvILs/8EM85o6kvsSZ4CdjJk2qjEC38vBVX1Vdy9e1inC
gsHNyJPTc/Dv0ci6kMurvaM68Qm3CnuuHh2Qj+yGU0IWHx9FXxAFNdlFur5dMfz6I09v1dFUpflF
qmEDKng0oeIjXqJGTaEyFMFEvnxuron7ymmHxjA+31IEEBr37y7S4SlMfGfIexAdRASrrU2gWejq
hFw7JD6ghoTayLTVFoqE4qZNz4op1qylIi2cwtrDRxfEqe/Jkh/mB87gzFFGLMU4Sw3B2sAQrFzt
sqYrJ++1mpJoyOYfqnJYu2f+rcrqugDXk+oBHUq81T98anAXiWbIa87iwQCVOi9mawd9z+d8OeLc
YEnZAQmFVCVKJAuk5GXwmf4tfVWm/LdudpmUdUqEW/QsdagLFljXS+0bwWIBl8Yn31ECikeSPlDl
U0GVDZPiVVJCwQTUPCDippN/jlPpYdGQSGY+OhfXQXpahfXScV7hQvkshdiD/5w3LUmIlXAUhotB
BbVozf/U0+VORMQhn2wrEsAUqmWlG5IRbHrj5ca3zyhwPrkeu0BUL0DSJnpFdmEfgvyXORYfFSdn
rjNQrIfvr+mYKSXFd1Ou7Qe8x3gjwyv7+IzufjojvneQCNtyhGXlrBuTfq9LdkBvBS2x5tTIb/uC
Jpzngf1MfDiKVkVUVQGuAJyy02lwzCe2HrjBCQKc1o4q+dGLJvm+Qj7o38NcA9iS7Vc0jZT+3U2J
AOCekO3ZwD/B7GpORREUM3TQ/0+MyYqiduKt+jgPxgmwtoXHDqwR6/g1/SfhAe7ksR6lMIvR++3O
mXnLMAJUO91+N6WXKwIoBxx2CpIIBYU4AkcJW8E9Xo/9zP2t5MpXqmOyDsE2Vempqs4sJ1PxHRqL
IoMTaAFwjx4vzrOH4Arl7dUZO1ck4/nZASJYUtbrEmfSJHtWBCeNa6iocTUc1NEUiYVJ88DGqdlX
divgKQRX19PIZ3yVgzzgkR088SEWE/mr5CMSXAIcM9ICBv1ytoPXjXnJeek5W2S+B3AxpnQ/S76r
1iLHTthkcM4OF7z2yW16T8/fKJK7W0LtpQQwrTNhQxD2TRtHehNrZGXD1hTCEVNfwC0Id3N0Kehr
scrVGGs8icvW9L9v9Fgjjj2AtgTuj0lqK5FYzBiOFaAPTURZPe/dihDRFXiVdHUkUdPI6QxPOdan
xMoVMUiUnShn7KllGlktl4rPKEBCueUbdjgMD9w9OW5/ih4VdlsYdFYhmtK3S5UpFJfeA62Ki8n+
dTPQu/4lX4Tgt6EngpCO6iI3zlGY1O+taqggLhiDxeCvNqZ8uzeKoypTwOqSxkbFdZ9zXDWM5ewW
32kqvd1uRMRzPgrfuwyfqy2yMB5MGLR3d/ulhwKwEqwZ7Zvzd2VZAL641OcUg0N7izejfSPl0+xv
tD8Jt9wkTlnryctAHadSqv6kfTLGsaK+/ITFQlOfi6GWd414/ZMvPl0enoGNY1DptxQLPZrV3ZLb
VqbfkKZNs/dCzKNsUtdGlMVkhx290Nv4Ihuf2PiG4dBbTk6LkDYA184KwJCeka0kt0NWFYmAthJ3
I4kHXYUE+OatwKtCBV8PMHlTRQX5jF3dBsoQNiONsmm//HPUDiWJJxF/pf4ETaXg4vS6lAnzUI/i
Xl+ljKima8i0mxE6fXBQlD9nXydRCUvhmr5AU4Z1O4d06L9z6Vrkn+XPeBpYYu8nXYxJQxnQaeSA
/VnnzbAdE1bZnJ9fDh86MEvVhEWznXp9gizHMpQ6d6+0+5NGBm6lub9l8lhtk86CkvlEYpvEtv95
Z3bcBORLWgdq9JTFEW2ufpIt8hyXyrhhLXPzUCyUCGVFrz26X3EIe9hGGndjhzJ463qv6EBcvpBd
dJgBbmCmm1ujA21R2ebzaZemyDsqFU+js2yjU4Lr9yj2+LK40s4rB7wXWJS+x6L7FYpWbDDMwInh
/DoCsSg6NseXLZZIVhryH5EYdVO9yl2jtlU3k9hFfklVbyNPp+V9Yce4hZgWPmjJgmB9Q/SmyLdS
m7U13i8VnS5LEdqOH+cyfA4LjDZr2wKa/utEC0XcOBnS79AquyaL729A5XSAvi3frJuZNO4p1ohB
yDeS9fwz4/kMZ/EDGca2p/fT8petMSv2sywCqZbIQehUN0l89UkK1dIcGooCZEZs6vKm7kvFILBQ
lzXwpT5IxeBgwx65cYdOLsGAX/3Atilenphu+/vM2V/KwHAsW3Flrk3LJx7Gh1GDpcwUmv5xB1EE
PI8jXm4I9sdVe8QD0S1oLLYk1tvQ7VIz78UuT6Mhbn3kEb7T6PSkyMAyCisdsbsN+e+C4pw5PkKX
s1QOZZrQqPr5i4Lz5wogQqNj9WWn4Yy4KhBRKY4+JLtKKSWSvew1HuOgZppEntB8/jJXa5HxbzqR
Q21BRidRcnjCEcbZb5gTI4wToQYI2/ONrQdmgHa9wy1ysRBhxaKjccOP4dZXe/Y9qod52ZZhRmJt
IZ6BliQJdFGc5qhrhWw8lTp99EEso1YOjpupnZJXGq+eNeUWmeeq6UXU2PxgL46dF4HJyq08b3Ie
n1Sqse7l6yMUEhr5Y0QYPFds75b1GfCa+lMj56eApEL7j3v9H2SVGzYEFqK/1PFeSnTwxQKw5jij
z2NdJYDYEVgn1JuCSLGQV8LeZ82mCfXv4yDvUBiKKWLvdgGJ/5ktleTnVodoqRN7a1FUV9z8YM6v
7sDwYq2aM8inGF/oPjhjZYC4nJS6hCFaGfb/HR8SCUH72adxFgtbQR+D7kTRwgKXp7iAfspN237Q
ph+AL3lcbbWpAQ3N4/yF42waBYOmSWsrPe1O4iI+O8IO3Xw9gzHaciV5nccZA9nhc/pSdK5fBX9W
p+tMkAkw4OZnSRuphQMEu2Y4iqqkwb70I71BaJabQQkLbDbNkUVGJrFCrTdSUYVvwoLYX6122xWG
ETGIG05pyOGKEw22Q4r75GPWwV6gwB6CZrhAYNXfPsmkL6hzO+2/m7k20FHVwS3csinP5p1k4bMz
4+eBjhcoiz5Mt9QuCHFeLW1DBnc2jF/2XFPqsWzvcUzhxl3iaObX4T+EEja7ft6GT3q40cGz+ToG
uQHB91HYpXcKAF369AN4nkNf2qJhzZRVEEW94PNDZ9d+G/ZYVRcHoQQzeYX4MoZXHV06pfrEsKuT
S/urmyuiTyoMaSjDXi8/zFop6kCgF651BTDc3qQT42S2ainyzl3TVz8HpoEqhR83+bw1ZsFMmV89
R3iZkKka218Qof4JMDUfuu0UW10L3dkK72VIzDJXTOgdkTXp6JTxPciEMWMiWKgpGSi8WqLztwvF
/lVxzYwz0nqQPLHsdIPZVel+5ZBpmd2t6LQ5sSu3F8hIyaCiIQR55STfSnJGqE2+BBaRoX6b3Pj9
ixZ/BBPSaBHqA6W5WDqvqZgHgNVsyIYhnp/SUdMYYFmFAq6fg5vicIezGM/fRqLUz1QpWi/1xZji
lQ7wzXbR2aMOC1NotFmD7StCPomP/5u68Zglg7MSFe6DzzeGwy1ToQUZr8Kwii2xRLBhUAhm7SNk
Ib3X4S/3smdIqM4SJ8fzM/fglcWnTAIDRTGxLcJ9FnCeP0U8z7P9sePKHa8UtxZFaIvJJCnHOs0M
kpPGDOy1/bY3vJZ5XXoJHEmyJhw8ySP1swC9eAv6wdzEDCZibU7CKiiHarBzR+eZVc3as2thJRzM
kN/0MDU/gLw4GrShUfy0i6USIgtx+c4mQ50rxC+39XXvKT3RWuRkDmG0vvX/E0hX0oQDEixh6vAH
zs+YOLftnKC36HlxOODEkUEHGuRZNbIMt6UbAl6wuy2+S5SQ44DK/x7qSGak67xVCIJ8+fBuxnQl
XTU0x3SQGmoYt706x7CUT4qZzV6Cak+qohIihhU3x3dFl5YvIpmgH/PNrklBEeTbPCoqQeWfMFKo
648H2pIjAWrrlWpBHT+OvTpufazrAbwZAX/XOv6/QHkDYNzEfFzZoIN5343kxehqtqRBONK5lEj2
ZY8pAo+Sm1f75jhqHSppHi71/oACiBZnO37Mc4LDR5VqCHxn7v5NPouETij9/SVgxtRVs1mKCM1M
mSGnv/BAkzg4a65ZfEX8sdArWNaq2UUwkhQXsflIsCxl7YoWNMABs/AhIzP8v5obpQswTNZb+JuP
ig+wLblL565o7CJkK0Anxd0NH7R1v+wC9cYYq+cvFBJdVbnowCdI3AeFBLYy0c1Ws+glwsQqFqke
mcBzGTHwQFXawwRe61/As2CdOaVVpCVtzVqYqnxmrXsm/2KAH/i6c2emVQj4m9wzSF3YSbIH5hsy
lN6TiZopvE9KfcqSnUVZi33JPYo5kWPjGbj8Bco+5+8s0ocszg1GTBFtVN8aP/sY+9jywLIxnjOE
bw5fz2FOOCDHUlnFijwV/zI2m94dU5+Cu5r2WM27GMR/ARMhF4sFL8HvfLWWXjHvvQrSjRCadDW7
x42p7jaBVRInhVATHSRWAFX0NF7YnnOBreLhOFIo4LrSEh/goTlEiYw994Un/QXKc3Uyjf4U8Hh4
N8xNZphYj/ZPWE2EanYD9Alz8JO9iMvgesMGLa+jaaX+HbDxdM3gbkvrKU8Y9RmfHRK0i1D4YAtc
yHbotmMwEzG+m6IADmUY00diBbkVNZzPUYVyqbgK+F1geTsMt4tqTKmdufnl7kOjffr6qhLU135E
YA6YGHQTI4SJsxK+fQGNKqSQp4oO6fnBijCLydIdF5AO+2ZjCPiDRsO0aamMU2JaZoU26io6QqDr
TuIUxylRqTn0eCEeyFCFBVqc06/pxI9nJ2EOQPVn8RNPl6Dl6//EvRy4UsZbV3iM8M5fqzJU+v0J
TusSzbiR5Ysk44rGHClWK4YKOZWULc6LxVwXgoWhR82cHk2FnEnCMj/unFnOAmsp4id8yxqxJvUg
BaQTTdyzoOBJjQkoe6+h69BL3F6/aLg3DPsLKxr1r/9AGDdIPhfLdkoX+FD+yOgsPl+ewuFvsZir
H36SZhxzEfz96sfSNnOogHxo5Ew/YWL+sDqzjzn8MNGe2gAnRorpRp7t5DQbfU1LVfSinBo4xTYA
L6Psgo6NyR44CWmtl/jEEnpERXUKoSObfKkDEfAgdcUBB0+YBVQaZHiPxVJgA99vf9JP6V/WJZXU
BBE2i4ECIjw3Bt+gD7lLiLTcmmRQadHQBYIAXgDJ4rbovZNdsUrLrkNPHe8yzJlYccgjwK2blSCj
2Kh2+eqAe8n8KrguB4TIgNX+Qp2bP+q4G4PyzLMZZFvrDdLtpBJxPkibs4Ab0oR6JVyecxRnG58O
mIkFCM/4XgeFxBiY5bSliIqXQnWULF2waztsSGnWWKtDe+gUnawP1s3RZL4RyzQ5FEtmRmOUrTzE
QCM4SNeppC2Rcu6S9HDz/hDsMTs1DGuHjhH3hKGDlmZUWahbthx6b10N5KEfxj4nh6cdvxf16zp1
G9/iq4X1IjAFGe6FfxBxyAurCHiKklxSC14JxNIBTasMtK47+kCqtpHEf3Z+Ae7Au+l6vGBoC56q
pp4Llci8qN3DOxvDqYygDCpujzOcInrxeUj7bNLB+I3neMrb6gnG/oS0TBhy0v5DGoT00+skpr9c
yx3m4pO451W2GG5Vj5nEf9PV9AEOJgu0YgN6J6ilSMC/D3nvvEoj5y2Dciwwv94ZioQUTKET3DM6
OMq+C74jYiCaEjzCaao1w5xrx51CFQ5MiEq+viRVtzw0ExySR9568RlNhLUM6WhfoPsJBxNS/P8P
8jpK9HVZORvgKTtBOJjvo8C+cO5UW4X6Kh2Lp72jLCzN8RG34pyZPGs7M8haIaQnGgNfVDqgXBfo
tE9BsUP4oqlVYXPaTJOnFDGZ5QdbynFTCKMdBcnmzZXCNfUSMl8YDLdby/QVgXcsjwwfLjPF/+px
8HGgZldN06b0RtFOCLFbMxHb7Wx6jZ2J+m73qUlNHfiWIU5L4YHfE+6+rfperwgwc795gLoQAL8/
q10WVk+IrwfAePqPv598PW4gwl1ByVb1ThMUIJEWm3KdeZGcHv8pDOPJTi3qQ4/m6+PkJ9cWByiq
W1Hf0+CSi6t0NFDkPH818RcGnlOViwBjtjBgxruGqs0Bj+UC1WUW7fFmhvvchyucUKc1K3+BZhUi
MkF9JeeXCD3B9xaOM5HUa88VlRJjENvg5kquWEzpkhz1AQIEi87Jk9yRnECq4lFcL44X4WAYRId0
XjzGLP1iZHMVzJglIk3gaXppUErDTjq9jCqT9Wmbzzipmr7WUr3YNoURN/6HlWFkQrs4rcTAuvgR
QA6t6rij+KU5Ehc7eZoHzdJ4rtPborrVnFWscHggk2gRcz0So3Xz0VFVBlgpZpLNKoMpx1l92Aso
8ZAklmqhhH32oR2yEst9a/DKKpdfe0+2NQXR2KEq/JOGkB93ehJP4yvfXupvdvB2OuealLTl8EDG
+B/k0htmSpO/t2VBpgqyVKZoE1e4MSONLWqCO/5tWwFffnWXs+cC1HC617VbpF+d2wqFJlaqNBEO
oyUJdE7EtOK0EQHqsOUTGxqaVl2RUk250F8kesTPiurmbiVAz6ySrHRity/Xi1AZpixEABGI0wmY
0ip8jwfrhoWgWUElMZ4Mt6pF5Nk/idVmqPqT/+uHIw098gH+oA6rY2oMTLsIMI+7+87OE7yHxhnv
/RWc5Lo+of4tlNajnapefTVFxTBmdrsWKh2hIFAIEbAYX6FapIrA0L2qiUsXWABCKUfw0Bu8hsJY
YqjGNZw+6H2rNCD1euCI8RnKI8T3B07PeAoaHqI5zbfGEHcYT5D1CHNgBZhA0KyuZL2b4HuJWlpk
Qe63efWKdvo309PwnWedpOvapMgI74kod3RnArgTrslPw1ijxFkke/QM1x2YL0nWdyFsmTQzLBW6
kjaGte0h1FdTPBIY0Zmc7lNBMmw9Ru0y4fZpn6RRzBfy0wKbJih/qkZKkLDD/JFXZET64fhcD6Oz
LkkPpjgHUMJf/k8oE2AgXrHN7YR+AjXX1w9vPCxrmC8HeVaY34S0Y40wr0CxFTmha8OcvdRIv1oN
qv8FmtODkZDAwbXQNYkpKft6WHMX79aDCifFRW2R1z9NyOByARr4uceqUAKiVntMojTpMkRwCBl6
i2W10dpEtUb4Lfnf+qn05+iwWz2bGcfpGThvz2DNvaXTwKJbILASFgR7IgoYueOlT7Ayrzz2IlDy
E0tkNxhOLoV5PDMVdAnfiiW0Wxx7hBesEey2zqknkb2eW6m1DQui85ltazMWB/Nj4L95v0CM297N
t0Xs8aDjZXzJwn2t/uykj3KxITkgjvxNzZn67J5xSrQpGyLcNZUepSRnCLNhG1yqJf/Aa7rV1JxR
YjzPEzhlE3GeWHyK4DXj/J2j3dPmfDP2ZIJkmVXXFpNrcc7lMlAY9CByCCN13r61X94M5K2YSa8H
p1kJCMrFwywhFZD1TxAO0T6Z0Vf9WdAYNs1WvmpCcFee7JdSBRZTuTzZ8CnxoCZ4uvgRV1ORrHnE
HzgxFOaJHtaJaEjWBmBdNRWizm422x8eEz2o+qeQIpYNB01Q7zLYqtbGdVHV7+RoHYjVUoY7zEnk
4Y0ej94xSj8rJO4WkCm//p1T/EfXFsxxB0xE6n6+sEBk8yrcPiGLGS8gfvuRPO1e07w1OQ7Rsjf8
h0S2a/QjDwn4RRMnLfKdHIoErRlyq71ur+sYyz6XV0RUi3iI1gleWkTpLm8/6sxHhnqO8b/zY8nB
egiFFo6eKmqyu1Oa4/aO53UGJ1J+1T8r9zXAaUthSFquYHrzOLa7ghFkqpvXi1ROh1BfxX0h55tr
XLOgPQ3YjRYsdxE6ck4txIY9wwSLO562YIqtkWwQxXBc1O4OaWdgMSsTkb0Mis8EKwhdTDKt3a3N
OS9gsCHHk2Buw31cbDyGFmGKQ7WIav103ppYnadZtdHrwW1kozTkWldmNahLVvoUYoANY848vtXZ
Af2/2CNec+quPPq+ru/RjI3osgjw/wXJPE4TRvQRtAWw/H0+gyNfWlWL+Pwpf3PLQ1LiXeDAcNIG
Swwqvw9P0g06jDPbNGkxTYvV/Qvep66E2bSG9etjFU9gOaPYgz0ClvglFM9V8oNhko2tMQDm75en
+R/Q9IY4LtNrOlwaksd+v6/SprPGPitNyjTqkflH+JkaRMki0xnq9g0RvTcBasRS9LcItFOa9k66
Y8YbdC3q8mtvbe1/cZ3WJP6gUT18MpRtNhNS0C1wz6kJKVuLYfmudhIIfEmCbGear3tb/4N7u7Yc
v1W+NM/zb4QdAgk1csp1p7coLodQtEHKoCmtqzOme/k10v5UnTTuqzLxIhlceiZLh00QbWX0ucfQ
GO2fq9W/Evg1y+7PzXAZTVdXDUZEKd6Iv1cVzxawyZMDCCsTR/SEIXqdf1hbVihjUkUr2Lk/ytBX
KOv5nmQiOhMDq7K4eNIrGLsKPyEQE2SGdoW4IRmAq43j8pESpkK8oFkU3SK1qld4TYgsGRHbtgpv
drhopE7fX2r3DASLvKuxU9O3wmX+Y+e9EyTBBS842j/DsB0erD+FVnqwkuRyfhpToYmhLN/FPTT0
B7gwgpyqoGR9GssKfLlVUXZcbAMgsekVTnfeRZmZmbTW/gb94g4sDMTkGLycM7T106OsIzBL5qyS
sO4GdXRfzV69gQXDcOjzEYHkmsEa+U7/jlAH8H7YohkZifYl8Lq24zczbaP7wZRRmJmCcPvUZzEJ
QeS7oiUhBWNxu7pGu97ILGZqbUxnWvUuaAjAdoxP/L3kYdULA8XjDfh/0eGgmudrugZjb4y+ja8+
dASMZWD8s/g/Tn1eNrtYohRGD/AG+yf1woU/3bmuNt4sTcZoBeAwobtR40tg8ButAh1HNI5QG1j7
kb+s2QxorZS8FBaJzOCKHNvcR88d+aepd63bYaTPn6G7pVOkomWNeGzKfdBI30Ql4GryPf9cwmWD
6XhIo5cN1RaUmQniUS2OWCdqcKiMYHiDhDrA2uJB35QQK5MH9YnCvOf7P+rvwCdZ5xOQqekq9tBO
Ma/CVOt9KSobciPEz0p+qyPcXRCxulVfTdLmT9hoG3DDIpGMgU4bOZjOS7FD0+9cpRY7NMSzBXkw
7JuMSqOCxazII6o5QlsUy3d8Movapvsag28pPRXB/uJTtxJZwKzp2/vNtrYBu8rHv4z3zccgPQim
Kb7xEaNH0OQgjlscYa3n76QUwf65A6u8xdK2OQRGLHy4PjdW4aCJBr+407mtxotfMOIxWMJs9Xej
kpoCV2w/qmDjJ2XlBUitPenVAHVKeCvjwk7d70MaRJqAbSzoOzzPG+1Qzck0WICZFAjw8SRGmgLO
+yearNH6k3ioNQg/TpnaTi1/Q5WOTSZ3UYDob3/qo16yWFn9SGL4wLmOoSIl02kR7IQ3JrFHwp9j
FKQEJyUXuv3VJvVAIki7sjOiLEaNVBZC0aFR5bSBbYk7GR7DtPijVyHnCVNjIf0y0HjM6kQ9kr1A
1CA8+Bz7KqwjHSRdnOJvBAtL90JjDEZlbVuiGrhXiYT17gwDxpMnR8Gjv1JjyG+Vm0GHa8FQXeDR
WOjNjMacxEMrw3/bKvn21N5LMXcfyRpFaAOlki+fXzoGs/ty88amxbyS5RwNcbAUHUbufKAzGSbj
ueNlbktTmM++D39I/5GBctv9Tz53fpG/4g4U5vEGMCHKUNwySw2eF4Zwspg0+mHFCj9sYFtQmKGz
k961/lFhjjfohJkM4zp/TUjcOGJm7J7b37cfHJLchATBIUwkVlS0C6JMVwRM1+wskV5GFPRuFjUZ
Cm6dmnzNcw42gIvWlEf7knXKzAg7IBzlDacjNzSscX++sY5IqDN5dI7SvhiMHWVurXrCFu9TZH/D
1Ndvl25Q2K+v2V/kr21OWA0NYxrdhf03+KdYSEk1nSSfiz2Ds2VCzhxGzW7Z96R1XcHkMixh7xlW
ldxojj8H+aLkdiR4YE7YNF0jbaXfStIIkOKjGS9SvgvxUAgAQ00+Ev6YrR6kMHuCSiBMfLZkYRW5
UVAgRJTMBDLyFQoaNzKQrkND2k/hWqf8iIWn5fL35x8I2Y+YDuOcAxiH34rLElxWxX/v5XV0D/1C
Y1UO9VYemmH+8PEbFnQb7vJocFMhxbOtpltvI5qVuhv8tsdIC80atoo5IC9RSsECniWzis1/uNes
2yV8FWiq4V6b6Iqe7w714fb0q68wjlzryWfP66BG1LJbq1IRUJM2lSjKI5nyJvvZXUYJFzy5WLWp
L16+d+eEmv8SwrQiPVs++IO+JuWp1GNyXqSXGuIRTSK2bcWECrCO+WbspOnhQ3pmyma/d5dKtz8E
G8UHhC44DjHjiMkmKO5SkTjPU0ae4Ggg7PUe5oNH4jiXnRwy1nkmm2mhAy05ZlrCFq/nRaycnHPj
i6Bn0VC7n3Blyjh2TFNMS+gXrZoUTQIDsCLSRu84cOaGO+toovUBDbk+tMsRllCrsAD5m/qTwVyX
W2KrXWw40KPQASbHT25vKkMq08yLqueEoZF/lnYpsswI5fXbFgj4f7Bt1yoWzxP0uwSkjBas4l3q
DqbCBYvQYn6FAvyoxHb/eXzrztQ2t4xLAz6shoTWSurDWTNGTvNIei4dOqcTa3NOKOsUMZoon4bE
jUEEnzBkpW6Zlm7GyqDzFcmxRnfzAz648l1pMER1Qd2Tq4ONY1UdGDVaDmBaIV74MEvK595P2JkJ
+jFEREzvzhjMJekDy0jLrIP+MQXFwgqaHza7J3dvUAdMcjJzW9vlQm+x2SHTFin3Isi75kc0oCjq
1T3KyETrHX5lIDmxAMWtoTN4DAn2NJoOsJmtPPYN9Gm0SWiAhyB9cw3iZnRzK435fSrZc6hfzitB
yZFZfaHU45M2rhpkPEQCbcFmHXFW3Sz35ukrhIyMZhz7etp9iI604vhQsDPX+TcPQXJsNdEic/8g
+bMkCaUsEuVK6WSsbfjqjfFxo/KLNRD2oWP281NDjNut5M3Qjsw6wad+Ef8LKaiAorbaOF67VM8s
hFxcZLXfl1+EVz6SBQW9fJvHvFhL5kbkAMCNMJeKkGZCGiyD9RyTXkSrZBMwWwYXn+ImTKfl5TbT
ZllahoYD0UfeSRgHOOPTcov2hU30NtsMfxr2DJYmac6RWxU8OYuEDFWZq2NbtJQiKUSQsS4byVzU
f3e20PTEQb19Zox7Gmx88v+uvJggC8cCProqfsRulv0YkmAii9UUWbjX+ANrkKVHao4UgfjPlz+h
fKeltrlDqVKoh11SyfPNE/kPZFTtUbSE6W1hu1zOqFyElK7/zq8meJREcjaC4Av4pIFOSecQQ40X
Zf4MIbDjC9MyZ/fDxG3Vn7Bmb7fXRGXHrmVUkRBneuOsAlIplPrpu+wnboU9Yi0h9HDumqKLc/EU
gmzOkujdKyQD9CONU8x0QnFd5E8TnXeJcGUmIXtFNUC+Sqc6f2Mh4btxqWkl3lVc9mtJNu6DtzXa
7DogEkGkPEFtztCZQz1+nVXlFYCbsloPEFG8tK80tZ3M6+p7eIL6BC/eFVlVxeS7ZLzXrUoj/Wjm
s3bMXJNergeijG6o6cNCJkjC44JbRFIc4CpEBm5RnBzNZ96A+l8KPx03pHZGZukr5ZyE1eUm/wvb
7A/SJo7zZEPb3wQwmEOhKg6SoCBaT2ysRayQTRCfGdgGDdYJFVQK0P5P3/gz5rjF1XuqKwB2zJrG
CCpQv+DagFR75YI51pqLXKYRXPCGaGeXBnhiaNiPju1HYIFYrhmrihWYuo54ZLjGQSGIdS/P/vdF
+1XRKpE8rPtGPBXESJKst0KzscQ9SrAhhk3jzm30UZkw14A0HnnltY0NtVl0L2Nj7tPcLOeREJ7P
YjIhPcD0wRrZHhYUGPlMo4nnuNbHZl7+9KaupkTt6/D4nhktkGkFHQ1iEh0rwGq0mEkcNN54ajcD
wC9n1LMeMnun17ky7jmWeIUDSOmXtAAQlk5EHmvhnWAenLiqHLs8OkIuEpI1bkGbmGjY/v8QOMN6
lYL1sJRnHFZVA2uBZhxwG2dtY5lPfpZTX25uo+sNdGsB7d0E7KhDQtPVv6yfrV6kvVi6N0Y/VKwA
EHGIK7NayPbuw0Zt277HNnJroo7TpqPfMNa3kpfPxuF1pOHrFW/9+FegGqizF4djeQGyGfzqrxaT
tEiO3h7ghFKLS508HeYXvWVw1GBHIyDRHle4SBwEioVLBjM1JUd/Xsrde15z2a2AksLzj8898WbA
hPp8rn9daUJh6FXOI1su2gVF3WQBkmgIegwMxdpewaKZMj/vRKx/m5sMGlXFwQtBOFPpFdWfyi00
2NHB3bRrL5jGIHFU2wKXdpWcV9LR7k+rQ2Y5aEH19rr7EJXP4rVOG1paVqgzS6YcfaEAVgjl0Wab
MSyCuZxiPh4yoQVvuzHv++4v2Q5q260/9S1cHQVV+sqeqo2JzuYaM1qN/Z+XQFiQGp/X9U1IXtKr
7c1PGg4DAoOe926udShLDSfu8p+9SCvqEZ6YdXlWgGvT+n1ROUkFqv4KnxClE5X0bmsqxUi38H/P
Gueq1m5MbLUIfHJW7NuklHu2jQc68tKNIyOYCJpTgd9SoPiftL+3lzZwo9rp63uPCYHfyvmxBv9I
DjC/aVNgnUTbtLFMzoMQdVnIPhm2Jxo0Of8KfIbonIZdABaQFo+1cdCQVY/8mZ/ZooCjTIVV/VDg
USO6ZQ/TG6+wZJ6zftokSpek0QH/DoqfPn5Q/+lnMCD0IFyGEIqTGJGBlJ+fGImHDVr85Hme3ib7
9ISByvX8Gd6K/qy2Fqy/5J48tgQ7I38M451BT/b/W8Ac7/m2YREO4omRid9fe/BjARtg94UrQPBh
rVCOMS4ECryFK5aIKwFJYwZ3e1s1bqFfyLRZ8HXj53tk7KY6z8xCoQJdNsu6M/9DhJFfR8+bbL7r
mzxwp2B8CfldBYp6oQz/n7TSKm61eH9E0MkyKMYyZbyoW6/1E9d8g9WqK5wOjyCmThIGxnFMGemt
2LxjcSsZkuILCYGynOwzZ97SddTZNbGTYPzQ88vdre9f2LIYrToNpO1V5oGSrkV2Co3+l7G/26ZE
9Cv2wiQOCj539Ltr0ZRktf+GpVoYuGv1otUyze/BPgJCTLskS5DixwI+0Wc9xWFxazMgwxdf0f2S
mwnASfUYwYBNlsVqDkWyv2wGqgmkhWaDsTFElBl3fsUjybmv+hJLimZdvom9YjUTUxCdi3fjypZF
KcUlPCUvp76frEkNdiWtpU0TyftHbR+2P15k/BCWwKnZruzobfWEU+fGlYY9fLOzMa/TqPGBYtf1
NCyfeUi5gu8i8amlHoU8OhCtCTWGMBVzic98+GF1SOjgpbICw792Hs6VWTI/7KQk8qDsDemTDzry
zoTTnor3e4xhQZuZIW2ZcaYUpw9jtStZBTTB1YNO4J16+W1AyQd4Tu0g81TEnwotmjC9jqo/KbTk
pVn+u56NaC5P0OJuNCOSx7BYVkz6GBuwZf/0LVyGU98FG0l336c6Rd56Y+g/DzNZqhCvWUO8y6+f
lCi0fK/OcIztjwwi4aHXCfM8nwlxC/J1VGE/F+IipjphgVzOI5tmRHgyFfzj9ymfibiJNggsDhrq
MkY7avKohtgeUStdc1wuToEnkmVtE69zpwB11C7/Ut4WHgABUldNfzpZMVPaQ5KYwJ6+PiuulLLH
LMyAM0qADBPVPH10T7s77VLQQftX7GpDvVkNnVj1Jbu8McFHQyLEkOh1MunF6Ssn/f6RW/LdgjJe
EuhG5HBYGSGtM+5m3DuxicAmCX/GUHRBz/7go3VKprUwqY2E6RwKpCxNVkadmeY1W8QzE9qqJuvo
cpbZ7Hl4PeBQDbNaC7XYRsKxFdPld51MScFJll7g3xyvbFRJhCf7c8X18OXLe14Xn+47Sw+M9KsT
leCUwEIefXUfi6XzgB6aHUVOQdN3cOh3H+f68HB9DWN/LvfnRDDxElODmpuuPibOKk6Z++ZBsXqg
2A8f/IEW8IwTkwi64ahGsamVDlZ5FcZl79mHhbCEPuAz7V0fofMvv/bihNJ1QIl0p2UFy7YFKZTM
rdn7VryGsHaHy1964KRtQtbyOwgCZ06yZgH/iCeviSZCdMim2j9SQKtQ1SQmvVxqO5MpY/sdmMwQ
+I9SVu+ZZRPXnKqwn4Q9xPusBGL1bCiXW/Q+94xjvaqm9uYqShM+NAMvESBp0e6yzbNuWmdW2dQE
7N4AtF8S5MQuVyjxanyLEwPrxhRFOcOFCzTI8nGtkaksG9tq89Zymm+T+mHPjmD/5gEUEhuJcsZn
20a6F1p7Q7T5OpZvF2HuOZjSqy+CiQQK9LneGr6JGUku6vSDYYlelcpf+L8azGXLjfcn+1Ernf/1
DT7H6vPXG+lnI6psWfUdOSCxTiz1bIn5BeNi+4TZjvRxVxfKnjZ7Dmoll2a4IJSziFJoWdZNiBf0
bs+CD3QgYXZ79OmSRRbIrJBce+sl0mYevRHHGS4rgFl5dDJvy4tKtFg8qMWCekxa+i9KaASf8CO+
+AbMkAawooeRQmFqYe/ekXLnljKGJxa+gLZEZKmvGs3GyAkJW0u9k4ftuW3Xj5KOkZdwKW/sEuIY
Q8eJr6yUHQLZya9fgZNYM3PRCyX8GAOEELkNCyugt78MfrEj52ajmqHyzLkNujugJqUe73rSsN8E
RUGA9bIt0MkdBSp4akolreZwHYuUZFlO4S9mDf9l5byxsfL4oiro4505JE5khbFO1MS6xxFiloIH
S4KAW/i9NuhCmHIVLBoz9jVCJT086DF59qv+JuQetmqBpSsvgNKesT87TTXE5SDlvAU2p5BNcSiF
AR2PsD1cWzB4VVyVhi7BYO6oqg3HrQd9EsVJTStqlWiRlFTgVmrGhdexk3CX/50RBuIFJyPx/LUc
9Hn6Dwt0OFPrS67+j1ZERybuTtEe+QB6LKIFB8lhsRWfDq0Ql1SkokTTMzVy4yPVBkTxURMVuAqw
h0QHc10UecpQdVJf9tiDOvdUFL7o+ZHUnjkEumnXtAZapHRrcd8Ee52q8acR3e59chFcrNVY2gDp
vZGGotzkFbJrBtC8PAdkhWjvKKXVkqAzj8gMAp20z36yq4EJuc3XACHg3Xmq9tGD8sNraQVB5M1/
FX+Ga0XmOmC/ScMQ6KJDdljCync5Un9kq6/UTQkcvAKtOsX8GpSvBHtEtBiQsd7NFFivLF1Fz67O
K4KQSvPLYnj63qZk5w6/3ydtEc9qFNGuSAJ7skbbq3DqDsZpt8/shSymyS5oqC0/degt8T4BzZ9a
KOYkEk+g2B73BodQLkPnIOuQsWE+sX8GNKfESxOHDrru6bRqA9mON0XEN/uICKQRX1GhxaO6xfY+
V45THm3/Ko6XSq04L8zYBD0dm9DH46NsySjXEPtwEBqZEmfUK7kydGa2RH+IBDD7kU39zUKfgc82
7UFddwzRckX2Q6A1BwoCifoQ1mUFmZiIjvwq3eLr2N1rBCF7y8cWReKSNwVI7hYwFyo1rnoRebvM
fqMwtpVHgzcFApfR313A9aAtfM+ag10tfcSMQRF4sAHDhsHata5gYC4fE+PoS5x+J7+xGBhaVJ2E
UqP+ptBcoUWaC15qEtOjU94ezGVI4A9KVLNmT84EeXBRfDn2cNitw/huOlT8nJCCoUQ297V5uyLN
nQ4JTuzr7YxT/6M4vXCCxMuQVlBMsI+lV3CBgmRmhN+KMFywj21Msu9/zQpshuHRM5iPPb4oiX1W
gwIXl8W7aflFPHa/kIWr8MBoMKc07EOGPfeAu+1AWO+49vw1ZCAvTtsU5wO4/ErZjz1uD4a4hxtD
FDQoDMiaXNqadKVbSf6Tg0Oqbqy7P4X2hvivLHMTTXRNOlsJedMtaiEZGkEDyURNK0p4lwOxT4Az
vOJ031GUEoWAqdaNUbfetzF2v9pgSdC9xK52VT8IN81twJ4ZZIWgnsXJS8CzA4epvcdxBVTKzOKo
sz7cfwXtrJked0xBvRz+rHmHbl1D6lVPsfvnhuvuAykuEbQe4qm3JNcTNHE9+kKfYF3JyR7Vskm4
C/kfrmlhK+Oq923Na/SmtdF9eG0LKd/Fxbq3+YL2CWcTvfuU8Wc5MUqh/Bvd1vz6oyx0Xb3oC5n0
J/IvLUViXlqbku6ClXsU4aJyGNxgSK3X8WFMlS6cV41uHI8++oBvTxZenFXzYsZ3sIAjwf+8EuRj
L6jnxWioqs/3TzJHsKxuMwwO+fJjjC0rjo/RvQ8nl4v/vod/lxremwE8o7IOe+VzkEXj/Jl3yyW8
yvNiijilMNPyPS45VssvZ3elpnkC1wJMIGEISvrI88aOt6BNDr9THOxn2wvXtjmNlxTFyo4ZhkdL
Kw48j9gWoMUg8aOEDEQqgRYUSK50ONOmAbV9QedGX4IlHJZSKuVBxgvmow6aDmZw2NGSn/Vikk1J
W0ghLc5gtRwfS0yj0H4OJrVzf9zZiBhEFHqljsg1grjS69BsBBmVnUxjNhj9Tjjb9tFCb+y5LSjR
/MI46x1SOPsPtC4JkYwzGG5+Tj/aZTbjmeZsXVHvLXGFh/TEjZHYaLSlw6zOLt7dOD4dzEwDtfNi
DJZQlzYFaWC0WRMSZNLbP+b6Zz7eUCI6NW/qepw2TOItA4s3DW/qfxeCQXNQvGWzfQKse6bcAtj2
vJP/L20dK4wsiAyFYXtrgsakh1KOHIF38/xfJPyKhohVVeSxQfzu8qkbW1V4HlRp4pbftq3Gluqf
HSPjrKwBWOAqBhUnJ9F8UVY5oT5n61bA26RGueEpkooffVfFQYVPEyHjVUl4PcNL4CNGFzif0w1f
FuWf8uF48oJTkxzqyTtxi62tEDOiG0k4zd750uTVVv7hLZkaeHw4AHBQ0lRbxUBlPgoWLFUbB59A
JL05f5X0xpvnForR2cFQzMoehCA8O5AD5tTte7HDZfGnA3ZVacVvTCUo1ZmAOIDJi+/GvQyPFqu7
Y985V7ERkl6bSkUepiy3rzuSX/c3PluJKShP6T8b/f750HvwOaEeuNSuE7UEq6vl2abzBXiyGuwM
owRlMzDPlOvLTFCeqcRclQHKNZ4Zap7PYr/DcecGqWRj4oxzDJGQYD7dXqvFGR4d8XN8cK7YWJdY
7y4PRWs8YzIgNDNBYQjPCpFH7wyzUSWSbhwHwOYoD1SNmNIAPJFcSglEfiMVngmoY4/XBnDL1Zg2
niL3MIgaFbwBF/004PLFecwSFx8PXGbe1dCxxBmw+8bmMsk/r/FyBNE6TcoZJhjeInS5Whw+kyax
8ov6IBnkfdW1Fslj0NDX0yaCvWxEPas6F44kTsfy+FjZGLQ5H3inT7xXUSShIwrQFpu0Vz3FnZxa
sYBTLNsvsAijZv1zjWV92O7EjyA+MKHqLGoYYxAKXx9ob1EaPbrSrkZGaIBDQIk5cVhClIPxgJQ9
Xll16gPfcaxJbyti59YqXtozP5m61qb8ammWV1w+IeEcAWaqylcNsNrKFTFTMvm9fM4PzBwqCtZX
KrBzKSht5arrUUC2iQVyQgaz6pidXQh5NcQSAkiBmYNuenEDmjufpfZZo4GUdKVbcHIoyMSCPBSi
zB4Aognn8htmlvlgeowYjQGzvApVOmd7cGeCyK2/rkXTSx5aqzP8uNFAr4o2SuZg6FwTTpT/9fIF
/0v0TSpII4OhDTCmUghptYCuVCc9Fe5dtni6x9IxYCVK+oh7pbUjfjRH5RKRzoNSAccpGe0v4mnX
wlOlo0IGhh9N105NHyfOoK/CKnJDis3BjqfvjVf/Melx9dJF8cyRDHLIwGKjqq208a9nFhs+PyBz
TBmaaAI6T7ioBstfJjqV0Vzwq5YcKlGD4vfrHfD63Weod90j6kIqWFDFdO74jBwasOEeDwv85hwu
4DznSlYs7kxF4sSsbBHacO7yioxSWDlPu6EJz1Oil7u94whEJpNna3TGp0EpUD611INa+tKVppvS
oSdlJcBQVtm/qhZwTPSobxObptxgzRt/OdaPr7RZVylOrXF78QrdZDKYuiZv4jF9kUAh5T2N0p72
MdgVwIQRLIwOn+jEAR4wpz8h2qDsRcbph8Ot6Mr4khZGzUNcXOUhZPX9BIvl59fRaZP0kaxgWjI0
J0XkzpuLVJSOfN/PrZQFUbs4tlTmfr0XqWbtv4apTMx3MzkwFuBZkVgiw23UzNKEkrZBDX+DFpZQ
Zhw3b1SUdIYBccCUk4Q3XI4ECo1sQW1HNRl2SfxlfPvyiCao31eSVs0+P6KLk2IzBux/6J9aS3OY
Sr0DFra/wMC16gyFJooH8Hc/DyuuxM2fPlXCZbre/JHyIAk/N+elT/bJ1Ymk6BmPPVE21k5u4e17
1PcUtK7amvtLYHyrGelmmEp+M+De1oZwGJVJUpcVkKt9JtySmNhCNv7o7x+cUulLyZY7+Vc/Vwbl
Aq3xG0ycMaOZEx0vjSotrV8EPbotyrM3djx66hLUMca4gdq9pdnfUg5T1CSUf9f9j2JLADCKza8v
JXfrpMgQrHoNFKhfgOq8H1RPbhewowoZqJ8u2esxEqYlxPjLlyqFzBLoDYXaMiaAtF3UrN4W2k1Y
iNegn4uEbEb/Bhssy2m00pgZjJE7K+AmzTrrsMk1uhqJNsbGu8t/1wv+don138XMQHW2GW6mx+9u
DUsSYceH1PjajtJHSToEiQBt97Nla/PrvoJT0mf8MM8BeCWD10n1XP4l1XtqG1cMZwGyHPOofLqM
QEdEjA1SsGgF8t9Uz8PZMWIXsdEvCq8B4n8Gqt64j9z37Ygv4XOTVIwvsfspk8gGN/GGO/Ii28pn
y5+zSr5G+pUjjmJ8U8LED5ocX0AvC2kvfgkHB8puU94nNvuv5wcwttcND7oL/sxV6cY5/QHfWf2u
PxJ86CBizQG2b9/mJUwAnZQ/qgMPIODIisTGgwBFRSridsjoKVsAoNZfRg8jk9WgUrsF08k3PTzd
4Y9OWNOs2GSIe71EQCGLtnRyaXIe6HAO1WT4PEgoj9LUJYLO1ANxV2fmyPGHxDfZHQKEK+GxKljv
YXcRxRv/SZCGZFhNQRo2KiPyzOnQKJByp3NmIafWnS0z1qZ6nvxMJRsQBlh24x5D7n4/9WzvFIPZ
K4Z5VKFw+JJMsCzdZMRX0MjGHsuWCXf1v7OrQVBDNwKXTnvUcafSpcimXdREh3wDezRykPJnkDTW
ZmEaek0PaVtIdhx2/5im3wskQiOVVOoSdW4J4oWoaQW14VGg+xZAKNL5JgYDXrbDJKO/94+xCPwA
qRERe33Et6bOFje7/cTXzqcTBwPInzjTjcczHAw1E2X3OcYmDIKGDx4GNNOASGTkhRVPSldCgsp+
afns28eC7ZQdAaMDYpja93fFqFbf7AFIBylIIJH4qkZn6GXqQy2aUtd4jnvYVB+D/0CeR5ek0usj
VnxiO4SGYS1Scjkbx1kw4ozni3hq59MxsVWA0h7QMtS5uwradB1rt/Uc8L4TyUBJ0yLoDMvOeHHA
72OBmwSrBETULthMWJCUxdhNBk+hMkPsRGnh0n+5hkR1fSH2koq0BMOX+biN7a2B2G/amcDUdHcL
EpcKQmMc5jMbg8/Eq49RSDnmfpJaMkdlHhzOmYVma53G6UBgDtsHy6FxMoaIClekQAfKQUsBYPpV
UE9RTX4TwLV/6fl18P4w3lhsA4WBUcOMmUI0G1GyTP0KKWx++p662idSVoraNopy0yUxx6GnoJXG
JMim9RVZ+JSJCbNdjQCE8Mas7kqFAKIRiDFO7iSIU5oGYxI6RX5VnT3gi3ff52qhhIFUwCCvm25a
LSDxJcnI6k5JJ4UbKf6Yn1639rh/JVpZYtjTTlDLa0udugXE5C0Gf3G0lkC1i4gporrOODvIpCR6
DY+e0TAm+P1nBOwn/QLhGuEZ8cJPcIg2XMFbND4QvMc9SMB4GzMNfbYmp0Mi3fGnvWrfHz4cQW2L
00HU/LNrn8JwBlTy5SjvNlFEL1e1ksVa19VOlnq6pCjwKnMKnOvFE4vMizFgGqNWt+T0smHO7Gtg
L5zQjirPM6ASvvh2+PGtZ8Ylix17pWYDi5uyq48aAwV42azLrhVaAUeBMH5F2Wz85eHxpbRkXDnw
xqRdncKwjmj/naB3hyDWw7yNWChho4fMiPelmbzpGSnOmT21+QOyksRWJCVKhaG63Kc3FNHAHQNV
To7zD6hLaxpGr0MBVDDZuBXyfvEXigqqrutttR7B2I4o7eioE9KPEiyeMc9t58G+PDmlBQk/IEIx
taStF7U6tWyqF6KIVBF3Da7BPfhKsefrTMXPDdVxdNC1GvIiSDPKZgtNcNelRRNFZ1p631xzDBJW
VDLVq2cYNIYaYVC5vA5vC00SRhBif5+pxSbsrF7MtV3XP+NleXTJrbOXE8M2txHXM+DZHcFXLIY0
4kiotoZw1GdGKypkB0DCOOb7H9C+9pmQOCD3V8DP0m5JwCyaCaPdATnUcClgi0pjLdKQTsOgzpzm
kupsxELWN5/N7yj6U3hassY0rZ23Xr01RC2Re9f9DLPmE8hjnZXNVSxTRNAtby7fQ3o8VTjMEUbl
27uWxhEREaPvyXvwkyCc5ybJbZHmy9KbBgWp+gIACRLqKl8Beat4RQECybSe6BlAVlFWLQLoqIyg
LmY6IXrVY+UbeErCRUCHRQxjCjavlChi/Kbe9wi6LJ/n5hk6hEIYglLv1SKpU8gEI3nWQywO8fMK
rAqtm1LBRMAZOqZDcaoxMRw94XCuq/Ve23XFHeXN51lhkZQIF4/uSqHoIH2knG+78zU+Utv1hOUu
iH/IQ/0riYlImYI2taIjOH43wu/NuVEBa8XpkRGgz/rcct2uNsMzpboH3LYwauwt5GtkDFy54hTd
D+rjDYp8JBMxUFKDoYGwuX93UvMfmlYfciGohjG/v2LvmOjVQPIIuayfLyMijloaWyITyB/DPqnZ
q3cR2sXY7dX1+TF0JXbIiH7km8mRINj5tPWXyRvaVXn17/Ad31xv/iMNdIy+53jZ+V6XsoVM99lJ
mRJmvs1NniO/tRCfG2wOarFz+/0h6xz9kIHmLtUHLTXF3+SKby+i/hPa4kAru3UhTUOPpezHfCbS
bGJQISyYmoZ0G0/XCGSPkUmjBFK4TPLednEtb7qi1t6kufVm7fxM/Q14jdwwelHf6uN/LiesSoeJ
3WijO8O147hMZZHAdro7qTu8f0fRPtAhpqxX4GqX97MztOzaRd/pltMnwSQ5Qg2BFFHyhxel8zrt
dUB8LDIKgXqfibNgFCcdUulvfKtjKm/sl5+Rg4+dPtLW76ZuzVIbsg/wKQlb74o96uZWqehcQosl
ZsfPMeGdNxkqR36e/94qBSudZaYFU85S6YLM8u+XraShtOntSKM/RXnIbvrqLrwK19DPAOr/lO21
4QTAq1gfLwt6JMaYhsZfIl0tGvveKozGHdrAKKaqwMP49y6QQGm7Oiqz1mkb7vDFt0eTOT+dLRg9
ixr2BiqxohAtXICT7P6uuRjjWyKtst3u26c423yI9IKqM7JB/H12ZfxalxCM0fiQKiVJdPgXlkyY
INk+a6wIeK/nkLOKm4hJ9MLoRGv3AUz8gPBmB7QSABaQX6vuqs7lBiwpHPOsrt2fVP0wKUuhZgcV
AfpF/YZq/MTqoRGkzg9fSJEa63qB37SVe2bOaDXbF2hrSghoGcjyMMJAzMYLBp5M3WxVv/jOX5dl
g3162HgrfQfNX97eeOjNyE7HcrBWw54GwC+pFIXBJ/SO9oVd8F3GXHDTUTCiIgcoMhZP/BcJSdQj
gNwU5tt6Wu5eQvnAyGm4FogoGokAbWVynve4XiWKwLXcY28FR6wWtWSPCDXzj6+3uVoPR6LW1IU2
KRSuFbAk3fzfZVcQEGpLroY3fsiiHlhrXWQvpw/THGrRtHMCHPHAXfJzDhrbYNAWVpEzX/jao//V
c0E4gAqJy5cmwTwJwCPTUsiHcVkS1OZhW5ptvJe6MNV2N+KpKSyjir9XrheJqiDGGAnmnw3taHQ/
cZrRm8h6MHHx17WngW+Io9JU+KNwA3DWGfkCvHtOYws3sB0cToxE1rqnMwKxNVDeLEm0UGtWynHf
jiDr6Q+5zw2IKmsv6YQvqg9C/INSfirdgzG8GrgUnhvSyBUqy6hPIxpZQOy+quRv2DILoX6itIej
Bpgqy0qHH4kf3Vf0L8Yf2XrQCI4pcXb8WxGgAy6UyrimRrM7VhZQOk97IxhYco+AqtDr/USP+iZ0
1vXBvrZ1a2e1YOdvM1LRJ3zZehMJHjkQulfRunXSpy5pPV6U2OnwPxRMy7ydQCm+6aP9na7eSqe1
kbkRrVu7DK8j0awajokDnjyK+cv1Hi2gqT3AulRJ9l/o8Uh5D5w5NjqMmfzntnaTth6hw9h2vwxZ
nArNaU/Nt3JoL7YgVkj4hlbCCeJ3zCqIrJibCh+cqqwkwwCNAjZFuFFaCSGU3KQ8enjF3fvK/+Ld
orvkPcVqWVszRcxX4oEpM42827K7mQB0omCqVpwetqhVt97owdO14f+ytJrrRmgzfAi+2yATZIQf
jSDvwq4ZlcZmcNr56hqnCOemepOCyT3ub07CzDyn3XLE9C6YPc1GOsKPhUXHRh8zs7MoE1+fwFXw
iOgvAGvl+v0u8ejWwPpPc99XgxhVgcVUbkPz+kFj4bzKHmzL59YGB3si7JTzqmmOV+0obWnURVUv
llaN68fKl0Cb8N6EVsICbPdvf4ua+qj056UWD36n8vY6QEdZDsisV4yZQ937o85wR6YU1baTvYkW
mS7ZjYmQL/UTWre1Ybl4bhkID/A9ctA57g4hOcf6t5sSTxyAnOSBqBj+cTNpEXX3GfVDSzQBH+we
8Hrr5mOtRtKNgud7JRAXBPUbmiH0O+2d4Kq0mmIbPNXMUCDNGJqsYAPImc1dRohC9EvKvBeaaVhn
t4s6H8B7qrDhsk3SqsBztsCz3k5PeBstp7NeCMZ+0ZcH5z0hjSOVVJgiXZeVfmZNsh5dpSd4Arws
53wWJI+rDVCfhkdD4qoNU7zd1nm0BVSFSXdAA62Qhk2qA9gNsZXM7/NxdI+hrsctSqZmlhSWeS61
hHQSLv8NxZc+2YSkK5spgAXR7MBCOtquem+4AKeXYUJAo+dq0sOBiXoPhSG2bhkuQXBqhJyFo86/
IBJilUo7WyIfnY/QK25EmbOK5yMtA5Kh4W5BDEAtkIiGugY4hwP6KgF5p+Na1UUb2+Hfda3PSFpI
alNMOwmstodBfjuhMDGvGCZlasE2MWR9zphozbShPa9fglDOZbLfctACtBMrDjeba5fclr1UD3Sa
QzOYQf998f05cPwBC12yfzujOxh4T+mq+biWwjyC5z8npHSOETpvNyGVN6Q5IuDqQb/KLjGFtXXg
hnm7GHOK9oIwcVdNoN8W51Fp3aUGciLuP+GpEDRgSQ2/rCH4Jm1xyIzMnsy+8ADQFDtYBBshrvac
TL4sKwwWiU2aGpWNa8eJNI7YO17gU+9WQrjMpm6f6hBUQLwrSIMSG2ytGm0EerjteLtAszvyqBBT
CDX3DaO+mpKPx3MFffTYh89dvbvpyNN2xL8KQVKScNw7zzZFkZPr1doO3OD4yrJANmm+yFWz+p8X
z2nOJf7UuVr3tEiJJZZzVZFlndGuUkDHQg2F1mYNQraY2cwQ0EA2J1w6IwaFUmdRzDQYjLW+zhIg
3jFC5WsVcBG8Bu/LsnUVBlqcMGkvLVVE5sVSI66p89KvNqSRuqFj5aA6FK+ZNtnUIvN28dqmgUKx
UqwWO4/2fJo9/l8WxVHaNKBBw7FA6fCILkEypgpX2LF79WPjpinVsik6WrKytCTfN9eskSpA68Mr
Xw9gdyebeDLgZ6Z02DldEnEDb0EbQtJ0QbEHSWusYIWT7u5RZ/gfN5Gw3sL2UxFyHk/UD5M77Tf1
v+jM5DOsIIF/dxD8aYcAcUmatmFAt7eZJ+uOT33Hjs2XfLptwfE3ui+6BmFwvOOkNLKYUGkN2zuN
gfFFBmqW/ObmUVRNOgV7k5hHjXHai8eA6GKabLOzvWVSZVHKnW00zlZtQoQAWpTFT1bm6Q90rMmH
uceoUSwmVi/TEVAQBVMznadKj9O1ZCebFuArsCA2NP3ICPa9ghDFUfIv8F1ozjPPvkhI++XpyB1d
XAOODQSvsyq0bnIQX2HtNflYTxN4nzPX/JJjITkWPN37mRh7Z7JuDPqyyP4nWddHirDtC0DZwTtl
l7m+Wa9lGESHnvO2LMXbyHU3MK3X3jqJIQU8aK+LaSK0MKt6gmRnM/SnE9AO1OSr7YJC/detArTc
eCKK7tlznTOtNGWpgdZhn/9hPqCvPrbhxDLhZeg/hMgzqY4JfbSXniOi8HTWjmVdRzFowBg8eTVT
UautKSXigQUWpanuffTL2+9E7pnx53YQdWJDiBTad/aLoViEOcyOFRcobaFMZOa78DWn1q0sBkxY
P0YGYgKhloTO7UuqauNA6qn1/EiBtEXIYSheMM72OLu8+hVmiUi0/ZCp1i37mqW+pWiM5PcdFuWr
F5Zc3hbnhot62UuZoX/H9wfuaLpNCfz6D8riNqJ4rrCvejsT2KeoILpJ6QKvFRxEl5grynIJfsbQ
h1mvL9G5fp8rTKYX9usL7aBZ6Fxgs8OkqJjXsBOIUQ0LocYT8BCgqNkLGa32gBp+VrIcEg97P7Bu
10egf6pj+zaOAas9nZTNLvxS8PVxZA1X4AMqprC9daeHkH5rGuFbZ+5JZR0Iz1KmVesGJvBVczx4
i5Odj+LwZKW0PlY4qRBuCFS/4Ab29/406FV0x82eSo4EQ5sR3hwktB08JjGGGwGPdT98WWihifKt
DjMB67d4i3tc79Ju+nTFasPhHJZtls8jziBIo1oRE+3PGautcSadkuC3hPr+tmo7qan6//B+jK3E
9QhuYkpNXUAiPcP51jD+FLaYG9ogzie4YBxSVwOkQfhHP8d4zSBK67Zo6E3GQWXISsMEywpUgGhc
g5ZjOdRxpziomAIxnfIK0rw43+I+XKBtwig5N4rAKZhD7IIz8AZvUUfpeKAaBYThw5OSaABvU8X+
ezstVrNVEB3TACFl0+HVL7iytHL1EScvBn3B/vYqNgIaMOJRPBSEcVc9BozfN6vIHwdiep0qnlW1
UybFeTTIJjMMSSCTJzpSi9gAz2iihSKpE9PAT3tX23wSS96Qqrox7ZSxezt6QQk692mL3lrRPWN4
rLfRTo0k9+CkbGRrGT1P62jvzVsGA/++kNJaN+gXfnbMH9S57Ag4G2EJMnrW2bT2PJUOnJaHrLdA
ckDasTbrUBWBP2s7zwLXluoYYiqxgZqND6JySuvTGz2C7ykubjKeLSymnMLyR4OuH+UuQtVwZVmR
jiW4gcyHBEqxC00DTbjF+G6QrqtZFZa8aZEmqIuJ/hAiTKC1gQ+S/HfvyH+/RyIzAfLunuZ//knc
12s/EcXjjf88XUj45+mFe33c5ElsftuPHAtScemvp35VcXovKp+VTD/SIjx6+SkSliidrdFSQw/O
AO765vs6hmt4bOQB673C27A5ce2P1yCf7Ws7IijsqiIS4YDJIBmQKdaskfhqz9SqPmbeylmru88g
ysxJiUT8b8jyUHXWIK97331YCa7rI74F/Du0FZ3/gXjSVahc9LHMURTWlEUSKxjHLjb87j05GhWU
pZQLJVD6FSKjIoFnQlOa9ExyS2hBCWxbFHFExn0xpkoS0mH/T7IVgGiJZZh2lhkleTdABS9TKXwg
SYh6XKYViMoiYlmmGSg9t8PKBxLJqYEZqw5cEYbfnXgZz3Bl0iSgc5bW+nr6E0cqarLDF82kxbVU
VNeUfG4ELYEMAKos40XVfmLk8A5Y1Jn+YYZH6BrB26X+o+fvf9cDAszsnvzgW7rDJM53EZl7DQ9n
yIy8seQAkHS6vfcPfXAee10+J8HPLPPUtjKlkt8NZkv0W9eBhrr0ookIEMiw5V6VqaJ10PDr56Mj
hazIfHrpRYspcwSfb3LXzEUuG8HOGClEApuBCnz4nFBsyjwWWsIgJ9wwLvfaFqOgvHe7+8uAUMGM
vcbwjLeHJ3siywG+UH50evwbAB4FWbrISmwXWqfq1FUJ20pqzNAo6Ltda4kQrD8EYdhiF2Fta4s+
00YGdYB3LMTJBP6HeKe/D1yUDVzmwSrBjdOfpIfb5v9B+r7xYCmoD9a1fRV386CyQgUjdGkp3ozS
RWmC0PEyhF27yisjC2XqaYUZvQFXHbo/St4jhZlHjzadVV6gScBnLCQ3FATUjzeQCS23xfE18ToK
g509512upztyC12WMjSA8lyMEFRMIYf8naUUZJ6DxhSOa1XI7wPTYPXsF/qfDaYGiH0KDUyndxeK
iV++KRXLDIkq3gIx/FZuYwbtjvF013OBkKourws0wu7HTCcvA33clT6Qi9Y0ycjIOV01vKPtDd+Y
y+o/lAyOl73CKiPRYF5qPIq9dh2si1rNp0gzc1CxxrR4BV/Q5tidfoFLxLLZDca37LPqiIz8fcTG
PYGDYXA2JBCiYxvLszdMlHnZzMlW6fN28UYQSRRaXZc3IK4liHDsDNa2PdpvaYu+pLfTuPxIeqR9
2BmiDkexgUjp1Q5F2CDAySwwBMsspyBfr4Zf9kbyc36IUvk9NfCu09qouJ1fijY+JkGnRlftLM4o
dMn0Jj5fxuDysrVlgqPhDIBlAhZ3WRBXNeMpEqkpCq681Y7+vWjw/xo4E5GTGYH/z/ES5fwVeeoE
Vor5wkBbovdVimPo2VpS+sMXVTCqL6LnPbXyLdK35wa7URNsYilx5mHinGs59M9g9bguU8u92AGN
lQ3Rhr4PFenEecW/nvG7co8/GG8jv2xLyQBUawWE9FDul2YhlhpNRmhoqjdGazxCV4YZxxEa6n/9
rNoioKBO7vqqzzKzbr6iIzFS69/oCR28LrbIMhAmIn3TjbYzGCKcd6JLEiHmcgwNUybfeu3klt8a
VIJSK22I5CThTX3V55/ij/qqiL3JUOj6R4/TUHpySRv7NB2y2snibhI3BC4K6OD3BosJurhWQmwf
5sAJXvdg/cuYBPB4cGp+sCX8xje2wKN0284dvy1S9D2mVTF5aVEnWZDXWd3A8xato4px5MUVH48G
N6H5Zz+BaCrfVLKvlVBn439eG1RlKoyzG0oi8xho/s1icqp9Ckn1U6mN9+JePDSLX6YNgwLYE+H9
Q02QuZVCWLa8/JAnR2dR2Q/icp8tWO5G3V99rIkl9nqHTP0Axdly9JKSbMNjNAmkg9AfRCNQY+Dr
mKTj3+C78q1eWtw15Svl550WpQ4hRyE9Bre43eJiSwYc/kqCsI1g1ev2yk+CNt7KJJF37MSYTIa/
4JkSTuL/TYV2je6noTzzHVK1JIqNjRT3IJmyLwXRydvto3Qqyc+NprY+1kJDfP/RGt5ta1HNlHnB
czObOQJGOuVWmFFnLNtIp8dpJuuqjnfTY0gHleEpeYg6bsE/QuYGMMsy+lNx/rCkJeRuETLYmcaA
q21rry6r9GUzXLxXVVReQeNwfbDJMF+G2wDX9e0ZvhOhnO9SjdfJVLDb4WZ6yJS3aCxeNA2E7RQA
pw+F68fC27j8bq1tkC8kSVbquohTl2r/ySQTuDSNMhT3BQlxBToIoAP3eZSCWVykevFDpoeAQqHA
A3GcWgRK1XvXGD9uU8YpAUiXC6gIK02MZ7hzxEPvfDD+JBlaHKa3bLdqqd02vPXkrVUIp3ioGTrc
zsiiQiebIFwEKI2Rc/lXQQuoFYxgqw+C+1pQUxnIFRyht4vyF5GPsiYIWcxo9M+u3iVw5vOkQ4nn
k5EYPPfeKsw+2Z5t2wNabmO5oC90Gc55wpIvWNuXfhjHvMo5CmcFvLZ+cjQoEQOZZjPlnVpqtDXd
46+6QkGNM79HzohIolDJid54+gzAqScg1CHd8L/jWc17dwxf431a/Ts1CLGDFpzsk4x/5PZB5f3L
DtFcCgtcJ/RcNyk7jPhpMxrsFjFEJTL5s2388bxj/j4M+yJI8IKphSPwPrCzklF1gPRT6KanxXti
k5ztXDxNaL3K+iFHl1GGPYeWqdhTEf8B35B24iWDal7d1f/d3dM/BOUQbGpB3h7kteshlP7VL9QU
2jQprYHP//fyE3+KXQzoWVpNlLSOnro8v6TduD0Ey2u1PKIdlmIe4XuP5jSSLbRhuEdpFNz9ajUQ
RYSa4kmQdLRwS7HY1WuWKVvDJPLIABL4C8wSlH2K/uFPpbz/xecujS40h86VhtXRhDvOY6Cr9aRd
yn4hF535h2DOh8qmFkzqfkPVQ+l3KkX1qWhUjnIHVUsd2L7damenhySM4wcTqyCVNNZY85r3F+gZ
ZVFVGIAuM68f0G9VxikGuxKa3J0lcnqIlYZg88L8TUnNMSjXybvVnXO9zg1b5y7lZFEN0FyyTfaz
DpX+4xmlp010sdbhSjY0jXlRcQzmcUtAiY6Oufe2SalpIYij49NZNREobxI8KhyR34rKamZLUNgy
DOcQ2gJC58MiP8TNE5qJacFzRXo0GPBrAtDgtj4WgzoGTQLcUV+YYruDhue+oUlrBMVBWEUzLv4B
07qKTxFBztY/kbyuTA3LzVnIK0/3wf1R87aBEFrkHYWovLxCD92DlKh5Y290WG0KSaIOTyJ8yr65
rR3ILr5XAQ68x96T3u+siS9UET/HIznvJslMh4gRA9FaWbQ5iDJzQmW5y5cD02Gdo+S5yTW1Rj3F
EykrZ3alysu7QBOqioUaFRFbST2iuqviwNANc+ILufWuqlehiQCx7rgn9ymVX7SfVx02p5qPxAqK
Y68kJL+3CC+rSjLV60M4jtXjteCWjKJj8CuGDkN2/ukoaO8h3xmC7CC3FPte03NY+KtY7pJpbFcL
z7GxnHjgnXXYm/SvSMhiSSK516XAJb0drap824viGSgo0h7Q/P6u5dzf9iShZ3QmiQTlOTFzh8PK
sMtuEOeRnKcVRXZ9CUbq12VLsY53qcXzmFDINhL/uGwiQsrF1THwk46f0NUXNnfEzB/CwCXVw2Sp
lkKqJtQREbfZ1c1hfXLUDmiKcpWF+AU2VzArkcGdBWGoxJia/bnl3PLYGaiBZDKfC4/4Yt+NCumG
PEUpq7lx6s+D6IdtG6919SeQwdAMVrk7YeGxB//I5n5vMztbN3lmJIPmk4YDYjio5FE4ZmHmz+XI
rO451dM6lYuwRd+pwyETCj4GQuz2xUQvWhDhU+tmkyj52i4ZDwfNvW3sOdJOslcG+V8N/Ic9uLod
G1/NkJrG+Hk7o3819GL9/vEm8yJHVZhD/MZEa4OtM9jVi15ft5SNnZaGuVbmV/JOPYFWwch0FX9J
M8M6YUuRmZdGu8tgtETwU/bg6/KkxSQEqSjD/wL+CX1TJCi+d5D5ibIU1MpKmuWCX5udqZ3EuEQa
pyOtVBs6ii2711XiK195wkuM3EIXVPz5NHe7pr9Ac2kulF81K9CAmo1UIJ5Gwuv0Aqpliwecu5SV
MZ4Hga7EXKoQG/xsmxmqjDsRyLOaz9MA8zel3aw2vPJsUBvR8Q9tYDHCYSxG04SSFL+IaO/v7M9i
oIzQ5YXDbgf8MpB4kGqX5+qZddDiIQgXjMCFszPRBBu09TjeKiHBsMkFpLPnkJ7pdCaX7lJWnDhS
gk9GNIHI8UVeD4GuaZLfhWw3QyJUy/hAkZAfLoVQQHRBMsloyQ7S7WWRppwyOCMRyXBcdyQhjhlW
R+BDLRj7vXA+fR7h/BwbgHSEYhiU1v6uljHME0oPeIEsMUrMj7ui5NOfdWoyBgHwfEVRo6EH5jzY
HioopCftnhRn6e6madJUxXyrBc3sEL4tJrnJTCVukIDALQ+FlmFb0kS8+xq35NcETEUVxj5Um/5T
zuYGXLBXELGkf1tNL3FMsGsyH4cRz2tl24eBbEftbv9kbi8T/L7Vyl7XQfs6hABwuvwe3v68a4Uf
7cBr8s5XObyWfzS3sIHSl4yyziL3a6QE8L78D+7rLQYTWRQWtbx06ZwJQlayvNpm74Mj5igFz5SO
Gnoe4XiLaYZZws4pTcoKtoqtMIm3D7hTx93zWnJgv7KCnRD/Qle8LojAzfquk8SOdzwSDLgZau07
MBMphtMjecgvEP1/9+VHawruEobocSzbcbsXq35kdE6Sj0TAOK+w+w2Hn6CcJqjXzF3tiIM2yox5
0QIleKxaMiUD94MdCsFzWGGTWZ1XQiqkZsTj1KzD9USNztVLUxZTqYfW7D6HGQIDFQV6bhY5GnrJ
BR90jWLJe0OPiqwBgqYhlNbsdRlF8oopDm8xEPxbOdglGlZw3xnwmPcvUULJ3E5CjLrOJ+aH6L8i
/QtxYU9HjWqCZi1glE3avF28ibWtEk6WuAkoXiW9+N2h58YaL5WFJIgNnEcTURTIlur7yj4ugXds
uDKTEKIsYxGXFv4J/OuxemBw5a64EGCrCNyHKLkovAOLBk0plTf45imrD/Oc01EXY/NaVbxAZFyN
DcJ6eXPHvlB1mvMWy5IRVhb46X7FJCmpwwH8ekTNwD4tBjxgH4eE86RxBlXqxhhhR4gZTF+jTaI9
3FkELCq5yi0YO1ZNOnVGC0gmvuCVFe7mJvRB86TbAzMSPBQHKf6sAO5GrfEeKjZDdR6BYTaF6vlD
rLn8q3iiws4LwxG4zV8U8QCg2Sdgr7cdaaf08Lwd65J32R0SF4v9dMr2i1lUnCfsVCxRy0kaLxfS
9paB+EolBd6VtQ8rD/2nJe5VGioxL4QMSdDRsD5UzxtYwQN/eoLYCy8GjhKZHnBOeh67ifnHGAgR
mE/RehbpvR25pqIvLJKupBYb8SIK3a28uZCksfTMdkySW0frv579iIEHpiDwMwe7XkpNU121zMKs
W6ysOnrBiLKVvnYa30I2/2P+Tp+yl6h9i/A+cD6VZFYzkCp6b7rzw5yJXNmCEs74zGIxjCAva2Dk
+ElZSL1aZvAP2HnGP7b3wh8C/bwAHV/f/9ZrF86hMjKCXNO6jr4vx2/4YlxC2uURgXA/1XVTt/cH
tecgBCU3qvjoQw8k9PlljgWzEogkWCfP8E6SXwpODfrYNv8aGiVuCaVru96zmNeBpu9HHkaAesGG
XvTqyipDr1611QHVhUkyzBcAiRmh+O5JHrPHiPbGLoqxgu4YjM/ez/icj+sv3iliFsmjMxuZELFh
zV+DhRGivAP+cKdD1f15we7oq3GDLN3PUabA3tTHd4jHxzDdIL93EjhiJlmEwbxfXxEdLJa2etPQ
dBAaJ/5i0RCiS1KH8Utv4DugU8bHXLG4U8BEkz1GBbUxBSWiOTJndoTaz/Pe/z8YCV+Kx9zpshIS
U6PpopVE+5ZHwPER6JhgQAcckRmYwWkDLibhdHUps0UPGfbLyccUi4Y5tl6z3ul4KSIKU3R2pST3
jvg7KVi+svRICZ7I1mfEABWmVZHg+3rHhQKrLXkuQjZMA388OmpcsHajsHnz7bAX6cZVaOEAYVr7
yDQ96VMdd4bQJsthH0zRcph2HqiBs5D2WDseg+pa3ODTqlvXpLon67HJjfSsYOHLRQxXZ90cjbIZ
+mebOxKgzAj8g8x9MSOj4jlNxFhLbD6f5bsMlS9lP8c7PKjr3hOKQQaFEqiv9BMiCWWk+iFGiOKj
ycrFoRcLaA8bIzDbFWb9Rx1D6gakHkRP3mXVzAVDK8Qf6fENnmRmK6YcxXhPfC09p3YVTHe/Xfh7
uSnaAR+pb23ioqlTsQ3g1tU3SH7d3B98XVQ2o3bXpxZACOXeia5sFTUcfXKt6PM76TwYjQPrsQq9
hWjJmBPEDGf0O9e/GPFw5O4aJTwzC+U+4uyjCflf+DO4P1Yj+mjK5wviIs4fuCTkIR2flbSclLjr
Z/1X8b6Eg6HDtaZa8krYc1T/taAnkH/QyJ3P95HbrhOstGU5+F50Pz4UoeuuEh9fJAOkqgbCAEgk
K6bW/osgAMwhmLC2dCeYEKZxC7oPAJiPb9NtSH+mpqN1GGUuNSQkiDXrLbXFi3LDNJX+GNUOhGQw
pbHUsGzbdsQufUn1FqYQp/E6lFh2H02NpfdEzPFcuxGo2Zw50eYTuXVXS5WnBd4eaMZqq5TIE4s0
J3sNjdoYN/rQDTPpwkaIcBNPD0ECMLkcHNCAMiroDsqxxlaqyYlWuETog8eCASel5k85WD/2H2qO
51jDoikfTcqwaQkQxIvjxb4umVf4m4vypjLX0dBSIoRwsXQuNJemfoIwninO06r4wCAlNTE+5Z+s
uSJqzw+8eKSDOGfROGeA1akFofSetNRL/r+iPPnZ0sFWlJl9Ax9wUs3nUQj0r5QNEY/ytvRbuuNX
l9vGlIwCdxYj40RRVqDnkwV+PnmHaIpMgL1tJL/aERqzZurNKa7LXJ5n19c3U/t7428vikH7UDvz
a7Z0moNNfITaedqGPOmBn2+0Es+E6gXq4uRbDCfxvNZcAV3zWXWPFxysoAQzHE16n6PTdSi6+VYj
6HGxk/fjS+O7F3k/zymspT63QF6f/pipRk1kvwfpNFcWjJ7EMWpWWP2PhMyElj+vqVJYsqYpIAv5
nnaCKJHDF3mYjEGgsP9QFgdEFXolMRkxWQa5Pqq8te0KsyJ7uehrASEw8SQkOCNRN/sPAdvEcM2h
dbA6OtLUsJj6jp8EPUcy+zsp+ZBkOZ6atXaD9mDAG9qgim4Td1QaBy4EP0XSqEE+IjY1aWj5WIGB
CCw2SrxmuW4JlPi9cp0opdMcZPlsK40AX57+ZWGz1gaONM7PoTPai2mMwuXsPuFv2gRSHbWBuvid
vzPcVsF9AKBE6L93Bu2q53H7P4gUyWB1NcalSjFkOSUw1fFkpd9+yCDPqhGVlwoPbvZh88A9qPBE
Z12JZSNEBf/aqY/hr0hFi8Rse6MB6WKmt+AprtO/WsNOx/yehv3JtDNlYMLfpzwbGAUQuPpHCfLn
z8JKlJ5Cd0bMf9iNeH1nDrmqj/eCgtvpq40cXZpZNUD716EwzJUvJao1/gIPKQ+Uxp7nhXFavY9p
jm3EmCGZ0OR8B7j3f/fZmxaXYh2ek+42NMt8YgwJm/P0Qn53d15J5shmJg7eqJPk7S+H3eLMNmFa
WXZG3FkyVNFKqU1SnG/RiT8dHOWgJ0IXrFhIfNZtf8CNIuyKM8e88/OKG2X6gqPf/5zdn5AUwB/J
ODcPCGN/HKddetpZYMaCyPu78943x9Mob2JwGR4PfX65XdevDZCm37KSKCbP2aW41+/Fk8QumVCk
7RKZgLtMje3ob01UtboA3juFIpnZq7Lo0ZcJmFIZZbIZg8TtqB1umOTyX659kA6lFrfl8NJr14sU
TSm7S78OZOKJNm262z6NDkLW02TCUzMGTHrMX1yllEhjBLuSxJ+n0v5OYHohouFcq68kk+3kcB45
0ojUcCvgyGYdFoQe1VMIY7a75hYsAbMMRSndyXA975OofMPMma0geM5ZwOKL540Dnb3lYoum4TvN
VjCKoRRTnBKfKzd8SIIT7F8QZFnMI/si99IBxTI6QjVA8PzAOZxHxN6p5Dgi7VM+2JRhIHwdHQQB
ZGLDO7Ncz8yArbgWPC1esYo4Y+0HbAckmlZWegJeilHAYoejjivTVrRtBQizD+UcLDKmQHX1fAdk
/1AgKNYg3nd0OR58O+KeWp+06C+EKkVnuldobkYB6ONtkKBLCPd5V4FjD/QYiNuw45NgKJ7lKAVt
vp+NztvfV8Qtb9FK9N+3URwSAefoF5hjgZLaPEJcOeaHT+EmvatJ8NG/0YTEMFkmIyHphVT0rWbd
mjBQqC06mrrGnJieqfCQrez6ysEOoWGH6wOLJKrHF2z/8MH9MeM9OI85rXvPt5/HCSN6dQu9mgAS
YbNExl7x2j/8iLbagHE9MvkF9zaEybCAoH+GFfP3nK5haH4Q+zbdIhu2LKP/N/GbtzsW04H+bChW
xDkkwGeotDjfsA71+1cHHXdJfasS3SAu82VblDC0CYZXgJrtg+gkktWA/xRHxLctL+LusRnqr+RO
cWNSoaXoxHxzyEFhFGb/VWcsLXac67yberXkzLUZX5Sl45qej3oyb2lKVBd4NOZeP1Vubu3VzcjY
lpvNNjn3awXx/y6Og2lJXSCxQKp6Xgd8d+G+VLGI09bKfdSPqWKsnUVLFuc7h/Am1EEdDx7xpEj1
JV1o/aG0H7aywzVK29edNXsvx9aW0UzwWlYJQhEKaFRpDnCPvGkUYuAyft8kKILmI0m/qFQpt87G
M+lBJkjQRIbY/jxIiYOlKAxaCMOPDcEaovv/Wuow/xEnp6AjyZEqtHPBMAGrhvnGsyauA7YMBNNo
RtV5uvsnAacEKYvlIn4YFOk0SIxlyFnMZOHYrneg6hr4KYD9aQIWq0zfEGdluNrOunQzFwoRD7YW
mJtrluZRsszLcFTKJ5xtIUu2BG3rcvBbVphIWScy7HR7dWiFBRBQMFRYGcgPhOJuQ+4QV8pErLRu
KlBJQhs3fHdaVqIFSn0KV8UTLJzEWY+hjVXIzYtIsBFjzmlZ/IkPuCUHWpynP1WlPGOywpdIurIE
a3I7vEi99s4abXDbeyluT5zTtcjp/apea0IlgqMEKSv2203vaXaqzaSaKutQqj8pZyBI56MihRIw
yJXVwI0HfKgOyiOeiQGN7JhZCrgk9Fw5q56K/w/Lg+hMHeQtRyZbrFATcdAj612KM4RWMhrgt9Yy
AE2IYr592QwhQduNBjoXVYzj4UpQn8K1m1HGRu4nV9DQ5gGg1KeQXebhLw1yYib7pJr6GElfQUwp
rPRdqqqBHds1t/6NolfKaS15tPUUaRpzqEUkYUDh7PKAFWZVHOWak2dLTJJQzFHrEHq8EotM35Be
R/KPzpjfcfgdFkVSjomLa6cBvCT1sw/Aa/CuJF64442ZJrLFxKwWO+6MDqaCBi7pRlE5L02YMXUF
ZxfmFRYtwmzaZ0JVBDloPmU6GIBt5Z+y3ZwRX5pOp4p3LLNbLYPCt8+AyO9zH19m9MW3mJwEPhzO
5nM4Qf8YrFaWj7Orm2JwXA8VAyIvpQ+cl/H0j9qYoe5pIv/QbBU5IN3j7FQkeBgO/IIoTeZ8NM4Z
RN6krZnqhiT5+94kbIpitPDWd52Ez8MVSSEUgZoZM2FXMn4ZNS7t9Q9wgIQX1O8o8vbdGUx7Zthj
eKMYEWHG09G8BOp9veNyN3ZWwsY5ds7XsFBWRPapsmsRSduKkm/jbEnpN5ZiIF3G3Y+deZBAFZAV
VegO7rl5AyHShHJQ/hIWi//uJqaM2akbgBQsaKfCm6QzcEH9YA+b32kYQUonrZhTPps8yYazIPi0
yL0HlcffvKJOktJzotg4TsxIos4efg28ECvLyO/hAoX/TxJ8A1sOXLehQGwssA54oLcDljGYzhBF
7z6o8vFBcIs3N6fXu7KCzBft1tofYW0L7UrcqmrQzNc6BDAmHYvDJJgG5N754ZEo8ZQUVxlsTCO0
/J2YVC09G6i2VN3pfePaxXdr8Lpst5izP/bkC56qDQcsQXFOWV4Px5B9zsyBCqdBBkBsfvzkMJnu
V8gh5llxX06cayvVMONO7XjCzKf8nkcIHiZeUsxlW9yc8GY6lcUxjck+BZPObit9lPCJCTR+ZzX3
xPJOd9pVbf0KXMZ8Dep0NQTtszC2/sUuLF4/NUOYeqifNOOF1zyA/pjSsIfx0ddTNS/DEDpMaSvB
nzXc5y7YD+sryCu+OJUjKZZiJmUGutvfYStaAR3y+9GXVchMzYGgqkXM95ye/AaDlOW+fhjBZhE2
lcAHJMGfIdjOJku9Ao1IfCNHRaa5fYCfJv4mayvd3XmJW8Zs8NYHQqiRTGgWMe6m/6n/26b8CfB7
BC6BRjby/n1+gF/nem4OqHgut7gR8khAfkQOjTy8u6xYVguEVqScdlGc8Fx8STTJY50QxgHiI28B
fuBerEkWzGUIs9lrr6MMcTpQ4a3yEojRP8zX12H8YhKCDvR4AcmezyYUxYBvhNfuWFNf+upCnqJ9
joaFVq1djRICoYsMK6VD6OdBxy46DdsE3PcBv8ABQu8r6ekDpGGKdDjxNuWYHQm+ULA3VaJusabT
1HUgqR4yoW+Y8gEo6TuydcF6gOTYWxCcy8uo+f/1Vf+uGF+K6RjOhJS0tl661sSSzvgsOzVpqeU1
9Jp964cTV6yXqdA7ZWi5MLvDen884Hv9tliQNJO4ztFkYAhyMipuks7urwuR1dBnypq/KTexYtb+
A+WxHpqudIqO/0BfOBpE9bbEvHr8Gwp1d362hroMzv3DLRFBac7UJUmy6NplEE8HNeOrnzxPK47/
OEZUcRpvVfB2w/Wl3fVKnkPCRmXMRTLXFB11D/OsBNvOxvcBSgBhOPp7qvOcZFuSBKLpJrIef+SS
XyaGOd2kG0GEzY4HT/I8aRtWnIiXuqyUENe5hU17MWVK87vqbTVtzc3IRAgylxfkY6nN1DTlG896
k/sRCQXLY9KoL/DYIpMpxh8RSDulIt5muB2o7Sd6OxdGV5qw3XCAkktuQ3MeaLwnKzb0I6esi0sa
902K0MRBIVpcELfrg+STI188feYGqiuZbkfxAJMyV7s2GubZLtp07QlHFj9om8IPJsDTwUcx8kie
ePrT9QrrULzdTEEnmyZYvH4bBn9QJ+a7HMeD+tSf7b6IXgRdZrwFueilFpgZ9o80Vm9XIfMyAItH
Fcv94oIDYIDpvFMsRtzbLNv4J/qPg0w3JnTxA/pWPYhBgKYBZH9YO1wey82kV9e7I8TAH1gzTE6m
Uvr3e5XCFIlehFcUMzzE0RhSDdVtii/wMpWATTwlYINmPx7eNh42a2bkiC6jvzRwbFFgConYjbY8
/nyyt/SRcPboAv6T+euMEQopcyw9A4WXnhPbSEqgE6zf2thBJaUqOVHucvG6PRniB4MxxWOxdrS/
o7JhPyruPz8Ju1mwc+XNk08v5OxmTU1CrwSefUAVpxHiMYuKhMe7pJTOWQH2RrlbAzjcvmFSW47e
Ah/Ceml8BWxnJspbDWHEhVvzyjBtrcDNNZ2WvVt0Qccm3/N2UWVZ7S4Hn6myLuu6l3hZjhNYCPXz
Dqq480pnVPFOpA8hJwARZw8KoeegESDibSGCzoezi1eZMG3/jzdtWmKviZ/8aalVELfPQnZU7Dvg
GO7GDYeUBqBiGpuHSMHqneexDsHawHE/fkJhnmJT0ON5yXIuvmKm4Af0nOU2o3eXUUI0K8FY9wDC
r5ynsMpMbgDm20a+JFttZn9oOzZQv6Ul3vSsjGiUv15Fi7CIcX4oGhkbOk4VqyDs8KrXv0X1E0sE
JT3/eN9aRWCG/P8Wso9k/JG5OKRZd0QSdc7x+TpMwWiifSl71hFJseozYhFIJdfVq+ltFKzHvzYg
uvgE52L4f9khFJyGbMlQ3sv5zwDuHWgUsjUG/OFRZC/x5jU6FX6AAezbcKUcseIA0XekXGvL6Ryd
iGLCFVquPViiMuN3mt0JSaWQdTJSJF4r9CqAqgXcxxmdRaFq7FdXR87vPor+UTca7pvR67xbzwsG
YjCvQngTNbs+F5IT8KfXc37yr6vvTr+IPLIachBSz/aE5blS/NgcBen8ovlrMyD+xxVeNviYWCCb
gA4Owz19mCk42I3nnjCEkqrdx24QwNQg/+w06hw6/aV7tlPEXy6itSRXUvMvFw2D8WqobHD/XZ5E
Sr8lFuuxugPY3cBLH3YAPv7o5emhSOgqAp3FJoUWSHtQHH1HXxPkwDAfF1x51sApTFqect/BxZfh
PEq7U1Kcrk4+UrJTi557QlCwUvft2YkHMmUWWkqbxFPQK30OD1R4qzF/eF8vfJcdf08ZlVsaYAdI
QUTnWsVh+XE4/vBvEzh4UZLt8TrJrhrbzwotr8u1m6GVVjwkwAgmJEGAMU0ZkHljO3FGHImRL9D0
w8P1f1cKNfM7XzHU+8AWC1sInW7wyCsd1mQ4JpqaWwha8RUiyY/JoY5D9WBpZ2efk/f5LJJxUm9Y
pdMbyEoGpdRfjVM5T089HBApm9GIqsO4IlH1Jd0+yi4uDrt7+1PKaL9QaNn47099jtP4oQE5IzUI
Ukp4LndOb2UqLB+KMlWMkoLEiWgKSV4YSKE6R3FT3lFITy3ydJIBqH3Igqwc/a9vQPAzSyI7sSAM
r5QJT3CnS3lGHKER+kzcp1jutmT9d+rYi3rMSj6yOcBJtpP/8hp7ULP7BRJIiPz7mhXTcp5PDPWf
XOWcM8s8itu+w5GR0z0UZCnEUfB/jdXaz1Wr1j3Cl2axMgwyTdjMXlhw3moLHu/IbwEeye1L+68x
a7cytzjkFrxk481h+91MEll75xhJiqJAVuDcKuM1UL8OoNjUJxweucfM2QEvYVk/UV077iUYuk49
S16cbbFntsBaiggE972lsGO98zWMtz35wHLGCyWVAuH8OoLOFW/c9+IACz+Pu4/b/vt/AeTHY83V
qJcSjHa49dB3LHp0SaSKzXQVr0w8StTOVj5Qvaievl59WZoJY9z3qLNOC5+hVZVz++BwVnsn+sbV
QksDVOrJ7vLK7bimmPqvs56LoSVX09VL+wjEHDvhtygtXdSdOUaRIv2hDn15PZz1QNArmTE/YNg+
Sfk+6KyC/QV1YxHOjMTyZL51vQ4I2hP8UjNOti+iX4ao/54w+omeNnSXOtOriKEWCddTJpB2Q46x
UWHS1brIpxx/3R8v8d80kErtrmFS9rQf7x85W203o5UEqhOekQXKNi1+DL/xx9hBuB8E+Fh69E0R
czieJbhqUe26qSbVIBPcc8+JCC6dasx1pkU5a7+O03CnUqMrAGguoglWjHQKEMTYzihPHb6uLRq6
Tej9Nd5RenixisjPyKNMyu/Ckiy3v+yoITZzp2mzSy2YHuEtz3dMax9i6RnQOVRVg75Sz+rKd/7e
h7R6kBSQ92UbzdyERlH0QKiskQWOMpITBVT2awjCeyiG8ebYKm5skGrnRD6tvv9BLWkaaUd24PPR
iQP+ibw7GYTm87gTnXt9+nUzr6RkqjJPl8voXslqOxfwbtzFdA0WvnG46bjoaMCk/gOFicLlOHgC
8I0HbVW+L/fYE+Y1lEp5/DTmRfZaak7MU2DbHBINkyByIOzU0/87xa2y1kx58Zz9tQL/bJmNBAw2
dkfOgC1o6AUgcz9gTuHnRi8smwAY+X8BJdx2y1IVLUcDFZteclKq17FRyV01pAJ8dRm5vll9PhZi
jbp7WoCLEqRXm07mGeZUG7/QCG3oD9rn8jCoqWyLarpHN1rmuRsA/PWb7xaQN2KCsHZJ5GQxiJMs
CvPP6T+dCMvq4WyeCI8M+tUFjr4sW1PXMa9yGdYR4vxaH1MaXXAIMK+AhhJsXif2t1raoZ1PMBhV
5iXpTlRZWsno8zuH2CADJHOQos0RReATN3xF+siGxVvb1xElCVoJaib/plqOEjE6y2yE40T/FyBe
663cQKTPIU+VYNvKusuVqSsBKtKsUp0O+Yx4yh6MnhJjEyURLKWBmlLYwQ8wBxjf5ytNkcMfndTb
ovwMbNb+cdigsn8qUAPEQx7HIqcDj1kXivPVaLWklUUCNi2k9aOg7ofqr3sYRK51/5Km9ZSe4Rjx
M0ENQFTf/Q9ed3s9aOSkXYCRa+NyF/WFFZE/+avCWPjeowYXx2XtjMWuqLfuaS8UVU8c1m5tY250
JGN6DhvyU8vuvMRF8AZ734uq3tk/1gg/HSKUi7Tasl9bLCJaVsVim5Q8NyB436d2iLIC76L6+37r
DXW5cCgXrennIPEIFDR0f777AzERBnmae+CdFEM2V3PDkI44aQjx2VWpHO+qUtX9hg6/leFkqQnb
0o+HgjJOk8uoXY/ZfiDD5pprrP4UERY9mXh+qPdlMKDlfNyulgEtWszyoZ2idyh3TcysJLAxTspg
3n1LRBRLNAGsKcC8Psbt6dt1o4/UopbDDdXuJJ1YnaCZyJ7/B6z3MP25W6GC0FYK8+hj+99A0bch
FxDZtZsw8rtlLGyfzyLZzsmVLqoJPiQzR87s9wCrmB1umgYYpBVL+RJ1oKuzHikimdN6gvqo6Grb
+WspnQm2STj3pEawOn9mX+1um5lOGRjiMdavaBEFldwhmJTJ6do+r3s7coJl3q4TMltTOicRNeMd
RfyhKrCAqgnssiw1fGIWxGDje3SWvFAMdiS6LWmf5rMYm9ZoSOIcROPZN4jIgmOhzmfG5YtD6/Rm
u90oxJYDzCf+Kf66X5TiDOXO+Bor3eagU5Bx0awgyWnnKHcgfXRd8LTDUitroC9D0Jz7kjrCPxEA
xJzAfwBcOcNIWT850aCi3FFhhk3GCEc/vj4d/K9FVKgvpW658pUVbjz6QThTq2ZpBm2EuNP/mSbI
jxK+6feNnRXMeagqK+saQMIFQqjjgbisarlWA/2jWIV687t0Olqo0OKgfmdUiAQxfaALoRoA26HM
Gdz0BcW4TIXTZxBtV8cNdMPfnjXRJk56FOd59OTDReTJShsYikFYB3uI2iOMX+4Y6/vkOC4qn7lI
54Vk2HI7rJtD4ATEEYhvfXtHRoAkD+fGXOFd3qwGWMdpzmTdS7zs8o5F8nMYdzu3uVxZa0wCcSEg
0Hxag63gNAEr+MIh7r46Prl/Jn/D98S96mMC78J7BaUWTyygXi3tgU12dpyiSW34J7L25RhZk89I
h1EhPPASV7KzvzRuDXeDghejDTn9R4757nuzwuc2GRccqhbb0MMXRnEZiRwr5wsoixf3ofvrIz1y
s6zn+vEVFLujQx7qjYjJBjtDVHg0/Z1YjSyzyvS1JlyIOEVtwRqJ9sRp2VexnopoynnKmHUrmfBj
toCHpws4d/8rgzu1jH7r6+ilWFkPxJdyQA1IHYSu9PXk7ZRemVasYq5VKkO/PX/OVzT+ZYIof2hB
gkX8Xzh2fJ+e6QKEoWN4i3TER8d+Q570UxXauoApc0JxHvm5f1QFbCH3CyrB261V2JcEpcmPiXAV
PUo9xaQN/RVbAZRdFdjgI1/PoudxvoiuUZMB1hYkHF1d1PbAH2pbaQlCV9znMgBD50RWFvikoM7H
9bL/d+MBaID0aDDOith2uHb4dPPW+VQ8qsD8c5G8/jTQL/yli3+hJtyXdAGSGNxyHXVC2mbifxjH
DFQeyLD3qiTqjhThIohl04KnIPACfg4FI9xAAkY8GqUGsiDD8jRvTC3kPBTHjBe0WVx85U/QUSTm
AALR+ekMwtkRhz9RFQ9Kts9SdAaw79jvbMTFQowWg8NEF5f3cyQrV+ADOyBw5C4cSI26YvUq20jz
BsxjkptZA6hTnhF9VUMmJxYXm9NYsSrGdgGLWaqjCDIQqA12ovwAkZQnXruuFLrBusHXW0rekoo0
HpFIC+JqOlscfqc2KUqe1D0ZcRSaLcNBeSkoL/iqwZM5po2We4trVcP7ln8cp0+XyHysYDIua/Cr
Egw43eGN/aUoWP2/5l9DJu9dsFvI5Rb8ZJLyKbNol6HjWGNXJ1LC0xjGWv0IfR4G3AU97xDaeoaz
lgLX/86es+ritWvkt23I2xtThD3GeyTFHtdLe0a28gnU4IJOGtuQq96GQym7A56So0I6hgHJVZsI
D+Yz9nTHtcbPiwh5uec1+GXfVg/lYiVVaC/GAo13G143j6Ik+frCRvOoRTk9mzip1UrRvrgs4Ixj
htgARTS36gVXagG+1mRMhUiGEfcGRp422ZgVCNL7l/rziJ99mz0h2n1QaNHRZbvpZ8eYbGHQ3Hao
XlbWa+fI5NVK8M2OlnxuNFjNvO2bsMoDv1nAJ07uiZ1jkqNAOE6kY0KwFIHNxDA5kiKjzCkInPcd
aLE88MAVPOZdbv3tFInY6xu/5V9qz8tF8JJrks5u1TW892MMBnw5MSQrL0nmUkdBx1i3XLKhA2V+
PrLHICI3A8OFSOssVh8IjNcDIS2W1ryu4/grxozLIZamADon8vYesggY3Q/DpzMY9vFniVzPLjii
mv9MfiBESN3igiNMHRPiEADlERg+afg++fcANIZ2HVTFwYotbhuhVqr8RYK+aIXDUEchvAdiEXLR
R0nzb3FKAII1oz6T05uRsFEyo9td3CfkiYHVkVj1SLiZ/N31cdo5KaBd5Xd7BDOjFmj8WHjNfSTJ
xhDc9mJY1bTcB+ke8T/Emt9TcUdktDgerbNjlVGIhQTsXM6o6A7u0NdyeJ7hAtc6NGrE8slrPHzh
KUDcpvic5E+yH142aXgsZDj5PVwqMixsPm1FapnabXZGHx1SDLUpOn7Q82MSt5CIPpsAey+CCtXt
HytR6ecym+urnxEVkYWsLq95mm5plxTNXsvA5FykKjKHTSsPx8FTAU6suH4yWR6xy6keF3ax4iLw
R6EsNiveKJNArADUEqpPgiJ3boKysKoG+Ldiu/0aAFYiCn9tAl4H3Bbp5tInQHZJulqm3ZpKkcfx
B2Kh/kv+ZMGCQAtemvWiNDpGboIBsOBN0oGOW44VD+T8ksEUszR2BBAjhtXmEftSC7OjMygt8hbS
5lAv9yIyKFg9gwwLvUxIcKSogE13XmpEcuyM2gAVCIQr3Jqlydy41bDDKizuFSHsE3xIgtZf4pC+
/AD4wWYtvw75MuROU0UYeHjyEJ9OiIhYx4XtVlahzgICq1Ot7nnxOnGpmLYHIqdgjHxxJDhKXKoF
KsplhhNsa20ZgthncKXzQ/HTKnRdfUnQWR1IfVxpncxYEX4qyM8lSkfYUcNA4dE595sDblDrU8rR
UmP06HeBe0ctfTiwAk/8137KEK2VWeg8LzFSADda7bcF/HjcSwZU6/5Mlf3UmzdsEnLVKeXCemiA
EsZm2PCGI6lWxfZbFpaylpr4Ofbkg2m1us5lJe++F5yP96Ta4EsfxTjJ6saqSYOuMfxeMWEpD8JU
4Hp5t4Rzed0fDnAOgI7feF9G1RPg//N0vmGuQg+0uJOCz0VSjS/BFv9W6HyaIHL/mNNHsK715rUu
l93z46EC6LQeK1eptgEweh8LVua7ibxq6hTQtRjUBYQdRIOsCJhUnj/9EhX+DGDkzVnL7bFiYF45
DJpNWK5CD4ehEwHcAlal2Exoc/nnWSmMwZl8cdeiQ9lBGhNhY1OFMnCgSPDcV2QKynfuMNhCBnNK
U6yYHwnwlFhYFigbZBD6Y/uf54151WdxnwdT2aXcG33Yf8x5pkP7CMFZPoF+9kkoCPSb3DDz0nO7
8OVEwhdFzWmgaJiacPeYxBb/xtaR1PVnOjVJFzUWuYFlKXYI8lMZ+VCFW5PEXKVpKRNVBSR2u6uZ
WlGpIpbz5hNcDcOVbglACQJ9PTQwxSjMjBgaU5HnIP23pqJctqRDJpjxUie166bF4y85g4ABPQSY
Pq2UyMJ41pI5wO0vQjHbIOveEhpBS3IaUKqY0YdXzPtUM4dSJQpc5wB5+64zfr6vblu0TZ0kLkqp
P+piRKalC9QSplyoDyPU4dXCLGvgM2Iay7noDwlDF6fCLGt013klxxx6fKW4pO/h2TeEdRoHyW4B
MZ9u4qz+eiBoFp24IOH4MlM18p4VC61hGFNLYLdrXkXI0bnuJRuB09A5CqngxPGUF4dAx/ZpZ9et
3J33Tl3udSWFY/2KXgp5t5ORaShgjDpDZag0tRWWGyonqfSvsyYkUw3pWuPcrY1lDl44biq9v6+B
g/QKspH+l1nKyNmFNMYo+PIdqM0IURm1fAVJ68KOK8IyQ6cP7mE39II+4l60hmbfAV4OV9Y6EQW8
GEA+diEB/8zKVrUZReKy0u2j1O3y16aR5dYOmJU9mj0ob0D7MFjs6+3bzmIPSLUHEjBw8npnVDiE
a9mieRALQikPTpogmPyS1aRNs0Yz9W1f9lfTFIeFqlke/iPMxH6jpv9Cj/1X6izsO3cjPq0tioXR
O9ti31LDxD59kS7mu63ZnO1brcmnbi/Dxb8bP4U4ruR8L0Vwby/ZychqrTHDCpxC9WyxcbSCuuUc
xKWC7rHxhpxnJYLRUeZnsvdz4SSiIBRwlEQ5URlpow8sgK5Y3ZOESSZAlhS5lC1EWKjiLb1lOTIT
vEdHH0BPjYWjhV1xYRCDkdVyKLbEC5tWaOvJAX1tIvVJzXRw1xOrfnUPzvVow96v6f0ypUQmHCoE
Xg22jx0hs6OSSz7ydSlp/Pd6BrseSMJ2uBhf3Ljoq5kbbY2tT+GBWM0QvUt6K4tluTfVRa4qL5Di
8S1RoyqTidNW8BoKAmuWVfExLK53NcLM4vr4vuE0bDP1Vz0ykg3ZumFbBuLuLUlP4yYjWoz9v/XG
OSIxnr+qcmQfmVQ8M7ItlAhAnfBmL2AiG7atka7gKr7OhBAifY34tY2AXLpqgDNpQHf1KB8yt+kE
2+Nc3Z5J4oPyIf6RF6sOnR1ZZeMHCfF7SMLxWCFAWWbBSf8lCutAbVTyAmQWbmaG2M8JHUVJO4/f
6IbCXf+DvcN/Pl+N27GoEJFIgxJmDJv7M22q1GLsjVJvErr4YAuDFAiQQshdeko1lRVjUu9GkeEZ
Os5sSll83L3etjekRbRnFJenl+rmbBCQSO6ACBMi6rAvp7AH+0xx9cJQRMsNkSfE/pe8g2NZvTyq
NVJsuTQEnFHxKnrSf7SeQFA9DAN6uhCk9gmALpk9AzyvGCC/9fncubfGQRPrpxSXKlBtCSkuxq8F
p7xYdWOAtHxvNDaxGcPxcBIwTG5fYWyhPM25Hafz0YzBzyLNdD7/dicpA8Vc8SbgExZDziFsxjg0
xaOeg57eeYZbSkoVNERQ3amwAakafKWHVLA9lGlJFTBWUqjSb86+bDofxhgoY/T65S80OEdFQYfc
hxrKrnuNykP6/kUg6g1rn8PQQ5tZ0E0Q/OCrEM5d9q/0EAn48NyYBtwwRnUSbXQfIXY6mSzb/b5t
vAOa34J+m0iHIg5LcijCXTZbs1NvbocHQiz2i96B8vK5u373/ijaIBLJQI2yg2sb3WLa6oz+3X4X
exHWUNnA31ycRapqY7dQE7GRZbJtE0NyWlbEu9cUcq4ytPtBzI8SjyelPbLMeVwXBRYJXZjsWEpk
bypEU2xlGahRI3ObawYq07Ss8bjBx9IiBrS9LaBWLwmKWrRU6NokWG/IXVia9fe56E718EOlDIVx
7GuHq5UIPWFLE4YtZvaGNmhu9ELwLov+DdJVrwAb72BK6jPDjKRXao67+tic5b40w45bgvwyvozY
PDrqVInlkGKADI522febJy3ZJcw7FgSGlC7T9FmNV1hSHAmf88zQLaLnEUZcpry0s92jpA6L5MQN
9ayJk+WOgepivzu6c2sEwseumQacdzEW+LnPPBRh3Edk5ftUZoSQJz7E3yUIBIgLJnzJPEogYdkQ
uwKv1waA+3ClVSL6RYI4nITTiHwRqrHzphekfpqJcww5J2qa0IYygl8LVQUWA+WBi7zZL5Ew1uiT
Z71A6XloOPfIpX0IbSE5ScRLH7eGPyZOKI99T1gsKuSz2ll80fo8NKKLZbgX6q20+Vp4YXxSIMuA
5s3k0xaGl7b1D7o8+7lBvRW6yljwn5QJtqjAWK3m6qSx/mqT/HqLOnR/wJXSpSojA5sxtJ/Fq8R/
4h2mBA+F8+hYS6tCrPTeYAeJa6MZAbYPt9ZiIOvijY1neZQh26mSP0UWuyjdO+dLuq5Y2Coh0uIu
/5vsQlpYf+ExAJTEntQkKjd4HyYbKeNbAZW9gFTTaqMWP3HHULblKhPBnQmBoocJAbonqqGDtq+z
IMnousoNbsAnp++OLA8ihNF2NCQKLk7WmPqzRn4t4jucrxLSpgwJOghX0XBHKNJ/sPzrfa7oQYzU
GihqqtFvq4rwbIfeYptSstQ9rK7N/zJ9ulKQNhIc3+4ZcK6SxNQv/rIrtobkPY5YvKueeI9y1UrZ
7KGPCQiNpuGDLxdcpUKiTMc1w4BVLS/HaIptj7aJhhjUMXip/7G58yeR8M82etvrX9MfJNh8bL9S
04kZ3RPo9ia64vJSX+7YxDimuoECR5s8p/fAtGRcfVlHvELvdReffaH09Q/unZY8jxoJIwpFi7Pz
5rhuyM2wFUa/gy7Ub0mvFP2Xi/oiDsGPiO3Ui+GqQi7DqmVsZxMJqLFvrtgsfWJgOE4ATIxycDUR
ChyCoP1z9RoWjndHk3z5RiSJ6PDp0O86Pjoua3AfnlktkMJ+IgXaUr0IZZpqW3V5VVX2jaPGOVNk
MoFmLX5bxl7NRphr9h+dP0ZEAGRY4VcmcSLK2ZMtlFbdLJBeZh44JHzumlMPSxxK4zv6g6+K3qfa
UOqKO4a7Jg6UKAd2t+fP3gy0qARbh/HlD96piMEmvrszft4Zez851NQgx1DrjOhdb0HlbaORhWfL
46r/12y0Z8S5nj4HhRsSvX+GGyh0RcbvhUPT89VQj/vjZ9J8tguxNVRYpwKrYaucAQqKdE/4xtM5
wxSYm0m1EA1e9OSjdI+H6+IqYiKcc0A6xXy3ugRUWINgP66a8gIzaaNJc4ya2ucLHaMNASXCoP+y
DEYHOlo3rNz2gK6Uy7x9DBdziYjIx9hH7NynYxwYpg/VMo8Ab70dQhp3TtBZTxD5q5YcAi/NeEm3
cEDKHoQzgpbRn4q/ocLTpodHXDSZml5MEXXLN0Ob2JhrsHNEdXtkgH1YlCU18SSaZCLfg0lXckxb
mETI+Wcw6vVspUAG8SaqVRZNMhuoval86pBUyCTqIPufuOUDZ12mfSwYIAc2NscsCIpjFq4Xt4cZ
PfTVJmovh2QhlCOGxV3PQTiE4GTqU8rS4RxJeGzlpVw3UEg0ddev7cfyEQe/OfTLD4dVHOrhga7F
dbrgabspsaJdp0CCpGL5Sz6S4ByTFcd5aadF4Tkuj/dtxPOjM9JrOavhWfEuUHmYk2ELVAOzjXF2
mkhC+PsZ6IGo8e6KEJ0ngs6oCEc4I7Yu1CHo1HeYGxMGQuzbXCLNv5LJev5Ax/F7lJKLdLNvC1fF
qgMVlXMfqsuSLKP0lmnqQww6Hmrl9OuXhk1gageFQRDJP2VEAsVPQ8GpG0wmDTuiOX4LrtwUuYnM
9BGC8ZRFRlCJPpFsbErqO8RLvC/R4WYwX8/ArmfDL3XFBRi6btQ0Eg0m5ZLqhFlC5SzRiKCFPws9
uufkoNw4kdzMOFEBaUXecwP9n8AhUZrV6SzUpti4O11brI4GlYg00JLTjG8lv2P7IdLqgokEYDa+
bTeBICtxOweL1zX1hn7ryThFzA1wVi32FeagE4K7uvuVSFEG5GJ3oHMOof3iObr7HFtJdA8WDnO9
CRr4ZtiDbhDCdElQgUVwOWGgu+ttIEorIei50unqZOqiwbEBgcFdzzVElrgO5Pbqy1t+/nUoCKAa
u0TzaaEnigUDTgHPnEBf9NlHGWv4TzkwzQEwVrpPHF4V5SasfACYBpeCQ9Gw0aH3DXJTMzmOxQtx
wQInwQvmEVTzw7UJXDun8sV9j0aZQedaxwcOzrOWR3LYmVv1YAZ274wEOC0fxNAmLL9DWoCmLQ+E
jQk2hTcpeR9El2yH5FQaS3PqkBHa1z6NFf4AttEjcS5o2gaHS+IyAA2UHR2CfwvUztuPNTIwdI/G
vmLC6XOzAtfm5kf4tO60P5OzpBti1geuULQCNE1yK84mS1f/SDYDGB577Ev6eSrdsHKW6FWuPfll
EuZrHn6+eZenlf7738zik8edAs0btLmV1l0YMURSp5tpcAlWmtPzDijwGz9kjcQ3eYxSl+D3ZTFc
h4jceM2UJQ2vLc0yQKnyFM+69GyuU7la9YkrM0pS0qvFDlHpIdXwQPPV4HlRacwqVcqGH+5ZjZv/
ncJCTn69q5whY2nF8LjGIRqXR3gkkE0LpJdPLFJk/1iy3SgUt9HMmXOLS2nbFu7lVmrVo/LT68mO
ixMgeI91OyJ1Ym/yr/2HR9ifvZRUWfOgRhi9A/pcTRiB0NgA1ELKkgh06sqrqsllravpQoKU3mJS
eD95pELXsFwfCnbsgwasxvxrhrC5adBBblYPc3L80boNklhJXyN/r40LyX3/yKAfapMljhKJ4zWD
3OX2r00eTe41ybsiMJrUredg3OCTm01eEFQEDOT/yUR/wIcQWBRWcouxs68QPzS6bYMrhUEv2KuA
c0XihS+ZUVd/J7DsTKV+C48OV148HPoQLspKC2lPZ3e8rpepwRRsvSfxkC5DY12H9EwoxO2x+JsE
GRqunSt0XckBlhBfzc/5G5lZFUfLkq9ok43yfkjA8d3c2a7HOvSYN4O9N/tqbCqZ0WyZao2uFM/L
wHIxT+h3BdhtjqT/4/zLrnG8RuN/KV7wuy127osLQ1D4XQ+35Nl5YWeBFSiUAf9Pdwwv0yOBBJAA
vGyhLjMLyHTMEijqAndlgFvGiXd6SnfEAZYvCAdwug5VcJDtL1r3aoHMLjM3HqX271BF5TX5Qce+
PZs4M9XddtgXUiZ6e0UwNnh39tOuSzaBoYGMe58Wy5E8DxHH3SlCM0k9rfDkRvGDML8IwmFC1SnD
WY2GJPyFmIK3/0Wek6+yJUwsCIHGrrpQ3mS+2efV3JLJcr6n+9q2T5sreckN7CvdynOcHbLVO/+g
X5OXEqRotNTpfXcHLTEJapXKNaoNexXAdTCxj5EaLxI6HAPM5NWxhxjpglbhYTm7pfx62GQ6MHtm
69iyFMOwndK3m/G6QCgajR31bopxpUIWEJctp9NiZyRWO4ga0Rti2mV1cKMx5VjBBHgw8Pq/34dv
mIyxmIu9NSdwvLxJFDNfjMLW2w3O7D4Sv/k80NwmovyaWdQr5jW9o6i1MiCLGYu+ZQ84vt07//tG
AomZ/wdlFdfYCNlTc0RdlMjp1d6/f0JTgcEcczcZRkuWHotE4wiBbgGV68SsXcPXCLWAHC5m9x7F
PCEB28OjBFIWTA/QsdnK4+h7MAqzixlWycgwrUSy9bVFfCO9wEFKiX75ZO5/W0P8CUrsV+9/tfeJ
0534dfOljzsBrzpojZP02kgVhVwZNQHfGRr60Gks63L0ULNZctMmfxhGzpJlBYNbhQoNil2+aN75
iS2LUEqVezABv1W110PG6Fnggk686afh9fG/dfSmR1DAGcA+u62fi3kg1GaBwptQf/3SdBDFluza
EIbf6bqCFqnkOEHQcgRrx3ALmvLmOMnnO8qv5Ve2JgeiXyIU+G3ifR3iMLoRYxZUgYOvd3ccGvy3
i+ncsyioFr9kheYjB5GN1AkkI/JJ6r6hbAhOHuGp8VghpQuluGLHB3hzYolVNigTvizfyIdWKG2k
d+w7VkAePaeMxVXwpwDe2w8d3bddA50VQ/tRqH3RuicElhluNNb2vslyMj1PVKpSt7sl/XXVUXiE
mDciqKqedbNZRplqKfZUBJgpi986HmVT7M03ZLn3NZC7Hhy860hvsi97SrN/zTH9vVpyxEJrAosX
tCdtzoWGDkbgpd0ujv4Ka25iZTL23XSvhn5CBaHva9I3FGjYl2ZyKQjohMn1VbCVxK4Oz31fXb03
j22J+pFgRrT69vHiNdy3j7WBQ3obmP5MfIRrmigdmYnnAqO5ozqmGbby1r90Xja4leV1O7f6afMl
DvWo29ELd5sjWH76JExSf72daaOabkXTsSqucpPEfd1i8HnuTZHkYfyphBMORy7vp00rBe30sO9v
3qegicRPc3A2hEOBce6uxlt10/JaUKGEcN6fuXRuloqtis871ThwkxJq3tQp2x+/F7i7+/VZ5kid
T7UFx0W15wMHoE1AMYDNT1jJO8Z0ZSTjjz9TgcCZr/D06h78QApD2v8STys+dlqsBK9fCrIyVSEv
oZRAsZrT/aNSbNMRNXTtDBo35wYB5RAnTgde/Rl4DB/pYOHuhLHCtoH2nw5kTuTHZY3Hu2FBn4wk
pyWurMIwMwE64aGJTXzPKHP7a4NYeJAXsNL7fAR3HMZyrGlgrCB3aisfvLTZBGkaiPbgLY4emz3N
kkaMB20tH7gjWKwpKcp8c2vZpyUUZeVsM2yNUJH29np2iwGHMgXjil8MCrXkx3WnucXJhQKU/lXK
+TRGiFrn2kcRzdZ4b+E5Uo5c6QMuw+nx4V8jPOXdN4JCjO75FEdGuep2fHF8TIaoYagGZ6hCSN3w
7dTQfcbGOxhe6ZDbKQXs5tTiH9QQwSDH/aflG15cK/0nvSW5Vr9WBuYylqVfrfZDBmeJqbZ3ESUP
UwWkL19PRwaaYNe3D91Zd4Hj6N37P7jK6z6U78Gg1qVgd7IDhTX81hTGfNB+YVMZn+B0ebfEWyIv
NfecBYtZFwGEcGhimGEBPDcHnhs4bJa8B5Ue1JhGKGGypp/yZu4gLygv4xpP7EfCvHFGMFb1egwj
GNAS+1o/liK7FS8G8XJK0ROvnSbAcielaD51IC767I7SznJhi9AkMRDdFjcKyvDiK0gH6B1uNCQf
BhNJLqiZd2us9G+JsZqWdTshybGJeImQVYES4HVaLQ75RcpWuO8HCssYVUyiM+o2DBuUBqKb+d/W
ac4WQqmt5W5A+f7zSExekQ/rUHz44f73QRXuSiB7Zo/NxCJfWYtLUeTbTJnvMAvgdf76whrwLgA1
eMvLcv82bW0d91IbdjALRzF20YlvQDYaHbqoB+2mK/EPJl1iQynr/Xae5kWue/TDZcZpEiVQUxnC
xRUfMkd6NNAOEYqTo1jsKkhGodAWHoX/xjSHpnkMwjVrotU1UDiqFqw1z7RXgb4FBABXS6A2GKiV
kOYCSem9vCc9d9asuJxbMDdaiMpEjtRRMb90k74VgVRozr3CagS90xvx/xTnm+WzX6T/a7fWu3A1
oZG+AHK065e1GW/sC+n0k/sOq6rzGpW1tIlDP1Uoeq9ZRQF5IvI+zcg/JfRL6IldC0xJfRyb+ROW
DMPLZTZ8l86J1sRKexmAakvKJ16Gxxf6sZagi65CU/HH5pm1ezDK6mTgMOBQCdzeiKHNKdHjQS/f
b6aM/CbvtsULmg37c2GG542c/ZaaHeA2kTrHZNnbbQy04gE/cjYj0db7lT6aAtXEnXWOLCbOwlXS
/zM5LRuSKT6aNqkhM8qmScY1ztFs0Qez60L8dzzEEshSpG6AC1cc5rOXfGINxtBu2GlX1Oa/MdBf
RX3t2en2ufhziKnm0xYfjcu4s6ubUdFUN/OADRRBp9GNdGLE6vNCsQrAEB0XXmtb4jrpSIC4fuCA
ija7N8gF+/Av+kdzEia5ke9rz89yUuOE+F13wqf3YKsIIwUbgPu1o3OQ04jWbdOpG6i1rgqcjVeP
UDV8vq2Uf9ORLBRRJHZHXcCIhDQZSefxwvdzicMCDkAXhhYnuGZzdgAFCP8IJPNAIk4dpoVqU1Xx
JWxl2BT2OWwE6/2kiabssKUKCpXUPOeDkZtUcDW4hCVc0SepTWo8kYWmfXRPlQuSMc2nst73m1pH
CW3UaFGJIXWuqIRU004RYnxH/mpgO+iPFFkQhwiuNaRBua0EL3rsMhx6KvdpLOnPcZPKBCTtIzNu
L1Yffk4OQ02EAW3UPVVGD5iKjpWjx3I6n1VYTYVpaiQIidEsYKjb8YwvWjGdSJSEfBnWqk8esGSo
pBmgOa93kT0hXYMoYmTdFTU8nf69IV5OE9z+vY51YgQzgk7/08ziN+j9+3Jj73XsAj7BM47yMr9g
I5wOszAl5xcmV/W/rNV/DPdvsTdmvG9buKCcyaUelXE5fGJMr79X3OTV6jqDCy5BLbZy9e3UAHxc
e9TNZpKVTrjBGhuOxlaTSdYtLDjbbfpL0VN124LonSeAXZglUWRM8Z6jlqYkYob84m+lc+VVj7SV
BQoo31d0iIP3b07kMY7z7BodaRRfA+bHWXN7JfQ20EUg2qHvecgxQ+llBEtyOD4ewkwyEAeSkfJn
pLWk7RH/0wwAhHGCfzkOJQhN/6mnINrBI/S6wKtoU0lNRQpeR/3h10wkUkrjwZdu3sdYEu+CP8Xo
PRFpAU4ORof1b7xGFIDKlxXloR9KcDph3QNeS5S57k43bEthRkRa/QIqlCK45Ojibjo/N06qezds
W/oY5q4bPKgLssPBfJ363axBidchB3HTKxdlFEeWgDDMa/Qyt3vj5zERTaFV1LKtS1I46vZMrISW
0BNhSiXIofT9NsIrGaBrKcni1jIWDbQYBw4qHNscsEwALUj/CJ/z5IcurPUBK6MKpEyQzgQWGu0o
7c/+jnl0n4H8+kKK5bdEI5QUO3/v0tRmd1enEoGJETEuB/gXQ2a3SKHjOTo/hJGariqWgnBqa7ES
bcXkTP7RCRzqWANk7LRw0NoEyvrIkxcDmi87Z+mDcYk1S/7C77K4cSoUsYcLB1TWts49nGp6Qrjd
w3cpdO00t9kRWnMHi0e8DIhjoCn/YlTNhTnAlTmbguZEmg2fSIVgk7ScKO3oURW3QfaQd4OxZ/Kd
nVyWGOUmkx/DMD2Q+1Lqv0IhYShrme+LCEyCbe4CIy50JlTDmKXCRXYwk6euiA0rp/HhL/M4RcpU
rz2LEUC3Yg4EsygI2Ftq0TWuAWcYPs66GK8K5bOWqN/X/cHkuF65PWNPqRvCgPjI0EK+HpnpDLxj
L4AlStugCleYC59WASlELioQdAXjH71/wiw7clCsK1DKkde/LtqgRHeB2PKg4u0J19zw6Nq3EcDn
wVZ9yk4Nj6xLmmEqOdUAoUGPJ3OSq5K9dvcRJYQUuAIl6GnYStSSL875+R2EGHPRznjjX1hlurrD
uO1cIv5zEUBG//mSs9rnL+QhL8rDuMYErC40cA9qJTJ8LWPWF7Mb9fDytFoGXey3SCIioVwvNPFg
gXv7JbQThCMH+GJIinjUcsN71rBMbhVNAs0z7bcZqAPZZHHxD2h6ymIcmgPUonII5t1EFB/6XalM
jo6qyibyTg5LCYviMWOeLCIyow6fEBU/akMdkCcKnT2PP06EDHT0w+Hsz5M3jE7XRYGsWGLDP6A2
XBQdCubpmmQHIuQS0TcGfrCgOS0c/y+IjtrRRuOprK58hMouSZOSyKNXztYFwnnGDLz3zCEm20mR
0osmm9JSXQzmaOViulyYSRzziHY6qrNzPnggadYZFLVHCrdnFIBYmyxDvdTtSCARc+K0x00xzeS0
lh46BcDdlr+4+0phZUwAkO73Esh77DZ1YQJQSxdKgzz1qV1vyOzsGQoqVMGLOeVi/0RvYckUhseF
2wNURFgSJjhNtWCMT5tMwhL4+/7GLVbRNDj5dzIBjnzLHvZsDhXEdmLfOIOpcdnlsT0W/PBFI9D/
4QPZ8cGYRnypwfl4euevN/vnygBSyD0oKpbNYsO4wn/2O4ZoIV/eB+6DOXh2Gaj3J10faSsPr30y
1R8sDsk1sVMx1kxVswMHtS+9zvEhEg55G3aTGbEaR3ZmFhBl9PlqrS0v8WvCeSu0wINr1BlujByB
yeROHstdaoujRz4pDwS9Em88ZJRgRwdJQZ3p+2kIOsR9WuBuFqNbBhpbQrSCMiJQJwCD2TEQ7MtG
7XugeHonjJmFv38nUdUtzUzEzZWeCCWunwD9KeepQRB9udtQmSn0lqyzfE3to241zKh1Bo6Au3bQ
ZMfEggcg4Lrih75AGWvpC/Ryp/DCYrpS/VX7uCSoYknk/tcSO1DFjYwfyHis0nKlQbVs7AxGkuZx
JEqOutabrFFvx/Aq/04iumUDEX9vdTDzCjxQAVEi1lFq255CRvvn3t0Z25birOtwj2BQtG8crj1k
eTHk2Lcxo206lBa85MrjZ1tmxQ4hUI0tsBRzK7UR1qNIxZhv9cmo7VtVqqz1CBpyqNa+VhceLlqA
Mfd+PT6OJ5cxlJfghFJyqllTGd9au+qgfRZUPi4NiqfAzox402GzD6JjFT83QJpsCAyvq1FDTWa2
Ru/6n/PD7O8ZGKHlomtQ4UqedekZe5OTh/VUXq/qa77NgqdgxJwxFIqfL3qQqOvc82/pS4ya+gna
KcIthhilxf15XzQAsVkzrwGUNDF5uQUf3JQZAphPR+z/K7c7qWuEYwrfctq7SVxWM2B24b9Zx8JL
B/iPtghHoeCR2OHyw38d9GsRG10EOoV/cqVYI/zhovCfOwz6LlrJTVYnNqrd+7Wpf4lWyUIDh6pI
559GGLoE4NPeV5ED7XcGB4gTscDjR+9wCTz1hQ1cT3Z63R5vAAROCAbBceAWB4Ub3qNvcwfjTJuA
pjahbHRx+/Gvc5NpXoBlJ2LxDOhkhN2mIQmpZbS0IPmWWXcf3kTBc1qYSPmUmhEdQ/pBIYBx4a5B
mcPbKhx4/APSEjZjbZDIKVkX0Y89hvHKlXn+mXmMIPOR1ZpFROvlOF/1NoauSmO5jSlA4axMFSu6
2QO2v+wqMTR77CnuFPLgOqLvItO5BqQdfv4lFl3mf6PzZ3THIcnpYeK7WqMP7IP7pS58ftejO19b
IeosAqB5es98PTQCUN2lkiWGa7GpThplEPDavVh9m4iG22IXkHuhPFOmYQ2WCLUlAUOn1mPlQ6BW
lmNwrZcfbyAS29CZZgA9Ps+30bnPzySiupDoPcryzfoh1cZbjhs76e/JBfrVC3f+HsC3mO/Kf2U+
uV/4T2MmufcwsT6UPttPxhyYV9AXFj5Jnu5VwIsz3oNHT0NGMWeJUijyxoIwWYoZF4qs3tzIpWTv
RlcFjGHnBiyo9rSowlb4LdrMBto9Bk3lJTYBb3J2pkEYpswOpMeSuBaoDw988jjPW1MuNohE4y3T
vRx4uA5XN4s3eWKZLsDkgoolpFWSbST9zG/vwJhuENHVy/YZZxnB64er0POm7HvCQmL4wyp+KUIN
aOklEGs0AQ8U8/SkRCq2iNs0G7sH/RFb3i4yea9sfcJtnymKvl3o2bBfcwuUNuk505jgzjDD8yWa
28xfirwl5wfDBsxiZDEmFKmUu/8kmCoAEcNbJWO5fAsreBbG3XFY9vgeo5DqgnjMrDIQJbhbpCIh
DfPK0HfUUnf/lp42rVpRvJnLezI5JaewAL1pMlD4qWljtyuhf8tJQ2S4QWRDCq6EjxCTmS60aeXz
San2OE7KcK0/FeEUvf8AALn1cmbFwbQdaI5Kw5HZiOENNTHeL4FmImD7rR3JjZBUm8NP75JzSS7x
3ZQT4b4bJBjywEZniichwKxa0VfeYC4YE3zB6kvnOKpW9i+3ce+oTiG9fk8lchDe6I0TWUjyzZas
uavk8Wimxu5HHui2AIdgXNPhEOgu7H2XM2FISxZYuRFPiZ7jJcW0G32XTQaZxqh1lIoEQZJdwY7V
wzIvzZK+azPudAyiVtc/vyGSAdlBBUF/929UvC3AJLJ7JuMy1QpcSYRJsXQ9+5RzKKCE4N/l/bqb
SqU68gr9aGMf8vnqRXYb3kjF7c4Rk7Pv62lhRsuIDqpZpeeudJ0nXAH5symatyVzymxJ5sXv/4At
yhSGkOpBU2mISrjLg94Znf9RoPotu+4xLqZfmqk7fA4Kw8PG2kRLbOiZOshTJOCE726R3vJvH7zE
YmvBCicmnb/82gK4N42T1HY9IcUOttuUCGQ9/MJlEpeY3zKYUe8gTieWQpnQbVs32tuUKpVuccyo
5KzOfa88hEI8D8q7MLAgcLiyiUkQkP1EnTEF397FkFmsBDcmF24eRyro4EqqWrrPv6XfLQLhKMJ9
Jv4hkwj5PcoGauyykWjgFM9xA+Hu9Tlp0mv9HgvhAy6+fdCwmccX3ztsZEyEEa4q2qDFPYX6Md1j
2pzHVz0hIOaBk1PMpqtOEecfQ3ufNtTf8a225L6Se1qqtiYxNAIn0K5AI/NM2HyXkSCoZTDwDtJB
QxSY68nytfW13ThDHmn18akTSAhnNJdgpNzL2/N7Nx1vNl6lIn7vcBZQzJdr6jffXUVNFQ3n7awi
j8Pgd/oLfpIitym3rxTC+0gpQhoS36jHYxsJMg7ug2QuJY+M9kRLywyF6kpjniS50r9/5aQmNobF
q5/C9wv0n7Gk+AsLnK/HbJMZO7MF27FLwvnHkqcLyr4/V3jvtEuArcE41VXm1M5erJYxS5xoQ5rr
Rp4eW3aInWo6MJBtVIk7CFPT2UeknmQaKwtCvwsRuk+fiEB31KVEEq6VmaR8clVhJIospqDHGtD4
nfj8LhbGb02G5NAydWv+qvm0lr0Bv7A8eD9r1LUFycGAUv8aE/2l4h9HcMPVRCRwY+MXcx6Hl/jl
/grilGNND+7xW+hHZ9VSl+VW+HKGHABh9X5KdGpBf6e/xTWRIuC4aKhQ8E+2DEjbWz+ZlDXIi8by
//rOO93Q8HJYVpsA0j3yHZY7wkKJuUn1vgRc0vsTNMtKeFu2bG5cHzpkYXc0ceIhcU6EFyp/Frb/
I3qavvieaF3Padl8BAwjopb0QxDCn93uL19vj0VJ7wh0nHMOydAj2RX72ah+9+coQvqjZJn3Yrp8
CPleAxrF3YbxwycsSWklzTlTP4pQfXiYG3gvJNSTf3Ip5soxdfNSNQSQgmrKmPmOef9zdGpSefuv
Xfoft1Sb/9vtH+/aVLYcTfUDOvtSoqDvqPxYJDxvB2Gi9vObq00ORnlTFXEtufUy4YJtHeq7jtPV
bZmBv2rJnOAQccEj5N0gvoFw8q0DtyanrDAo3xjyt0RvhgRn9df8rwMrj2P+1oXKH+Jy35435xMd
l4dKubV9Adu0cs3pPr8YSjemAdrlObkHZa6OgoE/b6W7ZqMFLY9gps6YgiMrhDNG41H9y0JCuFAg
KqYLdBYsLXsISJfWln87+GUVDpNZicVV9uxln/csSUcK7Xwr2yVQEzxyMp9eiXyU3Q8DG7OOR8vf
UICBNrgLplZjGL/UAmjcnp4uvvZoB0YILBwIAFMipHo1OGOgZBORLoiXejPjD2S4VgWmumQcNmcF
FZwJ+hopKkQrdhTRUl//PuuTyGk9nA+WU13dc2GHkiYHZ6mfMYCFSEIsaQAtAfS3PaARt7iSHiWx
HPzaKcZ+Fzna6i9s9Gs+GJ3654OTmh9usRBhJQMP6KZhyz0NfreVon+YcTk/sbz/5EbyoqQh77LE
9rAJgMXMwrXvYe3TtWfAQ6LUexSAsSiKExUy3BYv70cwiugyBbs4i18FeGSYye0uzYIujPAEf9Ey
+U701qB+FnVor3sTlTRIlKoupGxHb979qQjmvkQIvlFgGVF7XS2swSHok1POV38UpwpQExMiq7QM
rJfgzqUJY6cXrL09wOpQQXPmqQ9pgBYwGcPnK/Ufds2t8YBS3XQxbfNYqSeCJbJ2LT9tz3abFQzf
gC3lLnGPnXRlo/SYXNtbKwtWhGrEZMBsi3iq6zCw47JzMGLKK6cFZ0NjU9kt5D6rQrUrkqX9Jy05
m7TJ8RGD1Pk4IlGfmESqVBTmkRThcBzf3R1h/kUtC2N3QAbN/Df9vJmNPQMtIJS7XJDWODEbubrM
PDPZPuWUzDJcAPaYesoexwYaq4ZAj37b5tk/EelLyiURNswcPzwI/ipIqZOotVq9z4htVV4ex6+v
zG49DEg1Za0JNMKmnVMzh8GvIKpHp136zj41XvW7ZB2O2177JsYGA2eRAXZAexTsr0fHkYOPxSdB
dhzHNlYHS33MFg7ldKN84phkoYrwNS0DyQkyC+c6Z8qUFkdn4LDVPdWypfkkjEsHpnIOWg1c0Ct7
frIisP63/BUj5NfIwqkwoGx49Dw0SC1E9cBaT4kBqvVEy/BSPJRg1BtIQbHW2BeBdNd8u2JCcSqM
GxIRr20t6wCMbedEpgi7HHkJDIyshvw6YSHPz+dk1PzvmiCmdcQMJDX5qBbgPsIURIVDL38ftP6O
68Rk2ZXoAyL0A35ijOaeDovb0/f6oTXPadaTH2dgs8CyaEUGjwjzq/yDAaJBusqjvipMTlSO72WM
et+NOccfufIBcZ2/OyAUtKGujzVqD64m67K1IWBeLbSQmtcJriAaJ137wQeWOPFt0w8ogmHr/KVV
GNUsGXV7i1NPqGSq0VsY4UKemaV2S6i4YvHGAay503HXtZqcU/iGqZiG1hxz2RYyXr8TVmAupgXi
hnlGOzFL1jAYhnLjv69IoUrqzNkRBgcQN68kz8mdEkJ4UPhopsc8sDorzw+lTBssQO86WR85VyS+
JN78+mbHhZUsvDMWrwtVpe2tSs6Q8xbVoJwKWUjlqKsrxeKvg+CsWrUGNvZOreZobo2A7pm0M9ys
nd9z+11HCL6eWqQB5Iing/NdLrEL7QXC8gpnvXBqdenPorC0yrXc83JsFt1lCUUrF7VjtvbMqPcs
lp9YgNn93J/EetFx/MwzQKHeVaV3NqsHfVynT7sOYvNGbtzhlGuv87lgmzNeqHH8uPsB6amF1i9A
qVE55lasulg5O6HGA0raJGWPm3GsDljZtptBeCs2TwK2o0+PMU7+ai6t4Nqz0v5mUGK+rozO+n2u
QPV68RJ2qwQxxfJDEWOacExbha0JbcHgvInDf3T0ftP6fZuaxK06mokqQoW5RSHGElcJK6xhENFc
EUetvJUql15U01pdjCI4/QNNlBppgWfYD+5kNzXcPVHB1B2eOYvpneoX8T+fIA7FDl2rPnvkwuYc
p9GbhN5aWLrsQydTecVKLcmX8MOTAcipIaqrVmZGzWlsTkQiK1625EaJMy2ACpxllZJ1K706LT8b
SeqbblfPobBP8WmhhX9PwinmdAWYrmE+/AlDdLwbD7SevyXDr+Y7YspsO3ubDBrBYvF7KO6/plXk
+RZQqyhH9KrYeobYecZj/Wy/d6pPXmOWXr9VeBiTorQ0F3hUlFP+98t/ABj1d1gZqOC/AsYN/Hxj
DGT/T1xItNnc2OZX6fgmEwyID8FuXz/Mk06H96laHMp0kEGMQV3HE9Z5eycQY6FN6sCsGUAeN7Xm
31NWIvkHXDHD45LIxfjdOYu8hJi4Vq8kJbeOo/FHbGzB3MyYW+juAjbtybO+pEIhVHJQXurPU+wi
e8tyOWOvFiCh9lrHNexNTesi4cbqUUpV80O3knwBgpCURTg/lPLhDJ4H9rQuFmZJKFk5d1y0PtKp
rjpK8yv8PsMlg0KE79UZIOyDlFYBA4W2slgFM9MhdjJ5GIJZvXX6nSxQHnMqSO5N4maGcQxDGMLu
iR5TcEk23i746Ve7nzv5ANbhbSXULt7rLtf4+5nIDyRkZ+o44xJtO4gS5wCm9Q/xwJLvNdi7Dh7V
cir0VXvgAKdvxQ+D9OM54qW07LVmPic6c9498XH0naYTvQCcyO9USZ/l5LQuv/hj/Qr2EhFrfyAz
y1uk9JHVqWpAZ6KtGUDebYKQtATyULB6Tqiy+e3iJ+lDPoHQFjE1qHCWV5wCPa6hGG1yh7GxcREe
AYdihMIIrhAiklMSg/ZDwLnLvvwpOQC6q3eG5a+gQHf3kwRIPjVgdVKGe+UCSiRJQIT8OUplIBAK
d+tqvb/yn/pB/aR+xdF5APM4Yv9QXgdv6c/iFnZDnpqGXk6eww91yHlFOTUZJEmSUByAQTDl6GCz
z8JdGDMYNFH4Osgwq5aNHkn9HZuWZBRqVc+HKhZ0Y+OyRc6QqHKSubusgsiKCjNkLlW7gN3Qh6fP
I/UXalogmbZ74dmmnAswzg5Z56mZVQXKVFZDTIS9dbn5CrBb/6hfQigFgRD1knIHl56zsh6bnBas
B66Z1y4ogATlDLu49HJPuDjLh9bqrxsxZBIsV3AfvvqdL7IAEyahyxb+2iKCyYW0Zbd/1k0YB+5G
KnascxcLXkuRj6oWav+Ix4QPl6fcKfeYGjIBg68MsKwwuxTSCOlLsJotIMecOENyLvPXSU3Sq+qk
A37TNmfhaZZx0iDDgfKoU85ZBG4o3cF0ZkGV36wm5bOvEwwIweBLcmtbwnNcovgh6YCwDlvDCFni
Vp0N0AGiJMT0AHdIgLPPYhtOlCICBtDpwmYdsTKnQXFKlfsnNPLts+Fux8JGCkSrukbg97dgN73l
ulZy/Bm+L3plt3Kz/z5e4UzI3z2WAt5x56Dw3KLn2dm6E/8NMDW2eFMqfzrRQJOCiX7mVR2FSZQ3
Fbx224hdt1a7En8rRKjvsAWn9ZYBqRX3l8kyJr/D0gNBvHboYVFszLfWnXJyZHJPknq/N4h5KToY
sDSuAXH1ynVJuZZJZQlSlLUBhtqKWUlWXwRukzMOOppub7GyyBnOFdUZVbwbi4k9/e/xf0OmdNY+
sUMG6tIFQAIyovd3CdynK0tXxLcS8nQMJmN/ClQNan1Z7VMot3MRSscoTEhm+QB9tV8PGuwu4wMD
bpzEEpDX+tosD/IKkzXxNFeizaCDpKyBcDpPJ6Uf/+EkpI2UUYSpSjzl0t+QxQ6irKv5aKhCl99f
l4/li4N8VYisGz4gNT/kIvsA1VcgempzJVnPppUaK50Y6AB7mHhSC6zHHfzuIC1aMP6Ox3nx0CUf
VIGPPj6pwgE/tbDE12lICQ9h0dgDa5spD08z3sOD5NXSFpeWi51JdF7E8BVSxTWaiblOK2qrgJYD
e2znBCeZoR5qZbEKFUbU1HKuBoLTabs6HxRiA22ORlp3bjl3hRYd/l8xU38/eR/EalJTH4u4UtjO
LLZTRnO1rCnGLS1+NDZ1BoU8FIO3kp4TwASNdvsHxMJb2npneAZb62P33UoDQbuInmr3GBvmG2Dk
4VdyjkCBjvKYgUlm3E3KZk6aKNk8qV9tdDcnRjUAb2ZkyM7cQanYy+GngLnOgb77XW2umexBUTZm
WJ7mpqIWbxOQykJmJpTVNN+NPC6eXmUgMhkR+iXAmA3Jn/GqcuvY4/RBSaLJystReFbaGT76hqQw
ERkfYYL94MLLs7we+29jlInE1iAV5f71aKiSHDGh29vmijZTZ9Pd9rkorK1b9icG1shOKE7lkz+X
7Mp4Ug+2v5r5nx15JxXHZQ7+mcttIeEIhAmaK6mG7nKpPdcYZvh6ULH8+JBZXEVuO0rMEId605VQ
MIdOrYAf9qbQp3321NLSg1Z/xc+EGFnQnvWXQAgZPDyXFpqkNaCXmMWiuQZabdk3kTVJxr6MaDOG
9mTf1GIVqbpotXTmmJnsq5uL/qHmmEbZMKpKiwzuUMIYc2VwEv2DjrujYXCKE9pD5jHlqy85ElIm
IXvKbjHKaA/PxaPP9Mqel2YDwy919Qyb8MMHDkBRtCD/RbRs3TO4f0eFaj7U2JYDpKMOmDxkOfMu
IC99s5YX5nKZX2sRfCVF94Mf3WHCu/kCDAVlxL1dG8mpkqizNko3V6dstMZqd8BnToO/Qp1Gp62f
2xRKEjLQMA3ay3Y1Yn90rGM4nCo1OHXqurvaxwPCCDCunkiyr+HzKlbj+ujPaudlGhuJEI59w28z
nz2WyYGpCK0Mw5ymcaeeFF0JE8JIkG/QrsDa2jqyZkZ/rJIaYWN55hSzkc0By39ofKQ5r6UFgPnq
+1LtqJuGq6Jr9V4eI8Et44/NoPsSu5aTvHziiNMP7LZF9iUgEmQ7X2ttrQzAr5M8UW49SHvK9v4o
31rqFYtyHySLWbMKoG5WhTepVyUhr/6QNjkcFbfa3irb/9AT2Icq8tQeQojk3/OJSie2LCqxzahC
25qfkBg6UKZWMhshZMIvQqrKwm/W67C4RWZslFbTbNkjxubU2pe3khy+ltR+FtKnZ6Oje2nrSi4J
+5QekQvMHbWvzGgfkLyAlhb0d6QbFU9nJvy97TVVpS5NYnGYbVMltxqByK2w3MK4ifD7DoGSeGaL
/HqKfMj1p6PqV4j9R3NGDVd8q4cSCg43Wk3yreN6pRC7SgnjHuuUKd+PyUcYN3AI5AVdn+jrAl4U
TjwckWrAwvWzzoWclbh+sGzGARH7nldSmIRfoHIvwPXPPJwrHELJ+pKsm00ANQvyQZbwIFczt3tf
8lGU3y7250gunBrQor1gD7SsGco0gUqxcnUvRgTRocuuygiXd0MvciG1hBCysCMtokM3DJebG305
kToSvKkoP9TX6zB54W7OMHAjQamFoS/Gs7RGTL70dYDkyv96ipaxetSdhuUCJMLRZdY4WrzsbDS4
B0yPjgp84GQOPFmI+drhGAD4qGyTq94TqD2R9JeSTrJQPtBL9kz1tEleWQhHe5drkbFvyZ4U9l+3
W/8+igakR/drWNkYntCftoaX5uY6l2e/mqk6ziywAndbgFxV7Ra18ZDcNiumkRmvbaOW/dOicR3K
5uXPX7qXQ+2VM8mb0mZbQawseQEFlAvzUD5EE689tTCFMLGCI+dbQ7iDBbShLhr8PUEUlncqb2HM
WPy+y25czrmGlrKel08sHnbvD3YyMWrKgywtSL01lGMrfF4eRmQ0MOoJ0r28xaH+bgaO5TMsA6J8
adN3E75U8KR0iyZIUOTH1tIORM5xtTkZxfm6y07Dw+t/7aYBgoGx/Twt8Y8Fnk2oIT0n5CHYLiQM
I30e5eyBFGHfDBLej2PP4/evp2HzwFyXlIWOpBgal0tQdAAWeQXsjayc+6I26M8yy32evYA7Dy70
kwlSVAg033dJD51wOH3COE8pzQL3uqkqaKJayfyHsDwVLTrI+09H+cHa5qdeUavId119VBQ0bcYK
eQPez6lBbqZq+Y7/agQeMS7MltyDBx2ultQVjLQdXe0djOK1h91QHTad6exhnsnW0p4UO//YKE2y
XZw+P495EUXS4me6g96Y47VVGb0MXUhky+xVYPQKXInt31nezW8HLT3B/CwgmvH4SwGedUm/dGYF
sBSnYuQcPLkfumgsCmk847FYImZCJYz9Kylio90nDQiBrxifg1Y/Ze2d1Nfsr5Hhs+oP4sLWTEZM
y6V+ReTMzRhiOPbXAqX1XIUXvOK3LNg75Z5qsQZgd8scRyMw/sZ+yE96iN3iVCM6IcLEWQkP3oGa
e4GNba0oUZc0fiXO97anrVPD5vsCh4HBbw65RxDvgnd9KJs8NUAlzjHtOBZWzIw6SywSYF+bqTVg
Cps08i3dD5eIOnAPxhNR7Y93l8o9GVgZ+iU+aSC4F1Y3HvMlCO9Rz8Axx1bUusEajxu50OSHjjRV
sE3rC3yQpdmQT5HzLf5wtfUynblCh2zYtqkWUGNV1HXDwBEcjTfc8H8ZjsmMywT3zdVt5r+H/02g
blxB6sRIgekgNy9jrE/nT5V+/sW6/ULOWIRKH+yra8NEZ+STHKz6YjAXAHvtN2Exz4218o0p6Zbc
0ueP37JW0EMoyk1L6LYjlm0hGr49t2loZrScLufGcgWJzFRnB6u1gj8jSerCQvx/fkqVvn+0byxP
/Oa44pQ1aRqrU7XCQZoZDTiANv6WpnROWiow+Uo9MZcFevog3CBD6DO26372iZ/+2gkFPxh64J/b
GgUhvJTZb3XipDjL9+xAljc9ULwXGpGoFzv/aiOrGIKSl81foL+w/BDsHZkCh2G8jR5CSSWzGbt9
A6CuopSPd/CTw1df6UjlejDrVXk3rzqe2HkRWjFG6CFJ4mUCeyJeusaYNFl3cJNqkNI4y6GrLpdE
q8oxPBvLEffPqOuM2fjNoRpUK7/H1Ptx6DNkmcX0gsahxh0OewWArtiGEKMjuafk6DdlyavQdHnF
S8xG42SOGI4gF0JA6v37J+ceNKYfidb1A04sC/lJNMmD2GWSHT0UwMFAY/g8cgHK8lgrJp/83EgW
z9pKlHeriwDizrBv6CCEmCZNxU4pqNnjaT56zGj/IsYdW6whHqq7f7lz2wN4rd2aAiLVmIF09w/W
16z2dHGvO7k6gKntRduYynj5uMo0HDCXIGufLRh+6zRL0rkPpgHS+4vDx6CzxXW1t9g2RYdNsWfi
nNbpQSiJD3td7OxMfpTK6RhkZpTRIyFa3wJO/ozZIU4JQm8lwad6XVJmDjlNyoO3KPUlsLpwcUpp
34TXb7sWfI6R3NrikFhTO1GwtVVHSA4CXWJSHOxV0m7LamAE0ksQJziYWcJaHUwXddDxJHaSD6wS
RWsaCQPE7KiuHzzWUQDqAq525QtVo1DELPUpar9RFbrCbvm1JbVNbrX64GA0GL1r7c4wChZbULNz
Ube6WOMPAieIK9adDy0W8OTiAKFKYnYObaO7Q0OM3NBvBY+ByXBBtpRu0jVVPZn3HNs9nx5cgdya
mU/DdonmJhD+IOY6TTt8LXVtSZzkWwplpa7qxYHEkIgBP8n5CjVgvGI5tZBX+HhOHa3msM4tm6wD
FQ+vQ5ULPPLvy1aIIlX4pJG5SbGragPMAocE5HC6YSvfP0GKt69QKMsamvwCcANHMTZH1TcgQxcv
WApYzsC9SpEvHhHgGWI32galhlJnqJMzk5SjrQ+/KmNBs21AghAvRn/Y4OI8HJK9tjmWNiOT0fTN
g1WDnUbmJrvP1ktlHbTnfUk9V3AOF8FmPB+V4lyZQ+jYt51tVCR+BWrVGjRi47zB0DZg5GA8VgYe
jmaGcAwW7eFx/5uju6d7II4VRBXc8icdCZs4u0BNssxHUYiAxOR9eq61wNk1HA6S/VPY5bgYYgGX
7HSkm6CFBbGUcw+MsVuJ5LdqW59vTVfpYNoP+gSFZyvAMB4h+V2bLxVoHvgVg4zTAzg5PymeRTmZ
b01JnicTlwXjOa4Gzhk6WsPfArCZwglrSQAJSGpOHii692y38jH2fmtFRjcGS7UFHDANzkmcsCzn
7zuhv9wOCQqw6E/n8e7BLrzZ79W/plDNUgDpKlX+L7TJ1vRv7eg23G7iR3APAMLYFtlF2YXvEuiG
aMor2C3Ge03r+9qnWWNlTP1z2cfVXk0zujMpEIWbMye2LU2NB+bIg2SdJFhbkFWqcPIkTMXvqs39
EG1nrPeE29Xy/w9u7hzmwn4F+lTowHoRaQ3VCc+d70OXWDUE90Oce/R7Bj4x8veH+E4q1d4IRGFb
FPuCMq2DwVGqDNd7zLvxn4QiuZYkQrb9n1sxbWPhqyItVQLzI0wgcgVxZ3UMECCP0nVxeHZA6avS
v0Gy91goEFKa/hs65RW3BAfN/PCihgQogvMsLx2MMCSO9FwwHY3pmMw2sa1NAYKWmJQ5ITMcrYAq
Vf47DCz1gRpZn0YskpKV/elGlz1ZhTWRJBq8XbyTLlmfuSBEaIhhjaP6l+bifb3l+6BWVDRfhvLm
DS8D5SK/lG2tF7E1cwe8VyyX6i3hg2vSjHLyjmSDEriVHiWoGcZSBu54D7r2If4Yjdt1/MG33jep
g0ruDj94QFpJkh+90MTmFK7agorNc0d3M1JKc4Ej3zF6+7ulcmkNGrdPiWGk+xcRgrfli6toc8s+
2ZHvJ5+kA+4Bxf0yOd9o2kMHC7QeyuBlsedBsWCm+ECIq8ILhEnFUbrv/VahxC3OyQ2AnObfTZ6I
LarWNYCCGkjuSySFoJ9LBxbMODBWzKcYg6C+OvgG7glt5L4GAHT3HUQ04+GlduVyPNGE1fIM22V8
vECaB1ig3h5CLCuryNZprk6MeyCLbe5qAIFw66TNZyTxnrDykoOw9f25QeJZ+jLN2grOYwgsZtpj
mrKsB5XX8H1IQoOt0n4S0YbFa9Ng/WgtGZBtlfcPpMbAZlXu/0KJ6jnHeQHmBr1rPfelydUWUKJX
4QpL5SRlYq7neDLxqDfbNGKRXjPTcSq6pl6HOlgaZPKBRTVGgm/VwvLCMaqeGw2oMEgUhfihkX6r
PBLHZFxjwmTjvQmE4+sTc7VYteWclPRxjBCinaOeJkIqY7lgSKaeqBuHbksIeftquXCm8YvfBTfJ
oDlPuq4SwGH1m7iplt7BXxphN2KWCfyXVOIU3BFXsslH/Q0gOb+FaxxCVgPuz8smtJyI2PfVQVGr
pD4BWewIBjzoGH12i76OyH4uOGaSiTlb3UD0/Y2S7afMMtQGWOeVcBP00kIzoMtopEALhKv0bQ3W
o0kZ9TZEKAQp7qTUtmm2Qj5MXHyA6y4Gidf02uP/faY/y3jCmV4meOG1DdRaeekWgai6rbq/3sQ2
5T5ezbtbNYHe1g4d3phaiCmmw6s2yxxpEUf+OKqCUbLPhqXEdLEmIb6gLr0VYeONaMtEhCxY+LCb
vc2dY12nUPhyRBw8WxxrobxsApkB9Rh4NVkv/5C8E0feYRQ9DghK8568dOxfCxe7SoKvEhhoOkLo
qLZWmKoQSMuqKhuMuqMqTKce06FotoMZrVCdmo8CW3x/dEOTFNsYU8yTje5v0RacpEyNgc8ZKxql
7x+cd/kTlqxJLql4BkmKtnZbnyHKZabKb19ye6ZlwzViLV/UNac8648SqZi9K4gTog7WGqyJrb8I
OJZPgxhkkmSmd5CBJYhPk5tF4MYtoqGLriFW8EeU87tRxznlmWjJow7U84DrISxD8nCZoPJCvhLy
wvODoLmjVGkeg6IYh0HHayUvh0t7VSH0Xm501Jtd8GCwOC4vWv3Oq3LVLiVVXiNC7TIv9IDt9Jfy
vM+O3JhzxwrLgCaiGVVldN5bIzBA8qdUkzj7JAg5Urnqre1W1gNZnUMp8aeJ1Vt3f8kDNIxPryDS
RINw4SY6Xn+o/+M1dAFAobMLAniGGlDT45nbEUUSidOq8OoTb0ZEwJkeN9lxQXg2GrOWxkoVtCHq
xTyjx+b+87yEt9FRXd80srsoadSADGYyCY4EZ4deLuxTF5ihKROapUZfBveM+XUEpPj/P0SmGK41
XTvfTY0O+mS5YkOYPdDQQg/l3etbpy/CIR3hX+2KuPBIKdGxER73xrzTq+y4+w1pOnn7Xhl81zdM
nVa6tm2Pw3uRZyZsrj4u+E9N4qqat0P9AaNEEsx3+fk7DZj0quPV9B1NCyOSjj20nJkwWVb/zn6j
y6vPeB3Qz9dOEr2WNG675JnZBx3sLPK9VMu0E7lbaluaxin8ITZDZ4H4590gDA+SjMus/91nH/PN
q6nQgcKTA6bh6lB6a2SmqFCZI6ZvZLyT2BSRm21k1iyNtDo+ZI0HTpaKyxSBSwWVgcW3Ij94BMZo
uww8rmybjKMx55WF2UowzyJowZDIV973gdn4tRBre9OwegYgCiIrRc3lrDtKWJhjLoIZrZTXNhOb
JXRTCjSp0aRT1HXFVur3mILi0CrP42XddyQX0mE80/+N+nfCQahxBBD6cLybwHipsLFeId2ZCbSx
XVbLXfiRgQkv2uUvLbgtpmYm+HBYGuxljfpsiOZkdSK41Af2A/o3K6GXEDKmL31hnGZvGnr9UAok
SYJ/8At2XMWxvfuiVyhp/EKrxIfVV9uJPqFpBsyXMdZd0DZJAln6CQ1gCzWfCQFoCeWw8lUNqan5
vhSFl5u2i3b7eLbkDPBT6y5TNjvmMeMWhAiSBjJzueTARPHfD872LPcqIBS5sTEUGuxZY5mhGukm
PYQ4bOnjGUlFIg6+TmrSnoM+WHMRUdRp0oTt06Y8f5zuD8Qmigoy+9vJaN5BTp9Z7+Oda8dVsd1n
k6K6NBC7urpbIVbVAkpRG7fR+/CkhjdJ1KqnVGQUS7EmfVgipZwSGEivQuh+XJmVoBePtsVt4AvT
3j28pBnL3p6hZXkKEKLzegpwn6VKMJ+zldysqyLRQ62Km5DPBZG8GHy0qNGCa40WdS2k+DYpGx+o
uLo2bdJOT7Y3KkQWBMUfevICJlDPNqDMfnUefsn3+GkRlpHDimY81BFJJDouSEmVVbI7PlmawLb7
kUenqu3EzQIw+/06SpoKldBQxqnNp8LXNNMStCq8JLKy1RnSVS78OSYPOYPQwGJierD4bqQWHFKv
/6wIGfTGcTWjrPd8tYd8YMwQbDqyVNTTeHskYT0FvVIwiDv5NtDYFPA5dFwe6bHwdgQoz0hcnBA2
3AErKKSqEcdUI4foP5Ewlu89Djt0JjmZKKnHZg0vJNKxiVLHSrbtf4RUur+3H8TH3Ie1PP4IEgcp
eR8Hqt1aCxUWfqLOVrp4tlaOjIOH2ZonPtaXqZYG5TqelVWdw4AzkJIAlK2v7wgiBzv/vzN2JPRL
6eD0GCj8Xg0MdQCa6iDCTP6eho/87I5YlZXCFxxaZ0Kstplcfv1W4P/0xGEAjqN3oLu8IAu7MmKj
Nm8Jbg+2PAtZf/lVvlC3XRnjzDZ5znEsjnYNeU9xOPbMnwgokAmQF2/2Q/GQSXzNvuNyAIpQ3gHl
fs380q2zz3JsaZ2X99a7NFVP+rORfGbFI2TDzsZ6MYKfN0ti/s0mqB9sfye6sH//q4UjfOAtCAcY
DITl7+cqumYtioDxwL0rB1mFLuEJiyoNKxJlWiEdx/VYRZZsngSmH+xvkLsgxVnc1ZbzrIC4ogi0
n+zFWZuVfjm7s25nHy+7Mo0VxgZeOnItFGPIPkgEY5t+RIXkA+DMGkSPKuIn5i9poSFozPr8IEqq
/lwvb1Duivn83IntBSPE9K85ouSHuN+x2wgHSmC0ZZAi/wi8OVbuF/gOPMYA6gTDOCmBfycSVNur
JnpVi3o3M2kI9ntstlTK12n6fkXojPJeeB4hVWQ/doqe6+Fks/u5dOf1q7A7EntIRzCo06q39ZtZ
Ps5QQLzcrTMdniJ0gXZvM4UEVE5MeA2aSTkZt3P7lU/tzgBdZLY0bDT/ldGgo9ebrmkqW12blkwi
48jTDhDKgcM3mExog10/6ZYhxZaX//aNn4hof3Txsm/hIwpBPiymqeZ5r9yXzzOSt6qgmo3yc5vb
Gf0CV3aVHS15cr2n0arZEzvYPZJdbxlBTAVGw117Bvw1iMx3bBX6GxKE2l+xyHZ46w37Idng54We
sdF1RUmXUFkv6RkPYMJqwVwOoT3asNIZrhiiWJyAQc3VRF3NC8t+TQaFGLvv0egTN8W9/B5A3uBs
7JfLJLeuTHMsShiY53Y01xUhPbf0c5W/IOu80qddOlnTmpjMaK2ZeyEVRC7w0sUe/xcxgKVbQgqs
Q0E4RDfoKO0JYdZYcUbjkEe1zBtmMrvZA4Kt63kIWeK04e7X90j/moZiPrxVaBuWGF0YoP7enms1
PGhImVybMZ+CsfQe5x9jDZpWYc1h5yZts0TrZvSUN/Krg5NebxJJ/vntA0ySjAtqs9ufoYfBLudX
i0TT4Bw3dUIzqEWdyM6mt8jyZJ5FTB2HIZ6Pdj1wLz/W+vr9WEi9N4v5Rt/YusCyYNC9MFTe36zb
ncTDli+B3XH15S9cJqwd11LNKgPaXO5qtbWcr3X5iRQj/Y6cT04HkNG6ggFcpkXceE0g0+YTwxrP
IwU+J9S3h6QlS65ikgbY0URMOMG7W0qG7c8CJs4DQ9mDKOwNqkRnH9tvxNTwxaH5M2HwaGAWgEii
OeZ/R3ki7QP5JHPcIBebzxik46QcHpQNlykKLAm/J3D7edWAD+Tq/XO7ASD6lDtAPISBqxVpFlF4
ugLE3SFFPBeBugTf49ISDMgF+t3U6ZgSBPSMo+IyqpG+qy+fX54QoRvLFhZxTjCV2dh40OjmONMB
rEA3B7NuICjcbCvs9EbIqFr7tIZp7h7wJRT477bDzLtzi+YhXOycrYATUvChUp3nZAY2dHPqEfRd
PXW/kJPkHlImhkG6yReCfhskuQGHJTClKi4/QYgus5jxdgVYY5U3cLKSOnf4vQp0fXFju/p0rjU2
cYuhAYm6K4RLJOuWJ8h9R1kOYY2HR9VdA7Lu4Bfa2br/FZpygBba6DsRTqW1a27EzlAexlIxVCmU
ulHe1A7kQGbp1JkSRbSrIi9AiMoQiRxVl8HJfsXm8v6ATWqOhYxhpNhDluXEKbX3o7ET4XnfCB6B
nhf/6W3yBQ2PDifCIc23CgFfTSnng/+2LxVn6RCtmZLTsJRh/Wxqa6U8PdB8pLw5UWrjY1M1oPps
gmbBqDvcUi9UzzB8gosYPB+iFLEHrqyfsfmdN6g2/jAL/qK9OVD8WyeocKcJM59CcpNqNYzKeq3C
LbBAYNGm71JIOLRoTGi8tFrZd2PW7SmsThSCmwtcbuITYtHT3uegMHowmeJMkkYNKlPPgegSkIfG
CiQcTuRvFpp9tm3KSikNCtMb3nr+lJwBYnZ2Dp0rwx27G7WpnVDGknGqY+YwTKBu/4pnb3jRGjHo
bgKnreEYytfqphViSviNsTVjpSok7cx8M3nok/l835qtWEsDwRxacX6sP4TrOejMTDcppZswOrWi
Baa2iN5torL944qHUMtBUc8i81q/Gw1t5t4K4g+oIL0GbdS8YnFQ15qllK1o0nHG9a+FQbQWjnAc
fgJK1btGYJ5SXk80o4NkPIU5+iMzB6S2RwTUdPseKNYtMPWrWSkwHgdBQZVYS6bpc2xk7E5A9Zui
HEjSxx7UILlmz6EICfBhuzncoejWjDwS22ZdtC8rwgWdfNtOHT8QJVEgSSjVso/aQfhd+Jk1VdeV
Yc4Ippy2DOLX/ytgarXlidHQ1KyTCyTtwokB9edrqB/jUTqEcnGX4LG7TcPmF1TscxcLua3YOcyX
MHyh9lS3WCqgup3b+rHLPYq6DrM1agQEW9hHctcouZCTux3+ht/CSDHu0/cB7AXx8x89NFZcxHBh
xBWedpIVCE3qKGfewhUjNYZsQ1kyzQSCVsZw4A595KKwe8/7/h36T0Nx90hoCL3T7ohoCUlk7k66
AWCiaBdsDa5r2sHaypRMH8vNJt2w/po+0wChKpypB8qQNKwLwOJ1pMrtYeAEIX8XnR5walpT/yhq
aNdvK7mPF67HHe7faZOGbLs0XROJTdMKQ/Z61LyXFn5MsI64qBuFpDLSSf3fAjGwlMTnHn9btwBN
Xa/8K0/cx9BpyvXDG7M+PfUaGibnzVl9hgcTo/f4bWPx2olLA6UpVa8WVBJF0hNJrsk3PdakEJ6e
2iQqr20oq9zgn7lHEsxtqhmGr6cpf0MRX0Kuj1IouUn43eMp1F/iSMoJkozhJx7OhRGidKRId4XS
vGuEHCfGCq7/PnXeWhYloupjHJ93C/8N+dMKrr56d2iQj6zsBXhl3OtqFris+VsYmbPPhDv1vH7M
umc4OpYqDHb0ePmzfk2I8ij44qhwgGImkQymvIWjlgR902MwVX78Ouu1NjiaERz1kAA2j1T+pEpB
0xYSidsGiPGU2CJSgf/A/bFexWc5DTwXRAM4t85imI9bwZSyt1BreuD7OTu/z6BaYe6FiToiVWHU
j6Ea1RPp4FFcxSRYgDlrCV3vZOFPHuJW+wCDlw8J0N6WiJ+gGw+nWLDP5/j5cpY9iGX5JGqaGP7i
42NeJXIKzKccHepi1wRbQKdPqk8Jpdl5oneKP1Us6myWRnu2P0w83P+HzD/e2Rk9L6tfufUiuBD3
mMESPc4mAoXuRio57heszT+Vxxe6LN8futJSTnpr5X8ohLE3bwLyhWAwfUo/lxD8KuZ2roEIBypI
0nYSqcooZib0ave5VYw8GFIsat7uSI4bIPnZMqeEPDLwibfJJO+KSS5/NcLVIEwVTTw/JaQvQi4W
3XBfWe97Inowh/2QsvQQeJE0Lh0yO/u9G0pxtYlA8t/yLjyiZazPuJjsTnuwwA9HxRjtmUd0XfEP
oUywpIr3doM34QjalgRae8+Tgbt9Y05psiPf6uHFpD6wzfklbWgbauwDvHgUO4ulWwSD3FhKF3YB
Mn7jxB2c48dIk7qfbrTKLyFxckk/9pwDF9BCOiXWUs2bT5BUPcqfrxf5UJyMd5dm0ug7xxuRWEDp
LaPwK3+Kdybc9hHxnKl9eiopIdUnswe0UcPvDjmgNE80d2fkBIcw9uepa2VXsgsr+ZgRKoNm7G/P
VgFMUZRCCTj/a1MQMLH4uxCoMOa7k8NcU7XutVOjwQBdTaz0FlIV/fWQGHIpqJqwJ/wDQv7E2LjJ
TWZ11hMkn0EVuVUB1VnRCAWH/QmCq1XY4XuTmRy9htlq3jyyXMbQ1m0ZvVvoZTsNiwzRjq9n4Fb6
VCJcIXS4gVvtxoaDmzr7wIp1PA84nujZI1gfYtLo652HZs3AsRmj63+v3KRZIYqrgkrwPmlC3p1g
mFvk6yVU0YcGwcbi+Uc2NewTtiJSavDWiL4Ox1J4+06SMZkNUTCiTYmbTKI0L3OLB/tpUlEw1D2w
q8Dn9zrAcwyE7vrvqiaaxN7XxODB3iE5I2X4mzBtAL/cr0eWW4thUO5Ijfi9oW7r9JWghTrDhciJ
Ph76eVy+b5OqGlt8pI8ueQhBgzlugZPPO7B2h4TPyX+GHgaebqO4tyIkKSi+aC7/KwHeV8qjxkC5
tP3gnKA/DzwfCkV7TdJPaWwW3N207gAD0kLGAIpVbzpdQ0Xuchhntv4Jja7lnz9vE135JI6UzBeT
f18QpU3NeooPc0Zcy4F9oYOJKFYDazNZRDPZ8VfnMeVoVXstD6JwM+m3TZ4cH/w3NZCxhizDXNmF
cLz3Z9Db0I8KLtlvkTAOSd13oc0D5MgrSHkt3AqoIFxQodEf/OBbc6JCrD0Zs4hiN4EwLC2FHNuN
zqXauLfdy+cBAB/+l1rFEASWEnLn84izH7RlwJVP16a/O1rpq1yoxfQnIXuPVSuKT71oKEbGFGeO
ONJRghklxtmyf4Kv1XBjCNtvPKwdyLzKWEr9r8PBz7jubiC/A35W7gO8k7wnyYk+th9u4JOu3Sha
jBePqP6yYIFOS488j+cu+/jQxh5xBqkyAxxbW6MExcNvveUfPiPLGiAM/BO9IfKUbJ8Gc0ICsK86
ECtZ2XiJztnP31WcT8CKaGrNuJyoA6uriT3z6z+ot+GOglNc2c9HPuOgea4vQtaNB/rh+DCwSA30
0ByuylAgcaktmSVpzDPVNGwU0Ho6ta5XduEOVLFTKU1lDg0ciZqzeVqIDe90Ql1FgmpL9JuIXj9r
mhJSk8Rift+0WxoWEd96OAHsmH9x4MM4kVX0zVdqEXpMuYIrkEDFokiyspaKTm+a15m9u9Ra4mxn
E9HD49YU0mhXEcs2sCYWfV2JQVEcyzgJ3oxUDZRAQqq90LTixON6hDCwTSNg7n4e5GV8kwRllKII
3HUpoFr5qMyFrjt2p+0oTfT9T+PDkJ7Ori8gd5YzIgUfvVPtj8ojKlXfPjzRZ4iP0xsCA/eIyTzl
mCHCgGPDxvZKDrKonApsfHOZEMvJ5N846WQsmrk0F0fmfRaMprCmd27Xr9aZWK5dwm4YTgkYHTSX
YqqcLt3665J3V7O59b1U/qLkvtieSYkKdqWc2wveNDbyuj2+y+WGe/eFpv95yb4QIl8Tv9+k/CDC
qStUd+5HlMLQ8onEOGvEiJgEn+egVm3oTNQEzbgOQEpRnmbvhuVuUy4KMhAHqu5t6y3SbKe4Dy5M
YiT0MaAIngSHGuRv5LQxOcy2cPO2hbwFVkZgC3Zal88VMHVCHd5qrp9mHX9mxLmex3ijxpw2CFwq
h6VLcVScxOC35wGcG2kBT+Ta2wyW9yFnid52o/zkU6iGEariktH+6enf2vO5kiVjQ5AOzn6Vl6Nx
XTMIiz/KiET9hHOT6Comg7Pe4344cdqmHadkoTso83pjKFyq1Tenq2WJOTqCg3sp0t5WNWinHQt+
QBshzgYyspudCtbH0m9Ly7U93xco3Ax/qWqiU8nZO3OR4hauYzoSvBKjqVDIH96zY0ycIrqBwrKw
DO3+B1c4vh20k52n/iDGDzLiQRHKkiG5j0cuWU/YH6gluO7qhh30C+VoNd/T9WQT/hvU+3GYo7Qb
rQpQIpbAhlJHb924SK4gFcHuZiLGcTuU6fylqIv1w+iZkFVTMB85d/1m+q+heXrXsDL/z9cM+4nn
fFlW7R5eAMv7gtuY27pC3ewNzR4iRbHv6Q9SVXaalBCwPUCn3EjKVo3ZUPwLV+pwrOp5azvrleam
uq6srapoWWKqGMOTYitPvzk5E5TI4Z4S0KNmLvRx+/3TO/33+fBtfpUzfHxlUns/vhlJP84/DJMn
0+L2W3QvnE2EMdvzrXwgC1Dilm/RY9dtG/8Yqhohnz/CmB0KAPpMUnRRaSW0ubleBlv77VGXc+6V
sgRJchL9Per2y0S+EEolrFxlO4zX46dA7Np7VY+MerDh+ZPddz5PzxYC4D6kMGee9GUO+GyYnd5L
e1oPvv/HLwY4KM2OcO0dsxveCfeMQtmx2V63fp+zFnOqReoHOzwF250Y08zzLf4xRWdxEjTKQ8KD
pC6teOVjh4pkpP9ZrQ8Il7aC3p8alFcvBG7s0W7tvgjFfgGkEKHx3uxItpYt+XzRycWloKxSDI99
a8mvk0oEIGvRlInRZ45cb7w6W1j7Ai7R7y5sDT/OklY4WuzCPPmf432kj7le5f1pvh72itQ7ldVE
puc9t/R8S+fpLWVRtWwT5YPh+S60afb2r73RJLZJhC2WjeffzRn+p9tDhctwgRIE/52IdQyru/Mx
AumgBceG90UDCx4SV+W96gjOPwG2C3POWh09RHLlvHNTBk5rWIOT5zcDcz3/39URM6G3ASmX1P6R
tUqDosKjS5gu6ArhGjOUbhrw8V8iqGUxBVHSm1NusjNIecqbjy4+DJis2ZU+0jkU64JktJsN7uQl
tAKSbyxZh3fUQVpsmvYJeWpmfZ72wRKQlt1pYOpdieIiIBKVALNEo7msN8eLdV0M6+bg2FZLdgbN
B2XdzXy0ITbhp81FrlLteUUB5Hg5+1G+0R8mtYvX8Olaty0r+7ptfWhdQ8Na1PICF9qoOu2i0suz
ebQ48DpfJY3S5Z06MUj/uQqPqAK39YkfSz5dNP3KOVymzBHJnwJrkLaWSTZ7Vo+ZN4ArRvhMf2em
S6SMDaXLv38nc3gjM2Ds4jK711qR4D5A2Hqnug/xbAz3w7IWmnDfMyRnDVjUbo5JzkShYLba8thO
/IJ3qKGoqo/tdeRR6uJOeaSASMSbWQZvePSUa0Nt7KBNVpa6qoKZOZD0DLkMwrJamWc2IzWi3lNi
mhzQgBCPQGyOGqLwgcwyM+dAPk/kadVsB84i5GztYiLb5kef5nH+3gKW6R1VIrpFGBujEgcYR3xg
HasdsJiaRIAG1RjrguyaFFLtEMRaRDaCk+flCi5uwKo2/5MnTnoaR4r5xk7rVMVCj1YoFdymsK1O
7edatIJRSf0ScfYqqGJx8JlvzQK5b2oY7FARw1DRGVPUd2jCH2v5o7gBI2BR/IhAbDz74UCiSLow
GwZuoWoXi7hFo40y45gTMXjEftCVb3VsM37AErARm22pFlToqEmk4tth9Ei9zKcjARlHGvILXk10
zRVrLJpciPpb564loh641OfeJRlUIgb6UIbUkhFf4FqKrcw3slIC0ysjay2T9KMiwZ+RDNEiwQUq
Cpxi+0qMcCcYnGjpPltJUG7vtb1W3RGo4mHVJEMV1JHfgCgEjuuMIeq3OCWlwEFhjsXCdxDRvHUe
dzvSh5+1W0GOubhuO8Yy/Vqmy6lsu2Xy9IurGBtqTgqFfeIwSSgPdLis2UztiglDtXh5lvZ6qe+M
tXxamQ6phfoE14d93x5Y379ahEclnNgqDltotugbPa6CFuZEj6jB6LtLqZV2xvsYGJKw/oPpjdas
fWhawj45jMHHy8zKug2IaZEqbOWTS6M37g3nvxjGI4oyCpLu6bjs5n6KxnViHYplOaKeE0r4kFf5
9s9YlayAPY/CRz1vC3MzZphx6NYT6I2WoZlJBDbIm89tO9H3JAUhLeOzgKMtqMM2zAyDst45mYs6
LB4uizXOC1SOIBeZCRu3HVnCHs1LjQKqbc+vMS8nkWtPILy2gJ8bqhWAvR7b3tsfjJAO5kjKpjsn
HMZgvSAUXgBt1Kjr9pBXplUiZ6ugCSonxLSv7H21kL07ob8a0A5L9Y/5TzV6NZXhdcy4It6iXtI3
TNifUiL6TZ98WtEx/jBMs8UCoPr+w5TC6aHihemf2YyEjZDDEAx/0CWZ+2R47YaE6biZF5RNNuNO
MH6A8PH2dtzVPVoO0557QhSVdFb/CPICUSZHk3L3VMkcVTzOtnbFnYFbBbDgFcKiLM0Dj+G7WXQj
LNIPWzB1ZJcph1g8jZ6TvfXRshBnVTvj4dcPwAChNCNAScywBg7KTgjXdl1P8VyO9Vuu3zSFJAh/
USeKocQSqRVlgf1LuT8q63Wn9lxmrHubkouPsZX/iQvh8lF/7glx1ba+bspi2ugeM2G7BVnTjdY4
VzBd1XyHJig9Ua1DmXCCE3E10J7XpvM66tupMF023p0bVjoWraKzVjZRFsN9RUhqgja1ojzQ35PX
MT27n9Y0KnVtqCL+UhCdNO7x17F/6p8J/0zK2x4lDLNjMpfrxKmmaa+OWX/FkoAI4+rysJzDSc5T
SkKNUcfXxnk4TqZU3SZVP+fbPzVU8eywTvztFYUWjanb/50DyyuUE96ar7drzuc9YnfH+m7UVgEi
rlqQ1+nlSwMGhhcaIVZdwWfMGiM+hkWBpCGFSJNPBpVMm/qWUAmvNyzSK0w296jtMTie0aDwiUOl
TF8tIrKxpoTtfIlklxESCIYj03qMayyNrG/jaK0DsU42LTbT2mLIBoSOmOwXW1aNBgKLvyRd4H6I
oKl55MgfCHjdEtzR6Faeecp1fnwqe+bcu7WIEDVqinn5aYo4kQC+MTjCieyK1GkJWuILhQoxK+ZV
ub9waOg1u9mMd8rVuGCbY98Stp6NEKx+xjbdIpwxAzsUYZB7hwCiCk68WI3pmyD7ab/tdO7DBLzJ
KpC2nqDez5DJvtbn5/Aj5AOrm8aiJxuG06TqyHMmDA7EYmlYt+6ug2m+/eRQMUtQKq1leX0GHNJ/
SnXEIraGpYTRUfq0WYHDpVy6U8VJIg8Znd5osXA0548M9IhpoQGnXFy4lhQlVMZr7bjKVEf8Wyuf
cn66aWgD80EQFwXGv/zTN8gnMPETWM3OT5VfRtlRNSmTn3Z0Nq2shtoGdpzFpv1jgnqY2+DyBApv
qp66l7/R8SxVWvhZ80dqe4O779wMS3v35JJH7AmRn7mcughGbGvT+6BwrbucFCJEclMPrehlbDPM
d1Ftw16VWeJM38xIWEHenAsk9+0bGer2k/2laTmoPlvcCoUIKXJFsWkgIxhuvODtwbB4idJTRrD4
KBagR59ks7ImxMggOVb9bp0A7zywKQx2lY6H8e8C9Ek5ZEFyEjWhK0U7cwNwAbPfSOPwyMh1mUNt
UrrVaNT2aj8PJeFc53qJtxN/JH4Mm7N6tNuSVkVT9uJ5DmOZMJIM3cBAAggwFPmYduYWJ/fq1Bt0
ddk6NuWDKCxyu4ODHuWcAYxLpWFVxR1vH5vRpEQmrXKY9BCMTVlOeMslenSYy0GBBJOuPO7vEAKZ
SrJiGPY216ZUI0Njvawry+jpwQGrPp5+yuecFapjUaDJ2psLS4A061YSxW0i8zF6k42b7fX/Bj+e
czpANOJhrllmHOk/EACNCmP/vslgbbydGOMyM8WXq6LV8EZ443e1NaeOncfRXj5+EXhOPN5Lj10w
lhvajgWwVXvx9ghKi180WS0iJhiIHqBqCogW8lcNna5eO2zInKuFKxLDazao4KEZPeBLGEucXPl8
UYPCXvOV1OqqXUgHFepZAiT3iQ/B/H9yOoD3L7uk0Ct+931HDaz9w2zoq8GTi9IogMoSPSQQna6a
rpQpjXz7V3lQSA074DIRVNk+z0HSlxVpY4Wg2KLbr4yPirT9kvU2AlIumvSzb4Jx1/HO01xx+Yfe
Jei0bhB1EcUOuljRRNpAncDrsg9FxsNFo6Qn5RWWMgtBQdUoKq+npQNS2WT4NVZCyX5bSkY/OZHC
WFC2JsM1mrFA0rBhj276yHHcJIxBcVh3EpyThiUNEKDhXp9hu0H0DOxlFpwjgx2jsUxbKbEMt7Bu
XDoYm+LycjrN215WlEWQbDrAV0I2Uclhzi+EQyiaRJa6BiA7ZC62gmo0QbO2RAZJ0KVoYlQyovix
3ALoYH9lZfVWaWM4Q3NEX5SMVhdu1zVzCOVruWhpn/bXRG0gjhcx1RLdnWUdw94SfHUV1VNJaI2y
n8mI2PECnxMKYGtOV2okSuZyXPtdonGxbBeN2cXi8Rzk6v8kXEQhTRtXMxs9+LkXRgR2WMzKWHDE
J/Gx5J99r5ycJDBOVWpe5ijDz2o1ht4BEv76C17k3V7dseCdBFoYPNgjmm2nO9ukVmA2DoYTMOpT
EJOwi90Zl7ZR2dARBuQf8wBjYCkOp2rGC5hNakk611ZIptvx3uCZk8r+3i726guNZYrEOoPPfI11
RXCGhlv/pudqYJOmnByY7NCny1z3LECR1lORSC8lCaq31AqXRbHKOsa4YiEfz1TbGwBjJ6W7YoiD
CvCgpPZ6El+MOx6/FQS0S3rvkaxawFPojN63Bbif6CvMVD02XKP8fS3O0i5eBMkcazmZjNyAZFAz
LyvPVzzvVqSMdaUf1vG88jOEXx10KThGgNvAJEqOqtH9B9SkXpgZ1Y4koz+OuIgZ4tQM4CWyhEW1
vL1zKYlH8LlvsVTqZTY6WvpkaVfs3wdnavfOK5VnS8g7iLnfwjhwbDiY7lXE8biRE4bAYpWZTwmk
uoJjtiLB7pv1zDK+8M2F+J9Ebx2uVpiu+d8aZvobMfpetF3OUjVfvG/BUicITOMzTURzz1WhqRVF
tMtw7e5R91RQfMKJUfbnTD+CYCPvA5yAjb4iAAggrYH3r1nFl+zGbx+I/55LXo5jfQpeluwTXQFw
422Gs9TXo+8XNXZPRVhoyEobIVR4NIAlLAL6t5yBTb5Wg8SQOX8J2X7rQ17o6zSOL9qla5OMMu1A
ETgecG3RQgnt6sailRx06BFsKEurRDBy+hwLNBIak1yBxQ21YQ9/vWfZeRMljODJnAZNe93oARN3
OloeiVDzyuQI8IqMdfLTDZHpBN4Xmh0ROMLoN9NKQp+8dzGsjWCtMfMTG44/OMjQpqKGMYwEQOs5
7WdB4w6fl+eM5NTLT/9kRkGT0FnAmBBaasD2ZPndmlHu0oF7GyuXIcsWJUEgWVCW5yH3fT3S9+vY
CB+goPql8UDQ9BXSK5kHYUzZLblTsug2kqDWCUoLx4it+rR9R56xh6E9aCZSPTbEd5oYPYdlTwpR
rKK/Uesvv/zHM9mF5qHM5p6F0PGi92cBXmKaEt+62YSlsnBNctTTYdv8I5tPwq4kAY3rNhZhvSZE
kk9gEANCCiqL4wZt+zMzVcqPKcTRGj6U/u2rSLajzNvW0oJEeTzeY06zk0qAv+Y+NEW3prKq6NBa
5csAdJi2sgkyOYv8Dxz+66EGjXc8gROGlwVdKj6WjydS8rpb5zmINrXPahR7Qswl5fcDEwAuWcPn
k6cw8SKtpz2mU32rS5QJ2ZzmKxJjavRXkSp2TPpukdZ1n/sDd5uCbgF2y/slqgT16spVQfT6MBhH
HFuZTbwxBWn3bXPAKNOScs7sKlJS9aNgaA83g7A2O+I9Y69SpfEvdQmN2I6ecsbBhCYQNRcs8gKq
2EDPSdFNGJnoEtGKQ8dithERMFTt5m60HPMPNHs2PCprgLlk6ypl8DAHyHH25vHKrB88gTFBy7w1
zNhsZ1xjdcFpn5AiKs3VNEb9UK2Z7KVx6skCf9ejidpzYK38AG2X9vGm9kguktt7oM9pS+MW7v23
LQ1uLvfpqD/gxbkR38q503/xDdVyR9vabDRMQxkbFwZu/uPYd6HwoYVeYBCB3Nm/ayAVq1rd5MZl
kFMnNl/21abKb2+shYV0pnfHLUNMgaGe0Knfd8DajE1yajClvl7B4cbak659jmC7TalorP/3R5cX
9jU2+GCcWSnpnqC7UmCmZCVnWCpYo7cEzBSCQkVSiCKdSpg1/vuQAP/wJ0ptsgabM20NonpPUUYP
G0Dr0iB2Gad+oE5E3cMwajrs6drkNT426hoGmewh0ADvYDrQbDKo2PJmQqgNI6rN3sdQ1bCaXYhM
FFJDMi3esyjLW2cQI+A6XZlhhaV4x4Tuw0byeahYbqR4W5o8P0krSDPhPkcqCiSibzRCgbvlVcg+
dLt+DinyIfq7kRnhh2v9/pP1bY2H0R4Fllkt23LKk4DCjCsUNwtxVXH6/paXyCaGnz5itUSzQVAH
dBh6+PCZbyXvOje4MW9NxG26fD//KXrsLY+HVe0EhwOCYs/p3PZ8KtTPz59VpcogeSlvJ5i8m+cN
B1lm6PIu4fB2UIv34Dc15HVc01YxnloideN5fUiDclDWviLJAUEft67/MtSF7PmxK4FtqwB1N4nL
FR8UjvlXl286e++ONKeNGf/Z1SL6Pv+jIUXzv07F/BHalz/c9lxU1VRFbeAhsyg7ZFRXW+WPiAEl
Ha/HC0eV1BvFsbEPBO2Dei0V1DjD9mICmaRpWO+en/BvwSSAnZDP36ktYL/qJ/enSwKLJ49b1Ejb
s23BH1+a2OlTqwiKbxcY+yg/YAIlsBPebqXZ9Vvs0Li87+zcLQa90wwssF3Zv86QIOU8k9XBDjtz
fYSdJVBMarxGKGeRSMqSZM9Co5SwWL2fuYEuEXAm0CFag2eFtgOnGq1ZtyksmSrnjVZ+O+117F4w
XGSe1/yoF7a0JO4Mo91SqOzm3yXBX3MvuYEr3WS/onfA0Fgx7b+ZwxDjX3QHhksBKKlWcRCaQ5vN
BkB4gwMPzDwspHcSMoTuSoPCB+h30l8P9ivnz6iqaExhsDaE47+3GWrYZoMI/89NKguANdv7xdkj
jRLbFNxTjFnPdLt/ZJ3Ujo1doIvXCxm8RSz5BqwLb5MdZVs+UYgN467RXe+6GlMGbkzLVSIHRRzy
OIm3gV96ANpmgCBsmtJPLrFaIeATuu39PEIQ2tYkrIG9vfC1HF71cOT7SA5W1zSoGm67Hgekgi77
U8zVQgu9a4VJI0j5Jsk/vfHkQnSPvSB7VIe6THrppHd7Tf3d70vJvkkvA2EVk9vWWWAPWSFmVM1A
TlFBxEp7Fbc3igJfSgKfKlf3HsesN4u66AdlNqhHRfIKgYCqzvcffMeQQ3MEp6arypj7lVlOXgqj
J4LdbsJYcUNEfS0kFqS5BPVqIfqaaFi5ekoGcAZXepF324Ye30jmccWRtpvgBSW+876O77VPzpKY
fCdTzFchSCCOVg/K4JCz/0ZzdmwBBBBYVP3LIVnjR2cwi/+Han9tHxDnp3HNs/wvAixloDCLuNYs
7OVVCRMLXgMCLXYUBznkkXH7AnqAepCDkcM2dNmdvTEiPbj6jMNitzFF7joaQP8gdNXVzBN4oGH/
6TRVsuV6QhxE1exI4stpBbvEIiQBgLH0Wkc3/cE1+huaMA0kgr5tdV2TjCwWAzK81mW3ZB/i7Avq
AiS8umes6TP44DXyz1ewmCB8BYkWXhO8pqc6wlMEjOsVWi6XPaOWIQ/077SOt++nWcZscZmzo4Sh
u08vDBRbonWwd0oKm7NEdRc0rpg7yqNagSfNwR7ydAQQyYgc/Qfm5BzioIY4FdsMoZ5F8lyE5UVk
xdemhFH0WpaSzny0iYChL4ZHlyQjPFkZQqEbjavlUc7pALbeoDpOg2/DvpKIzRGod4vTsDk+bxOX
OoptBXO2DTU8RjcGc3Nac7wiRRrE6KdY0fOwBPQDt1n0pHzVC9YDeqGGkpOheZWAeaKn0ZNpd4wz
uveTcM9wog458ZULJhSdhqU9el2ZGJUsW/vIyxF5cZLhKjJaF7BaBnawv1bx70S9JUk6FWT+dmEI
NkYzOv7TrdaHsS6eA1WHzadczSJ1GoQYni5qvQukmZxxvZ7rXsVBX3EK8IxQ2rnEbyZxcIkWGB/1
oWU+Z31yBkMrc5iU5b/t1duWaZ85NDp+bvvwTeG+96INUFQ+MYuPgFMN3SgV0/ggIKaz96lq0/u8
X7u+SSzcRimrl5Fbh0bfuo+fJCNbP3paHupcyU+WG4ub3ox6j0lYjJk9TPqrCSL6F7+GHTH5s8C9
TzD0HRIly+Bfd297cqJKYIwVY1vPJMz+6Oru2TWIaeXCKwjHnyS4eubicje04U/SELvinx8Txavn
9YOECc/TPnZM3tUQXUhJm4gWHyU3wyowWRWSQ6skl/+MaARgl1MZBgaqcNzJSyaWmiKjSeX57gRp
XHtUtI7S+iHyljFf21FlX8pwPk3EmNg8lLmj0qoDZ5MHy+Zy0njRZo8Sdfz5epwazTvnN5YEjoN0
VSKt59Zm3BUGEbzGo1VobliFXJgnPDRSboC5n7ZCFnsYwBJWBz72Lqqkw1+yLrPsP/kxvfJB3b5+
/+34iIeXhbuGLOhBtAZP1GwelvDc2ahMsGEUImwxMBgzjp/UgRYYBmvxHYEwDOSyiDZ3zPzPUANf
zIpvnJT8Ae19j9njXsmhWiATHH+ZVmqIZhhKTBlGtX0lrE8mGL1NcKmNXUbtAo6W8FRVhskaH0Hw
JYzGIDRyWVecEaD31BB4dClXoSo0IUYUaYTzb9KBDQyXjMx8lpMipSB8nwwMS177+4iXaj/XqizB
ClsyhfdGvtpuSNpojFPpcpqccTvLSFRudJHJXiFvkKWd1ttKrI8+GpK3aEnpkoNh6pky2xUC0eVz
q4u75r6W7q3k9ge9ejAzcFM11pWNyQLFpppmLQuUgTPDghfuFsai/8es/uTxFtZmiHwayUiNzSZJ
lhPpVWntaCwjok0lWAm3k20Dn5esSdKMLLgHozWd49Vve84+35+ITCO7mfh+DI/AwU2M3EnDJv0I
38ZfP3cLJU8Y06k6sOVx7cbIL2wcJXD+4P+ZyNchAeoJ1yuxl7ErHLOZ7K7wHt7VjEyDpSEfQgAJ
T40bvC9Qlo/Q6trLugydqICx/XH8d63BkClh2P7hVUIUpgye2m0pRx5r0b3x4o1JVWbS73gb2AnD
TDjPntfX2GD0O6rxPdDjSaZxClJ5smpkWktO/0YAwWJ3udn+tVjmA467UESTpQW6Bzm7CXhV3Ivj
7Gg+Lke63nC7uU8Fmbl5sfVRWgl4LTTicNEChEC21GEcRFP+S2bm+zM957kjS8IrctI8nTdiQ8kL
hfyNwtteKPr9CbWU7VYcU5UR8qIaXu1OOBeGusaaDRGuBTpiGbpgmguAcihanpJd4j7WlpIKLlaG
TLqlmd3Dc8odpwhkbfOp3qGkJW5goKuWOUvyDeqDDQ5xocO1LQRLLaRIFqTLkRMH81IEn8WxSQcX
lu/LSZl+nm/6IaoGfVaIIsEfM/yDJQaliObajjId2R8udrMPHMLYAOsVcFv1yB4xrU6mBlzn5ZwK
DaWc+Havlf25ETqROAg1CJxTuVElA9WUUoSAxcnlSxoA9tuLkcSKTkfc/2EEmbpJRO9IFE8PVLg/
IteWePzzgYEhhOQc/3jnn+FVCJwXBNZZZRgWf3LPPfb1ugjPUoOMcbJ8wxAZWvkT6FQPwt2hGt8r
UTbb17w9zXI90QcGRN8yxpPT6i/uSratgNSVxF85vcotYSN8sD5hWR/FawMEQ5XCNZg2bju1prjk
1EbeVvI+iFYFY70Zmz/pP+K4SStolarVBj8sJCOuiNrwVuddl4Wp2/RblOlaq4rmXIgXbCVkU37Z
Fjx6DqIeei/8KqpiBbHod3uY3TLMXiRhmKDktc/laQUjclMOcqhrbhQBf1hqV0GC4ZPJU4uu3zYo
hBcDhTeEHhDeipFp/wOEF6YnzBceZI3AvoA7SZsdpIi0F2Ji4Zc8jAwqMksqF+VtJjR2wZVootMk
HBhT8MIfvpfbArHEcVQ205zMIGfz7jGQF7CJV2R1lT3xyDcM5jWtNCuSgUVs6zIatKxEcOIbPQGN
11wXn6kUIGukvQ/zBDGRC6gtG7EK+erNVTDqtkTFsPAOOw2LVIw6JguoNc4BvsbsioAIrE5rcSmD
140JYIqX3FHxQUDWWEe+tVT1gzW60tPxZ5lBjuOLvEr3PyBiDgM4CyuE3lKtHbcrnn8TUyj1spal
FUgWA5EWkgkfHQCYZU5smmWw2kXBuboX/2W/noYFX8mBplvbw3xjnLb8hAYD6TMofMwCigDWDTCR
tMX2ZCoqjgbXaar6NmGVKZ0RNneXAcqfxFsCQKMlKCYFU+c/OnO6jfe4o6INHqrzCK4BXKOeggm0
0Cq/DIU8iuLy1BJqKTAsBj/TG9/ABioNT/D4yXrYJC9VbBAiOlXAS38avEJtyq+9putMP/Uf86WH
c0NqY/F/ia/hRiSwPLXMEBaZRJ1AAK/SVRgHhmN3B1aK2+MzQ7vkmnlQy253Yve5nR1CjAuFITJN
b9UIMMFkbRDMQZmeu/y26cdqcWg4g3k+nWMfTSki9G/WQL8RhUDbIRVg4Bdr/aFfVQE5ihDIC9Z+
k1FPGNO4UU5xCRKCUZSgRYIzOW5LDTfeLU/doTvUrtGHAnL6/VWbJpNt1WjfD1D6wyc8GGPKwcfd
ytq9+lHCjlC15DxIbilz0nAIaX9B2Sze5k7KnjXtSZm+dSIyk8xmfrzwtLozHH8u9Foqpi/h8KmY
lcYsy0QQ4Do1xuWbRuYj6FApr7r95aAENtHT3GLbptANBkilMo3fp/5nMy/cYxCd+z1d4GYQk1hu
ISHc0LppRM4658tFDEntkzZbc1kx3EdkW9mPnlvGCmK3IsQms6yfDBODkc9whGO0HOaNgs7OJ3jz
Vm2Et0ryOdRtXvuQIpiZylQGkEXjC3+j7ZtvfmDlroqbSoqDOt7qwxD4pPGEAT1dvs+mUiglo3ED
3aMfk8g4k69HL4bC0R1sNieoSZnXKN82i8GeGDZXkhKMCCPHU+ue7uAIiwI+enNV+1DPu3ozvFbA
n3k27J4IOJBUfLd5e9lFD0zdjMq5Wfxc9d4q6g2n6jJoFOOT0gv9iV7WdXpFiD0Zs9P4IjHqFcDJ
jBw6cxzD7ukykob94pMAI2u2k+EshQmohhBhOwHvqC+Xik6A7U+NFmhQ0Y8u/0tpWC4sKJkXIaqJ
F/cjAxLwN4a9GxrgtHnNmPexb9UuB2rVcGSlf//htouCsW1edo0MosqLxWow05KSM4i5r+DvhKxj
tdKDPAC5qHmAWh4C3+uVW3yDm/DbGDx17sXR5NEiqEABsJ1JmvHmi4fYQwYNQct40WrDmZwxU4CU
noAHVG2xvk6eX3msrtPhpAkqE2ltYlWN81Fe/FrRqir7go8g0UXYTlVdsXzYiVYVbnkYbmExmtGD
k0ZubWixGKiv2FiFBNDtBzHwES9ftTJg078bIHB6ASFa4KZOXSvkjLnIBIUOp/vi4CyKxRwVtcw9
/LyFkXiRqpj+UaK2EkFVjjRTifBTvDh36L7O0hGC2qmFksk0hw7EpSEKezMvsTvcRm9cldClq76k
xYAClW2pXazevwuY4/LUAojSAo8DS823E94HMU/yMyt4l9B3MMptZLypPUTBATkuHcpGnffHzol2
5xkqRKj7tOmiKjHQBetalk/13CzviV/P6qTCLc+wlkBAguIADKbyFcIkBRYKx4/RbhFdz4xWUk9y
/wjNdz/l7lL7Dn5t05f/wDxqCfr1xvwmeq3/WIWNlLJL108BJ1zxCvNAKyuaEbT3sdCyR1rNuHlm
LBzzuOM+4MYtGpTqKb7cpnTALQAM755NY78ReT9P4w/xTVxFxflxNLW9rc7wYLhqq8JiQCVPO//r
IzUh9IjomyCzNlUG0MHEwvwSs+b5vnv2FH6wkEn03hArREs7ijHUZSyhrQQw0wDt16FABJpE0LEn
UNAO14jKMDkGIjijR8qRbHpt84PdOHTkoFMmXfqQn8hJKfqd5oYi0hdBzHvnor2gEGHVrgsCQg5Z
+90+NpNJ/O5SDaJGIf5f1VSyMk8cDfCebSDH4bKe3KPkvJUOzEZGFUtZTK650d/hy8aRKwoHH37Q
7EFsUao+pXv57+keWCLlWsn3z9GdhTP7Qwdv/6EIpO/Cr9tHdhIfffeq8NisGnFjtvoSA3vYB9l6
5Em3smlfTDph/mkBVCOITtIQK8VJmrS6yMUABzU4wfM2nD/wEGazX42IGfzkC7y/DuU3D8QRVkRN
vM59Lel57nytzWmVBWeAmNFBbNZV0VSkJ1OdJuHU+dkWhAzRYTaeTWwZ1CVbYA0YJrj+hag2jZZQ
YSJQjhL3BgL5h1KIVhXiuMExRJjLttH+crSztqgRtAXobcDxKL5O2S4AATUw0tNtLmH8idfjBeMK
QWyXeNEBNpGwJ4FhKIWMKZgqBADhmdzD+kMKk/xAUusyVUyyLEu2+giJaz+0rJtkhWF/AtRvQ8S6
lRk9c5ycojs0lD1IV1rV6tJMQPIUYTGhG/G2U23d0UZlh6yuqRECmCmyYGOra37zjZG2vP5O2rJ5
9zPdZKRB2q+2IoirLSgIap4rUnojrkP1HunS0NIHdQqQHQKWPid5zlCIDex5GL3t0c/IjAktKNoT
oPtnKsMwqdFIOfMz9NCXPLDtvJ2+RtAo93PTtUYkGmCdAqwSJehiYs4FAoGAPUhCSdVfXdJzq4Nz
E6eJOJyZr6Sdvg63iTNEZKC5Wd9vGVBzA6/tBfs/5erxbRqemaalO8fYgxPz+HnTmAyWq6dpv/Ux
qEJtUu+0SjXGMuJmJsrKK1WEA2QzWXM9eixnr17iuGNGhULG/N0gw9wO9E4MQW0iOmWr3GXiqaVz
PZhvBTBMEK+oEtDkTGBToWOZxXY9j6hB/GWnz17dtkhvcVnvhcCGmcNnN+WIcv4KZ4veCKDjp/n6
Tg0L0T4/Om6zSAQCTt8squ/J9ALUD6cu6W6Hz070F9v+OpuRLxBNCJg5s/J6u0D1aM/Cr9oHKOYg
HFDdHSiXtZXMAlfubTZx3HZ/izKV1+TY5+ReZia+672UUYYG8UrK+3JwbLN3C21v83ezeYggpMje
BY2NFJn7S5yAAxByNFH6ss5pQqJ5RkyuEy/iZy8N4ifZeetCIXwLgGBzw9mpz2d+FstXX96vwGT8
on0eOJ2aNhvSuS48yUaZnRfHrMcSKJh1gLuZLSDIxCfALKYlwj3ADtkfd+BEVTBqDc3AC8fIcyJe
JW5giZWA0ikuSrYQqiGlxAb4ry72oAk//VX9P+g9qvKL3ngC/KAoIlmPRjRSxue3/DKUdfdyg4t8
AuZHEUjTu/UgNMVEx2yxHqqUaiUcxSmk5V08Cgux7OonBgOEJ2+V880FMCKmEwGkUKsa9oVW8d5m
SoB+uE03fPPOeP/qRCaImEtRaWpTwLUNlZpsYoVUnnxyvs4ixxVosSRTK9xbq18vrSuaEHxvJkN/
JAbQ9bJuDq5LZ7pUS7xgx4Ww5FC4y4DaZl6A9PEJJ9D7nSKM34Sy7EZbhgX27MN1G4YisIb0efmS
WWxmWxNnshCuyajL63RsX1yM+AkieNvtFDOhoiweFIsukUvIFMVXgrN7uCv3+FVVbhur7Tr4uIxe
4WWBdYVhPo+VJseUDmsO1HtRyoZovEmJ/35XDeoUHA44eSYchd3thnvnW3NcaPTZdL3yD4L5kmfd
GZmg3tWVud/NZWimpHyCjsjLoOdYE9nyyJPg+l5Rl9YXdZg1FnQ5NS/YHnQuP8PCpyiQ8BzKbiak
mQ5bmehR2QQCc60ylyqh4Mb7TQpow7gk6H3VvsuFmTvc7TLHTSHy8KY9hQRSIglnKJJ0U2kSTeQT
1t75HgNVCh/7PQVFQY13SKAG/TBHd/Uw1Qjrlug9uBZLTivZEyLH3dWjcrOPFOF1hqO524bFk9Kl
y9AV/6Ws3lPpWJNAN7q5ZwVHLd9quQMeTrp6JfC8zLxuE/m4oZ/L7OmWWoIw5f7RRlbm8Bw4/Qc1
kUuzhEWGAcQwPh0ZjocBNHluFiAhSQPCJYdTHPivSdIlqAukV6+8Gtg5WFvQeO9aEQWQ6lnLuyip
/vWKgmEBXVFrUcNWMU0717bGBoj6c8/X1oJmF6RpnGqbQV50rGuQ25rLwXe7Xs3ISbFPj8VdbxOc
yb03FxQbJP43hacXnYl99kRRGmX7coqfHCGTDWFqp/iKwDJGtGu0T+cJ91eI8wmdNd+CLzDQmmnJ
m5j9bFAPl/oUcT7TZozrPKnTjtT9wIingYtfH/sbC/w1FfzI7QgwujZfpahbjbqjvfgd3pffEODh
rKE79vwwQJ3oC/fkWTc8C8GZ+ohMUEqbMXHl5QAZ2Xv4sconEmMbh3mW/ulywrLO6IOBfluJdPCE
hB7xRJ+vCMR7niXbFm2qBLxo5+jzDxE4Y5E3YhiNZpdCeas5iOBx6B1G6ukzWcLk3R8ao/MGWZZA
phi9+4AN1r0CONrQDiuwvMC+cMEWo8zIKY1u8LrG2MQ0/arCMR7WjzeHRFLZSTZmUXRAffLcBkKt
izN4pwl/pZd8CHNXDxyltey0XienMSrVSwRwMjFSsy/FDvsQM/iOjFlmHMQ9YQgsmiMsSlcsLvcG
MJAyTJkeDkcrLpPIq3OHIov23RWSRSd3Zfrz2OFSBSUmH15VFy+mGpW3nxPhz9u5K6Ki35mmv3Lm
7lZ+gF3IG0b1PJEXIZPMLMT+Gg0z+KxsJoAgrhehfPOK44eIcXVGvEkWeucw6+aGQSfLAafmM9LN
REe/tWMJGFCCfyodlUogAuf0LolAbOSFH/mmtkZqjTQcgHPD7Ut3lxMhkAye7e1z1OYPZV99Fc14
c00xpQzRdIfC8+QIUX0gm8OGX9RZqn4cu6eHbcZXg7QCO+neCl7tkL575nvawvCOdYX1l+gh5Roa
0/3fZDGu3ZPGJH32OENXdtHW1fYaCYgC6zBoWxZi034fD8FMye/SmqzQ4cGgCdvlKNE9JfPhkVYr
s68ASts8+3OzwIcTzJzCJKYudOqZXK+3jyM/7C8d5Z/z871cAimKElS9du64pO1kFPYMGaTHb5bt
hiFfCdRYdF0JOKnYu0Srd9tKxtEDr7uaIUeqVeLkpb+UsfpHJVCxBDHwqE2u4+tkgkp4U1OPD/kB
X4rMzA70Z6w8yPoP0VWGWfbQDodMAXMi5IxVpgTnYE9Q4mvrlDC1RBraPRX43tr80tb2BXnXEp4Z
P7uJKdeLwKlyhXlboMD45zB3DnRBxeY+JzV/+Sku/qKnDxQ4XayhQd2PpbbQG3JRx3E8yw3zsgGi
Mab4VcTcmxwCr/vDzvhn1fsrdCJ9gJRcrYXOZA9j0tzru+2+g5n3WGqUCvuB3SftcY0oDIM7Xiyb
hRo5PsZXWLjGaA1ctAoG1cSJirECiE8IbGe3v4VeqsepS5p8rymkzY/ZwVOMOTR2GICuJpq1oBtD
cQF539O+EU3KdtaaDg4YbdlfqK5EeCJBt5aMy5Odw3oP55dsLi9xqBqZPz4kyVcj81oeBRAyTmWq
M5vRqwI3ICJwi7r6BLDrxQxdXTW5yDB/VSgNV8dv/jt9gWWb8OI9tfg24WU4FmYVPcSaB6znaf2A
qRo6GIuRkmV6qjOPxC88Z5pvfk71RSdFDBZIRHql5GKnW9Bq6nWLEWBJ5IzZu+7I6tASBPoltOVe
wO/5w9o40U5zwh+xizA4Rc8T+Zpg/ARjWmDGnGbCgQ7ZIGEnmFlII+rRujGnouJZWVD7Pej5vHfO
/NK6Z546X6jquRLsish8NqxduAUaVDkKvkyqtGRveoQaquIvLbT8BqjcwDUECK39ZX/50w2bvg7X
iebBmSR32IvHiSQVIf7tquMA9VKrZwBf0XpY/IS1ev1oanCoyKGfN1D6TccNUV+XonsFRveFYJIC
0iyycQsq70FKjc0nhVMkEsJbfB5s9SbtlJnnkRg4zysovLx4K116iYd8rkJaMMQR0+tc/3i1mjF1
pzvV4u67tPtTCWvqdycNtsVkUetbmqR/AxDJoN5om3bsTXPAj4ir/RjiTbAaQ/IPcm7yj0xZ2LwO
1Xqg6Z10t7oydGrIZ4Koegn1XHib2EeoSrYajdgbdtuXH6I6SaQgM8lkTKsfYfuF9R+r+fWNN3tf
OtiMfY0iTrPzCd5fhqlMDwA2aV6FvtQ1J+CmWIopsg0oiXlG5v0hev8pt6l6xV9a6QT07RnkRpEH
VNFef+SPGuM8eRpldikTf7dvfStBAZJ5Qq/H2IDh7MZ9ePu+TgD7aCiAmgo6AF05xmxMa22u9cOA
AATTr30sK1g9/X7W0hF0bwog1Z0c6Vla6urYH3+KbRnFRhiKHbyw7nRQr9E349zjfTRVVwZswvzY
cg1PLwtfaxQjpF1jJ9qmDYDO4aqKkX2NWlAV7X2lMOLRE3YLE4JdbxS4NAEqe218QaUcGOihYQm8
VnVoPmERWZqbReSfHX8fNV4fkE24989UswZFp7EQzhsh6YEoiOq4osXc1JsrcCPCS5hCUXc4vzuk
LHBEeu9DCsaAkgDsoz7aHXJrtj5OyVvGjSyX7xaJn96qgyBhpOt3yUsq0R8QtgwHkTE2gYssWvIO
+RvFnS1sAqkZ8C++1YnVD+gfJt00PHhdW6KIcIFrVTln3+XPePCVopGzXpcUaerCnqHRejbOrpKe
kvOJjRYfYJdi6ddg0y4yTtVdaXlvgxVf4gViVWqcnbMw2coWNhdtU23q8dbYUUy36/v8aXoawQiQ
mBx3+IC0xIPodHzclfVLJOFAGC7TX/thq79dwmSbINDl2XC7bVpQIsTfz2eUkjGsjLrGQedu2JuW
9kwdBMEsD/EUPzG+3+x7fHe5dcStz8cTnCotTkDqxdfy9vHxgniXu+0FTZ71TK7eXPmfdCMXR0/s
34uO3KWsHVBT6OvGTjlXwf/21wGrO5a4dka5QW1R2+8FMMjOgke+rnZPiF5UOvHWyFO0LKF7sLBM
qKxEbcE4t12SFWVMbl1qzkzYuxeY4CwLmuQhk4TAMF4jxzp3tZX7JUUIShUScfrDxfuL2ucFUT4X
Ved1fcZZwPgkqqNffDoPvS2dLOZwDtftbNAjeIm35Ozog4k8mfJ4j9TFAqTS0laBKUMKVaXuNV4k
D9cAtcpJAsxp/ScR7IcuCQhTQYJly4RKcVVzIfzTZqmb6PsCeulsaXHIoL4EHo8L7OUeJotmUrna
lMHMl4eBhm8MlI06BChZ+EPB/WnJC9CbNdZKlSMKqE0ceMy/E1xUPcRcf4KKAXCVNKLLybMBmM0H
mUkbqkSeMNDSbyDWnp9bH3uRJEMuVP9v0qHbEz/7kB/oHb8dFcUmQMO3uZQArJXRG1z0LTyiX3Eo
S+LbU5OCK3l4SwmS/LU+m+LZbosN8jGBB0R2sOs2ih/9xtDKc9ISgHcVANGrAyE+eQrsQTMOFhx5
4bj5RwHL0dVvAWWNqm/fCTS93ragdWDsVjZYNADQkygCqNIt7My4ZdGhpqde2ZYssqSp1nCXlo3h
NRu7WZthEAJutOdImRq8Rc1yklaf+CvVWG0Xy9TazETCrbZMmzKlNxK72Hgwns3zkJM8raRzO5r4
WeS8dEGeZJOkzSsl4wb9OJ4w2zdLiBump2srXdegL5hXx9bGWvDzSTYBsSaEuoQX6mEQFxzHKOYe
wQ2V/Y63olMJlaBEHSLc4zNKj6UMuzdRXcnGklY6Y3xr6b5XXLMju+ug3JMFTBXZdQWt9WvSwUWm
IjjkWI8dhZvO/YR2boTmUKlxw4alcfu+xUOlbiqhv6OzA1lObFnEEb13LqWxbZYrxfi2YctrdZSd
YAyiMOZTB/whP4iUk1Xcct5zjAdrTAByHRv8KSp1fDsnScpspGKqYQTbaP+aMsuP4URaI4mf0H8v
qLJdISf2qCvm7coNLaJiJAEGY48bW/jznLuzlY1wm0U3/WWRp0rH9E1QPpJ+bmxPzZ+c2+X+BQsX
j3tjNHQReZDLyJnK5taF+AIJzW7NY21cuy5wObJSbat7i8HQjj5He1eSt4RzqaCQle6vL7B0uSI4
3WJvP8Mtm7IUAN2iHA5iodEFnRaodOIlWTJknjSD8azeDy5bsNQE9sREya12rNJM3K3Apn1Ci/Du
hoLGHbDCGNkU/nIBk1MaZaNK9s0TYGiPIsOo+t8yDHPGO5/k00h9gEfmtscgvi+cp2lcoSju7qA9
KvMehSecK94Jk3/cxKJY3wcomyGGpTRGl+DovZq8NVY3N9Y0mkicY1qE6/S4xo6FdnEuAAIuNR5S
JEXxX/EyJplyrwQFuSKSdB3M5RaDRyvIfOiD3l36mpTa3bd5PmV/q7SgQ0jdBu8/KB8Xi0p0wXSP
Gme3M2dPvEN9REq3fYld5aRZwOwCpTGBfvGwnWfL9A/esiH0z9aY/42c5kPl+jdTtbVHcXpL0oo2
O/imjskmGk5JfeD7e8h9ubQRJx2o1iE2LNMRVn/14tUZm681NxKBgwSn4HB+6eBQsVU1uuq7AvTZ
VqNKf0kfa3QzEWpyZwbyrbEVOyd64ly1JUHeS9JzZNqaVA7QjrNqIDwKgQNzjmSsBP6thoz6vHaK
utJjYJeCQFp9f2L8qW0nxzpXS+RzLDAIgpn51nGdDO98F5nXeh/GeZD9JIJWbnw2XbhaSTkWpzhh
Tki74PRkL+/4Ro7+mQ1qH4+Rzm4OFApFxxi8rIZup0q7JaTM7b5dILgTi6yd7vCNQDnTdA8JLEWt
UvkPLkfFWVmbWhJh9pakJh+EeKry6Az7PUcLw+Ne0tdvsUNhHpvXN9LBnyF9Mnildo0/gDd/Wqyo
yxXl7Yb26WML42BufF7gSu3QgXVUzZaSXgfnWu9wHpERtmODTOnH6AmgWsy/hDJM1YaZrtgVS1qf
9V2XHGeFK9MPK7yXJfq5cGJ3oGkBvzAEF6fEIisOMwgHuw1TnVQu3tWU2OcBxvBCV88/uaEzfjHB
2BFG0DDJjSZD3dH426vQ6UjQpV132XWtvtZwH2/sQlMMhm4AKBiUPqZ8PdLoBpHals1NNgk+YOer
mFLgcpcmrkoEaDz72Bktcr3/wmMmSirTdH+8XIVsBPhFG22da077+n5wjgFEni/ycr0tNVo5s4aP
crFn8LD2lm0/6+AmvJZadAfd5tQn4xo+k2m19WEOhlQgQISENRtO4jw+GEjTWTV4L42jZmOM776j
b210YZXgDpESG9P8GUNarWgz/WRlTs1uqBfy3CrvWcC46dKanCfeIzVN7e/k4DHyzX9MYfvxjeAz
bhbfFkvTeAgVwt/TvlheHOAxtm+AYcLm1GDiq/n65Wk0eEYoEYlhsscfwQwhFxlTGddUfmu5OaMv
TDlxd5FenasGKNVjbtkokCXdpRtMM6L+apq5hAPugb6I4KuJSHxjiFv339WNcGjo2+bq/jIcv4Yx
8JcqsMBRqm1xGXt4AYdEF0yHtSDF/PkmAifRtN/jSF7Er3FktaHnbs7j9bcazn9VlcKV1jWsWbfl
sNbLu24Fc+Zt/MQcimZRumAaYgnLuGauEz1nJH/uhdLd9sMBndz3OXOUDDaAFaHh1TAgriXruk53
o1/kWdc9Fk2JWteJKHS5QHFu7HkXj7u80Mm4ZZiJ35NN0OF1Bt7zhMIL1LagcQxSniSgSNg5oP0X
Wk90AFLCehLBFK1lmbJucUS6ErEbs3EfsCe1/mqnHkQU06RdNXdfjv9cjJkvMUhUWULLDdaS1qot
30Av5W737RnLdEeoGch7QnI6ZQFHgOUfwle3d8cF9Hxkw8mOirKb/Z/bT+cD5Robg+IQRpqCYSvk
nZuH2fL3fLIMINrWG5Lkai9aTsUiUu1zI47hjZM8AmPctVsLtpPFwZN47knaZgncDYoWhMEORAu/
wjknVp2BaN7jFurVLmBiil87j2USxtzv4PrUEYLhE0zNluD+XxVLYgexA94Tel6fXwE4GzVCG/Og
YML+pGPQEJe9A9slidncg8yNcXxeM0oDkxCCpwrmGAs+mJRiot7EFMwZX4tCZWujLmCmAMfcPcky
6SANPwQhg0joOCVUvqWTF2g+uaCwpdXDoQJcNCeruXhpsP9URa3Mc6Kqu7AMyVyi+fIdvcO5rsUB
wFZ0TiaHmLB4rrVRFdxPvjwWVcSf8MhoDreo/9mVTG/c1oM0S8co7kVP9+D5/FIOBav2kZE5Abdi
fLWjbZH1YLLfoN0y9xy79iDVafwng8P2iLLCt4XhyzHHSBmSRsaGQwhgTlNyecAMRUHX3yBeJUhE
EN3ljnfRRpXS3K/6ZEuQV0l0MzFxTgXP2fLivo8Ws7MY2yfjAEUZYjvLfOoguo8AIzG1XhEcz+BF
oBuh3dHnDkxrdvpzoDOMWWUmhV1U3FhdRPl/GDEBFlP315m7j5qmJzuOdqsFCal4atYdvyOVvml5
s7xCY2t72WjzWa7aYCyLnH33JOcCNms6/NQamQwhXajxuDLfRhW5q9rcId1gvTJDNtHkdTLetSfU
9j57NyM0lhmo8AzQt/yGENYNiSfZiuz7x52i+YcWnC/KbB0ju5KVcDdmXESRsUv3Wp0TC0OaqdOV
KrtwxAsyVQCXcB6Zz72nlnwPNTSCwZDjwsSo+9gUTOf1bcXak7rZqRU/5dGu60TQ3HMDfiOvBvSd
YklZQKb1rU1qaUUVtyQwHcfpGsrWGYmCCGbScsgno8ZQzUOevCBhUiJPJS52Ucx1mCjNBvf48UYx
He64bN4rT7iOoDDyfAYuPlPzpPIHj58mtdnWoCVpK6BwgzEi5wZ5Avf6XctgmSuOjQkQw3pEkf1q
HuRymb2eLdaYnanlkuyuHRgEZXUXAXYn6wNeLYg6liRU4kpjkknKvQKio7llg5+G47TNl64kfHFP
LxVpsC/+WBAI/fzB1nDVubO4/kT2DBrsA+L+fwzkJWsZYiOCWjT2uFqwBmsX9wKFC0YPdeaLCOvC
A//C4GYV7DjGOiBUxwRlx/HOWolG/zXTb01LpxEPXcNbLHoNoI+7Ofw7ZQUjTgfOxR9uh1wisNko
O6BjjdnLaw+EZi8BqZKWVBibnW5UolNWeUnp7T96+E/zqqXcDeRcv9FmEyHfXt9g6VUudwd47Sxk
o9Rr+aDXWspmSmFAkvxmoOPkbpS1LP07cHmovq0cVI1UjlcglDvVTH6fxI9i5EV+S44CXdNH6qVa
6CQYacCvbr9htdSK9Vqr0uQpCdPkeIsaL6udtkfiCfW8taAoSOq1fnAUq+RBAlwPac2gVx5RsOvJ
Rtr4uxUCicmK81eIVwI6XF5uqOdsC1toHx3kYZCee8R4ZFsXbHtoYhTl2LNuZXpeAlXmJsw7txXS
4qWtwxb36k560Oxd3CPYGESdtHfFD8j2hecxbQBSbesYp2IlmRJTSEoZQx7mv3Q15EKa1wJ0jizJ
qIYBUh9cvmz5iNaqdmCIQeumr76slm/pGlivC8dUq1xoVFGQs/NRMaGCVt+S8ptV+r7T830HlUK9
EFilvtwbkMBXmlRajxvg7A+HJ9JOZmLFKPYatibriubTLYunzMrH4jQHQK7HBRjatLLmiBy3w3nb
MGBpocygAAPH+ujxV6GoEXUqXMuMSKST8mLJbvY/drpIiFAgeX8w2XGlZZjno1JeCavnRDbRPGSU
dXXx40NogtTfVjf5J8LJryOCdjuexK+38NyeXo4kXNs5zwhPRC86yRkgNn4J1JXlp41L5xs18hbL
lV88RouRbuStg8meJAUgyiHvsPAEAS0iJObqDYPWxBi+/vIsJg9nL/GpW4F062n1gU8IhTGR3TLS
JGUxCNa1Sz7MhJbgJzLgIyF7OZ3k33hAUL5MdjFSffO9GisXE3FhI3o9XiX1lZ2L5wVR7RI5DHPZ
Jh1t9oikEPeu2sTGmNbr+J0SbhqHXu7ojDejreXIkmAj8VrTE9tTuwyBjrRm/XAE8wv05XSHRDP/
QkQFpL0PrT3DlLz2U18d7NY7jNaSjDCV/rN9sjVbE7UyWw5+9XDfFXnlHzswuhSuFbXOKbE0J0Gp
PcJqEAkkJpnRffspo+5cWZ6/GvkDUmVXCTwjRFW+iex9sS/2PWHVPa3VYnPS1dQzLOjqgTflQeMH
IG+hs2gKVb0QpDOWOG5XjJRY3j4fD0pyUg6aeg4Zx1FxDcMZpoVSrzDOaB8R4OfwQmcwtBUIt5rK
VBFZmjUiQUROQrktyfssd4cD9Kl/JBegC/zfSaiz+UGdvonAv4V939tH3eyV+GH468I8y/toYGqc
rM8lQxvlEW2y6ckDOLglsgCd3x7opxJN5uR1dlzdZhzAKlS8nStA2iIi7akiKYp/6zOjL3DP+cOl
HHNgyt8+nne/+/1SBABDqsrZBFBDTxhOHDjZlOMZWFJ2pivtnhbKSYr8fXWeb9/2IpFxREqeQKOE
6AdYZ1pggGoz5N4hLw4CQh0ClPBwmAjVJPDc/pB8B5L3Er/bVvwc4p68uj6tm/CIGF5URJXoRVWD
NIiCtX/Gz/Acs1yD1uOv+opYgy/UhmETuZl60MEk+RQLytXZkDj0nZ5ZsSGIJRwaRJP2I9NStF5p
ctV5M8zi9d+Gq1xZ2UunKDA73p6qsIh8T0DD1VC6k8BludKbgoa8eRJOLbCodw9nz1uDgJ9F1c8p
z9oJp+t8L4hZcqC6+s2UV7RNQIBeBmL9AugdyV8lIJ4iWUk9dSjSR/xHfJiw8a3cktCHvTeTpYFx
gCMRIEJgCochYkGma9NKwFMlViaQE8iYfJgyvrRLfxG4tc4j0/5ux3oROLPYn1OQv5ukUKUBoPt2
KWA6qdBYcjUIGMwam8V6ewC5XPMPd/ElQICAth74fXa7NIwhitJa7HbmsHOqKtq5Rpbg7g+IVl3o
f8ZsH48/Tdb1rmmzsoIVJttRA0wr45USisPX4Skp5i8CXXJTXhdhm/ANMpnx5kSohxWRRTqwSnWI
Wt/vDs3fQmfrYvwmxItwoUdlSw37ZfpKH1MZnnWbknkrPK2ZT750uqtnHjiq6J9mhI1LGskEftqN
Yjwedq/fv2OTJnDwYO9KYvr4L7q9Iz3KYH/hWZcvurW5B2uCVh+GmP8s7JXFJoQMNECya2KXfaOB
DNgaXcUFYX+KL5HEu9nM/bIDHBne/5sICFpttHnfcuV6GJ05vw7cHNkaMgyxKFjf6f98vtG37Ftj
5UkVaCpOsJC+J7u5W85AkN7w+B1hILn6zXbQjtS5J+RpMTMFdy8FmpOlC3fx+imji/yZzIqgPNbc
LXON189UTXeaUB26nncoXsoyVgORl69LqoHDwS+nZNTU3SrzrGWfiJ+UH1+Y9hfayr3Z38aNnpfT
QrgFw+XoVG2KwA8vvzzGdoMaMMp0jlOFEg7sdbOzdChw+4Tgjdl7kwVKL3yLETuRbrSw2mkR2pWr
Ov0tx3fkBeROCfCYGC6Vhkccw//BxopWOT77YYpST7Wu1ZUJc81RG9IvUpc1iorbTkXBSlt9PKsw
d+VGw3JMzV7/DsLTNNpyKS1T9p6+kKySZAI9QYY47ZpjIUJVtjA92fb1Cowk35EfgYM6OiJBdoiN
+zNhBk7pHltZjakLpCPxFOR9KVqlV0fwWXDPVVwobVsmJtOiLGBNXIVCqkt9C/TTeDluZKVmmqsV
KUu8JH2LPoSw5rHrznXEaS67xg6Hza20aCN8g1M9FbCWi3D+WqLwXHi1eFfTECVzFguqIl1LRFP2
ZhJPszUL6OS5wHMBziBOVJh2D9VzhTAEQzSClTBDg3Z27IH/L8s8cT063n1N1B7zgcZ3sZxOE82+
adB7KiOmKiXR+q7L2OdZH1lHw1Ec7WxH2cdL1vo4ND4QohFUYNxjGyvE15HFnwb5SP27bXdHQkL8
z8zcn/614iR/9khe+e4KyHKomdkj3nPTYtzMbjaaAqgr0kTZpOEiKcuF5srbmWoiAG4AQMWUW4R/
Gaepblrs2bnlo8A5OtSl6r9QZLscYYwFQ8k2dahKMAl/Rh8rbYHSP2awcEqkOg9ObFan1KqZ3BsU
diOzbEbnRRdxPhGxVptZ6rpLrWjzKLLdtvQo7gvbfOTBaI4KAR+DyGWOgcVmnWJtiF9XCJ6pgLFS
lfeWn9DRpxGoeCszZJDCABynCrRzOYmaXezLNYQe1r2I/YnFJ7uxbvahiLr3EufGWwKWGY4Gy5vM
zv20h1GWsiEFhHenkCkCLGd6QpE9/8NVK5TlUfZGaABixUYSfqZ1s0BSCRFCL4Ts1tW9UODoBwIR
se0RRyIXtIf6Jbe4pVa95UvxjqK8KNJCukght3gz4mD8E01g7Wlp/+HMtCCGYsR3/TpyBF3f/qk0
9rZoZ7z1aeRHER8rFR4aaP+3lIjnhQtMEo3IpjqE8CbXPc8zKiiN4NREfQgAl+1zC5u3Bfh2Z2FD
l2qHh0uBmGs3xXtowk52Dgy9/27fWPiD3R2lpOMSJBXgHecR1DEqz+iDLwPc60mld6qPVPmrAaIt
dXPrDod3cxRuuvRnotsv0rUbUDOJOasn8Lc5v4E0xmMPXZDJniq92aaTyYxJwQarqcYWTtZlArfh
gs4z+gqUiK8otG7Fcn81/QGoByXghHjIWqwj2O5xwRX1xx5Jteowem3wVdoInUedkt4JW6UibTHP
BWnXnfI1ICAUnOC0xPCGVhTJsNQd8B7htrFXyQVbbN16LYOTkoJLTm26ED3m7elVZkVtUJaSqVlV
WfwTgeZao+RXs/4b6YAhxFw3LufGiSVfHhqsRVz/3YwqOFnKckpAaULKhPeLd1CyO+H61q7O4tzX
loP+GMhasA+v6dH5c3tmDtlnbOH+U+CcHNXs858oD1WDpuv4FKBjJKAcPTiMi/jtXY99rFK1InPK
v7byX3JbBc3bGgmumOexSbMBcbHgqPTMc7dZ70IZOdHQFkSMBP9/B6XClgQ1KXCnIk/ptkc78Yby
Q/gaIozbOqmubLiUE5kp147WyDWVUJI4XjpHLjYs3AvGop1JTY1MDQ61p0ZN3xMFAkwfxG9Nyzep
peiXbU14nPj7AhguG7JXyN6jAQ/oaJdLJyWMNLI848DFHrbdKeFDkzMPq8ty/uihHfYYTviX38dC
IENT1nmbkRdpWgBDsENDdPMH9BjjmB1xOBVr4JMT3f9xCNdC0iXyXKHceHRL0am6X0BaQQNHAUPT
WkGxoqeW/NnhdnwXfDg6yWiwZik4A2gPeY1oD6z1lPzsz+sFpwQf0prpO2TVexBKGydES4BgNfyw
dmyLsHKAzbZkfzANIcC9qf0JQKsy6EOaELrH3FTm4AIDgChFiUc4bM2226Ml4c9DWsaVdeFH5ZAs
IIQ8nxom5kYvDpdS1C7Rg5Xe0Tlce4QUULmk/FhKAyf3lc5Vboss1tMgXyQeYwDeiQUE+K9bQcO+
58zaX/7c68PBmvcQv0BYikBuzEho8vaCuRU4zvpBAnl6mXd4afyPM+YszgGJh1OpqS+X8p5LERiA
Xw3NGMhkZvG+oov1vrfhXBG4CzEYpVPiVNoVZea4zrVQM6XgXZH9nluii14qpmrjGA+GzBkUpNxX
/9+DqEMBDscUWFoQkPGW1UfiZ+OnqPMPQNrh2QXqYJPVebIlYGOQjK4bKDYc1aFj2EOeKI1WHumh
VD+c+5zlOLMkfJRCyns6vxfw6Rypkx5clWhD6fyda68FHSOK9PuH71qwhUrqowl2beqUnMaHYpHV
UqjxC+GxNzzbY5wgva5CNO/bSINWZAxfHdzgWwczZixtfizqb2CRhXe51fNm3kLkUC1ihtlpvIZ+
OUxM0b34hK/EBzs/UDHv7of6VP/D5urbzD7TWFC2TqTngcJNEY1PwY82NdpAY98FJ3Kij/2TxVvU
z4igKGyolg7bLPdB2Lf9L8K3E/BgBn3TZ0/0eSUCkO8goBWOH/ecGZcuj8AUBxdZOA9tt0dWteCX
0ha0TXqd47MwAeSRo/+sHHCtyqw4Q1j9nDhSHBh0uSdvLO9Aw4r0jEOhkNGbAcsbZ6sCCFiYxdc8
JWeJDlcDw4PGCqS7sHTXRZ2pRs8jv3LmpciwxMQDyZ1edhcHDs5LunSj9zv6AmBbAt6YQG6giEJj
/dmSs/XwTHbOd8LIwYW2XloQT5AfSDwCV/uvip59W8MoLlw9Q8KT7SRnNx72mEMpgGVBEE9Dbsrs
XQKy98Oz3YElx9hAQNYj8C+MH27LoG6F3W2ecLni9KYxut82wHtlTi4itYNfudZeUvWR6utQ5C+U
cQJIndMWKaODXGKhCZlDFLT3btzkZ7EEq9NoMtoPdiJY53tkxbctKgNGsbhvr09vAhxonMxr1H2r
R+tOcl33peb5vvSI9UBI1aqipDQcznPtXojFrYc18VsbZ+35t6KF7lOlpj0zbouHN/l0wFtTlnBc
gMRRRGJbYDdXMFUgmM+RjRge7Xy0eeuF8c4BTGB3qi7RwTG6zjgyJ6yTv9/aK/i2A8Asi/AFhLHI
KSLXVaLr8igd5rvtov5L/9Ty2eOdeWitet+7phtG3uHTN3B3LT7zOC+vvkui1JXCaaplwa49tzK3
RgVrMlXA5cpWSN67lqDV8PGpvHoUcIkIgMO1oy2hzfy7I1GwTk18oJ08k2cEVSomBIwEgMvnuqO5
3HzXCQ+7ntl8uaabOwtKn/QwlZKFselxnF4kMIvfZegWjLGBCe0D34glrSk5p02ep40m2n9FkSXm
fpZQ4H7iROA1TF6bxcuLPsrlfQEEhNCgfA3h2Hw9Jq729z61W5Q1KFYlrcU9rSFF2ZcwevzChq63
mrgpZBlYvB3LW0T83y0jhk83Ev/GhVgSAaGmHmfW3aeS+b0ZV3it2cq7oTo0vW4FkaDIx2ifytt8
avTu8yT0vbuu0+gymEO0tgNm09pRRNc/ejkQ2IvnD22lKeS+Jvj0n1ZYcTMgyBVGwc7KhDqYEQr2
MeXGm7uelCujSp1i0ypHonXr+o3PiJv5j0TXnohHoVYDqRCkz5RDR02fHxSyKxxhjE3OTsmWsrKv
nCjuUnJWuMdPpuECygX4PiJvdIcixhIxfE0hhhZYz6829KzqLoyCHabJbrUglRsvsvNkmuXs+7Ml
ECP6QCknxUxqpalY6+Nq8ecGHB5fcUGWBa65WI2izMFJv+4eugS5zU6Hab/h+PaITPQGzN7uGN8W
To0gH8ciNdLFzljrF44Pv6iZcXXG6Iz+HVFC8Mo9MvfLK62uQKvDrynrpVBArxVlswYAqX0idrCv
YyOArRDa7GuK5tnGRD2dSO1I98HUqCVElApbgiXiuqEsUTwtmkdyH/JPNbaJjKSPDc1c9ukHm21V
6BhstDkfSAtyoH/DqVbsIgdGwsdKeKt/JSF1sE7Zk777H4lPHDC+JBhyFdcdX/eZFOmTDvjOuBpS
jbPkloe9hESTG2YFSh2fwpkgNIW6QVPFoAY3DdhTfa2PCQ+uIqkJELt5MLAjLJahioztmCu01I2q
GQgqevQCERL2toBhKTWepbo740VoHI4zagrxuQp3mHkDtC+iYvTHZZUyQ/LZuRWlg9xuK7bKB4Ba
ewIr0sZKMgiWXDvP7R69vgQY12HMD05z9BlD7Eempj0/KA+VNitllor9QGIiUfCt/zMPfdi6PUJU
z4E6n6X6z5eBAlGhA0+1/LhqFf8FhCpPSbYgH3d+oZ1YMPIC0l4lHhtzob4rK1elEHuIrehjBhWM
d+72a5zOWpt7JVfJxbJnQUEQC7iEJqbJuZra3ict98TnUNQ7M1H5D/rw3xRHwk7lX7HcR6FL5GUm
mHlLbGI3GJMaayKJLQy8SCScZt5WIkj5JQ9YHKcrKvRH5dAnXI+Lv9kjL4D6JHtGRVBco9EUAvxl
tagbVT+8gEfaBJZUaD0jmVUkRh3Unx+AP4tgs74D81Bfckdk21sIV91IUm3JGOrXzlSY60H977Ba
CgNWfbA+AGtt/mTB8vX0sOLOz6CpROmmA43Uh12ZwmJjKQ9JCM+NZlNcssG7R8g7ERTJwHKJ3+z4
rVWJhniBUcM73C+JYDbtWa3+5OEtfNuU/S0GkNeTrEVWIUZ/92vo90BHJGRB7C4e1NGKYrSBkKmz
J6MS56ofvZM9oUzf6UhhbVi3O/7qc37gLwiqNoyYt13NyZIsVyyvQSDaBuX5ea56eSFhzM8PJJot
xjp92pAMjx6OLV73Q8LJogheKgcy9blSWfaMOw+l4oyD4G0PhrXcwz1fqpehbrk9gy5skh5PkIvw
Yj/MeSEXxdJxLcynjWT6PVm3fBadaZmfv8vPsQefP9mzGvHnQiIZV79jmFukGoj37PG1+Gy5awFw
ZmS1UI2Ws5Nnz03o8YIcXhOvkifeuKtxSR09v9PL2yUk6r2o/vfWylrCmMr3EcvTzwRxYPlb5+ZP
K1/wlFLXMYoME5tp0nNUIgJr/8O4HA4lo/6h5NV7cE5j1k7dizY0Li7eLVkm1PqgaAVR40ZdVMC3
qc6dWfQ5Npi1zOdyRMeTTMkVMmyO8SkHi3obAfYbAC7rEE3jc0zKkMCH14YCGXMPnlreHmtFYjlM
3ihCs9OHscXVWYfvxkR41MhnUlSWbOhGatrtDAl++nZls+uRZRWnyY130ZR3CSPN0XLLezNJ3FyD
TMDbux0uZYENJ3klz0+pSTMiQgsNxZYYchA6fN1pNh6+R43ZwZIOsG/aDZSvptkTg4+4DyEbuSaR
1U+qHaYoBvkpNH8qnSiUfLwk28rZh8sE7ejWupqQXEJ7bJ1JnoY2Ak+nPi+TKkq/Off6ghjJZBC1
fQsBg6tzBJah4o9LyEvCAFZDePrmxgZNLruwvCUcG3RwoUAmMO2GXJEmMhEi5TDL/HmM76dzofc8
0Id9aPNI2V87o9Qfp0km/6TX5hc5j8DX5psliYzgPGPvKYHNk7NdYsVdB8AJwbpMES0/muJvkGKR
ky0rRaIBdpmOjuGYI8Iacbz80tRI2nDKpsKGIE9mUYf+o9nRVPlsVrUwvkJgHKqMjhRNBuG0AYlW
Y3HuiLOSd6Je6cL+xaORccK63d3M1uxUCYfjS1vbhvOkhiQt/tTRrImktz+75h+54VJ8kB361c1M
f3QQTJeu6NMI1U75739nXaC1+zVjGAOdnFzWypnxPoK0Nh7auB5ma+Nso7hu1Dq0HUF124Ze6NLX
bwNYHnmGXpzoM7E2zLvpOAus04O0tmHmZcVwtjEEUuXfIylgLnwS8ho55idFkFBUTMJ8Y92039ZH
6tkDyRvbOf/Asi8SsTTrqRZqLLFAHGwqyzEdvqJarV+XyuMiQPXGjJRSEAO9fySWLkoo7kjf0b7c
nXZjazlxmwAMJAGb9f6UsBdQ2TfENls1y55cnypkl/82u/8x47ipKzUv7EAoBylhljs/VZ3BJbWe
sFwlIxA5ypqrRJBHMJlozTY/49nOO17DTKHxX/LSBRPsj9Pg/1LTrfZ+C24sfD2Q/zHiN204pz+0
kvwEn5YEO3zKakkbW96WlmrDoYyfFe2SZtHeO/BrmgPntdffPkMjRAAymBgEX3gC4aFNCl9mpCwY
PzGxCVZCJpDo/8eaC/SDfZdpPSAa+O6TlXdF3gSmgQCjATF6sfI15buLHbI/QfDKdtKsG3x417Zi
1szlJH7lAqxZF17NMBPIrFrt2MhfHGFZH48A9GF+QKN03GeU2x5MqTAXSvoIBnVzzUDBproG65UR
GlvY2MCjcXMXl/yLTcDMqneXNCGrZgHA+IPgulenqkSHo1U7+Hgr+iFezNo3fLOMdCHy+Pbn/6d8
5Y6dunB+jXJytVMRV4DAcI0gXc4LapampMhxj5YOn6sOJIm2L7RcYkAjlI7yPOvn8Pa9VxD1kbPn
nzat7wGl/gW0vUzoC8rGxZ0ImzuniQCtDZjtS0VEYrPl8ejeP5FgUjdAaqdNKwMtfgwEGPukn9oE
zb4RLf0n2ao4+/gmJc6Pmw2APtAUKahuS5LX1QzlAbWJP30Yw9g8WDa9vSPnsvjat1wuJ3+62RDT
GXremlZEzJR7ccVTjA+cbzhf2TRdojk35WqG1ewIxEtdVmedNlR/9AAD8X6YknnXi5IRabAXz+rU
Vce8aB86a2cc61vu8WOvXetCOr6cNWP5bozLWUWqSFVEHBSQUQUtSyb7ZmPzXBEgEjsQrn0jRL0P
Nz8JRqnW9Mp2utEQ8Xm7bymH4h5YZ58pz9feO2Z0EFWlcUfmXuC8mcdPT1Uf/WO3uNFxnyIqQqvC
3vKmpZ5TvwHWyKNjyG6+Nzj+DHjzM11Qz2r70rH7/7CNaefZzkPt3WG5i5n0MkE5EAlWa6BS3xhM
svmAT0lA0kz0AoChv9P347cLXb6gffMrgZC9ZpLAXsD3E1aSCmnx9aRt04Vc9AJxwBns+0T8cIWm
6W23HXmDxjRxXh4EFs0ie/6sK9OLQrc7nEWR17AL/ZdgrhshZ4oKCUYAMugLQurKSGVIk/a0WHRI
elWAvq4Fz3rjh8jnQqjOwt4rYDnn58OvIFRnlOeKm7kp3+tt7pAhWx2rBiApHsipJPyTEeuGaNNk
a4IeUVPPmRsVfdue+72dj5enhL17u3AI5tYpuqWrZPs7TsGKpTtPX48UYZ08UTFuUealN6QK4VZc
LBL2RYfF5jC6Pp6n8t8hd5+2dCsLCaHGawgRea7O0M/ucg+22AO266y7Qpa3l2Zv2pjpAqu2Wm8A
hymphLq3GNcHe74WNqoe+xUSqXLTJrG4NS7qKqldZNrCVukLSfHyjpi2bO3Y4tjHIkO0XJ0KcDOd
OXCCw/hsrJR9gBeIyuEJeZ1wWoEdLwJSB/d9/sPsmDhd4DW+9cD40zVIgHMg+yust8sn6Rmv14YM
C9nxUSj1pM7dXn/bOXYODHK5eJb5gYN7InCx+IHTk79VkAJ7XpF3ApY5MNNMgpS85aM+zjlJ4qh+
Q1zjjwUubnQONYs8O1JPM6n8korO7qfzm1f/6rD9aDnZhwzxsRfo7Zt/xDhoVOKj91r4DJL4HLxC
Z17KfM/Dx46yPFsKLTLIgNdO10lmo0xxCMZXgnSrdiSn2IDhgWPDdMS9G60chu1/NH/5tLkE65Q5
uIIJO/5MSKh7kEqaF6gHo+9kWPDki6Zh/59fsBXksWJf64KvIytwud8hq7+dlnf7aaI3fb4T756X
2mmHXD+3jim60xP7kVEiGhZN8jIW8RW6ZmcemYiVI11i1RbJXMsS6wcU4V0tvx87IOVrZz+uv3u+
XWn0IOqk3msT8rgIZ1TcGeeV0VVGAY3bdieM45MSkpPMYZZnaC8zH2q3/ZDiQLInG5E/9qfM6UYc
sj3WtwYBiHtDRUlcEIYu9zFqVazZv9eUVGI4D4cIs5/4Y3TSw1Urpo3c4yNK40aX23/guAOaDEII
IrfERMUCUgNigFNt+HtTbGPGTK9/2LU4qkGzGWmgCgxvBvHS5V7RhVmRkwCriqAJRCVwNYsbPHfu
Nas3SmjgvaHaVH9q3PDsZpkgATyDfaemP1vjiRFmNVZMied7ERc6afILE9zd1rQpw15kiA5JLmq7
RiHuOlnqIVoRhzZd6ZW8/D8tMjOyzywpL2kRNXU9Yv0TrPCnaNQBUGjBwUnhfs55KlXyZi15Kssk
KkRzDrj3bUI/QRnv6//CQYNex/DOd86FdF5TmcIwNW+c17/fKe5/R3aQnt7uD7rjNHPTVrleq9Xo
lQ8JsId03K3rW0DmuTZgEi1apd4/medz3upNX4fIFXxAEuRnB9IiSQqItSBpqgbaoeSiUfxp6TWl
2nZamxuAIlrhmyZ/3SWtpYO6bsdc02tqAIp5ekhkFC6ecYqDfEfRDVcKGYLEY78zBWylgZUW2OF+
jRUQbsgorD7SAkBRT4kEIGfEF+c5lfE4RnV27SJ93ClWbSKGc9suL2ffbZOveP+0qmUlyos1aTt1
+pzjKstT0zo8iZlsqWk2ZZAfG24mR613juBBKxm0ds2Zvs4voERyZSMo356xq7mruTXWMOuB4KKo
vkiExJnllRPa/qnltFspnil/N8m/s8hW2d3VktPLeyv7HI2PSkqfqQDXohlgNF2rFH7w0XxYCklZ
UhAGAXCrzAj1sG0d//MwYtNn7T9VJgM3HEvuMB06cgVxMBeAIqb7eP+kZPvKUwCGzQSbWnE40DmJ
3JyYnmjCvJ6N7eD8HdKubt6FezQxz1pu/dF6ckfU5HZwfR3vUtAEPmQrWMtccxoD0jsyZX01P57W
KdVyIQgcPLy5CHZPpGr+JicH2E8JQMPRSQPUcR3/ILRlWGbMRkHL8351+54+tKvrlysN6Pcu05IO
M82o6rSBiUsU0D9gOPysBMlgrB3oYD4nD+0cw6Wev/cHEZcpYztwWt1pDOfWVqtLJxMRCFw9Rxhu
k5AcHz277DKFo2bZ8s2HXkkQJR1Uv52hQ6nCqoDvPJB0DlPlmAqHY3eSBQ0rZVBlfzLzQpDPNtkH
J92k/vpZ7daC9kgn6oSLoFl7oK57Ef7cP320zynor40jHpG4eL4d9NyjRc8UAyHtel5ngcSICZ3j
2bgMUS63two1nGsU85UH+W7+rsFUyJlwJ1WL52fJY9s211ofcow5b94vL9XfWlsxcTxLEcAmlkzZ
EWz43Q+jUWoSpeP61mItidVMFQeli7r4FcnkFyIl7Lwhb2xilM/MFBNtpMJoEdN0pOQjByjG9hW+
YJr3UYueGzwjCeDC3Ojt/SPApHp1/Pp8rrzRcjqI2rrtBljwyzeK0S+gXX11xCXj1doXOjGUchrU
MfMh+SzA1q3dx5K6wCIb16sKg9mj2jTBC7jLET7nu07Ed/iJIWfS4lXKDXmU1D0Tbx2BPjw1Dr/K
ib6rGXE8Q/mtBxbsps9MvchJT13hBibHSDRCYCZFRL6EHrj3erTYo4LCTFKKmLIAduXLdioGvwil
Jryk0qU2VyKzKO8c/CQi/LrxoNSKVq+FbuXBfSgtsGOFnBzSbgbnxIQMY2yK7so2novCOOrYu7+W
K1jaW1nPp+FWzSht5SzkXiRCllWAUy5NeQMFTBij5VHRvfjQKQopvAA6OnQGFK48hI4xa1v9EEtK
faRW+3aZ/ph+x94sJGEFXiygnhMtDMoAQi+yQpXw9DOT5VzJ0Pj5MN/yqB1VU3ZVS+CZj8T8cKgD
7qUS4MWKV6ePtDxT9L23gGta0cSReKjSbc9JQOi8vuNKLUSMoMT0VFaH7rbhnbRUV5g3WH94akj8
7mHr2jjQR+Vmw+x9AaAoLQ3fEAjr/pHKB/9labJzzeBXhj8x2Iyk5rg4VXYHPq/fMymoKTz1baXg
dtc5mgKai6rzS7ftzMYLealxkZf7WCQKKhhcTs43r+IIJcR9lkwno2C84QIfPfVs7XciYGsUF064
ysiK/UfjOnvZfT+LLCnWwh5CIja9IeGAS687fAPEZD7i5tn9R46eoEYIga/smHXGFV1l3hLB44vm
Rvr0sU7aEJpzfhYammoL2o1cxrkzSWqmdQ4rNjbmi+cx1BHfKkKUgDUc++vbhZ5Aeu8i3ISETj3C
v0tjT3Ba36IUFMoDA8HYBasBOimERZtD8QfxqP6+V1tOW8Emo6Oryr2FJWA++AiGOuz0/Iu6YLn9
tbAP3VGy7bCXsgs8yDsa/azwe00o8kqjfJV08LdIRseBI85/MoohN0kYBvrP4zRnjplfmdADTLUR
IT/tnjioSS7U49ptY0eyGIP6Pu7aDVJ5G6GhkjDatM9WREkgG63n9lITLK8j8cpuSvg/+L5y/WKA
k+g53xLpULk/XvyE+JM/aZNN1Bug5m9dzACbJM2o3fbBU+BTPizAoUSZ2aW3GsDRivy60fStmAPH
zVyPcPoP70khLIUHyXNcmFQFjXdK46qOtqzJGpq+sIs8DJNVBxurnhkuTu+ugpl79VM2cz6YIpjr
2DLfraSnQH/WDrURj6niDw8/mUxBGUFX6lg+bNevOFCIVhzuaIih5DObw5izwmEZDULEMhY6FJrS
2W2xgza1IRYFwVvqNTXNdFrUEMZ/gHlctCR/q318iZlLzZc2k2sM5/L40OGr8YplKMlKDeIUPVPy
gEyZqdi/kGuZul6WhS40SgIRi+QmwIdE5S1nanOBZiy90jmaTCdrTLvDbH5knqJYC4yPWF1trZIW
oDsdCpvOwkkX0wx9MqMojOfnwD76b6nsl+K7C7lDRBbQn+iwuzraLIm2Kg5+wi0SzaWTP6YKSIi2
fXzODaCX6d0fe+P6eaoWwNH75+7/ppdKkeSQSArNegt8gqodmvKh/TzEDTSqfj1GkeVBG4TCK/hx
wUKpw5Ut9O8520OYI5qLfYjjMkwwCYr6BR1uqv2SxO1Zf2OSfq2ThWWvba4gLMO66DjDmCQZ5MGW
EZ299eWvnAZQfCUGmwXPM2Uit7U26d/2lZKFknfhokOUYMLPO+jZcBurper6ae7nQs5JmLO5mO4+
2ud9Be0zWDhezBJRdk+Ea+99GBioCGba+H8rIy4tgUMXvYigELnWHjNmMj//U4qu6A6C6k8/UTo+
z7Kx0MV7bQmEohM47c76gVbkXQMz7vwMvUKNAQQ5k+lsBuhdWUBW20k4QnKMkF+cN3t1G/pmGANU
o90pVYKQ1d1JRVmxyxjLshS7Bx2tWuWpJAhpsrut/39ELUtlylskgHCnNmB3SuBCA2aP89EcFe59
G4ANisVjUrTiq908z/fwOWAFkGyvCipbuBs8e/sovBy+OAN5wgRvc72CUkW1ezRhrAi9teHMr6X3
pTo9Wa3Y8+mviWPi95sa+rhEJdTqOge+oyP4gKTD9O7r/PQQIiTV3TM4tpnNBEpT83Hx/Ab+4TDF
RxfDb/uCaMrL8YyEuXvjOB3aoyk9TcOkAb/Zv+4I2safFS+YX5fAPx8ojit9me01/EWgrlemSidm
7/x30qgR+3G5uncT+Ld9sqRJHSG4gAAdBW2NeTSTOyHI82YRvrHH5cUg2g1GgKNV4kohe0Fv50Fg
7KfKtaqlfYEU6pxY7UnEvMd2LgCT4zsRm38+QY+GWj34Gwg+a/P3dpt0wLhhZ9vzsJ6iBvJ4P4HN
0uNylnvG0RbN22qL4kZdyG4RU0q9gboNUnQzqU/ve8UYY/4AtrKmIYxSzIQqyZ+xNMxiC1RQ31og
pOl35/Wco52vdGIlJprokHMXomxCRYJc7+/iCe80Qgi7UnBfEN5IALMTa5TUVtug7X2wzTeW8VBo
BQ/GulwW9tB7b7cJUDG2L2PLu62NsSshp7C6EptliY9PM51GAGeXQWRfsUqt8FYrl+WPVPLsSjyQ
ggLgzjzRCpVdR2YlOw7nnjlrJbbquuCqJ8gVFK8yPCQFi9ngYcXPqi0b754uE8cacZuf+XElGwrS
GV/7O8UEN/GFhiR5UqdnmHbkwfBu63Wo9S6EvF7ifc9bW8l/7/rNdLkv3X9YJIRgtS7dRyyWfObn
WGMYtmNZuJCPahUrvullkgoVz9q2X8XX82t5bTqiv1Wfn2hqAFf3VWwjUWxesCT2tkkChUfFHfxh
vCzM3lfQyCNN1k8/YEs/uBi+GwT2K0X7S30hgbDpTTdciWMKmWrnLEVXubkb7DiDyocod26ulbmU
vXkXbFLUQYApq5foFHF45ltjDhJyDoMdQL7MnuIUYS/Ue7dqD7PY1VQs061AhJYmQuIRyYu7TmDl
6Ldm741ptOgsU8h/SZ6JjQO2/0pd6Z6PFzDwn7Nhz8OwSv9rAZzv5aMcZz1431eBPNbvkklbvPEx
o2rSm7RUGlMfMGqE3kS+92GSRb94uI7ovqtf3Tyt/3VNXkydJosuiONW97ChEGB7SkxeK1QL+Mhj
hAgPPMmci4h8A/16KbVy1BttQs3qx3jB/wUZubFsIdscnF/3q3j0YCiTnVZRJLCFN1+rbSKeDAJv
09ckdDFomsY3gHatknYev06Z6I00u45VSQZYQl/B7DeSyATxbK/h+RXRtmo9ttTHfEmQtR/8VspW
FggGXGYOWzAewAsCRltvtp/Sn7ogS/PAlY89VyDCS9ajBd5K4A2ZZ/ot8Vy+EhgGHq0ciczE/IzW
t1DAImBu4ice7VHbmUPzh6B40P3glwaZxQQbjoMqi3vdSzofMiK5UemSP4eQ2UjWeHvt+z6AC8q3
GI59tp6d7kXU1AOaJjHWaILQ5bPFGkNEX7Faoxd0sQ9oXeHk/j1tG1JJaeH9vKiljji2yhG4ErKD
BcrulZJxjaPie9rmGY0ls08r2nY7Z7OyRiuvLUndaWmVVzteFCcvzvmjEmbL22Rsj/Vkoq56C+pB
weau0DcuEwjCbmR9PyiCN9JDedwkA5Hok+wso+0zQ5DWCmMWPXQOHk4fiEWDZM8r8anbphq6CdCF
SG6vwa3/srtod1cBXSHQ+4pZ0zUKc2tIfGrgA4RXTkHBidhGz9cEeoUUYXMoa3kz/Tj8Bae/667+
whQMQiOXTI5/+1b+n/Gl/y+KGjMvXzN0ngl2H3NvayXVkWH6w3JkoIWjrfZsDxiMTjvjwDf1te57
F/JHGs8Rv2nfZVRtIHAJhvaORmmFJnhcLuM8Mp8uB6l+0u5yMZDbQY0NvmIK3BsOuVN6NqJTDoru
LW+VwCsvBDGGcGsf62zQLDwISvC2jFCVf3fQT7OayFpgrRbqqLl6C0H1/TTQc2HWNpVzIietsjYn
LdS+okqsNOScFyVPKIqxiGIebs9IeoN70AN39NGibSv4f3TnMiE1sj6h9oC+TLrY2/PWgbVzR8Kt
2MjA07UmhdAsS7VHXfR9MhGC52y5qlHR4iBDH2115DB2T9WirPwDGaMt/WlnSQ2WWEyxQtEoPdgr
3oxXB2MAEkSaiLCrQRnGTL1ICyFkwvWfjdITsTnmMIj14m5NIIFHqXMl2EQrYU79hYFf9UxenpRV
sgVD4zX0l2tFOuR4ugS4c5KL9bBPtWdY7S8H3L5whYCWkkcTYKS2dYyg59tV5+RzggLwBbcABYdF
/D+DBk5gK6sYpRgRk/05ws2jCO72uRMr7u5R5Nihn7TsvLx7jDk1N0jacfdipCX554QTCiuiruP5
ct2N8F/JLwRaDgno1Mitz7Lu1JxC1I6pxP9HIGF20Tao3mxV8AqQR08/90/aiLO7Dv0399fFDPCr
S/Z8qhGXHIkSpMQr5BnHLdnOZ60/BLpQRa8j/q5IQTXMFCL3qtK5FNc6p93VtZ2XMBfOaIHo8PDV
abpETEUagHlSBglVKNIPREG1e9xhNJs8UhRz0iWeru3yAic6hMkKHGsJKF40mnj+AkuJuY2PkkqJ
FVwISFZWIp3etaytIeOj9ZfiM+LxCoyETX4SckcZ/HY2jcK3nQp/PBxXCyAKbhrdDiEb/VjuStu8
vDC3opNoxrDyZ6K+RHgDbp6o2YcoO1EkI6yClwcaViNbELRyknpIHDT2H3uZdmPznFlFjstG2gwo
qbFcP0G3sjifWPvH8/rpd9WtvHyUbGWvRhQuqmC4yHf4dfbumoMDSkshhcm7zl0dzdpbyoQ7jxdf
oLJgwzXDjMXQ/6Z7tAYxl7z6qbC/NYDFs8xX4xXVQH3RpFFrq/NWZ9pCmSik3YFRIBRQxMW+utDx
+LN7yqyNEy3qYDVrc0Gf5u40mWHMDiLDyuOGunhBJdsc7pXucKbku4tVBr03CXzLHOgUjALAUle0
7Rs7Kv4SBO5dDTxMV5NTXQ3N3W2OlonMPIVO3B3+I8Oo7sgac5l2QALKnMlYy4P2+R5nVLTN3Zl+
tQN7crCl81Sx6vKdt4dLudBMjySCSLW28u9x1lj2CkmYuMP5KpJOu2qmiNeJulHXmu+m3Sg62TJG
lqgjUjKC+BcjoFmoVRF4MKEgfEvuKaTILzPuBKVnfnqpmqnhWG5N1fiseKPswrZq1oWgEGbT8iip
wNs0nxuDiW7LbN1ZchtT+N2JVs42RT8mK8HBx/EPd3+3MKXeKbLI+Q6wB6x4zuunSyHlstF2WF6Q
4F1Ytqv0oCWXBbcamm0DcKbkDIvLj4EH2lXPkZc5hHt8RTaT9wydhEuAyE/xPFJ/icWRNtpI4OLq
t3yrIs2j+V3XRRaREKA4MLWhImMHKAeemA1CcMRWDNkH77+dRft96ghv7eX294bTOG4O+se+dGjW
LESL/71ekjdzbgqCCcP3dGdrb1Ldug7G3WnnWmvvmi+LuVJGy8KGM7fMx8j2b11ZWOPXy/rZrZRw
CKuCSbciFseJb6bvcy/KDJFWWN26Kica+kDuucPCtL+N3yb2angRGiDXkbRUTMfTB9775oSN2z5c
bo133mPGzB4L1smpuHZcFI4BrzP0ABCPvfud8k5oSh6i0MqoGGMbs3V130Q5hAFfM5ZrCsGRtN1w
VOsKqRsqNwQOlxfy9vvjZtOCzJhB1tVnYMmLcseZpyGl4CCVMIADJ0PAlmP/RqT1etABU2NPv3VW
CXCsnLcyRf5v/dVByurtMDpBuZzosm+iSUDApZHEkrsABXXaj7XANHaw5oRKQpV/2IxTlZ/uShnM
VSopL1FgQ09Ge4Km29ZD6rJt56F4MuZRaLND37ZPxbDwjI45E6VhXMWe/FsBS76M8XLOJ/cO4EJV
mPMDXrzpNOHQT5AaloAUFidgNtgXNzWORIODQ82RWVTtAzKX7ZsYodVwcb0TRtCc3CCS6ppPve4M
lJYuGrlPCHwGUJJbu5Yqj9FP2ko9qghNSs6q0haaiG4w3Jrgz5qSD7gk4HdYaswGKQQeJ0hceGhh
l7hvGviFD96U933ANiJA/Kr88j+OrN8L4HK5flrnelFrtGJFt39xCPMBaHI8afq/81T/MtoWKWUb
A3ZAQlgqLuU06+JpLTUY3jIj1tvWDQxpTvThB20G0MVGhX6MTphbXyT87xL2kJjHbkSBUVfgqxof
J6a6ZJTjZKOCMPlc1/QqmgU28Q4yUKKEyTns6CXtxdsEtTZCIqn/Car/X09PXn0vII6AlBSVkOPC
2UU8Sa8jsjPqrU5e8LPdI99XL/1HyI2V7/3arEWThe6M11HZJI0nTd28ASPTz8LYo6qareEGXDLu
xZWTQhTcLbyFJdeM6Yu+lV7v6BOePo9wkqnoKYlXpuxfRiliXROeZmwH1j0Me2hZF7SU6D4c0DgT
NrKerxCeFdcpvrPArTUyW9Q0UPIQ3ARXKIsJ7hoKQNpnizGryWg7WrjOVDQmldXLGnTAyg3wnQDr
XyMO23zDrWCIqX7cCsvXOC5hAk+qyU7uEw1eNZ9B9UaolWuLk96P/PZwolpxKhYyUXasPKMdJTzk
ooDIGsVWsqS6uI+ZpByWq3GWsf0Yge+EeNwX4LpSXgRWOQY3jbCKEGLuDHh6O5tqpORj+wbD8EMm
POKlSZNB9BY/Mv0ex5ddcPjnorhslZTVCiK0Ez1sgnDb+6Y2XI1+aEDgoTfhNqMaQoN37Sv1ynpy
ajiWKFR8WIkdHqn/iI0KaRtCTbxlqXLAmP5vUHFZbUxZREyg0ucm564kV5tv09NTDA/Ah/x7s/mp
sR1KE6KEFpbNrtCw7WFNjtW/ShukzTUwsrmK7ZZBW0qXXB5xBe/I2PPCR2sYwKKvutytMW9/9hQW
FwUxD1Kny1JtO3qPk5CQvrgIfPY0Ep9f3ycajJDrQ7LNWjfpLx4liOS5St765IrFZuYQI3PisLKl
qX+epfus0lkRm2FqUI8N6FWhgbQuWjRuKBEaTC/Ux3jdsp15gaLzP4fs9wVShkIN+9+pm5Pse0TG
qT34KQ3ygcIjFOrYPnLYRo0tVhE7bx9koA+0E358BWohEByQKNpP22O06CYdQXNQ7NIIUgiGtzNE
u+KNMRLUr+oRoqX1gVyhLBtL+heFUVzPLBsyD3lkFEC3clV8jycAHzO9P9GaSJDw116FGYfvitbn
ZyulfWO9b8y/oyhIr2fo2aHjBFYZK59mlAKLjnsEHwBDw7tw2pfO0sqP0NlhMpQT+sG8vjscrwhA
Ht2dIq/fsXc1YTftcI2TRoejoqlcs7zsgq9/uvTAyx3+gGk3+5wX5IMKKHpv2X915R9FpsQ6t/9f
xnR5M8lf1TFkUqe9xU4LYyeAjBicxl13OFA7KMoVhCZ5EKd6tkB9KeU8SDPJzU21uShLdTFuMXjn
Z+WbVPK86OnC+HBqtk4gajinQKYkleq/V0uYjb8Z62XDcxcNAW8AyiG+ik73TT3XEU6BYj2LStRk
h+/yeollwQxVVGc9y61bg39ohtUcmFacKq5AqTEpuk3WP80XaJ8MP/igwbt9NYCYcCbKdfbmC909
ccirl1pLKlY+rh/perdoX10IdUNOLwDxneodw0mmrjArnpU23Oa6X6GCnh3ESEqFrPy+sR9LHsSV
dnYf1tw6hXlAj6y8YICsm43BguD2KSHV3nxLj6gtAPsDTCwi//BGOjKtp2fW1zi2gfe+W+eCR1CN
jVC400GxZLwnPaxqyO9NVUdVKZq8nvT25p/xZNgS/N4/+wNQXhHZvseqCcPFRys6kcRz+jGUr6fx
fZPS9gDXE7Se1xsbLC88UhJDfnZak17SpGKF35BW9MmJjzqewZB62ic6/81x6BYuOhMUykk7Jk+H
E7IGjGhEzNaSAjNZh2OXwmr4igQHlqyqaQq584Awdk4izjYSNMJHQxcG+f4oN+3NUz1aZD2r/klQ
TUx+cTm5FNz1jvUOXk4foWqUyINF/gHU6sSYoux3q9kSLPa0qZMpn4iGVPPRJsVYvH3GrOWfHhrN
4bwTJD0fRGfedqB7o7A33A4O7Zo/aHfgzte1NNwrZk2CySl2d98oM75PUqhg/R6fVotW6LxN8H6V
4QZh+xQZSR3f+SpsMy1DE3sCAzL+I6kXSgfY77k2j2Iq9yA/qUKpDZfgsbN37KXT3TnUhMypZBjd
JZQe5LVZUADQd0RpJzUfKtMA9Mg4gvjhaMPIsTF3+a24ZJNJvjth+vrAs5N/IpZTVZHYTgEfmiH1
FwLhlqnv1fJ/D1zektnLbid3DadTTKEza9Vwa2juPvdsnLVyEYGUj5YilHMPeb519CcrqasL5k+A
NEXD19ZG4Hp/U5KPgd1jScToXunvTWHSGoh0LL1hksbLGFKGyCcKcC+nMX9VM2t9dkthNYg40eZH
jCvSt5vjAKc8kpKME9G7c4COxuKZkdjnvLrW2/gR9H2UTi7HXujWJJdMZW9mINWLYhz/gQwoR27S
vgqtmTTvic8gPB2eVvcZkxltTjs8WRZJnW9sJJ1W6fBpj4/uVE1amNe+fxLgww8gdxnLOSZumjVL
2ck76k5SfhxE42do8pT0HFN/gFuqBNu/rb9RxaBnRBLnhAjSdIoNUvLxu1nScsRON266oSBYM6PE
e01jHX4KJVnp+GphGnoxEX3wAIfQt6rGuwxScwRz3wLRNJNzXgOXD1/PjanNd2f1jWQAuyggb314
q5kgE4oHhtJ77IPxS9xxCH4Og0ZwxWkMJYR4CrTXRAxjYHKM4n403XWMHjS3tL/BD6BTOl/UJSuh
uvZAdknL28iUWFKs1HGqhoSl8KlLG03zmcKeWGZerv51RxsRv/XX2tQ20pF1a3Zc44wKBDgJVTrH
Eobc4MeBo7VWy9TkzHpPdwn9ieZMF5gy3uDfPGizpOThavDK6rMNTwJaCNo87chTnQJEMECn2QdJ
0Aqy3sVRYodL92Co3vFitfrOfFW17cag6rvVtyEkW7Fca7DBPpzCuKxXqAL4bu/SrEQEXjVApM7q
f5CdWNOBD4C+fn7rrI1fn0KkL0YZQsfG5eFke2Y21Xh9EXYgYXUFndmhFGB2Yq//pDuVm3UZkyaQ
T3Wsu7Kctj7PjKehpg7EfFE5VfJwjuQkBVt+NMgsZvrChGfAmMkLsISLBGfJQGZkArYCraoZZham
ZkM3q0yK/bE18LIUEW6BHVL6/1L0PoQpAKhO2tk9QDLWC6gUV8BnOFhxTXupVZi2vZrgOxn3ObwQ
OqAShCnp3dRzTt9Tsm5/cRQLH/jiwOIUuVwtU/+IelPHI6BXrWOFZEpiLYUkwf8tjSJNOueeOOe4
Y/OfBP1ujUDZs5W13zHgSgRHhGxat6jng41unPhKtGjq8BGHpLh2ezwQi+L2KsULBLjdzmThWo2x
N0ntymt3RF5EdlbbJ8QBejNcJQDUHCnl6m4Qkj0v41tP0NLVkej72sf2G2MGNjIS3jaV9GodSGmk
i86pFw5mwCICN9E+w1ZYIjQ/o7QPF0q/bl0IWWknSrCrI6WGqeFvcbGgGKwNz8wDImtx8rwbV/Hd
BAqLCqd3F3oqjZHbCsllLRSc5cywwVXp5/ptf8ILVGoT6AgseXuBqftAu7qXW6u1KYgKHs+hnfiJ
ApmBm/1iCYYFX+2Fcm2KIuacPIvCL1LQVfcRUUs0zgiynE/4gSOi95Nym78lhqkpJXswZcafGCTL
sI/em1FnBCxfBu5/4xsppWb0vbb7gXOWN35PuwBhoqfP+csmDBD+hi0xIla6CjsUPgjDHGxZgVO7
9JmPl5D27v7BHWRvTQ++EXAeZ+1+Z6vPY5hSECFicMREwq8ZpeEXY+sRzZuGbubRIFTSiLlxj+NX
l0AKrWIaU1nNC1jPhp1iOdcnLYnD6c64mATEPGUCVTKoXUlhsXZIJaYbdAb/J9NCv24zbqhh8VQ8
vVxib/Dxhw3duKgX4x/P7OiGCYXoOxUPadihpalkGQoRI+4KAIb95njNM8JUsdg7juloyCHPG+o8
ohFqGj6ZJ8mIoxT96cBl+I2EKUUTqSCx8ajGWjd/GprIXvhA29uS6DMugxkFB4yZBy9BwWc0HvZl
xtOsYeyRH6DSZuRtNEjnFWFR2BYkoxK/PlosRiKAIrdEkk74BEvSfhIwX8HJ2YCuekBX1cV/cN5b
aFBFRKQ7J+hi/LZN2BBIV8cMgfq8QB8yTaKWd8Ngp+RWbxfCYMVio9jc1TR+/NUqu3NBPT2wswMM
0dglkQZsrHUlMc1LggwTwC4YPvNmHCVd9r7FJ8CWv8YlkwPmWRiyBcmJJLtx5j+OCoZ9xJ7C0kRS
sTOFXHvdhGtk05OMcPPH1eAcLLkOqBG5o4HH21LWkJdIxDrcAcznirPHt/LjaOWZVAeOQxWzCav1
/adcCq9c1mrM1q6Rh4iWvl9MTFSTjox/voq1nh83CbXeC6WZFXGgJ/7OLToW5qCUnvMJPdCifUY3
gd4nIqVi+49vqEA4wTlxMM2FIK9x1TkHpbsfmapu4Cv61Tv3o4ovG5Ps59UPDp+Nk02Sp35KKgcA
34vbTU/qxDq1w1GnSV3J2vJPIyFb5HBrK/6XJ3uoYoWyUxHkK0fIrNZggeQB72f7eOBkwcfAiG5a
EKFa5AvxtljqXtqZHTPPm+WnauK94mKJR45ssZfijxTFDG+ONumawc90WUCF2+AarfcEeTWRFfcN
Rb+WbBIICH7UMssOPZHcrKqkW67wraF7Vj31+Dv2GGEXrU93+vT/B0XS/xdntgkBSKvJ9VH4jqa2
kp1Gmy10bPaya7QmFeRAXeOjPj0nNDrlMtsEvDXY9ABMLwN8Z/ANuYEdSah5OQ5KN1vjQ3WAxned
3zHwtvWJIPM/APGTptKwWAp7M0leHD13WJItLOKwuDxVAJCRJzqNafEMzcCaRFgbJUgpk7QxHmgm
kNeuxwAhmaUPASgx/hwv6abFiKryuDcF8IWWkgxzqMenkOh7b/nN54saWjwiK92SIJ+57YkLRqEk
LNOEcdoqrvDFVfJMAmtcTaj+CuexZYu/s0GQo9iUNK52gM2nhSamO0McEbYo8JmhGmlPrwTV4asI
Wczwx5w2uOMg6dhM7ASfPPZfA1Uoi1v5yZMRYIVGFRmxjK+ILGcJU01Dgbq6hdKKjGU4qnvqKQMv
MOAh6g8dj/ac6h9sO0tPoNzOmUy7CUDWm5maepbcbA8gefsXRmf0kS86MXkbI70PiMPubJckvXkV
KPQOslpvxE+By550Qqj29xbWM8RDvTG1y2zFBh1idN77CUGcVFzRD3WfYksMeDVYKqyJTSZZQtb+
RfqSPjUptLRgLgKwx9j2g/HsPYHv1uUalyBbTsQFEdcirKJDbHyC2bWbkS9oNAEw8aaOe7ZLXwJL
aIoiueEPBCU/cnZ5nMMuOTgUhu9qEogSQC/CO5CBByOocq5QKmX6qBwt3JF2FHILP6NHxyY6aapY
w+4WrQXk+6/tnd9+JDrSatUKouR24nQ6xCog0AmzKMnso29y8ygI5ef/fT0o57f96CGJrkiwL2QA
PrMX+Upu/7leKYozwM2Xfd4lRCpGleXuhl9gVFcvXrbBYMmSX+Ap2f3x8WOcFrT5ZKWPjH7DqAit
OqqW4e/7VVPfyZMiKLOL0d365M+VTBbmlEQ7PeAJuSQtK5J2ujXJKkuzpoMAqgfOJKFTWq3xm6Fz
bj7RIzKGqPxK1f3bHjLiUM3Qq3Z4FSZgNMnnr14n1Le2/0MuyXjXVHhPPRtmF9pLyjWgAvi7BInO
kbRIBChsseGc/lsnGsjeKDqPJY7mcLWdHswxqfZwJPeke5Blednd0GMDuckzyMOoDkXpuasBKdBI
/95x38xiHjZIWV6biKvZZz+oxP832nC0glhoU0BXs1shANvJEY3+GuM4Wdei6QiUjdZO5EZesGES
HOq2SZGpHU7Xv0RU7es7xFVPwlcXZHftbiPYFz1kWyVwxmHoLEv41mRbh7Qp/8Du7FBAfi8bXYi/
g/z5vYdv1Y+t+VsUI807fz/EwsbKSGIhRbWjeLI3g1h68I0fPWVSkOh8HwpTUqJvlMQ9Yx/7Ks3B
3NYV/vKgfN3XD6cCOH/wyG6bs9uyHh+q6eHzjlAk4fstyRSx7NJZQy8ENzvbMEwBD4srese1w4rR
JWpMGbn5D+vvKqoZcDUP8M2VAtW+2tmZWappoS1Ty2mcqqKEOyD5LtKR8rRJUDiFE8IsTojxwKx9
kdjqqbiGGlMbONLEE2rwtJx6pgIzg/6aWS6CtaZE/WhTUU/6tPclfCGAKtg0Qq4ox7io+1QMLllS
FtLNxykQznzJOlAudxbsS5OUb/eGebRe9nAtLNHkStI6olZ9cxr6Hh3wJTHCwU6nG16e/LWTvJl9
kf8afnmxhxZNruxZqqxMpBpRHKZVyQlreq5wjYXjM587W2gb3VMUfRW7Hzzu7epucL6W516FQ8mL
7/OaZTMruxFFGOAUbbAVtmwyJc8WkByAkZR0NKQgV8fpJvjN4zzNLtzFGb+O0zMl1h2eS8jtEVsG
oPXWGjn7NNO9jO/ZR51R1CTt3AhkpwVYlO8FiU/NFk53cHfJRKRpl6vugKIlBXtMgOLOPq5cAz00
Xx//Nm4p/JGAKPyFVEodyARuvpVER7GhUYa1OSnOWZzL306RFrPvP10gQnTKvD+3VYvhDtpBHE/I
IqPlbnRNDhk7FGxH1qnBKDQOSQkP2ZqOLcKlOn8X+wQa6WN71lZn2q/WnTf5SSlBCQerrewugp0M
hauQGq3sGcB9MLT33asl4VccMh1JY5ApdYUN4YSHmavPUWmpl2pFgyfpjuBcWe6Ni+2ORmKE6C3y
qyon5UaxA1Pz3ezEnkNDV0rz6okvOVD8guhOPFayW2bP1m3YMXNtFvu0/FXa3wGlVBnfjqt0fomr
59CltrUU+9577GJ1/RgbjNn1TgtSMC0DFvQlkKt0OVfmURsYzXy2Futjmx9OnTod1Pk/f3vXp06v
B+lepf2+EgE8rSNNK+PSG0fF/7d9+pTIFrY1caIdMWIWHLSdcMZCx8XUWcv2HmRI05gjEJtnLejx
9n7CGpTUR/j3G4+2hxGmqmH0bOWS580t0A2SDa8yc5g5CoSkifpFspLHEm9zmXiL6svFer6+bFov
Jldm8vWTVRUFCVrjVCj7haIKCMtkZHWlD3o9jCo/25DIglB0uFUtQ1EKZ3wf/jlj5iR6pC8wx1Ho
mpmgh3jttw3AeqFZi4Xytnt3m49AmF/XscgLzKtnWHhVECGnVpkuisrFR4NEvs7M7LO53ItiD6oe
MpJ3QeA4wd409aQBpWBc94ClOf8ZlG05ARpCmHfGwGLBcRbDWMeN31nGS6tKcXYqv27BcEEpH7Xd
51eXJ0G3eqg8l4B2bd22DbivujZ8tfz7b0KQDzS6kyUJLnFYpV3fAEf7rJoC21nNypTmyZcZ1oZL
D8K6Fj40B+oq0r88rwrIa2jdCxY4/suo2OcYz8QLsyol26b8Em/Jo1QU82ZUYMosPASSoq0dEWiA
RYJNPSPn00FcjZEtfkOPANb9j8NBgSq6VNdh7L9/AD2G3vXkU74kpnV+1DSWiNwZ+ED3kjnXH5fu
l3mIIo2lNjD5RLbVQiRQJ+F6VOWDGj2QStJ+UzdnGSiw87I8ehCLu31ySa8xmR+ySNHROuFi4ExG
7N9lMqnHYeZfVpxJxbnnOn9cYXaLvx4WY9rGYpEI46oxrCMUpUUcpTP0XXM+i1cxUQ4N6vTgGAgT
kjh7kzjBMAqrM/u7PZRFjfb9lizStipqTcLutonNNDvRGWHph7oE/WWcQIIeOSOWNRtgbwtaDS6U
oJrVIYMZ0uOmbds1xR0GnH/G5mFRP8BRuiDefIqkAUQ7ugVWARbkjqtdrFBFCDOSDVP7pV8lO56v
gglildAiS9TnMVn4BSsP+hfIYUmEjW7qXzkpjbaWQrF1FpPl7Z3LsIIoHaTC+sL83Szbx8A6BREC
fQKDU18akocgofi1M+Za800lw9KlF3ndf2FFZwtelmCgulx0UjYMUAUMy30hIFyc8IwUOUJvYkzs
wYcUGCBtOf3uW1tRF9K6n+r3O8GZ/NaUl/nvSs6TtczvO1q1M9P3sT7M5jfz9+1PgnPEPAdXSeB7
FQFhFFBKgM0OVj+RDicr/m2j1iWvFNAQMNF1bEAYEBTwPZKfOYhsgxZyOwAdwAyNSLmY5k2mqS8Y
JgIgDBhJDWLEyWpfYM2QvgO2jiXBnZUT8qvvzhOBCCy3mAOIJ075E1/b91NezwMAn1dsCRMkMctq
y1CZS6hAVMsjmZ6gVfvjPf0Zz4sEwNSWSnmv4FWy4Zk+QS5Ppb5emEGOG5IWuLUCEcV1Pc0d6JFd
Dd9+ieZQ+7YrxhlsUqL0uiEr+KiVLgm4qfdIujSXy2yDroDwmX5YB0fWOrQLkJx2yRlT1CRZMLvo
Z6VOd6dWdp1PeQcNXKdChCHr0i5o5OcAaZvQWs+2fTaW82m+oBGSECDEyVNmJazY0Ix+0GCgsZ+j
mTnj+2MObXhElWzMbHfMFbCFc2F4kdnRCJEtoZL0jBmablwOXiW/s83zeGoYV67vS+fjRx/DpNnM
o+1Iyndey1bLc3l6dJRKil7INi6X6NS4KYyYYWwTlZjlGP9CMGJma9j9gKB+Qpk/vrf/BiS0zWQZ
G/XXMWdvQYmO7K9YVdpXOyK5lQTybV7BUi71FpCUdlXFNRUjzYG0gIw5G7+xwNlG+bUDA0Feyq+u
6Wwu8CEEJMssVVIAEejc81KZTr++OUyGU/ib1EXAEaOEacqRMQG1RGT+jGUDg+kGnM7ek2nGEIIt
S+uKlY9Ur0ZOwQHBWXi5Jj7SRzqnTw46E6CaE/cEusqnSloBUGNCTGEzEneLxrmZI8C4zuHH+f2X
/fIvEy3YS/fKSK3mfPo9uninZOEyTNyVyGOCkY0TdYQBrdEedgOtnIXTlI6NwrKLRQzFJDOXXzu2
XFTTZh8PfCboP3SGN5s9yvkc6HO5jj9ueKsOWz6DEWHnfVDXtsan4CkuG0/10TNw979kqsI4nhgO
SblyVxo2po0BDjYSH4ERAhvwHvhAp82ja50SvgefW069DDJI4KGjR5AROJlrYnFm63gN8UY1TfBv
Qv8RA7S/a3DODLiL9nADbliCJJgnHqv+rI2ryn6cMrulNq9MIe3IDsl+2X+bW/XD2aV94ohhHIIy
fG8bylYoJOYsVYFWaa6LrFnZLuw8P2Q5d3cuU/+n2J3fTV+XG6bTb5inxuVCIdniuUQk8ks5hWjW
P41BmAiohKfHK2c8NJ11nSxM4w3nmgqbh6+Rpp4aWLSC5X4LrSrwn7nUtaMHcao2hdlnYAqziXaq
/Xlzn7qsx3lKNZXeNtaiG1E/5O5EnGmGKYo3WXVWccHxhFQx2CEVNy0yb55jRjOb/wET8HlWzK+E
lIAJzMiyoa2O8RweJX97caWtCQhbKpe8GwLcaIHxRiHeBGYDW1k80tT51D3bC/3R3KuOqHkGI7AB
UX8vTQfOzgiSFzzRUCvixk7DYXMkvnF+5fKHAVo45dlaDU635VP8Di86YaKQ+5Sxws6V8AeCNW93
w14HFSav8hWYeQ/qcUJfgCscN8oeB8IXbpZHz7lpuZl/IiwdPMWJ/PbAN2uGryCLiI+zRebWomV1
sUlymZIsWl7UXQ9hjNkUz1P53jPJATztbQ5Ze0Imggk0/Q05Qhd0HkYdHMqh+l17U8P27+Wht29V
3RQpPJKlgC/kI56u63x1/JIHCizT6vO3WRRKn/XPm6pdJA33ZQXYDwQEZ9IDUmO4Yfg4WcUmZ9CU
4wALrRdQpcMbXAyBDGYw69T3hfTHzCKvTCpA3B40Uw2fZOcmGQrEl89V3BBKct+FjLGfWrBeurt/
2nIofE7JvKiCtiWrzuFlmPakmm/IgsnpOjfWaSoTqLTnyPK0HZzIuq297sMB6Uv74JWi8GB6emPX
kxQb5fZUYI+sh95RGrP8d3KKzV0ch1Laa5x0MTz7KOlnlgK8DFuEJcfnPzb9UbzvuS2cY0Yj7euw
0KVTq3XWsocRQyh2TrY+9L6k6F6qtWGPJ76hCOPCS/A3MwJr2q5HbtMVNZY3tBkYDynalL/IXoy4
bWrf5cvQc20HnEoxjlcO496O8DOKGf1UWK1J+zBFPJgT41e4EOF5Mp31CBQapgr2EP7II0/wNWA3
Af97QVeM5uBuxSYG6I7A0v0M2A3B/Wtuo3/v95PbvfMpLS8bKkObHG08CTN2CrmdJvdbg4ggRv9H
QpQXgQ/Vs6ogH+/J6fvZqNWgMw6AoEUEJLcc9OG348CRQ8p9SuBamC943MBSApENcxChqyZ3cWL+
W45Rz+Iqu0112u0rzh0GoLBPH0UamTOEMLL8epbK12HujbZQ+UbLKYlTX9ZfCL9fxs1Jkc7ShCAo
iahVeIJXrSrmXlLR/UHZXeQ6A1kHijjTHnyJ/GxMSymoZLZE3sG/U0x5D1Y+Q/PlGub6b3m8hIWT
l8fb1beq3eUlhwUv1uS2OytThssaMoX0sRci+uzkQLqPGxsqF8QKsGgxrZTzLJgiedt634FtDGb7
o0EYU8aPrVN1ON8pKkT1LV+35EaIxkAsoyVfHbo618BoQft/RMlNe4LOKl4QDycwgBrLmsaT9YS7
x0iZfkvv8lgx15Lb+QaiON+GtzMT2OSMjuTYDos+VXLP2W724+deEIK2n3ZK3gfOcDol/1d6W1n8
J+L5894KY8bguRmax9UQW7nkZ576X1ob6MaIaZbf4qYXMNO1kAjeOV7Vf1T+ASCqR3XMeKLaRo0K
Q6EC/88TWNFjNMeiYXQKdQHu/W6bEicAnsuyRj676K040n2PPC1G07c762ugzcdgqVJdXCjazuWy
6UZQRpc5tZK9IbZsNvztnUw9+EjFTilsjVbmLCLg+YlvWvNOqtthBDmonPE8SRyENUOqFBM6BStx
RA7O8D6y0WrOhF0QQRqFzehAyWsUm7MSbn7HvOhGl64CJzpQRmIIUjfI0dIwHa/B8sPjbmx8GGBU
IkKgBx+dc77CPJRmjhTUqUvvx5YqEmZhYjqt1F7WQ+cjgu7eiHHCXXHG/Z2gKmB+dPmhEh7Yf/t+
u5N4nEm+notx2VTr3LN5X0W1FbB4Y22dpyYi53eyv5fJ5CMYovyc7FgrFFsKOBTfleFwMF3PWqjA
NQ6/kM7JrBtvcm8idOF2/Gdaq8GrjVkR69u/VsrDIjn+YEwKsBJiN6XQpHqRINuu+dmjIMyGFoez
haHcQTT+EzOh+FBpYV61gXwfVMcAwUM7E9693jrc8icTjr0LafGqAxwXvcLThUrQHu4pqbNaKGUU
kjPjo/FcxIZErOBRuGujlHmK7LNle7v7n/qVCHV30f07zmp6IbBJz0wnZYJ3yEh+UFPYtlfztby6
8DHKMvpEmV1gKaVwiqJAOvLHyAiQ4ehcp7O/0bV1IuBDZV/XqZkdS7qzZF9M2/ib0O36zQr8hZsA
g/4bqJPvcCTO3bkCRAtOauc/FQ40QX5OpkM9WChIihFNg7K6PBTIx/UGYMpVjnYFVoBtJRTu7UwV
Yb6YLKFxmTfIqEYTT44oalBLhIg94d1b/iG8JVUf6J6XzveIFSk90QCQgcydFxADgSgEX9inn0fZ
B7z4w2vUkMXRcFzurt4NS3VoknFvctuW/ZhoiXT+MEXI0q5KWNWXyeJqcX+tqsW7LtL5az0raKu5
YlZmz4GVyuvRiWFsQ4A/zFA3kdZbNt3CLhz+AFxH0JJh6CfrTUeEempkFjP5gcGvMU3pWx9rLv2A
EFlwaBey7q0mpwMJO1+0lj93caSwc2s62V668yjnZR53KuZnQ1IDkVL1b+tUGq0EEKXFamES/6PY
crtbNlRHz9yqHmx6WP51OT0hu+uulWPF5e82xQ+GfFUjL4KH30mYLD1BJ6/gAzLJe70bZarwGG+o
3o3tcN9Zg74jIJckD3y7HjTiRfLugqWLoT0S/96+tCNF7IatWQ3srHpKFHCnjQmGQV2FuuKwekF1
bYDwEALtcZeFCEpdLnBc8GyiWbgORFAo/+SUoti7uB6tXuG1OqlqXPp8Pttc0zDiGCbAbBeKyS8j
RTGzHnPGsk3gwR1C2bFKpJUGFiWBDyVsrlQbJ6GvIqEOYQBm/nFD3ZT9AJUSWIXcRZp9cbP2tDOv
WvBCaU8veRYWlF6/GUrQj046JFLMBW+6jWBCPIdbSHwh/roeIpJuZcI214XqbWlyQFzIEmiGBzfg
f3tot9qxz6jC0L1REYCizp+ODm0bHpQPfR+wSGR5rVQusTevgXmeOmi9Tz5Yu44a4Vd/mpBeTc0n
Ova9Nqwwf2qJnqlUaXRx9e9zLvtdgJBljC1s0j0Na92kEDUs1yJIYVPhDCrEPRGqwVSN31Xdm+By
6J/UuVnyrvUpV3N5nUoi+pp4RDcTtdbH/y2d3iwXarlfjq/6s3SZRMo1LUXpIv/pyaz6XIAHxZm3
KJxCa3R32bQSuVkztE0DdQzidtJD2Bn8cURfc8VpxSrDSh3LFbk7j/domYTFdneF2lOTe/azSfwm
W2jzLv9BAOv0GrHNFEs6t8pZ95zbZSEkSXaTh5WP+knPc5zQOPmbFc3+54fLZAXq38MTlHmXZxkJ
ZqvYlXAqf+l0xqvcU22t0OKRQ/A/eb1SR/zyhHuUJ2kjfLBJ6LoLjzz23NVQ+rEDmeDy06wP5FU2
5re0dcXltdPHVdDn3Qg2kHF5uqxW83THzZziI8je3U91d8Vwi+GAJmYw7eL/fbnw01O2wn6rSMa3
HOIMh+n+08tL+3yx7tXjHEv5sTwZ2TLBiT004fZBP9vP1Fxar7j0OIpeybzFpe1NswOKhHPJ+rGS
Cr3nbo/bn+KzCNxNchVGoz+LsXYQRDMTqzLuHHXny2kKkj+NtzulaLSZVkwqdP3shOEiHvRxXxfI
FMYOOvvkEd51Xq8DE9ttrIAVFgQeIlsShhxhXnWZmQm0XORhG3TNDpUhH2JXCvomEwa1VHEM+oIG
7zWe0fXgOOaANMXCW2f9WwKjtPNr/ys/WNSwSlcdTPDxiHYSTF5zd48iGIv2j8BW9TUInfrkFTqd
f5/wr2VGhXgwxC23UqQfWCwAVQNNp+9dMrZaI7yDDWbtvqB8o9fSHVvicMNpZKx+hGwho3qfqNgp
Nu9sR5RYy0vmT7FjdXTFCARyx7GERwQRvYYm9RDvQvmGAwFjdurfPnEIqzlcth7VLOK+nbZWzEAg
norbf1gdI0VZ/U+RmyGdd7Whgj8JRvK5/nCrVH+lNa96JQOohpDDm0FXiCOYgrqca+vQEkslCA2G
G1eHCG2L+2aQq3VBKATLx81QXLHj5A3VuPXx7k5VW2pskGgjB9qdRZGL3SJcPH1bYUvtCSUxT3S1
Rqn8ct5dpqMUPhvPED3Vk/BT6MOEs1zYrcUWyVOUFHfnP8oPFW2HSK6Gd9F61wBKisCL+7k8SLpg
QV2/5UrRr6JfKy+AHQMbyIV5MIeTKxt7feufglLUCFAxZwypzmdIdf7szPT8XQrAldkUcGPHFCm5
9lBYGp82kSevoOQDlsnUx54FJL7v9ScWDzUhB4UZXTmYHuCEJaf5rbKbZCdJteBX5y3C1aZ+QDgi
CA8MdzY5J2djDgyTXxyudxkgRC73PxmhJe0SCpdJv/6DvkqlbOzQSnxBDq6eqDeIiHAsV7raPdI5
xePUETdcqNH/EZbmYlvO+/13o4qvXfyWQ6W0b4HTH4Bu0vTFnzE8ky6wdlBmOaHM4t1x3I9iCb1/
M1QI13dWuOArTl4k9n+r02DMDuaBlyLCtWX3tYHFaPdY3wNMQgaAzLs8+Ef2L/1UzLRy8l4F6Y3C
mxVlj/MCsnX2+Of1nQtwk+Jr6XdExBRHeK7kWA2C0krNII950E6uJKo3RIdENn443oci3/g7B6ub
qLzeWBvzIVwM2G414D9FK11bn+7DIyNwKZGpqrnIszesoUQmR4ZLtchitVosBuSLGMtnGDn15you
re81UaScGZvvsP6wSHAk1Kec8bBEJpF5l1qJw8HEcVtyuAdJWhMSY39eyNo+/LyAGza56ThlPpu0
9v1XR9sEiLnSgNjCfOlSB+zXWNIxT47qINeotqGKst9xQibFNNVL4ffzqvQul8723hPXooI/a1VV
0/4JWCqNK7P0sUTq86h0/3Zn90NiZQjKD7tHXXg2LuEsdm6E2mrYKTwnSJicT7IukBD6Me4vf2wk
gv/lOG7H2A72z+S2lMq5RMO2FTWTxUtMDvD1ymyO6xRSpCIyewy1TeY8Rj1b6nYpmV00/rPMq1qw
0mcOy4GgZBN5V6kWp+0YejhZbNyhBGHqCOZIsqQT8uyKpU2ZDiMMQFEF91Ec+UT6KezUN2AVY8Ex
see1UPvGQ1zZyQsct5k3OgkbhQJJXhkg/OLeYBbYhRtpk/c3INkXJOggMzWmnruIYrcYSSqdjysM
/imPDaoOd8IuwwQEp02f7YSnK7iI5IuSwygSzjL4SNloeVEACMctGLNrf4kaU+rOqmxXptxi4Ivv
4VSL2+2l3Isk3qZdofbR1ruT1odTV/JbcijuATGW3G2FFN/bl904koS3j881Rr0snCFW3zkw0NLm
U6MMecgjHJ20HP02+BUNw2IKeyqmDpeZwRzwD8IXKXaFm8Ft0hcP/d1ceVA5Lj3wxbL1hcmkoobT
pP/FymBWgyuY5/Q6CnI+6Z91NAG44M4a+KQC2qT7WoDxMxOMpa5zV4CGUpiQUeGkLdsCRwuYWVna
Sg3DSkrsenb12nYxRvukO+4f9xBuc6K/lti+gpj/BLqgyB9h5zhED24sINiT++D5Qs1TQA5XIv43
V5F5fTe4TkYukLYVMq2CSNBtLxzB1oE1GrgU0ot2cWqyY8BwQmpg46bccmRYLJzCV0qk00M1VApU
8ZTT2XBRNmouYWi5GMCoIcD061sc44jV0ahSDBfWoAp8aYsmEgM04VxvaRDgPjZtZFB4Y0LgclaK
H9eKOZAQ3Mj0LSish7VujRN2U/THBeLA/EUgZLhMBvxvvrexgUAqbVw5FwjgsoC1E/1wBtYH0vQN
Wbr5oGMg1+KGuUfS7Z+t66CHPgT/BVLWL40JgpUmA+b+6Ff8CrlRf/WxsdJ62vCsyj91EOg1XYs9
SCZ3n3P8wfEfZcsobt66zbsCY9fs+5jPoepvJARRJvRByl+o8KPgA3fhgQlwIiGOi0aF5dR9PUOy
ItxsfQaBNuRzCfCF40eQtihZfr5g/6DANI5vcumfnbmpFwVuC9RRVuqOJ/e8LUH9L0vh2kTxT8v3
ZQRONz4IVKM5pBON53l5lBELxSRQ5btpG/Qi9wAD8kEMlFBrPqqMuhVwIkOw96uxG5Yvqf5zr2lG
/d8Dj3LzVU4QfmNXLBtKYldZrA8HjrwgH3uBRIKa6P9ecSpgAaweZhZHuE7Devl2PM/jA0R68Kxi
n19I97RKmDFqCoN1KoIrTCKwFSa/OFvqCktbG6IzkYc6mtzIP8iZqvmRBrca0TAYXW2eueUkPmgB
+bPxN9J3GrdpOmx5+5XFqqYVCNn/X9hZ3CzrRQBX4vpFC0jFFRlf7DiOt/RKig/Y2q/sIImM+BUj
X5JuGJM1pXtfm20PALBFXdC1wXOB1ckTuC2jAlWO74pe4+nWXxeUAevH/cdtShJQQMpvCmqGESGC
T5k4NUdIriSv1w+d659CYhxcDawEuw7j0aQ2mDd8l1mkZBFUzhCeZOImN9Vd22V/fTO8YUku3es2
vsdgHjrwtbWaRkSh4/NSoOqVRyTQTZTQw5zXaRHcWngg9sjoUwb5fP19ghZBaMn37HpK/FoTk2E7
M3QcLmvz1k25ekYFszja1xNC/ifl6fW0rYI08BH8dyEoG9I+M2VJxfMscpJi8pZUQzt1VJ1n9nWW
bAUYg+1DQq2Y0CmvKJeeQPfkqs6A08GdW7UpGHHvJrWkwpt3IjcLw//qaVizKeGCT64QKRZ7jGx1
dhZKpZdCxwJCD8w0YIafeFE9uiNPKhhWhsvemOaZfr/yqpmYVa8TmozabwuDccrrAsmgy2Ivlthr
L/3YdsnXmDQlDkY22wSVkFOOeQxJ87F1fneM8MmB7/CpxlR3vyw6pnFO7Zr6paw5YIL8V1LTSY5W
1rjrXUlv7Y56nZzYOFrtV8b96EI+XppootutFuX0RiD+7UqV8jUgSQe8KIg3cHa5BQX1isgVFUyj
ZIu4KtsUJkXhrIAJHHN13g9iV1SMURAp8Gtj8FVscVckAeDnRAD/ukwuztAPaty+gS2ehS9lPr+V
6gk5CK0FzZWHXDmiJ+KNUo7qaFtJiAc1WproYdbxJgCHm2yiDH2zLI5Zqru2wFyRGofseln3RgSH
N7TnVSzJHALdZvLLf9m2bP5OF2yAdPIbLnl5QiqAsd4oSZQLDnLoX8EAtkun0HAyXQtWP9bElbP0
myEIaG4/tGq49zunv22zEjOFKxgToV+ACNPlwpB5d15wmz7GL1x3UaOfcRRh9zUXwigeORe/qJvJ
OzW7GvoHumpt5LEXEOhysOOsu/I8CXBmiTsvcB9lgQDglIyoc67mkJzYx8YuL+9O2e17rX1SBKI+
naApptpcTqjJoEUI32yk5OVJaOZEI5mO6GwVknNkje/joI88Z1zyj0le92sLVUbKW5jjR2EkKf7t
SVuJ1X27s7RB0DJaesCNCRa3flZedyOGFuJfPZy3aovyuGSvdn4oYP79OU4d7drgm7yas37bvbXc
J44qx3FCObgbh8PhEvTZtmOS+dQuJVkW9xCp+VtmtKSmJg8sAlKtADR8/o4GO083JdSgc4oumcXS
7vXnl6zhM9UM5szJ+Xh7LXDaVYh01qMP2+ToYN9JBKr9VsFHmV05BbrahCScTglwy97F02oWO2YY
zM0DatAuuYrnGqDk7I301T2nXJVToUEZ1LjCNI0gikZ6//Y0l0J0NiXmMC1T7iJGCEGOh81oW0Vn
Z7XfbrQ6U9pca1iRaYEk+ViM4wiykGD9IAAa2Nydwj/lJsH3zCAOGldnip8N/hIbdsfTYzWL7WwX
hB8UGXSsvCwUt1PuuJf/c44f2WXNb9C4jUKSVoBzJtpOtWwVGLUJ1yd/QZ5U4fUGraQO6uX5M2se
UvD+WyoeF5SGobf8w4M9OEI1V8dLfqtYDLlLKkccPNmmskZ6/INUrXUaW0IoNmrDvscrSYP8gaKk
LLL8e7FyQaFJJ8Ma1PhQu1a1szEhA+dpe1Q+eS6o4Gs8rBBWwJMurJs5/UXUXWgflNw3IM2dW3xh
dWOQ3BhYVnzDOOOjDl4whM1U0Lvb8YA4MRTnBYW8C0Qd9sL+lt7l3qclo+ZWRx4IVEEyUcJm354o
V7we1/1tNAW7Y5GKsmoHzvItgOLddK3kImICAiJk1K82Q9E9QzU13+t4DtY0dC99jizvMjIKnC1u
qPILNthnUcBUy44FUc/7r3LAyVIYLUMW5WRy0WbBJP7G1X+T+HMPn+uw8E/LAj5SjfmKO/uMP4Wl
RddM6Xr+83J+a9R0Fq+GIiC8D6VXCUkTFoFo2v+1lh6CXJsnKe9hvUxMgFhVOAH6gd0tdCHh3a1Y
MEy4W45FSbNudpL68nXFZJaoidq8DKuo1XvqsyxlwF8CM8/30sBWfuo+Vac3zIVEpzf8iOhg21RY
8fz6Y2P4wgh/FktfBB6jnxZxGWTIu37iKA1aesqKUnbewq+MKRTu5LlUFIUuQbLuwT4o3lxD3Pwo
Y/4INR+STOwgIyFSvh4A2AgYox12BvRRH2YJeztmg0F8ywBxPi1eaYZupPLwF5PQOMVrbiaWf+zM
Fms2WvlQgyIEbSo2P7LcYdT+Mz6iqyYjQzVAYyjtMUB9oyUlYDkDS0C1x7F3y7WJE7nn6//s9fJm
LYlEG/t/kLYKY3g2bTd8PmQY5iFUN2x/bt4B/viOFdf49czgpfncnvlX5qocwSuqkSXvdAPmm4xJ
yqnVe7PaQPgw3F+Toiym7T1t+in2c0SDC9b+ivtSVo1Yh/ZSfb6uOd9S5YzhXULWvsg20/Ip1rT0
9wCEG40CkTW71nxdddJRXQ8ZZmsFV/0keKR8nUsy2TsN1X4FF/w+UJfJIZGHSjiRqNnMVVxcfZBC
6oKmMwDsYfkSTjXBp8SxI7LahuhS1CoJGZk9+OXprStDMcfsnWEkWcg/z4doQmisFpZFqgFjTSZC
HeZ+SuQdRXgJ85GI256R3I5gFnQlS88ZHZ5/xxkpa3iw8alDx9Lf6hvXeXSfSuo3e9tzkPEi23/7
TIiuI+1Oj5xEiSbQJj0AK3U/TMo77YjR/RNLu0TqB1txeBkq9GoNajrqQDyFNqcEVU4n7Q3oGigJ
e26GLqtBhuEL8RRwnDZAqj04H+FAoD6BMoGJgdj2rJ1DCCT9wZMnlgusfaGOG5Dnx+FiRY0e0qCs
Ws9JTW9eDdbNYw9PmoBaN9wRyALCrM/J9E3OqP10oFeXv+fa9MWctEbyxNq7P2LTud15EIh8NNz9
NkYEEF86BdDSxkQZyVTjblP6XdEF4gSlR8OQUf0/Sl3jMncjZH/UbKyxYULRGcg73c2lhtHif2lk
jeGQoKxNdwvI8K9zV29rOsOBXUrNRMjZBrGIIabdNAL/4E9m42gGvP7mfZu5t5fJ1CGSvCXXpgHj
4gWVAqAyGzs/pXVLI58753eKHxerVGkCacivCzIRJ4EVudNfvMeU1I5iaaazvsvsoRJ4BSIngIjQ
1/Ka6BFQJ5JTvQ4qFMI3+PcDbJxIQEnK3/QyLSYxAyj400/k8kBcbTARHlmnFrhNglLoSqnZylbm
8pCnV1Hw2SO/1ufW0GCSNSj1fpHd3tGAa0mQUrIEdDPU8fStblHO4iZpG2F5t8yFN5d+BOQpRcFJ
lSw2+p08pfNKVgDcihiDso06WX2k9nf6gYaf1At+Wdv0RGfhX6P+QGFANfFqeTBacXq7guyK6GpM
4XMdoc3dto1U09kZrEnYnsG+D8gNPRqko4SP7Gybmo1kuTaWvxWoHTFfK3/k9cgjgnax098O9e0D
AtVWGtnHsEKUBGuq2UhPQPXSebPBdztgySt/8G4FjpeCxmBHvA9+UhyGOsyN7v0IjaqFvrzsu9G/
4yQZVxBlgza2VnUtWwgJ9e1Z42lztGuRbla4FtZB553mCw3pyFB4y4DomaevcCT1sjXWRAABjypo
orppossqEJV+eO66g26ri5JDB3DMpVGStmPOZyZ7aXkx8REn33X7AiBDqYI6oawp5rIT8h4h+kMR
Ny0UlGKc7NXlfB0Gj6qLShSR7VPtWzH3q2EP6QtZ3vI2hV8qzmGArgrX5YLZI+f6WSBke/AnLFop
WgFClMz2G2RZZKclvxcl8rHt7w399c0RTMYWjMEf07c/aCthMUTylFjWDWT5zHURKVOjLxzjxtqI
CcJrOn62dqbs/55HWHqBIXgCEsY+CLR5wkUMcJfd6gUAWTsH4Jyr9fHXMkqyDlL+9/tj57YHyi6h
2yb+2TZtEezG1SJTgpbMQgKgf98rOl43PFTPReqAoQ73ttShmYxJF2hmD2Hm44yyxA5dhGOt8T4U
frwuZXbRzxJDVcrtl/JiKBsv8dU4rTZe6YRV+UuzPu7VOyRMdGoe/+0GETl3jFVn/El74om/d+hm
6WyeEQkGEdSDGEXg/7kEAwKBIZVv6PxKLI2SwoRhHbh7SoBqeOVReGWP8mAsYSlb3OpfGFKN28za
3LjRU+beLH0Twsc+03Tj0y/oa9JZTCZhYLtfx6+Fy8entQeE67S8fVbcXsp81QquNe4WjvDyWc6B
qoWw+G0b7bAXfNppvqraUiPcArFJL9BGFnr+tJS4W5tKNsvmcNVbv+H3135pJIroTI9A+ytsO99a
G48XAkH5YEDjKXH+qFvxxpaPImQG7jQ3PjdT6hYedpZKyJoMSBFrUZ0u6xYP+On3DCVo5KLcsOqq
/vtjs9VL4sEmY/oxI5xERDGPg0Nk9yBg9z3M6/BKJhHPyFBeD3oL7IwD3ywmSowtTFpSQUgv5A7M
QGRVvaQJC03fvbCxT4aAP+eFiPinwwqo2sV+Lt6B8RM+RFYWkngKp68IcMR149+cu5nzQaX1k8P9
yaK+DlG53GXsNMe7xRyUBsbYoTp8/N4IqA/SrCEuHXvFNTFfTDqt8VIGIo0pC+EBhHLOSENVIOmw
s6aepnZSDVupx/60wnBwiDALdE1ZrYHgMspbsiYpfMx7abOctvuFT5cxW6jWUKc4YxXte++KeZ5U
QUoGlMI/gII5Uy8zUsihTKQtS2nD1SxsDDj1CPJ34rCTav/FVx+NBtc2Oczebo8mtaYM/J4IDmqU
e3CfBio41pcioI2WTN8LOMcFZVd6le6VHLC4n8N+B3zKasQvuQZahJSIKt6IxPzL8DByEAOpi+il
fvbp2GeiAWqJCt/8BxeQdQdpECrmtpfdbMNk1dJ6QpPnBvXpxa3MSaiBiKmHqzONlx53DEKLcUoh
63GDquFxq2JezRjKrc+3xB/akIlpu/4GiiEsyn4ZGd5IHzfQ8JFiddvkppz+M6zAxzZp7v2yl2ze
VcZ2C3HbJbsh9OTWnvvl8rSOOZiQvz4SOw6k/E/XMooa4PYs3vU5zohCMDeF3XuLBgK/2Lj9S2dX
e/cOoHktjypxZloLdTi9IQd4IX23vkdbh32qy6eannV78j79Pofa9PODQDbTvEDO4uFDxMLLfFlj
rTRiwnRX9XsyfO6VOfbNr0Yrdz2tVXDKvPIAqZzTldmK/vI/mrLbghS8teFa2hOb1jEMzkQjBwTF
DruZqgk3vYIjmYQ26ElHdDj9nWTnkpdaeJkV0rNyVGVxYkSnkmtIyX5WW4WsUh2q5Ko/cwOxW4rO
yuvE/0lOJ/lRj89ZvtC5mt9f91R4HLU2Jz9rtGtX0s95+OBmsnOfRGATTYJ9MxDGtCsFpTMqdlfj
4m5a/g24nIc5sQKAZvCPsYck2/l6YqKp+8G1s1YW6qEaZNEnRsxaeTMpuQPg83hjMNBtDswBA7uH
3wFSFuBd8//XXpUIDJZfygckDR82m8S5BcW2knxu4suOJj2AD03xiEb+hCARTJPU4croPQskSa1t
Ieh+kEQ0YrFkc5D3zfr1ix41bxiYYdgypGmWGqnrIz1iOvBZITMiMCbteMEXkBwm8b3zUDaJrsvP
2AP3w86/hl+Xso0K1Dc0fjjyvT1Ey3tnwA6Ld8nCchYFV2YWkn4ecYaxgqOjSywZ9rMmi/KKh4I8
X0rkthvuu1pDhkkWDnBLvdj+XWO8s1shA0a4N6W2DqC3fM1z4pISwPXbzhZomrRnVBEkY2PcE31b
JxxA64IuMx/nyJk8OXau4W46weBIVGMFoyuEljXls4JmVNhQD3mnlI6fAgsmSSE0YvGdNg0gciV9
zdA7FPkLGRB8Qsth88PDa/eh3uYqkSJ+bbhjUC59SpyOQidyPxjVarJdtUAopvnyrBhYbVZ4sPhQ
N2PmhM89Z22CxfsEgvhuWHFV/BBV7YjRNGJub2OuIjMCv+Ax0P42wiBXN8B4DKUyE/3/qKvUjABQ
uYKBSTv2Rdb3QW1GA7avaC208I7IRZHJMFW4syRQfN0DMfIxI4VDKt5ZfayUjjyUXRc8vr4zH9lu
a8tphPY0zyNeEQZKo7RaSU0U3BRY7Z6jEvZ1JfuaZ3BF7VnEHp49rSasdF4IJmBXjQwbjjx5Xc0V
7QSN5H5WToQXEVchpWQH5oHObYFeEtUBFfrJZ+Ga47lLgXUchEh4vyLLr6kDPuTy8+/kA3R9tA8i
YcATITG4iVMliXKKGD9aYpzRw8JkECs1OAAfzuru7vsj3DIJGApmIAxk/eRuz4OB/iMzUZhXYJjk
8PWJHG/8C7CLmICWGlwsj1I7XMyoKv6pb7vYId6zPgIVWC2mgtlyOxy2Y+ighC+5AQmsRUHD/CAO
sCEe3Omk02vRzB3Mamc1rdNKH8Cs86RZSdvo+7NK/RvbZFs2bZLG9/ZpV4RcQfuTKkTnrGP9roqU
Pv3kTGVSIij/PsvciiGX9Pq8OO3f4wyGjnbQPukc3p/ZmNMOK8+iEmjNJH/eezLzTsb4jA0Jk3tL
mT4QEXMi0hy17i5VoL9JPZ+Og6UrDHWYciR0NJ5yxRx17/IDR4kCfiGY/hVC7/RxjwAFxURZ5dwq
IjW7swdhQNy4rtkyEEmplpmenu8sLPIrUs0gqbZgYuGX2CZ3eS0CWkJKbOLyFtde0kNSsnVj+eTG
UewcmxlbpzYivBKHzJq5h38U/QffexzBp06QxoNFYz5PS6RQgRYqxu4wNdbpPwoVgmxz09Vnfw7h
azTa9LaafjIMB1vMNIj73Qe6CAphoH5+0NNhUNnyogbNiq+OK7Ln3Df7g4IurtWyo++DkHMSTEy5
Pnay8+jJyaJynkUiLtMKZF0axy/lo1QIruruRJ27x1cei41wj6jfkwPaKjC4y1YBv5TsoyGH1QTQ
TBe5CrH3khhoYkZNM3ctsDHNaThPHAh0e/6BMu2mBresdm5QkSutUbCeAPwV7S/kjzcDT/4XNF0Z
2Ea+HSgvj5mWyeapvj951I9YK3VPwL5FnH8m5fR3upG/IoOVwkeLno23Sw7BhsGIIKDZr4nqWTNX
50yPpIBKDDVZ4okklQ2gVZ46Qwmuiu391pDU7SvHBPGI1RWkzxsJXYa+lUO2tDGM7+RZtkMHx0MO
qDbsGAMVKi/6XDPAAQ3np18jsRyWlhSCNpZ07XWr+PSJd200DY20kCNyw/vGVBupoFMl5gF4ouZD
irj95pJHyLpt1rnxKyA3nAcr7uMTjePOH3VMpihaDs1nVahE4jJhcRjzn28sPo/tmi+TnlUz8zJK
u6BPkcWO9K277OvA/Ff9qEYd50bHZw8wYRzYSVv51NlHnYkcVhRsevj0dYm7QFZZwAf4/PEkA1kl
LewYTWw/QQix6O6wLGqUOd28P3jFe+fuf413xAXUPFPRY4zUY0oM8RTe/BNryCDj1bNnpnBSzpUg
38ge0+7xLGShF55DoVS5OHyI4PGVY9OpZrCJaMJ6COhF2MLn+UpdWSCSmM86crj5iRwj/dnDNIgC
+j3oed6MGyZgiwpjKUT5gp2KtfpVe+S1oenp7gIfpS4PoIfJDCP9pSZDByd95QV9zA3n5oGXk5cO
9JnzGaC0EF9An7oxZ9PPB6lXML8i/xN8VyS+lcDNT3aHdhHBSj04JNIjQP7HPlcyPo4i/vuSl0OL
zgecFJMWZbFzy0CWAkB3RSUqc0iQToWBRBFvKIlk+EFnQ+EzWHLSgVuFK36xvGwqDdpZ25L6R+kj
MiCzUf4Nqcb/5k3BTT1DP3Hn8HDV8cEtnh2FW/zFMJDIAbDF6Tjkp9LpqwVADhLR/pVEZ5CATHwn
MGERlB5efewfwYm6WAPbO++xMhzFZYcNAceRptG/tdg6+ciW8U7G8mevMHJgtScXxQnaRNO78qLk
bYiho8WyxVw/X6CfHS7gORHI0UGk042I4h5MMbdwAtROtRFKvzdA7/CC9Hj7O6L9Ujiuzt+CZ9cm
fZ5lf/IcoS9KKijfXGVidb/grQwYJAxImuwd/zQX6Hbq7xhKTnPpBqmHOOIt+DypebMoqGkkSvFj
R7aPzH+D2o24J+xrTZgqCibE2WCyfkRJGWi3p221caaWriVCm1WxutBCujbsAiP+en5U8hR7jsrn
JTzrbfxLba6mrajFTqWYrmuoA/2tt7G2XON9sy3LzPtKOTdYfFm7s5dqBCJU2ZMpFAP5A8AJ3QEW
RYHlVlef3fMEEjG6SReIQKoq2sTPuI9hRcGSOzlRWjkROtCz9EsRNjvsQl3w+DP7++FgOZJUmmcZ
LWaWB+IGNcuXORMMY281cdF3+is7Le1RpaRhKfHWjXVVvGQSr8+F8UWbW4ujN3s3tC+7dwvbluLd
aEaMDq7R6d5ZR++cXKMKUtmlHCIlBnBGJDrmwMNvWIXRDQf7pQGHnwDFfC5vmiTfFSGhvBzt+BlS
6/x4+rHelvoOsOnCRE80BMgyprYU36qnKoRKeXsj1s6zs99WIvgSy0QMgM0qK4fr1uRnrWX7W7jI
/hjQ3YvC2bDbJ8LHuz/XKattcB2RhWtDr7G1HX0r/anlbQQSvds1Ec7MtVQfUpaEMlevw3pqdT2q
3ywZwwd86eL4j7joKUHzC9Dj2hFgmPXN++AiEs/60SQ+4b6MpVyjqklvFyoUzW/atg56etmg9Pz5
OfBgRMKL56Eptw+F0BEAcg/KaTVsp8KKlFjI1RT+vkwcxJKX6IJrGT+JEjxobOmQ5yd7hyneUDRu
jEoIkEfiZITQgEOMXnHhW+hOaYuamNYrNuORiBQtP5FHYe3g/Hr+o87tGeBXwyrFnj5RZQwfXMUh
B9M/2+FodiQdLhakI0YBRbcEUFq6/K6apAoMwBw9kE19l8ddK2LcATupr1F3/RAy6YxWR4E/LPTl
ou3Hoce0MrE/ewbQs7Wp49z/VtzmBtLIvPEuIAcq1Hf7TPmyusaqhRn+MIJMaK73GSx/g2Iq1F0R
Y3cD34X2FF92kl7jOvJUTomhHNCWB6uQtD9/36+gb1WKbr2+zr8N6mqgysQ1vDOdBUY4bTeF7AQ7
xn0elm7KifnMRQmBYKB4REOMlpn7eU+H2XG+f9I7VTF/UKgezo3lGgFb1Q7StfUjxeFmMTqB80xX
MMmIE20ixdC2VsJdn7oDoGoHyzGxlv38SCleJt3V0WfNlP3JQfoPuFVjrfeG6ZyaKGY91tOvBCnl
2zEAdW0YuoBrHyixCo2dNJBFI/shy3oyVXLxMF+ZHuhUjA3HQc21JN4cZYDbGBf5RpSoIXukMMXg
lj1xIe0kQ6Xb9PkggxWxujTjgbfWr5z3fjm0ne0DxLPLVz/b8b71g63xgoCDU7IeieLZ0LTSIc/I
wMgjED5MA30m3HNRLaXOCRzkpH3sAL3grQ+ShEsZiVdJfpwsqmgJRkYBLp6qedGE7P7PzxtZYHSX
es0hDEk06EGfsCsKd/rzqANeJ6WHcBM+ktZtCZxOYkhhsMXt0d4psmnfUnlp4ytkhstq9zIc93+i
d9fEJxsCVhaSj9962Q9/2Aclr6nDAioj/hcmiDNK4/oLy+o1d5wtGQAJW4Ie7nAbIKlCsnAzaPGE
vFa3Q6Km0H0KCAFCM5/tz1tITJNIN2srCuwqaPxT6dRRaILIF5oa2++/9HgrnehWuu3sjYFrgCnU
VnVcHBmV7Vd25t9XShraNcE7U9SEFG00ddyzaRbXEkimQH6OBMa5PIwNTgztejmBNVEjOhleAxqc
Hlsd9qAEecTi9z6U5mruKrZGrZ6dwWg/Q/hijFePZk45pUCgQjpV6v4+5ru6DOMywTOFMe6ZnMJs
8uQqgXO8HSBmiCdYLgphoHdMdWj+PggBrMxc8nZYiQRdeIsoSv7OCwG7xi38qL1VLEsw6xueB7kJ
3C/xrxkDC+Npgo3fGVB1X8K9jX8xTGfhV7MS1Xin4K8zheT3lNqjkBMb5LgGVXG5/F+gMPGjW/Wm
4443hkVqYh/jw5vc6eYODwPhyd3nr2lC0Ucfwn5O5hwxARdYMjiPjkgH5TS+ophpKNODnpzh/FMg
JS9EgjCaWCb0Wh6MQSwaYpFi66UToLs5RLXgdUPYc+cnxAVR7HWtWHhJaVXZ6pL0uTEJEOAfcXsI
+s0EUXzRXnVfsDDMcBYJRLSgTbSRFm2zm6ipjfC44VmUXV3mBHGghZi+R9PTdzXs+QDaHrObZNRB
jGPvlG/ev4DlEtEgKIpDxHaSyqYACvWPLmw/tA5w7UFRdxOLYzeMXMETVSd6gPwETAIWBWzoB/Ev
d8J6Fz+708Rg7BKsG06XoCT7VpRbdT79K+dUQccAhTRSHk6gy48iEy5zjU21gMzlaj2DuCly/N/C
iE5C9LhQGSpVHowoU1NjM4L12xhHRroapwRUuENj+Br6pRExMLf2HiRZNfBkgxEVMiXlYOU4GXeZ
ZOgS/C6eB5Zu0zHP3k8o7NwZj/FQiV0iIVePuwlocQ5riejdMeFklMCmA07bYTkOXrQWDtAb2V4q
fBDRxopl4ui4JHVVYqnGbXKXHtSDuj2MUkjnNzLldB5hTg3vM0UnQ5JGFTZiJReVTz6/XrV41XA+
wXrR/3rFZ4tZ8Z5IYn3wuLU7g/88OeACpPNYxJ+1jOzKdYcE2AizOxVD1KQgvQCSWJqdSrLp9q3+
nI1q9g4T2h/cv6WcfqcPFohDg9jhhxlqwc5YRcOO3nTSlxaZUuht6kzWGC4oH7U2L2KFIFv/ljv0
lSJc5IcnTUEQonn5A8J2wlXA3OXCA3hYMvcYFC7Jo1+i/HkqF99BRzMi26IfxEyyQVbM0eS0LX6m
dIzM1Xk+Qhsm0FgqFKqxoKEmMJHdC0sbjsPjplw33BqdqC3tNAY6MHQlK/Nk8YRYZ/gaYg7jACq1
CgGEIVVFOo2crtiLKqhwGUxZwVm7hpJtK6g7OVPshvBZ1viogVDeItKQP+EITQxAM+PMlP63stR8
dkdkjaZ0xscDMM7xFb0JKy+dUhag2C+CunwpbvWJZpQrpaq9fHzO/ZwlX2Voz4n/UY8P3HlUf54N
ImhenFbgK73hRVRfIMAAnsqp5V7RzLNY21khCrhJesdCV9Gl8+OUpF5+l8e5tKZnSVAme0fjTscR
8FPnvfVXK7Yl8fomnO4BpPR4lcZ/BeoYux/HV2OKnem/MCmZ0Eo53mhR6b7Yvr2hkc74OrmgBkLh
nbE5x2XeZZ4KnbMY9t1IgfrI7SAF9r6WUPkQewS94sFJmfkx6Fe+uuXU/hxVzuskY+YlzW9SRB7f
5r2aQM91Gvo24X42RLYJdAc3DwJTM3Egv1xQRSvIqq0jiOlaokgnOORc8Zg80A/JvCFwLE5xhPnV
oIkkOJnEnvaI85i6XDFlNLz32gEl/ox5XCZWX9ul2KxehiJACStCkUWvimM45GuGRGCPLbBqNR/B
6CFCbauJBoo9d286WsdcYOTc2H/57v/94BOOWDmM6P6kczbBqIHAFIJIwhgdFkYdIvQ9PSHB21WG
0J18uyzB36SEvc8YsO08l1hCsu/6OJC2uRIyFUPtR+zi+MHrQk7+BcTrUGAB98bf+bP3Pu+fH7pW
tw5tgSIPymxUihxXWdpAR0clNJSHLnLjl8McN38VEavwFGoPubdyaGJK/67UGa+7pckSYQK1slm/
IoNtSZbwvTYG2ux6mM/3//QlMnDCctQ4AfZigoSPOP30EUSXj7U8x+2Km/bGRZNXgPIzz+08A5Q8
AdHbL5Zxa3wYpjNOxLukhvA3kXEaUGBvDhmwap7kKQmeBJpRHkmJ5cjjox1+KrRf8tV1dL3h4spD
8bivYM5OgYQxRBnhlt+y6qHqYRdLrPmCaVdugxyhfNAdBLxbaTIaA9vLWD229cKDjaITOVJFt/sR
+1CMWBljfYy6WOyD32j3kQnWtotZxwSA/J4f6qtdeYek2DBzhcbgW6fpW9alAlhHRQNmitJ3NkKY
LQH6b+RQIw9jkMzhUxSQnXviW9X7g95Av/xR9hwxUid0eLzQnZ1ESWx3RBh4JeCf2pGomrxR0dUS
ailDxeD13aaFoCn0iP/g1LFYBZjTb7jTZWrOdXClZaOlCQKczZgnmHqfY2yWRyfnmkyhLXsYH6zR
3/wNivoKvsJFSMS+8vzYYmoyCTlx4gzDgLrR3Bt7iBwGU1swDmkK8GCIiOGh02VtboOwCWyAVj3H
IGFSTiRNgpCwrag+Vi1PygRS8zY3OH1sebsL2eFUJVAGFpy5KCbHGeMJIjBN7AgLJ8QuBBeIXHpq
tvuihkQtv+zVLNC4WzeEeQos+TPDYuUBlfkWF16q7Easv50N09MwWYL1ACiMn8B81cOA5D1fMqDu
N9CGlgTG/pt3R0nTR6u6eO2jmT3MDvrrhIn4TMyXikOq6EPHJFKPwpyzStFAjjh6rnpN+3H22afT
SlbtTO0OAaW7gAV8aRpX0ZucCIOb+wDL4skvMeS4V3kI7e2kOIJnVrLZbmTIYKGRXjrNzJffl5za
+YJslcJDYGo+6RGahtZdTf7+c/tf9YhbIqsjbVyLj85dv+F2qQT2dAzW1S1ZOxcZdH6o9f+rrWO+
Kz1dFJsG/ZDR985tmEqfvREYxc7S17lQ+CaHtRGTXH6GvJRG0yl2/W4jlIat+0yWlmw6q+7gA0SU
JhJrGWgU04JGbol6AXwVRivt7x9HiWixFe87xUpZ97aPdFmxbGnCsa/WcbJzS0hrmqW35KrV1u1j
A8cKLGXVfXmThQC2vJ+Bdymm/YdLiJyL7ngUs/WnW94KFJTqW298k7wPYSqucalORSCkPOqFm/Bj
QjrUqqu5XbJThGBKLKKR983jghTDZgQD+fboyoEsvL6/UlMWAVGsQ0XFRmpkcePeBC+ny+NNs03F
FSDSVgXydeIJPbTGN9teeDrIV1jGpl22sHDmTXzDDhZMB27EolIJcvt8cRIPrVcxGkjE/BaCtVDD
z1PZRbdkBPL4WDPpIDNq7th+tUc9/tY2Jq3T6J4kfZp4ooMwx185/6DhSWx3tdWl6f5kxbQSdpyd
b1aI91HORN1zp8vY6RZOQBqaHXyz7051KS+LEVYKENshzPIQ5AcKwG9hauHqKn+3POEL99DjEjnd
PvMyYgC721hw6zrVH+DbksYSEb9Bw3JpbPTfEdqkr1r2V9wHfsIlRrHXLpDcHqyQF52Nt2IdZa7t
jcwl7t6qj2KfQELLPK04KriO5uxUWPJL5DTFYrRAS9nqPRzxer+mbSbvky3PXKtZyCR/gwxWREFp
VZKdFAof0/PJBQcsXoUlOyoPl/2cwppKd1tIlaoK5ruaiZ9DUMRPioDMbt1KznpfQ1jEXBC/fWJh
uc7x7wcdLzSxBh9mbq/DAIBT1Ir8bf5yUG5WS0+A+6tZXY/5twB1ZHVbAYsRC7qx6vAc88I45LSI
6wU7IRkR7RQb9z/ONjv1tbe1sfgNkkgIh94fBCr4L2QW0D2B0kOUMYMymLM9yU/+ka1jeCHafLJV
RW7qIvcFCuvHP9Gf4UAzSNWjftWFR8PeKgzgj8fl8dmB9ePG5kP1aNmjwJ9IgXhCFyn2Lku3SdqP
RDga00UEM8XANMT0bIzZCa6FEyjkrHVAU8QOFRc5bTRq9H2R8f9Ce/WX5WvVV7+tE7/P/G8hGwW1
smXknXohDjO0EEeFa7/FYjXgjZHrfAFpxf8B8kXGWGNcLVIDJ2CECWdkxc6rYuJy5hH3nb3osVf2
/m2ynWvSyj+kPHR+0G0f7M81TRHwn2Pma8zR4nvpwaj7S/J61bcg/UH4oqO6ABq0LwBqTRwWm+vC
FNy0RYGKUjj3kVAcTq0r2RGOKt/9h1s4TdrKDSI6z4Y6VwZDLQgkxjhpknt2j5D5XIh9JkA18vgn
TgorcxXyGxdk4RF+vPHDVDfOiMMvAnnWxwccEQFQ2dlegyG4wSYf0DtFeyREkMfxoF+9x6zrmON2
0zG987eDdZM0wJEj3UPKQmlDlEi4Y9s6xEZvSNn7k5SeWTsg+4jhGH3Y3V6834/5y2SZAMe7x0cR
E/IkveOplyWL6QNTOtoJ2L74tD78NHz9nDpg0LKAWEuv9aWgokPZ5gIymfIxbXo2t3GPD1Dq9QWY
U1gW0E5Fw0Y8tNAbCvoqLwpWzugIijGr+YGC9BAfx/VY6Sd4yPbaK/pUzxS2Rj0FBRW5vlxdg5RR
pgRLP/4SO/G0lrME+FyDYMscEY6ZsDfCoDersbBAVFYk16Bk47323uffOMuNid+BpTUdGeF+T2qB
mbFFKwI6CNKyLV6Pcn8PWvy++L5Ci/SHkqkz2mvL77dZdh0I2g0thhbFQSTvfU6+4MuwlGE+ZfnO
kFdilxpkjnktZvx7jc2kRB++bBSnH2aawEeWn5RcVKvTMiKLVELLfZlpfvz7mlowGY7DtTVa7y3/
HFmEJQ7lEkwmM9Ts6tZx2SmCZs4IsQ5uUPop3+1Vb+eqiI6EPQWO3fMpy7JwuyAASFeyvZFhpE2s
Hpjx3V5WeKWKvsK9aIxGq1ccWO+xbwH0Ku8BMXWTvHAhJPzocJzdr8n2kUffMuilyY+Se/lPm+z5
xw5xh+iylA+cPW1HQ8Fk53ppEs97UWComSiMy5HsrRgy3MJi4/tpFOi98271YyB2hnrBeZjL3KUc
aaKzMGpdBnjpSK5muNmB/1DwscrqQDCCYWLQIE7Nr1cp9IwgMg75FbwyEL2SivXI/Kgm7aKQxWqK
1km1ofe2pwqt2H7SDK18CMMRiEj4yv74CM7AyA22BAlhQYA2ve0HboxqGC+/N6zxoBRoabZCcP3G
KkTmo3wsp4m0lqxhO2403u1YKU1Lm0pz1n0n3uOkQz2G+KyzYFh9TYggEgCoDVdcrb77rr3dws7g
8QY0mPOQMn9toa7709Kf7lZYRtPB8J2dz9bILCqa3WC/K6kiD7gPPk0uFw8efU9PSseF5tNJqTGv
zbMMsEWv1nO4dCPoeh7Yy6AW18H3/vtENiDL/g02mlKdMDSS2xa4HnpdER6KTuYOIjsHGOgzH1K0
c25/98imxZnycjxqBc6GfOmTEj8KNra68DwpIcK9I+Wj7rVCWTZBRCJfHrehOonYVIKxfF2t2A31
+6VRs5HKgCfwtSdb8VSpWtQP0Wy8Xz7/TSpIFiV+JvQnczMTE+lQGr///uKlEPs9VIIsfWAJitDo
/0orIPjRtadT3+iQBb3gSw6XzismPAOkGZI4R3+IlbONr8KHusbzSrGHyHFrqkV6X8+dxNVh1mFZ
oSoi4466BoMeW8eV9SEsEw7bC4UOcdNM97ttWK38yjHHOetsHlyG+RJSvh+kBLByP40+CT+ci/+h
Lb+QCrMfVGlk+ynjg8MIQ53bstLzT4Z6DJeCpYK4IdNnSpsH/RS9HlCBqURSiYyudvgP2vEYNm/O
CJZ7v41wTesqvG1AgChs6L0lTz+gkS5kgzSQy+rV6Ahwh2rBbRuJSPdXKSyhsYkaCN87CQbChSa+
9wCk3XgxZv9XpQ4ZSQ2FLh2Dl5iV6HJE9aooCO5YMUmzO+pVmRy+WpSRfI4ZpGEIWtbDKr+sWx8s
ojNIyqbBhTmCZGD5AcPnzrv6KTyny0BZmkqVhKUwr+6OZwrVwgoAyLKdDQFhX5C38l21yzj2IZwn
nDvMMm7PrurECtpfaytRCDr6kjZ58I3SbAB+ToSjQSlBmsmBzeF6mprlAVxnMvj2LM3wYREQQSRE
p86aOMv00j84t+K5OWdug94BjC5rSwL0BxywSgC6KNf3kuXmw0m/midnbGLeoJx5mYyJX5JVPDgT
CIKQ7o7OCKv6GHaH//fYmm0UKeYrpjD3xTRczyPjhLtGxKg8yiZGAP7MaUoYagIlWilgyoe49m+h
Ngk+Y/kOVeEXaOQ4x12Vzf9v7RFyMxn5y12Fm97UAMj4lAM9fCKmVolKWKs//ge/satVL6igz7ih
LjBw5j2w7pmly0zfhx8n1yqzHH5T/+83QbCyhKbR652M9QChG7e7I1umFA2XbyEY5W6FLxq3wfPu
/6JPDtZYL3I1Y7g6qQxrlrg704Cmq+hlINcIZl0ZmNjlw2mr03uzvr2NivSuX64D/lv6f+u/DtVD
AoTSZ45kHcOxQZA7545PMaUY13MAmjPMDgrolqzef5SFhDv8nqXsQxV9sxVhsk1VhmnsY7aBwMSN
eSHIc2zQYNLcK5dUM5/bkInoaX6WRnGDvMD9QMNe1PGUzsyaGiD5Bd4jzeiv5BCmVRGMwcegvRM2
JUwtFGJCUJIEDwtUznc5ilvYrngnDnz19PBe9uQluDCq44k4lx1Vnr/khJb4Oc1b4KCjObapEVDS
qWOY9Xm0V7Mqfl/7xR24kBm2crlzrOzZWmuREbiLdxmOKb1w6XPHd2sNgJ/NimO1iwpRC9E2psMb
IM+e/4HpQuPFA2Sv3lREcAtNel/K2m1DjQ02FEpNu3RCQ3dzSz4xqoJCL04ARBjDPo1TadE9SNiV
Zous8OJ7zIJh6nFLX5FGs5KeAoizdynhCpoxcFfI27rF0adrjye4SvWYLzhLI+KEx12XNBGAaGoD
yt4VluA9wq7pzg925Mvlup/A1sdsxrD0ZbH9ic0YWLYgni4wzKOpqc6vL6gDDV2orxnJeJ+dy1jR
83zFgynJCaithObwHUBWbrfCdzv0EkYNuzrboLzUNOKv7pOs/Is5B/YyA/74xGQ2FiVt25hWE6Rs
alxcoQYpPXm58hV1zkFeumpxCAR0k+s/fzRhlnwHW0YWwEFvJ1puh1ivjezPlZ4UYvwnNUPwVvva
zwCGv3CBEt8w26b4BCU3k53Qyv2Te9wmBq0O5nX1UFA1wTdptDk1x03LQXYT4F1ASLP+xraPQkxU
hKDacfTqzVg32YOlSB2EVuUx4ZOK/AG/x78YrNqk+NplscIQHTgu155Y42Qk8kiW9fGIDI3PSNhk
Uj8tsvugOUrsV5zusY6cUA1fVgr4nqg6Wbz+g9bh2ChqaODIH61Y4QlvDEZlL6d9ZmHio7auWc/3
XKO+cXMkZ3EOCUd0hzNPMloCMT3MSXbrKAWh6LhRPgmpsAsQJMx4XlEzX99gsME2x4N8H0pImtDq
1LMvknuWM//qYf5wJbC2UGnfZpdmhUOoWzwXYrwUCHp6xq1LFMOKHX4Ov1OBSpzLiYu+YThQNcVE
JvZcc5SixzgBbYWiODamNBXwT3TSqbsxIWFnIoqV8tXIBb/3M9Rjq4VeBDZMv9T9tvD+cWB30y2B
Z1KYEeaJhHSOLSBwFrLGqmaEDepCqEqwtxNELNCt7Kp3MnhCWvgvTgiRBkOe3J1YuJm49MlWzdS3
2YWESlP271s0pxy/nkue+d7dovb99ToW1Y6AzHhk9uEnTj81iYYqpttb/C29CnD2m3HbnE4ixbSc
tN9F8cjvPZGE8JurT9dLBQOySPycWf4KSJyeZSUHfAMUjT3NIlaDC6EE7mmYzXCt4pa/9zmjTorT
C9DqczDt+JIQDSccrGaHuCCRQy/hZHi72NGXh0UmrPula8lkzeeF4StTTGaIoU933OU1gpPkGdym
eahbAM1WBoAn7xM3RNwi4Qrlyqk4TUvGu3LpxO7jCNpvkQRcwKHBwKRojNP6unRFyADKF+F+KYWa
Grp4cS+BeNzbJuaZ1NL9M9n6JjWSuY0KI6h/aDJw/IxGVP7CiweDv6g5inIJkzEXkYIc5ovsuqW+
xOzgCE1NNynFJmyFOz7dju4OmGbxx60UQ9D9YpBlJ/ikPUA3c/f28xb6SgL1oahSIgv+i0M77gH3
Je9J+xCoyC058sT6azH62Ve0CIMTZSfF5DzIiOmqFWFeIQ1UWJE5FGgC/B7tX5FxbqBDoG5thSAJ
nLwfzAjHKZiSQMUWUGLysy4xggAHq/ffTEGmZEhHG1ppZhFkwwdUtv+7QUMQytYcmuoC01HA/F1r
EQef4EJ/I3AC9G+H1/l0J1FR42U8UoYR4zHYcxyovITtbrOs35ts/UvdV6F/jzF7k+IMtToKwUiO
58564b+YyQ9naLJ9BLbvTikOqCM9PaGzVPNrKI1qUzGJIZT5P8c//6rSFl+kKOJPYaG297uqOwmn
ZfrvXgDNECOJDvqx5b3liDDGdmuAli6SR82HFfIhfsEeto2J4FTyxAMXI8tzY522Ni8Rpmd7Dq0S
XVM5T25HPKLLnx++av0DhqEmwxcnuJrAuWBcjXBaFHwGl/EwFSrrALr01qF5GRw1HzdL0eIIbPHa
OfpxjOqAkTUM+SGSQxfZMHytQds57tVpcMNoqDJXThfGO2Y8kRrqJ1+z73FPZ+Kp4eolMB98linY
uVYONCUA16lpFUVm35MPo82gqfHpL8irOpiC247VRqcOubz36QfTmWN4w/EnbDkKUwl1JuGeeWM5
i24SmaB6Lg/+ymR6fIwu9IFDxiFaAj1UeadOvevuGsLbU2SKbkvQl+Cy72Fy5qCptS0wGZJE3DbM
2k+uqZKFdrnRb5GlUEwwORYP3DOYm5c565TIwYA3gYCGcTqQzsxBoMqOnkT2fZ8MA2EJPW8FEVkM
H1vqPbvdRUQUoGhpzn7SUR3ceYzaAryBbR2IjB/eJsoWw7XHNTTcUQUc61bdEgJXTD3mksfvFHmJ
2h0u3YdFUEb9kRMftdjhfaP2e2um3vEsETgbePBTVoANLIRhqDv16S0uFkgUv0iforIpSC3Xbd06
YS66uKpvOUXLxUsQEO+o+PZkmf+Xa4J/pgvmnsBj8IFUfTywR5HFQ8lk9l/4S9MONbKdqo71MQDT
Bagk79ErJD00WD7QvhIql+X0bqHDR1UkQJ4P4RAfUTX+h6Bxbci1qDvEJTgWtQdQalf8rFGHgQ9c
LBYgoekYFZOzMriyUwWW57QaAqmTgdvaTHG8i7ZCJY3XB4tUO4IokZJJ9RPvy0eXwCY/inSyMCMS
yGBZnaeNqDZpM6m7PypXPu1krT6Lpey9XDvAtccFxiMZWb29axfGIwx0htyTra4R7I+sD8MvPFLB
OWE0NwkyGcK0Q2Rwt9cV/oqhwoqn6L/HcQKlywLBjTeMcWoZeFpfm9AqB5z3YV6am+pkAxNqjD/o
yy/w+cDvQHrOg4IRrN8bIRuw9dvXgx/jPXugvQM54pP17QQ+9RLeCl7zdlWUzjPOyR6j6SlNOleu
r0oDkVfGpBWQk4370o1N6qsyB8R2eTwPOkhheDCXWnN36S8P3KMYmJ6bsJqn3XKxEY84M1qYAyCg
GRYU2/u19JNmVMEMxYyI4RjlDn8X03Ijh0X42FSEVFVE4ZbtG6bAFQ2LipX7G282YTWhMh/03ZyH
9GOAv3nBpRMOKLxs7VH45LizHYK3q+abOSxWbHNRpZ8WqK02mnbc+XJqfx1Rxu1Z8dNUO6nSsf55
Sa3IdDMR4tp3/6C4mWYraSmyCIw830YkKIMyvaTcLUcQlvqsssD8liqeM2JhMLV1Lay6mdBhrwiF
m3iRB6qVWxGKde/m7muRLrCukg0/XnAC/uoG0vijMxzjoJkhcmXuqP2Fdw0coL2ZYXKrC1OydHXF
H4kSUH36CDa2QlXiNUDunZ60F2fxaZLzozNkk26M7j/QtvhT6D6aQb3WqZfrJ7Stl4DBw0CuBZ7b
uSOo+SwCz6NHfcSszq+TDF8Hyy8TsR4/eJnAsK8/hAxJlMCLFe3pO+Ew56WdOBnKCmszDqa7ImED
mxdjsxB1ZWgqM6ynyer9YQXlm5n22Z1fR3CfFffxLvKQ21zN6d3YOlRp//EDhihICXLy1UxmLhSO
KdjCXwARs3a5ZcHXnbfJ/ZUzkPkFCpxeR7i8pSzaKCC6/C4DajjGpfCxeX/G3Ts4n4Ea4JP+o4uv
fuGeFVNHRCIgYHiCFYqZakH1PwG+9EiOzdic9PjDRyFmbm4MWuD4J57OO7sRn5waMu+TWu8zmAx6
fM/jwJFsxW2yTZP4AIJMlK9X//uNFRiYviFcE3FfHWEn88cDSUw8GVHTJg/OhnwGRxCZL9L7DNrP
p4iYgQxuhnBhE2+60RkTr0he5KlGns/3vB3DpCG1LIJjbEIxushQ/nhMjoqmlfjHvUbYXz8twUE6
KQ5wQC9WXw1i9+ymyx1bPLSs1QQo8fr6RMc+v6LehVwasZcObDOvqnFTnjaMAfN4xtKJ2jI0GQTd
32AlCYnHjb1MKF0qHe6zX7BMLWs5RawRx+CXuOv7GM95EJvj6pjBT+1fhgp5+aMDfdPPqKRNhGI/
A4n4GtNKRZD1j4MqH7mOdIoFPDA/WvkqSuZOn3BM/se0QV3B+/lPkuZv2b9Rsq5Fc008ceVmpAu1
Sd7zbg6zwhFLY60UJFusiQ6O3Q0ra6ch70rDjZ8PAU0kJ3Ph8KndlvYDG4IR29TtjcMVJpz8/TFU
7KZzN1gfNscldTKi5xILK8YLMVE7+WauRG7kHCZannxmQuzE2gSc9OOKnFMzaoIrnWoq5Jh6WFIS
/2IOuX5yqY60/oIY4PhoxF8jkqik7LmsO7EYidDSoerDDBAnV+3aFWaE3kUmDAEZEP8YpvzhatIP
dszFb+7kc2BE4zLPNug+nVyHiSEBFd/XiBg0nRoLDzCgBvGbsc9HE9m0EZoYBkT7n4lFxyzxfAHN
PAf2romHigv17Ij9CI7oBsTFkTI+/OKGG8jQ7yxMrTERmGhEOAXcC9uubloHd6xqSbuhw6MhrIIm
vSL0YFcQlDwHEQcI438wY2KrvrVEzMQnT/mQ7jjNtqI7WWLEVXeCBQcIY0uGY8WS/zIq0VvTKYkn
y8zFaH5PWy53OxXo0jrSVeSk+tYse0Y78TX41EvZkrhWwOdzvS8PGZEqzEyVqj/FyCda+gsFGxNJ
rnqWhaQ/RGKUR7meBkxwjtVV7aaA0Cxi8LdeZ/edUhZyrYbFcVNVTOOQuxxSBgfYvDvESTmANHax
KhyZp//jrpoKd9kOtB9U3isMQMlbfXgjFmUZKz9uBvvy6CDqpkfBw9UsnU20x1MYdDGhvcNfqSDV
9xQ56uCtmX513CTwvbeVilW+T1dIglOhwDvNQSAVpSvYZTosq7bLSl3isKvakP/oP4bVc3EoPO/Z
yRzgaPqebyYz1rcfIFgnyzkXvHp38+7ESRHi9sa6FkmtUzYqFsdCj70LA7mCMjMUUyiAUur+K1JX
XrfweDAC9EO6hoIWxLjRMxR04+HSHqKyujoZ7JmIQ4rZsEdfYa6h70N/3lnHzRUk62x6o1udsNee
kXLiYWnsUwB7XnJ0B5dMcfts+r+o5TZ1MaDlcMsDZRwfYs1I47M3wnQyCUo7XWzuaFVfjuVni0lu
6hpupb8refQeaP/mzxfkrBj/mumx/nbVc/r7QEOKwuqgWxDXp+0b4kKFhaIP7ESD0gKK91HxtyNl
shJn/nwmVoBmWgG2Ac5W+jIKg9F+NxVHMc0Ip6XSPSJqPPq3OYA5/Jx77TvQyPFSqut1EqKRQvHN
n/+gF9nnYaZIwDhetlX3FQsauvtjc6icM1Q1Srn8TTjc0c09IvfaVRgu+G75yWdkwK3r/R2gPv2l
wN8r/lhthgQkYf9v/qDOqhPjC87rqkl5EmOCU2HQ4B2HyCW/iQPiOQefYzMdcDcX3uGUcQiyBPp6
qaGtxxDGMD/40vpby9AtBmlxCMoRXLODLfkLXFPp5++0MVaCumA8dBJi5xaYnN/EjF7E9Kbgwwxj
xVrtIV4OoBDroA873qP8LJjjpeI3VRUeotx62gufybK+X8k+cFiCzhuSIXI8W07X3mCdeVXDybj9
o+AVWoOEOWSTj6/K6Iq8vdy31+c0ZicNnrXxc2c+9kOoMJAwy2mKkq9YmqZqQfU069mmjKaRYxts
C8nXj/eax9N0byJtk/GsjFNJ7oaD0mu95n54+aMdunOI+G06bX1MEXs7m+QrRVPOBppkBdj4eG/y
HybPiRkLkjtHT8KhG11j3YhDXQ0mY5O/L/vQhRNAJLSpB1crJwKw4HzJcwCVwEgkXF89vLaiPvVl
sKgE3LAemq0HSk/NII9GgwTiLyp6L6lNBsnosrkUyENVhLhkWai4sblL4e45l0/6ZRzaHKynvOjo
xkw7uxMjMb99G6c2uBAFjHvZE8hnn0q5oaxTbAT2nW0Q8NNg7QB+zv4DfvNBkjN+l5/SqKDFT3Hm
ibP5HpayfSAGxIuB7Nqd1FgCuznZZbQYzmqO+zk9omD2kt5eU4EXbCWwKkLQzlNSyJUZZ+Ce8gz3
Z36dFi/LRtIcKVYJByozf3Bw1zHDvGjEZ8bUSASCdvzlEmrs0lJ1lMjgKxpBRlkx19kTT5SPwmuB
XWuiwYZaVpvZCOTut7lH6Y0Ax6egCIZMUB+FlWD6eBPQIVRCE94E+5oFcsCPZOioq1ICPK1BR8FE
pyiT1UyD4K4uf10KI4URO8OC80sCXLFGkx4uZHptnFH9U45FpVYAVO8CFyQbpIZMsbCPi7IPEGN3
7SeUG/1clsIcvmc8iz2hKn3JWYWH+mFiMK0+VGqbUJR7B92BofonXiHE0oU7Lhz5ux2eyack3g8g
GcLfELoT7Pt5j623LsBfU6OWUnGqEAh32IZtOFElDLG3cGQKDo8L0RULzGpExEEDPxPt/tOh6t5A
BHJPguM9GQ3I8MRV+EARK9sdvgdaIWhJeNvpdtmwA/L8e+qy9VR4WztedfrReDaaGolFEeQpiw06
jf8577sxkIZYckt2kzIhJTJhHe0VZqmcL8MJWJahsYSAwFhTBJMsmxvKGQ1DYk255eeZLQwJ0Jrg
dxpP1haBRSVrXjMh+XXaVYIVZ1ZFMtXSGRlJ5+ExtvRs5sNCKbwr+i7KbUQDosRnibJqTFdyA1KC
RuEJ61vSBc6MgS68RLmzpGsnUy62JM24M27Kr2vLh0ZUro20ecENhhybmeME7ZyJoyd3ilh1HyPu
CfgXnpNZfMLy/DQXrPqLYECGZNTKkAKSpgO/j626ENtepH7d73cPQvIoFMKDvTKhw+GHK/BhONzJ
fCAjCYPqhI5emR/AVjj9Dg0M7UQWuHH+krPxBuqXMkI1tywdpt9Iu5s+gr3DFYntV4WKFKqrlN6a
yF1HaZ+AJf3mBUFl6eXhrTPJ7xTTzrGB8Zk5GAFnO8xRZvOFp/WIzgUjyO96gxxjSTWLiR1uneef
AzyiKqS1hArNgl1AXBvEGR700gDi4S1HRM/c4cQ6/p66aC3cDTFiL+pAkU0dn/C8pzkSy6PevTVD
BozlakAF8Zj/8sWnFqFNR8Diai9maoAZ06wFQXmLYnAWn1/KvvtixjFIZ7eigCp21WyySPs57EYG
oZr8eP3bf8wbAhR0bqC/jL64ciRoBFYcTAW9lKOt4/lV8r//dPkcDBW9Bj5zMkJPD7Q/0uQTcw5F
k0bZyBF5+iaeuDJ+kTpujiku/vKF2TSnbgdZOe2hOR6LItonPtrn+jqf+VjttbGFlFXrnEfwPDhi
+68QGkmKuzVYCrpxoiON+RKrXDjDc8ZQ9qlKwdwAKnDJpIYETOTo89HpiFm6t78dH+esh8dD08SP
THar1MGCeyBHAJxYnNTi8F1sNHydoEwVlySO3SmjyG02eC2gc1mtMkDXQSETapk2GPtib4HSWXaA
iXNpj1UrrXuMJCtGcxXqAmLD0x4gA+tPTbGCNcfXFOHzua29pcKazT836ckGrv5qugh0bwbcNAGu
tC6fxKEztUuI5dnFYnn9kSJS9stLGG/v99+pJFcMHw1eq6TykLqLQoKUCMEZYEYgq4GIa5xeET8I
wzHXXhhfiwRLtWM3PdZm/1xR2ckfTJmiMrSKUzSRhhZOlH+dp2+rkrROa0xvMBCr2ww1dqGnBd1u
cqtnVZfDtHCsZPfBLOezCSMl0lCsyVw9lw4kHjlObLEE7ak54Np4yt1z6kiwhw/STXxXoiKYrT+S
22+OeGa2j7psUoLCv6oqx4Car7Q1OLNPt0qjXIXTCIbOMqfqBSeBDiTu6FOzmjQjugPzSCJ+u6Fq
xv+yFt/3byTYI6wLzY/gG7/gs0TtcRIADxDkI94QacIrE30fRn7ZDdLQd0MqT4bY4yECaXxsm+YV
0CZz7g+lIJtO2PgxcGtYCdHeEQnnu1DdNsy85LsNtemrBLEz1/fJUWFMR0faZuBEsavxSQydD6Hb
Baa/9OypH/wMM3cguJZnfdAa0e8/QRoBs+6JxFRixNxUt3Jde5tHNDnV4wqBievcH0/VGA0/4SMb
MnghXD6odaVEwa5anU4EFMurC1HllHpsF8r+ZI6S0S6MOg8ld0E44GTdx9lvZkDb9rPnlawuyFNi
1cTqk+dEyQWtEcAllDh2L+vsxr9QziauM6MkAjsusyr2SNA2K0Y9yCZRK15tdydyrKIQ2RLpuK2i
UwOS8BsfjZ46JIgA3TZI5xgDpZ4qItnHUZeEUASLcC8ZCHk2QzJbmquudYGeWzbv0VkwBEN2Ovlz
K6nkpyrAwB76FWYC9fFLmuoslCZbXXODaZilw7+TBFDuaOdM1FlcfvwE4NczUhlrQFqOpGzfvvgH
HpLQEBPPva9x80AapCCz017R0dVBGcb0bbUkepJK8nLS1b/jVI/IrDxgzkDFig1FGmc4aZ+pC9cy
vfH2PzRlTc/QCyfnI0hamVy0R586c0h2BlCDEwlGeH7NHlZ11jlPT7f4mmX2bStki//dr9tlMhUM
zTNtTgzGXzL80oHGL5F3vRosxOyQAufR7sJw24CgLiiNjwHWH6aIEFP4dHZcUhPzlSt8aCOpelZE
w2oPK1ioUJStX0tmExwOOt8pR2IP5XR0hzerWBb0ivhvaduWgLhVWsWC84PXr4qYwiIaZqi0+k/C
F0HIntlYN59HvsOA4P6mM80EpzDwKnbteeU0uWrKuvdWZPoRuVD64TKf5gZlMA/o8J1DbF41KcRQ
xadtrqzykG7LxctzsdV91C19NDAAIK2OLFE54zLLGITbYPaBA58n9fkSWVXQhntnq8winnHtRrFB
kv5vWhd6C7Ic286qi4+Ked4SMXA9jVXwzMGb9WOV9F6KW8bZUY74+PJ/L/JBY14bXQCF7wIqxJuB
PMYGRj7NnBDsexhtebRRfjIRj3lgjMnOTfghVDprDtRxntlfV4u0aNliCWp/u9x/3MIUrmL+Qkxg
FVGHxkAj7MgYlR7HHbKMyoadpwj8nc6i+PkEfuiOaoBEsJVKCxFeU3RNLwNt+M837iQy3HJgaL5n
8t1tSjlHFise504LYKWk3yCyh1z0bXvhv/4W8iGy2m2Y7l1Gg6qvaYAc6S+DipJebPhB6uTWoyDk
tHUQntk283M/aLGXHOZ3jI8URItdiKxQ/fZS0MVtMuERhNOW16Sqb+C5UV1rrR/5sKr1yfWgMqsp
B+N/n0I8CApZ+Jchr99f+8cI87mYlqhw6Cwi2tpcgp3En0MzllEQ5ABbABEjI/SKkowsXXIOH3LT
FJYAoSawXWMMVe4Qx2zOZ/kvajR4B2ycBG/9BI0OqtScleg2tHHEzR3GyxpYvU5Fmb6xyTfOmB9b
Z4+Hf+JxU9H7lnK5gBmVBzvEdRfmHIk4X8K9hiU43b0cAZE0csjsIhUdxZwsyAsXbPwofCa4OtZp
rVeDO79Tjvhh1fId0+DpcmUXTOYUGsTUtfOYpTpCUC49/A11Im7N2n9mtp1WjKqMaQygE8KH8478
y3/G2oCn9V4ogDkx2++1jNxtmp5ufGNqZ7nUrlk8EV3EVAMKLdf7U/5j2sd/NLCguItiKZjTk9NS
wDvCPwN6FnEjI1AVaY7Wc4t+8Uste0Wi3rj+qoxvKx6dCRqaXXp8HKU+ZUfmgQxjmhD/vHPbTXyu
tWzCN9/wagBgeHInHt1hrLNwDJQQAb6DWZiaA18r4EbHNJAgmf6SaERyytCfYfUdA+uwlOqV/JBr
s6g2j2LuYBORKopqs6H6wrm4fWylITc56apLtIc8aXJ3L3GOyD2VmwUUSqjhyGjPwBOQYO3K5sEU
UxlSSbSPyPQHy8CBW1KvLWdSR7o9tZ0yeu5oPwA3Mxzd5OcmvpT6qmRPBJhynoBPi2mbaahe4A8K
1Bm0e1Ne2ddoo10QX+mLNsbZHVXv7ypmTtE99rXxBF29pLE/Xk7vZAvDEog7tVXU4Oj1UXoRxXzf
Zil3Kjh0xlIb5anCxoRgu+VCRkg5M3z60sk52Lps5LLOfYHOvx1RiWjNpfK4yJH2DJqg909/rJeV
tbCz8Ke2ch0lziQvNmVopsneHb3gP+N5z3BvMLXNgznKvU21MsYZGuLjavmM7kOYy4oQfv+9q5LT
nn4UJUtMWoXK/ShEiWlj5G4aDOAMlks5An7ByG8qYi+Xu7xk8N8fmtMsf1TmmhtgvHOiSV3wX4EH
ds7UKMRwpSm4EI7xeIL5V8zZ390/HABiWt7lZvPd446GoVFzUZT94tGzD4ZQEU2g89y2nEouFcC1
k3zNmxDvQDG6bTTkTQe5s/lK1VCxKU+G+q7xD9mvS0AO+UHaJBEHWxk1BKEoxLZ6MbjYwS5bRCUN
xggXR8K2PVO6R0Fzeay+STm5bFc7foPiFSDJ8kLE2yukHw/RM3VKkulgP28q3hQnWyhFymx8e7Es
u/7skP0bztakWjh6/FV+VmoMVdVVFBjUEZeaRqK54bufVT1ccgXedl7tds+aaI39lwQdkQ5B5rSO
/YHeHx5Zqrp9Xr/osg7nx0hK0v1nEHNjhEjajHxf1aw/dPftSMAqyv+04uTlTTTAEVCixaLJvlEk
PAOqdkFvdZIpOVRWHBZg3YWv3rR+n/89uNcylRXRQIqY4OGE25SdIeXnyrJ5nA7J8obwjubj20oT
9rVAKrH35OuNEf09i7FWlWT+G19CfulB1WKgDQSHKrp7GqtGpFrvWyYW0LFaTyN4pX4Pg8yolLK/
Q4m+404FIZuDQiHEwbJTqKBtvP9YI14JDp8RThLN6YnTHarfV6lusE7w8bVN7O6iGEz7OWDILooY
2EAVLy0JoaPfuIfozivTn9T1PqNgPx9UTPYctAA1U7TxKVIgMENFzOnQiTxfDhv/a3E5YFRhDQ6B
eL1aRpVVdcI0cvlO4GGYfy7bc17CHNBQ/XhjPFRFLXZ8/cnKlN9iz7CQWLmlyo4d9hUGTKBEiIzo
EV6jPa1jbg7UMF1xYaPybFrHTS26JZpbzuc4OPp377CJ7+/rik0ie4790YXh4YJHEGY7blhEXRgM
k9oHxYFd66wHTLLzvMcC1pC3v94bVfaKl+igwdLZy6yPouQhV0HaGBC+qn5QkdRAArhKsGV4HD/G
RPpm8w6ZVrfxKB9prPTUAqYC91yq5VvaHiy1JeRdhs28WBca6g2DEosiXcx7TAMRjCGYFJ9kQM/B
ERww+xUTdJsgWSfK9ZVfJp4pXn+gn1svYGLTgL+PfO/Nw5Se/in1nc1mf5Zhy6nIiKyHhog3DLUw
SCdJjnBxUfpCsEU5TfX3zo0egKwjM7c2j838tIjjPpTcpKklKcsotZZ3SI4dT7iPRAXFdn9wG4VW
N8/E6oc2kuaR+Mg7pbFB1h4vOqPs+VmwGtdpN2/rENHpEn8lWuYXRkHVy6yFgveXd8LgpbO164Oi
nZrbhXmxip6iS2MAKHDrLZc4oj434LLVVAHnAdoZNr34LEYETlq3woxrF526mJrgt6FKaEtKQmx9
1Kk8DLn2VRZyH5MgG4ds60idZwR2lMFrTnD8BlOzFouq/8MGi+PCG3FIl2rTTiTYrNjb3G6pmfig
UkEJB7xNOFH2J51fA5+qRCTIzkRHh30Ld3mXUY5dBLveqGnogfu88CUaenp6qCSjKC8u34dRPJlp
3FpMu+sbqovb6vw+u7dTCG1q+cdcbPCD6PMsjCuPE98SCnMn7YKroQxpI2UC7gUrqXnHIg6D/2i5
xAXJLsKp+qC+QL2f7liZkqRiPCymS+Z14TfTvnXaVsB8KDH/UEGaapsRWuCUdy2fnk9R9b4f8fRr
q3oHrBF9t2rUbneryRmmMCwSzo31/CWct5FjU/GeuwGkw1083WghjtB26PUP0QP+wPWFEREydmiY
XxIxSF8dkF5mrRXSrqghix8P4HkUlxbOjKpjrj+9tWBVBfFPepg9amQsDPAJpijS4g020+/1nJa1
JXpLyxeE0Y62QOOYT7MueROkfy2wrfs+sh7nd41JwccKTqu89DK75Y0siRwqftUM97e0GpH/3HgF
jv7rIpIUDp+XOPNBNH1AfwVsWEo/mnw8porT1mTqtUfXAHginlkR4ziFpYsp5epcW36Vn9jirsHj
vCBELgIPKmRD5y1UJxCEohjT309CDsTKL/z8/y6lfE9UCBSgUrX+hcbsl1yLpKmSMqJJTAaNe4yx
V9bDw0V2HuZ/I+qL6UJttCw4CUvpUWUNMgRgZH1cyIlysRCuXE2Y/jR7KC2CQG69jAlNZ8b3kjJB
hSAtF8SYI9lBhBtsFpX59ptkmONTkQInE+IDRpWdpsaX7UstZZnFCPqou2VShWCCJU8iHlf+ETNI
6bkMi5Q9qLAxuRsrYoYw0ZDATwzxRY5LMCX3wmhdCsa5NF8cOY9i+HN3M5gKKkWkLfVtlk2PZgYJ
oQj3zCUq7eeEZlPv17yZuRDUvjMHb0BJJpTfhzFskawEsK3v3h+GC8AZIbTiBM04ZIDmmmk24nlO
uwyVw3eXRPfF4Ay0OGTMf01J8EnwVGRjt6pEetBGaV9lQOPlxlzQVPjc2B2kYfenWw2+RabFuyRs
2f5fymBgkI59hyVqTjp7ylzH45egK7CDrHurhR04UP7lsG4ZbqbPwCsBhCXcVuszzCt6oWziLiyP
p4297uBcTXJ/Dt8PkfJ0JBB5ROPDRn50ZvmdiK9g+7l/D8z4M+7hoTmh5TZw04Lu21cliH5bMDnl
8Pw3nE3U0mG0deIt02raaAQ72J6/XMn0CsYuDKpQ2t+AEzv0BVfrRTJun3F4RmrmmifC40gg0wNe
OdVyzypcwA9T0xFaQl9eHURS9fmPIIbltYbCRStctb2Lqi9OlqQ3SBr1PzjDvv8G9hcR4S+dP1ze
9Xql8zdeG1u3oXbaOVxTUSn6sucze9zWP5th+dO4aH4RkH0+sBm8aKQUrGojh3lqGoZ4vsQgRjXz
jHyJ71TWwq0Yr3I5TeF0brq4rPzbWqtVa5cZm92lBhW7HfF+spkgENM6Xh/o+9myLoxRDfS8QofI
zLQFRbmtF2l73TDdBwS9Ckiw4LqoC2lBFOdsCmAeJKMv2gpIaRJBQI0SglGtbI5/LtqDL7kLq5Ux
sCebClg1cdvimBTvOFwGzrVxIPbkUvZnxjVFeuenQV8iVNvJ9V/yM4IdV1+DQNdRClVPzC3C8Z+w
YunvL3ui4Onc4knHfbcU4+ci3iwiQHB57qGwB43gZ+zql58OkzY6F4kKtWsiXl/DHhaj9dshtXQs
H/6nkxqhWtDLCXXrmJtHEM27VyJZ84u6y48+gX3rCamIV5TNFu0Pt7CIbbRSQmTm/Y+XypkJ1XNn
guMagAp3KZyjfaUt2WouMQnRsDbYRsIbdB3Nzrtdlx/I9sqpb0ga2vIoI8nJHWIUrDrDMw6XhOaa
xCLJVT9qwhxQB2rTDJszwtE6uV3lJVgrHF/y6jEDX6GEyncrYldfhf6RQJbjoq2efiTCE6cNHT5K
/LEsNzF7y7RHf0+LhaMgrH7l8WgoBslYXw/ePuC/w0HnLFwrzYIQ0F/xnPdBLHZCtDltOE5G2nYz
kZeJuKFxlueUH6eTT28RXxIGuzCEFBqQbJ0D5kOLZ/IYjN/rX2E2UUhT9Ptofj7TeMFJdOM5YAwx
N2Xq1E5g5TvcjdE4HxYw1ZQRJyYMP+CSg7srlmsQZIqD80aUR/CUbDgB/f8vttJ2fMULM4HvL0vk
aCJCvdJklq/tNfHoZuIwXQnFUziNvVX7sc39zZq8V+odXDE3BZzUzgHhAqvKL/hyI0iSa9U2hnb8
/cRcSGry3Ux11GgFTJVomEiZjFLVgHJ18ndMisQZJzeN50w3ZL2uUroP2LKIBdD4YTWAa36lC3Ls
PWLOmMApRU6EgYMQwShbjiRKHBjJaTMxnbYInkMDXVoEV/Ad3Ge9JGUbBoLm5R/UUcHu1GvjfAoM
K3X13MzsQaTu1WBHD/eVDQfpfING7KcrkvbPfFoJQ/enyvHdCWBj4+GP9e3TON6u33BhLUns+qVi
mkrzOJmhbCzewxPcUnOJeRlk/vYQPMFft3nScJdUdbpva5ALVlZlspyBgTWtbmHVL9COWn8UI98d
+Sny5Hm9YA453Qi4TxZ/xHy+gxOQ56HB81jTAymGo5rUZzssSVkL+C1WmRVhn4vb0l//VFbgFlWJ
R7m8bQNbaKe8DpB1GE2OIrLH3g1JCmNnPcU0E5h3JCGIPg4MV7YKY+zFCdyq0o2+W3xnXqOKFIi8
fCnT9on1/dEy/eo0kJws8rxCaNHrPpxiJEPQ86MQBkBSHwT1gmsWhCHGqOuuHfoposM6AVmU8Qa3
MMiSqxQzDH7uJ8QQROVVkOE6WfkhQvTCXrFhuZZJQVl/L/d2c3m8HbqEfN4v0QXqUJKhI+ypjHSf
dCLVXg9tSUsjqoBw9Pb3l9WdLP5GCo/UhzMIfTor40935fqJ7fKb4IpDdqrARlgY93AJwk3wf5yD
KeULxpBjusLb6eI6ThvXYQiiEFAiRN659hDcrvW88lJqZnEAagW/YKIqjBDwaVitjVlccvp71Y+d
JZdwgk7TU2S65KdeA5LRQvxJC16H9Ud180Y0LDu77uf7GxBSz7m+j1HR9mUjmjTSVCZsanrZdlQY
qkp8YcPac15dSuQnOi7FQBFovrAi5gt1Cy1Wc1D6FljuCJef7D2yNVv3SwmvGR49Cyu9dDNuhslt
rAJwuw3QJGhgvCW4ETGp4S1YXgJaXlmCqI1sgs9qih49wlTStUcyeLC2gqftXTGYXMJ6ErOwcttd
gnEHMrgNpGH97FiT+5WlOzY45KuUXz2IRRa0FGjoHqd5YNdsPNfwm3fQDLLOOXG6t+vyVz3qOfM2
VFKASL0NO9qEqzTMdSDr9QqwzAhN8w/0Q+Fs2VywkZxxXmHTWp8uFOTVi/q7hzc3y6E4l2cuWRke
9UsY8EPkFsjemc5LWlfUrJLnYNMF796qpsgG0kdHK8v7F0ePkhs6bN6yWd3kWmLlFWaL6GJdNhSI
hFvLJqDk59/ndx73TOfoIACQzJT+14loN7MZT1r8DUhHMvWdlixnPM7kycwyet9TbGFn4t3ua3RF
9U1jlFfaiJO4OEF8C1JAWp8qtGGgCGSALxHjwOmVW7EBC/ugRD0npMV2eItsSOO4MRdSlu1gRcCZ
N8Kj19oVdBTQbZh56EX9qqeA6YmGhWubMDUhh5tvjmuVq5+WYGVsWyEcQfYmUR8/CWVkiEy3/9+6
FG0iYerGRE7afH4nxBbB8UzSBybDoLKi5rOnulXdiXZaNZRA8DnvtPwh2jkktPxUWKmC99u5fR7u
qlHbz7DDhzzG9ID9jRUswzUZlJEQZ1LXyAlmE8S68QRU9f+8k4k9qu8lAyyDqYHprumb+eMwxvB3
DggJrAPECFjvK0YZEuUIZESeFJseEmWp5/5mukxl+hfIo6JFA6wJUOu8llh7cvKE7WI/mIrSKDSx
ACK/DzDv/4UFdoNtT8+1sp0VG4N9U/YVtxJqgJuDU91n3ytdNM5/JzjJRcE6nxOSXCu7AyPG3HIm
HqIaOvOfz39qPXUYTCIF6Bx2rrE+CgzD1k0W54ngWyp0Q1iFqaWlw13AWDe9WhPL7LqEnzkOvg4u
/3VBr0YAZybvlINCXN6dZaYBuv0BG8HdL1DT6GmbQYCt/hffiKkkq9GOnZLSxHNsS30ecmg7e1YL
LpzTDtIu07g31+j4HmGIRSNEZkWn+w6TgsC853GvEW9m5/LNd+2qc/RLtIqsAZmYMILOM+/QmfAF
iWCQsyh4qkfaEIOzkoJOrb2O3Eg7mSNSI5/SvCtMWNgMHDGE6xnMVNbiJbSS5frLprdlpNxl806x
tRIVr27vKV8w6YjgwVonoVf6pu4cHBtc+eLm5mSNDuuuEN2qNwD80GcrVnqUaPjrmknVPMW6efzL
CRJVQle0oWx+286xDxgYlYbFo8eZIX5PTw4BxlwJjJDOKp+qLMYKtlIhMT+vKco/pexGmUhj4Jp1
r7QH/I/rcilldnmQbCiD/257cKgZhrsH/48X/1xIkH5ywnuUX4MRagnvhtdUWB8LkZNFzEml9Gw4
HvKDSyMYBegliwd1pZtE8z6bOg/BllFcYW4LqIv0z50oZoXp/e0LZZKSrgeLxr3TYklm2US1uc/7
1CncDMmY0KJu8yo/Ny5AcLeAAr6xrDXOxdDegKxtXZRUnHOoYb5YpzSUh8GATWpkKToYRYdnPnom
pd4s08yZeF8U98KOvSoMlhzTC885ValFwBAZQN8DqiKFdnVZ7GzT1psnCXKHxbGdpbFvQFSOX0MQ
uofdzbkuLkyCD7olaF/TBakOcYhF46CgkWiCs2kh0IZeLKKtAPaRtAN8tD8ixhJ/b9Kzrl25RuJU
k9Z7+TaYc0LjOQOjjN5tO+KsCG/E2Jy6pUfy3qQHSb+au8qIs+ZhFAjoSmbtbAD+OCijmy8DtyTF
F1QJKpPvl7vURE6OFC0y8eTVz1f/BifY5Fd61i/UqjWeep7oq9xP6go/vFwWFYc9EVCA54nPDN+r
WJPm5mEGDXlyhhmXhG4hT6WW8yPdefmvb5njr1eatDnxMeFG1h16dro/NQ52wMnCXznuZ3tEJ3eA
V2dVlCzwEeCPGsR3S2TNXB+imD9KsI6oKTdyOxcXlTV+bvw8zsK2/FJn2Ly8sQMoZI98zJ4YwoRZ
x1/OKyij97BCeqayqQOh0qUWOzTjtO83PFsAsexJ8d6FZfh0i4QDgaZoFVFX5qzeEJyPZuUWQGfN
QU58TpDzw2Nb2wowtLLbZsZhnWAn4fsHoOWeNBYppe8m9hweN28TXRuHErEUYOo0OhR17YclfbIn
kSQzIggZYEzaTXVYJLD+Tf7PmS9nfqBt6ixZtYQRuiNHV6KPOdC6NyUKR6Yf+g9UhieOxAZTuD5F
7dVuG32RGRAP7S8yv+sHx4ip6QqCYuIOeF9EkDRH2rIPjt2TiY9X5ZFKAN8QGx0U6uBf+AnKVmsS
KQSMTcOIefijmYwhs4nnCr0qbWRhdfHxO2AzIb9+5UO5pGN9P0b3gMbT0egBesJCriLxP/QvjPsb
GpcWBQ46Y1AbiBhtBTdZn4eHhpX7bXfpRLws+hkhjTJdhu7YZKR2ZceZ/xWnHjBCT8Y7du5o1EM6
6WC1aSSqA3OgpOvNdwCCyKYHhXNx8VV98hZ1BfozQWNHbszCuWbU/o+WRv0j9Jb3QO45ViBuUwbi
rBEnBcYi90jLFDTeyQYQDLKAt8/WVQDXLLDLGdWb8XBUNClzbJ3B1GsvsgNt+ttU4L8D1evd+WMr
RINK6R9PChRgJiyNiUTAdhXG/t11f9yhtQRGgA1c/lC1aeICWnVxf97bFnv73BrVItIBjz7F6VPi
Hfa38anmahWjScY1+ReCYHkaKbz/FfysnQ7BwK7EhZslAJTOP0p5xyjkAz+wfhM1GKaPK7XIcg+A
THhhaz9HZ3kz7LQH7fMcjTpod4fMB74k5BzJwYJfGARvvOA5D+nAqITGuCTskjUD2nMeFImHSw71
C722t+7YGkjrbArg6w2viJvUAAV1BMMAzCr/in1LBCVtcsM9yP9IiOFWPRTpzI1dPydQdcO49v++
bbVRfd2Hg/VPMcp2G9UysQIkhWdPwa8xNwLsA9KE2U3/LrM9xx9WGDiWpKxhn1Vg4P5h4YutoD2t
z45y30z6z/sIPLpgCQuZ8rZnS6ZmE61TjauUlufPYQSCOGz/wKiE7/Sp46epE0zV4V2H92gUevZi
6NOEm62trrwm8/SYaWUkr6PzUVMVfq9jrd7YPKuVnUa26qiNHWRiS9z2ofc5oycG8oBoF/888WY2
1rhLkyU/Ij/zouMfsUNCDtF31E53OIYXVzJG5IU1SLNattjI6kk6m2VeVYuJQ5XdJDq5YD9hlXJk
PdZqRvjAF0FtSj5e56Sauvz/rZ7I0xkkL/IC13ZV8hC7sjqK8T8dsOMwLUdWvxoV3PyACjXyPJUr
4cQGIpXixrxPuONPwPA1kICPSEaefmLT+GRciJ17lLJxEsIdFPcWMPfKIR4A2jwP8fZLgcA/3d4x
twEHhF6Nf0+fWdg7vu8x+oSL/MtT+D5L+vcOOE85npiopftafwdt6hxOpFbc2bAZTzVdFJPJaUar
0EfNvgCFAs/F/7BMeH9VlHG6w9FvYRTay+SBer2MGPBJJP9GwTusbTnLs0qW21ACWIazbyNSOpLn
kgxfaPAfRvP6fSolt/9JqMWWu0px8C4fyp16hH2VBr6cKuacn8oTkXOJE/CNPwwHsylN2OrTNOc/
S0QuRQ1Ja3oDn0xyg+XrvsuOO9UOBuBK6AhoLmV68fvHDAnF+d8+OFYYb+iwyqdxY8U/NyUr6g4D
ScxNkYIRXfX3E+nql9dGcGqpGD8nrps7GB2/l/uxxaYyc/m8bTuuiCvRD4HYuvuJDqSdGyDwgqEF
wNvwehWyE8+97HlUtXamCCO+rmnjMX5LRUCQj+rX+bmGFMkWBuKDmJXJCZg4Jfa/CeHxhHT6M7cB
RSylQoWNywqIXzjA2z+S7t7ntmwiQsgYAgYPt3te5xUNlko8xJr+jdA+jSuEmxMzn4RIl/jZhRic
ZE5WnZlpJWfLGeS+cpERBuKrjgE79GYuO1VXNYHiIg1llbXERNzSfyvTDxA5VlZpZEF1k+09j2yf
sPtjEybZzduP80/iWq8YJXY6NsLZw8S3K4pOSJ9jGptnJJ1COGiFhSY6rzLbbozAA35fz1ll2kK+
ZqbloNeBjRYTV7B5aFZNhqurgcMhvldfSaPtFK649SUMhFXI6B+wKMgLBn/3othOhuXKUGnjKO/0
z88o80l+n0KkiJ/trYEVvHCAfSWuHvEJtb5f+cqkHT5lUIj9OJOuAXqfPB6824R4iHcwtjL72Lo8
P3Y1sQkss4o8YNWrc3vIlhIEQ29h2FFweWVvHB9Y5fiaXFaed+L/ayljgycw2vLagdPj69B1HTRc
dTDqrvxYyG1SSSC0Cwd1JlZNmRU4564mKPBbWHIaRN6jBD9wRbNdzddJorTTqEommSCwBdEOwuYW
uFvFGtDZ+DMipN6W+2HxuNvYfCt9ur+xG4dScPx+8zz2LMSaW9vWDWYywAmEqDGcAmdvDJcyqvsa
DAUfz4cwcBmGoRPedp4wRZEDvaL2fKtJA6Rs+KioF67Lj+/aaDM11M6Afj1Cf4gF/8iGsB/1Qbuc
L4EJigoG9Iex9lDxUAaFY156b6115UikjMRyfELLogxBwBPuq7HG908qtrI9Yx2wy4n/2SwW/z4P
WdzDNIXdJozHe3P332dtnn0tBMiJqtkZxSh133EQzTwlpQ8Yjdxtnqcr4VkYEr+oUG09FpQCP59E
LLY8ytVD3y9xgtPdsqVL4ZaxOiLZh1405ug752Ih7rqR+vaY7B4gxPLeg/4/kijTltLta5a6h9rV
CQo06VDyMgTJpHIyl75VUa2L5ry0Kho/wzSYfLfySsNAfN8ad3WJf08TkGPuStdCZY/kLlBVmsek
rz03BtOAl5S2oOzydEOi4ywGICLa6VUWzCRtEgn3qc3v3sfO+NHVt5fSub5ee0Jr4ekxjxeEBUn+
x8Mcskqam1e3nJc/WbfZPW+MRsxoKRUWK8vBeD24LiuKfqjfnxXFdirpwvaHEauk0jAVk1sOL3+U
ziJpsrHR2vgNkyaxAjuGa2FXneRyF/hO4BDceWVm5m5J22T491bccYn+WN3xmchG7xkGLgVT30OP
Le/NuUOuwUGm3XtKxABnpdkUBMP4KIFGtdhX7a9KoSV2vPKhjERQV1UFrm0jz6MOisOJ2FzGeGyV
8HVbv+Gf5YGt5mtLy6sPUyernVjYAlvWaqn7ED2VRrAd6z56WgLI59KLIx2BSK32EF0i9vH58Jsx
neoB6AJX+k1jXe1pF4Y3PQTZv9BeEpeIz1FnrjL85smehk29f8Kk+tQTVEQWexmrXBpQqQV6xy23
gLA83f9qD5VoHHooepqMLrQR/BcjJEWhfl6D3j80dY3ZmggB1tUBybNJnxst7QIfT3DiKsynZnYA
Sc4KmKAnUfuItWvFoDeH8N1FoLK+nOQNN7OczSGpFu+dEKriKOx/GVFJWEVVf2hgm8xar+PERJ/C
JuTN7lmGe8+/LHlPwUA3zC2KdJ8ahHd9sdjRaSuSJEaZkBwJVxhim/KsCt1crGF+4KRvpSevNA3H
AQteeLbkM4n5X61xI71Tlg2pZLfEndnEHUpxYwrRJMv6ivnN1ir8oLpxGzd0spmDC36dRwdgVYN5
HeQYQIPSemxl2ZuxELn4TPerwdEH0Z/k9wSRiu540+2xjsanxCh1HgU6WkdDZ1iVwmvBNSZHmD8Z
bn2h84HiAJ19b2lDKUgY/WekiE8AntNNmFax0GFoLtnmXxHW6mc3ApRtzN4JhJnB+JDBpaz/T+Ae
rhGlBPlcmBO5948OSW2ClehtxFojwQ0CDp3WHC9NpbLED6SpYkGY8fbkXg6kK4aj6W2LeOxeFqWv
GiHtAbCS3hEGYUO4so2cUcdDJq1Q8kiQgVhYUHUhhoCdBViegyfpTFBfVJbPnCTkK5j0NhHWqR+a
a+wteI4ll4QD5H2E9LxfRC//V4pJeCfTnwNnd2ti5LFSty7rHlgxD6o9ahhoU3RERPUioVAiT65V
66FNOil7Y7Jgpgfw1MyTgFwoDsp118HpWWKrT6rAYLKjoWQVkEu2a/uh1xCn+8xzFQVSZmUBCmmm
AQKbSSoCa3k7tFlweIX6DC6wofTUgKi6iht7aG6Pl6XhETpU7tu2jJeumF52LFzBWd/zX7EVFRk9
GKhvVxdddPJZvQz5CkwJCHvJofFro2/bbXWn5YmuKuwc/3gGY0p28GFdt8sq0TSzsqZoeI/efCKk
FRBnwLRCS8lVd/8HKIsyI+RaryfQDybFQ57e2g8M4Cq7jN5MOMwhrktjqOa+9ysZ6MXSeKqzwKND
AB94VsnnstlXRmaS/SvohHiixaE1ShhsEUmYnb5uayGkkTFa0jQHPa9lnFenPBRMYRVdTA5FmFa4
+siUYcbCCdzywOte517ZpcgDv6FNPmlPvHpnMbpBJqfLt6aY4FgwvRihNzJVm2NfEVlXOEbHOpp1
mLSOoCV3CmdZK6PUugkFDoEK9ZhnLqvsWZyDwND/nkranIrLZ6QZ8KlqShtkxtodadHcT5z19emP
+SuUCvlQc6dDwBZIkiw+HXhiMaeXJOGvYAwXzlwxB4WSRTKad/ZUmYYosxuVUnYze9Lh7b+Zy5uw
3N6O3/m6jkSZaFRi4/i6XmmChNOMUlwFCJEQnuJRTMaUj8jz3liHFFFw77Ka+feL/MehiLboNycv
CS+ui0RMdYoJXdAsJ2lZO3d8J4Gnd4/0Zs+cnGk0WpVmpBPjgIeygvxsnmjIjUJmcbfqsVSkmT86
oAPjbnChFAKdR89JZJpSCWUVwP9b/wiE+h/imqDUAUtauRU837ZTMnW1arSb1XX8NyvMgaQemxwI
wTKx2N5Tvu7Ek1wmvnhyyE/0bMHMjJ34QZ+8QE+Ik+dZn/aWU9DeK8iLQaDoHOso/RWm8uoEBP2l
e+Wrx7FZuxVec5ED5ahUGmzy2HsyLnpio4i/zPEnkN9Mj5ymzvVRoAYfrBRrj3u5XLbRkucmGEy3
uTw16X/fO4bOzX34NN9QXXCdyVtewM2piqckdPHBLHMLCHNAiIAEpJdvVUO8qo/qt93whuFejnaF
Gdqh4+HNx2/6IHMehM2Ug9QMnqYU4FzgJCq+rYLQpK00YrKW9/LXGozKHlSw43aNISA6l2wPuqgF
ZRNVac9K9ojQY0lYRdH/4in/usC75PUwjwF+pL3N5kJhpQpytTp5EUrblBSRwFDudNliUPws2P+b
B3TFKxjbqv2drSJ3is8YUCmo4RAqyCfvamOfSGF5WQZe4MM0WDVS9sUZW0zJp54PTg2MfiMdYCx4
fcCrUNT2YxShqg9PAGoas4v6ab08ZjROaGdjnl4uSrFo4W8f8yzgoOkOqtuNE4eb/+bWYHJglOx7
9+QG5bnvTQjmscX4Hc3n0/50xbzMskvmlRWOMszoHcTTpQ2pXSPPv1sdvC/dohowiseFnVqM3ecm
SEueoNAXWEsJx65OoquD/H81idrPXj3ROOmXnbsOCHYJ3+YVugPvW6x0YGHHyOoVYTiC+ZTJ/1VJ
6CdFDd19qmpZ27k4C47mJynJtfPNZUyBjkBclHk5YttPKdOHSprBNHBsSWAkT1wg6mBi/85JXCCb
yq5IbwDhPpqnFxqD4Jv3fJCI4ZH23qrZMEw/o4Ql4uGEFxu0EmR0JgCcORMqj6xZ6sksd5+VCgbQ
tO/TXMTA4ikImFkVaPuvadqRX4vZ+Ev8fbC5FswNRtIIvXxWA2Kmb99PId0uMAU5euhnq2hwk/XK
3lf/a0Fx/eB9j85CBnlbt4BIrn6Y6cRPjymhILlZV99P8ZpLAFmmjduFYTuCW8pa6Ycdfv9HerVo
SJSGdkn10H8VyCBDJDE00lYM4TbZMD06Zn00RAkreakO/2IbzZZhu3cGWpyVV4Pc+Y8kmekom8jj
Mn7/Y63LE0lmY57RFKk8uUU1xDJCQA4gZs0ZuA9YDyb2OKi5QjRgw/DQepsd4nLVhpV/WSqrVxs2
CFlh0kO2lo5knIlDQEopmeSMuOiSaKH5qY34ByF9IePX6reRoSOUW6YWp+PWVfUjQ8HsPVnkaMDH
o8BFct1fwX0qnTlCokns/9Z6QeR4j+yd2GOu8uxhNVhLgXmbmrL4QTpKHwHDdwkHJQfdHVBPpSNe
VGDXn3sXpO6SK8HalcTzvcZlCIVUg8Nq09AQU1NZsGwBmnCVFOt7TA7g1jE4fpMOXW8prNJprqru
U4CBe3Pv4b2+fpqyeIIdpM620VpSYwbw3ccteDDU6cYhIxBwBv+QYTT33yODRn+bQp+aeGQUSVFP
nT6KK0e3wc28/bH661m1i2zNdMEpCtbHsm1oRcPRn0YZ6jmqfBhIfSsFkXOXXxsdUBQG5FXwxE4I
PowQXn1ifQFx7LBQNs3T4uX6/NLzwHvls/vsS9mMZpSTfMvDt2xH7lXtfxZRJ8YISLXZUAjLMMpZ
a5hx+syt9oP5RpqBHA/xlBu1ZEeFBWWtH1cIOfhF8LohGzzeLgvJjp4B6rJy9592s051BuNJE2Bn
VZhZh/yLeQCkcf5t8w6XTmU415paelvIMVRBclflT9jgc6obhPMuXYVpz/s5Lqo+mqpBmiiF2Pv2
vHkUCYkWuJMUr7X24PFWA/WQx8dD22zFydOlJqEqnL/F7aDAH4/wzvj5sNODkRrCVs85ryTrSR5r
mer4FopMm3LREQPMrK/5FVg383K6KTty4y8edcW1vFbG2Io/6Bbx5w6OsJMFSid/J6nGymP/YYXy
IZUi5O93ZEzEYorq/jLDD3mt/N5FaD7ca0WzNGXihzsLWlaf7ohehjBtn4FTCc/KQ9YW0SBHxwB/
0+7o/cSkVISbTdUtpoaQPg9AnVc/UTgEn5K5lKtj4RvlY6UfGD5pLlu+q9NPL+JtXhdXrodBjrmG
vHcC9SAkS983TzIQnUmtW8Gn87mZIK6v1DtOeLLxSTSIF8JaSo4FgWrbXQOE5RABSScM0aHTILEL
GJbo2Uj9ZgWUxPjV57XhvdIVhpzBkVH2DVsfndkiqVLiZZTvfTi/c9i7fzBBQ1xHHe0DxZ+BuuwA
9/wsEgNAGo7BvWIqMGAhjBBMzWmFk9TrnrJ+p4kY2K7RyEo5e/iwi/ofzvPzqOSo14W1fOErdwKN
rzZ8gMKvnqiu1wJMSax3vF7E7AS0pMvV1YIh4pKfTtORPF7O/KgUhEnyaPxX7htsZL8oOApUxjm1
YuCg6+yyMpPfPPRpp7jiV7YCZQGZ/6ABLS1/GbgK88N8CXyU7Vdy6nNNdzw6z12M7Bfd3cItV03x
6veXldJBWYOGwdAfwkzOzGNNhO+PSDMuVagVkyTSrhdU2uNqsKR8Ti3lITN+1NfucJMrkro7liDN
nDE9zsGXx2L1scJnLbkn7xZYdxQ8CGdrNNY2N8A0XMZCgYm/DiXtLnvOGPjl+BWGGCpVd9e0bb98
FecUPJA4wgg2VNfFVRcFlvzRnaj7nPZvX4Hfo1u3rLQlGQR/N9wNtY6qZ98Lna1/0I6zKBsZ6hwq
QG5pzf73FiKPb2hHEpR2Uagr7OEzj/yWTrOC6rKTb7N76D7cuf4fhJDicuFQp4RAwQNKaXCQMlrM
R8u3naPvPVwvn3+aBIPUCUHHx+mruEPxDDrgyo5UygpII4CTBOCSXswXLyoI8jyiQ9Ct5H0WmSpa
b9IVJG1ZqShr5OHVhWc3jD5QggFTu1TJw7e2LgcMHnEji5YOgZWQoh7jDupDzVLwiysLgk/OdVsM
b6728v7lfmDdE3UpwCYp3eCi8zSsNDRT5dRIBDb8+/SHEvDdYuKe6710eXgI5CUgQKjHwQtz6WMT
5IahVnCHmnE0Kb85LcgZX3tmJLq2k6GncaCja9K7TuP52wOPCn8oNXiy9NF9F9RfiLYh6ZxP/nKg
xLV8U2an2c6Ufrm/DMey8lbJBaz7L81liJ/ywqmGSTB6w6fYkistw38N2tujFVOMubcgIeo6kllI
BSUBEO643KXM4dqxlU4Gonyu4q9IBibmWu+MC+2DNy0krjFYiAvBNrQXTu632eIuYX1WpzwqjnH2
YG64U920Hd2aQWNv5bOWlgf8xlPXYEsCOXuisg0vBjImSiS95xcPL3Cq6HsXVHYjVCfjeMxakWFw
Pu+gE0YkR/pMg2iYNt1L9BN5vKjI17CppunbOPadf5F/gwAyzOrYkIJsT0rmAo54uM96vZPc3Yqf
MqK140OoIHZWg6C6CvaMvQOKnYq44m7tcWZHozjCCOZba9YptzZ+Mg+KOOXVdA85XXWCPPz+JaOo
cwaetu9rRrN0hGtYY2UckgYp/CJ57XG4ZuI1lCtQRzhvdzlX26rqHPbgD/PoxaxFJfpOHRCdXkkA
iFL7teadi195lHEo6dhF6skFkQVnMB2sa/B+T6YrOpzGFQ7KsLvc4qDGD9f0WezOSYBEgWT6Bdpn
C0XZuuddn3HLRoFwAwR99jpf4CdAUjiwUfs3O9cVdpKSUbOCrzApLmGpH5vMP3SZ9usO+kmfdd07
DxCGhg176TsqGtPwHSNbqNhBrQaMPElgt6vvADRp+y7TAVF3HPFjxB0pedGeJdhw+Wd4v1am9npY
wVdibL8Jc9ifJwFQBBH1bjJqqYrjNHtlfSERR16U3v6CWr5J0f7ahkeM/89HOT8X/jwG6Dxitrp0
J0zHoipQyPn/3NiQEk0r3QtAEblXJl/7aFWmV0rlSAk09EGgTVGK1khxVhtKvk7wm7l4rzD4QauA
QqATMv5Ks9DfibuR2D/L1L56IPhZ0HTc69wIxdHd72XNSDd9QkTnKrnL6GyElAYFdk51szzxXfrj
eD6pM9AhsZzjisbQWJMcZE6w0DR0N68ZCd4qAsC7nbtP3DwvNmNPwIUrJR8VsDOwQKzR8zZN1+En
zvhhzSFsxlXFQp0JyU7Ki4wrTxgjbIvYBUcOsrEGh0vy3O0mgYNeHAbtmIpnzJiTAOG0unRskidK
mggMWTIX7tYj/AUHQ2AVZfkrfzTNB7fZ/EKCndYTq3ZVjopjgP27BHqMUMtb1oBiQsD9R2EMlgqD
gIaBKNYch4ZlFFMxYtubEmB6RoLAcic+XmyfoWsO5YEokkqH93PDTzzD0vqbMLJyz4Y0dov+btnO
BfiB6cZRHl7fob1FpSsU63CGTHFiaOfdfqh/ejsAOEOFszc6W847zbASpqfyf6S3jWCdEfrGaoAz
5tJv69QPP6PIKB2Kv+FDwaWesSAmEk9g3OfAFYbhR7L9/5HybSpb0m9QxD4bYSrlc28t1cWL2Vnw
LmPNru8eeApoV+IVEfaOwnripgawy2PdNEWDnYakeNqvoMdqthY2MNrn41CF5FONfRFIOrR8e9GA
fTbWaNUCmgd4nUrZgEyjxp27wYWqbIhhR1ZKat2wGU7q2hEIRX/SdQMQkFM3MliSPivGeLM0qstI
1Ac8mzAhHfPfF9IeYpudQ1bg5MoLex/sPKY89gcd5aH9Xwgk0NyksnPnjeXvAhV8gXZF7dUkmP7m
ptcaZp59xhlVmnR8xsON/5dCYSdBkLxp/Jc7d/mWizWlAKUBVx0e4ytJOJSzB0Xd/BlCFhktVRxs
Rpuzqgp4WCSQVE56Sijkyg7sXrIQafpY5MbR2de/TuvY/oZ0GcgYArYP4+RhqoLgtFzSnMgBPqZZ
TleGdaftcYuLORS3Xo1NsOcu5ATLdY/GuuAdMgYFN0XtqntzSRZQ7M1LxxhUQMwN8ishxgVVvg2s
z2zBQw6s3/DoqyHILLDohEQKIZrEJmB0KVL5GYXhip65lh6mAdKII5dLi5aohz7+YDLHWkOOPAB7
syRxV9iYO1FRRlM5vR8aMOZLg5NtpWONfEIxus6isMZYcSrw1D9W4ZNHaeniFLD1FWCqU22xWg9N
KiRKMzxSbIGYL28dN4IelPVvThhcIeKwWV629YnYXui51dnMYsdD5re8OEAmz6TZm486RmYHGDRM
tRGSqxUYxu/plAb3xR8pltxKdJioD+kRxC0zngr0VKkuphdHS37LJ5u3hetjfF2xZkHM93tuP4+m
ZEYeCMpwuPQ668q3oPFkSQ+4iFRniHyzEqbKO8nYuNiwRg/asKvV8Aj46x4QFFxBAjirZAb/CQH+
1ZeBJKIo2FF058a5PKqpxBcaNPhtarqaD6K/eQC4y3N8bcssqRSJ6BSqmOIKZieAX0JWSdcdp5yG
ayd3fohfNo2V1SLNJV3ZRt9UR3X6NCrn1XzS44c6AdX+63HVNU83Qjyy9nNHk1ZEfvnhxlzkmpXi
Gzht7rvwlZ8c+5qOWLZWR35G5fBPfVBrwwBX6PGuveCLB/58fbQjQECzvGbfFQf1KBie+vMp0wiR
4OPcFIfCOjjdoVWcelubuduTV/IBiwPtD3L197QxkGxJsIF/b70s98dz7ZyYJ7QjwFVeH8xqvVwF
7wXQkEVzvxRCUBT+Glupb2+jz3gHy/CXWawUVoihyNfgJ2GUQj8FTo3hdwToKt37Jv4romGppMaA
KQLsApxDmrbH3MojnmuwO+lLatU97goHX3tdiJjiJaw8NA6VBhqju7aOInGOxOqv13U9rHwDJJ4i
JpVsYoFnNK/VAicC7GExw/M/qZPQ8TV8Ra63ol3DiBPRz2ozvST05xWLUlQays6k4wjS/i7U0RYk
l5w1H9CEyD1n24jLvcj2/z3EKaOJB+6LdlgYycLoXdDGdLTy1bAcrDC4zixj4PUoeJI43nmX04IX
4fnPZts2SjnpVvb+C11fY4Bo1PY1+NeM7/7a2KYPMdd1OSFITx/XQ+2BsyQvnj6SCltePYZWbOk7
sYMX0EmQL/Uejzn/RoCKGoE8bHjGS0jl2rIvxjS1A6s6twJxfFNtLt8L5Afv3qXTOzdEIjMcLuos
i1GkeCBtJiqtYYgw5pFu4zS4pLimYbgrDwqdNifiaI4gFR7Klq0Jp+3kr3RTtsrseY1S5I8xtud5
D5khCMKTT+p9r4NpN3xeiPR0trNinYjBSa93eijyvGQ7KBnZbI7Ov+ccnHdTjrYdO80eB1h2/qid
+ZAmeCjzFk8zIuMgGCjNM5pUv81rfmQokAktpPy3r+HkyjlYgyNTB07jZfpOjdz8lMHCIYKorQ5Z
JyE9GHXhswhP5Tn/3j9znQdxT2JUjBYHbNp4PiQ7VPb2X/j0wc8fZVDNW88SKuL5VWRdzkkYTIGR
lEApdkDeahB/DQfaFjnFrLZM1jqTJsjzkOtotTdtEMSBVLzSpxUfuSoZOkj2WkOzbOmpTjhRZk4J
LHvgleuwj5XBm0hipnGSTkJyp96u/KUXKUYrKorw9jdJiOZ/DuHAiK84eoPUGP7i/PSLXp2uakGU
dRibqgrYWg8pXKsTzZTHGc63i4PoTJamkK0tqfIPo1D3df96quSNR2eQjcHRpYnR9YNtp2KO4PU9
zcHJdvMlmkXkICKJB/0sEQptYdA8eG0DTDzNZvEQ3wICiJO8GjWxIVXliCjbNmmpedomcEN5w1Qm
tHitA5081LutbY6LWd/L3tMle1b/HZGwHZZEgEH07ag1l2q1FtKxRoKblZlmCPevlIiyl2MPxgmu
zFuvvpQPD5vsv8omU6Ym/UO76R+QQQt6R2o0dg6rF3e49xo/lQJmcLSmUFrGAcC1EWEISinqizBZ
bPxvoXCvl4BBb5bIrBdJYvUdNvy/Im9FLWLAi1P6TybTnMOu+cXVrRKFkBzGYhHbKnR8RSnRyvPz
30dH/DMwQRwKScbnAzKvAi0Zd4kxtfKXRs64irFWpuqkLGd385KKcaiCb5aPBe9dr7UANdwM+ZnX
zxOjtqfb0d5F2LeTiHy/c3enEJFgEjVtFjqeD5dIDBkEAiphFph3fTFcWsSWqZhuo+QZxkhXQrBl
4fqN2vx5fN3fpYJ1uiEgP9xic17Itsyd4yt9Pl9yIr1lWQ7e4MSM6gfhYS5rlPcqqzGpezET/RXn
tCa30mhEr34GZGFYD4BHFaqzLiMWFFhWf6m0nxGbN9Mt9+q3XSdFsT6l3gO8xD7yXff+sxNSWxL6
oMKwIB0LaBPw3x3HYleK+CjcY6aKgaK5q4i63NXQf0eFrHetsFC4XRgSJA+ib/kY1LOg4oGMBGEM
SxWeROpy4UtO1dyngv57wNgbb3TelpJ0D3snLMM9ySwZS6c0FWYKYqDuGBpcsvJ6ExN+Sv83xCgH
5aG3AnYZUDNMw/W3b50xrL0HkmPVMB7j6/+WC60dAESphxIW5jFFe73HoDUjxYO2LhILskwE10QY
p7cyA1K/Hd5bEVWBYh4r/FgGFSO86hmu1yPYtIeC+d8CazHky6QQ9owHab/qP/0g9ZwnQ4ohTBQr
p5yro+qQC7fF2rF8zP9KFsAVPM9mUSsdFQVNORpOZygopeGs5+gZSWp7S2wnmJ5EESaTqW6z5nmX
qJaDyh8M0dsBjxtUpon7Mh76SOyyEaN8UeATU9cxfK2BW6HnD77p3bNTHjp5t6grqmUrq1sXkq0F
PLPRKz6pgFYf2uGufyF2rVBQ6G8nUNYrirj0++pfDC6BgK4dEOXoXk16QUbexgjH/lTm2ovAtblM
Zp7Y5yOVf8IBn9CCcuwFPk3d21CZopJ2B9KQVM5qzVJaChmD9LHbkgKzbK6ndYfy1d5W6TcOkJfb
7gqEl6jUsjngKCp6a1uYxpJ23aHJG18Q7UsalgpltQ/ULtLFfs7Tusi7WzvHKnY8WaUt1jOjiYXq
DAvStgHkT7CxS4xJKqOn+gxbMS7SGYYQku2RyrSZHweDeO9jyGkoi84bNb6kLvB1BUxRXsaP2en9
gtd0N4nFBD2iDi9OkZ8KLfQ1lI57U2T4ftXTNwzsC2De5xC2QLRSx3zTCTiSuGoh81k6MtzSPLYt
5GTKdaemvMsj61otmVlSjobzoygkJkphgqjAwHWLLQAfYAslJEEz9vJibKsNXGemHQf0Yu9sOfww
xOuuoyzmkGO6w/XXR9QeNTUNdnzNG5mzWbPtz+pLrhQT246QRteGLWMFQHyFOcmNXAb34rK+kIzx
g+B6ZdxCNfAwGuvuRjbeRXQUgFTS5tRocBP8SECfyDIYN6oBf2xvZNBr1+5BF4Vahswen4cXaWBT
gp4GD7pVAzxS0abhMej78Rl4KuWuUFRWT6GBRP2Vq/sHa8ciATHl5goyyX2pjH9CzKU9tt6qN7Up
M5d7wmUISNePz0t59W/aDqPKdvYJ6a6AN4vkJzijLj3pIUEcQBtXHiTf/Ejj5M+Bh5+L8SzPIaOl
1G9c8R5TV5u2qFUTza22W2X2CYE51fYhsXqTCkUwHb64tv+iWcvi1Vlq4lACkQqPzbPjPMrC2GAI
y7x8fjAQO8bHHRjM82gyQZQ6DRyJi1/KdolC5mml6Gg2ZFbV7nXEClQzuNU1+K3qvqkNvlbrM+eW
g4KsBeyb20kadG07J2niYmX47Nix3xdaPs6t3sHiDOFi15r4+225xv5kgsDpksHSc94HOzWG4Puv
p9miaCCLHPoWn/2vPhAZmVsKn38Qw496hgp+kaEIwLDdkNMt+xCOfahOz6mZBOe9IHbrQ/NpRG/B
xQgVjk1y3CIv2y5Mgro8XxAjQDZl7Whx8ByARahn32ftwslvUZjbqxwtcu0tyDUPocIl+p+TGGM0
/PIleVOharvI3ZU2SlaX5xy5Mz99Ta5Xh6zE8fsw5WYTJ6+n50MO5Qh2yip56vPEvQwDtnJtpOkO
T80Yl1JEDU2HAK5hHK+gGn8Xns3D4qIzb2jYer9/58TglofrH9Gd0sHJG05Vi4Jw8S8bloLWDGD2
njd8/NNHeusoe3ZHhKqlfTTsWHzZW/M+YQmcImu4WqfjlF0xzlQPxlx9yePlYcUaeYV9H/Td4TDl
l6he4RPPHnNC+YiHI/9DuzVmWHTxIvtzFhhTbZtz+UjmXYoijmJEsMfRfRjIBJ0GsmguomLsnV1c
DQu2JFD6n90AUmRLkmj/F8SRasu2KW8GLzOFBEHDjIpn1KDJ1V0BKTKXBCE6zDyk8Ml8ih9XsrK7
tZgsziijn+7CU1Zr7RsXaJNyLwnZFlkcf3wQBePVH8cKbNS3183EsFVKaSmq7wRunpvkMuv6XqyE
3DxnBhm47O0a0YMd+8QtjIUVoCf90fj3wnoCHOOyKz9MZ3Y9AHCI/51Doujo6BJXKYcigqPzmVFV
hTWYHYbS7QyabLMBycWcJsqpwlKsHJIamoz1SbNfP+TtEv+saKqiqs9th5UreOrTokw7rgQfk6kT
N9w3oUr4iprdqnuCx/1M1iSSV22qCmjk1zMh9QhcBP3ipRRMM86wx+KXlAlFSPgBeYjdPtBJgc2j
ss1O2x7x6a6Msm305MjHLZaaUK5jNqkDy7RN9j3/NsvBm4APVCJ6vOgCuGMsDPVqVWf0jtPaKk5s
klS0oShq7aAeouWxmVbDztU0XthgZ+lRYMp0ArxxhZHgXSgxN4PYPahCDm6+4T/3GV35DodCSds2
eAAi2hKbXaJd4xCb/5SoG9QUuuF9I5cj8o06sX6GVlhPTSVtoi8KB8A/c0FBDEhsDezY/qerxK0p
yehFxfk8GhPRgGe6kRjfcypQgOcURqxFGFaxnVqdKPPclnr4YyTNRSm1l5KHcx5YB5/43+VTBi75
tnk12rHinotOL+rNT/W53qUjdv0Fh0ar/PgqrPV3cwUmNv1npY8gWBR8OmamSOpFumrIii8Zr9cq
++jmcn4nm8/md6niGcSkGjxKfxvBjtKP2C4pOiMbgr0yJZ2gR/06UTqvtQnZUM8AN6ATy8v68FS5
EZAHBuzwxVq4zoJ5aup+99uTkehJmfH5JRe40PujwFUjTMKzi+0dvI0iA/sXJRFPL1pCMzlIlmGe
NaAfOXhbdDZbcll3lgYA6GgBtQvdUFVS8EPbeogOYRMyQTUc/tFRVZMq8e7Vbt8Bu5ZvsMP9OnUK
Id75/w3QCwc9sRCUQXaPywOU0wEiiEjBVpd0szNFeQd5zv3hodj5D7ybeNbRHoxS+pyCz9hjA4cc
XsDS6sftrLnnJRWVVjg8pF9z3EFMwUMTLq27naOA6I7sDfJ9XYlpVq6wK9cdKIDEbrqVyEctpjWo
s4l1aVf0ZdaIENkCa0p+IqCgloBbKPeLV7m1Q/+6LT1+FXFMW/sKUpG1HcP+2yNckpQUK7SRm2h/
77fbTpxx223H9fdtu1Sx8VyBAunjv1L20CO8TQFo80B8M6IQj32uihKI/46qLjrhobsRSNh6Y8dG
t642wxpWZ0Pnp/PmR/vHVf4A7LxqaLrF5YwVb51PQHxAVFIomdHg6oFXV/g5/lTwt0vR72kO2TDo
4evfBTjLRfK4XXdniq6F86PVHkMaDkHKkr7k4zTN9lnznHQjIWR8ikPoKpMUlgpEytrVP7Wvg9Q1
Ksgzg7BX0a6kdoQrjLYwolVvkOhtu6CNvUQdHIfi5WOpxCCDRLxVEQtg/ZuLqlLjop5Sq1WdhFE8
OREAz9sjyICFKK/3yA5fmCLuFro4gJxuFvCO1wvCN71dX7+UsXbYOXYQ9pdWxTftGlJaQSXiGSSj
+vwRhmFX5n1xoa9TsY5sPwdHegalFmwaf2txbLZ8n9dTkf2Qy8rCTGHeN+KqmMWfsC1RkHdpAoJy
9X4KmvCzMvtbs05dyT3OM99lfLqZ5PzBVCDXBWhz4RJ4UVRRQdxwTN8OMQXfsRnrP6S0fF+FAhMT
Ofh58e/j6LAVqNPRbhSFS1D9cQ0t6L29uQrVgoXWR6B1Ct86GbKJlIJr8ecSRFaVBsokOdN7/7XQ
8t66FLlyaHzLRY5wdVUUL6TBmESLXX+NBGkwlSwsT+PO2+itvIRTNlF7ngWwl6FSKQmRnFry4dXM
zmob+HjBugDoCjqBEo3iXmA9s6KcoKkxKTwPCNv3+ujJFbsH7YjmbZZP7Af7VQOq7WInSJ0O/FX2
blTW/x2vy3KxUpOaCA0/ZroOsusOshp1xHsJEMXTm1hIiR9iWdI0ItPPkI42f9eJACtiQi77jtVn
WiTrzBhwaoo6X3hO/SgTa6hAaSEINDgaFH0XO+7RKliQ+kgtjTzi8rA95jkEkAdQJg+ZYIlo3AmS
hlD2LcI6FhCk8NkQUgPM40sGRDExSlrmYolgBDWbUfM9RoPZr4SfJgj2WdCffXW5DzW9obXPk5je
KUTYMeY8R4DxC0JU8SplIYm9PwNv0MxIjfT4YD1ewVmbZI1J30qsd6rsWM/trDhoOE0yEXLPL7nd
kE9wUUnn7Er1c0b5jSgPoZadbCOSEuGlo3mxiWiuRBr6ZNXVX8YRGSGMD+DfCQjoXkn20AIdiv1O
gFfsHk205XqlRozxj9ylKsVkZ6KtYV6V0145IB2zvhZFYfZ7OzQvCitV+qbB/zDgqy2XBsHaDEkg
bBIX+oPainiH04uph4hePlcIxCaXPeG+5jB6LxAuai4MPksdx+dluqAm9J4x+RhpgIhtZcVAxAPW
ojqe58qlrA1amw3UxOuXPk6oboe0OzTZxhFuxlf2f2vkQUInetmGcB0vqbgOwSThgfZlhCj2ILjb
SVirOItNe4jJlbDX2vZntuke+lFf+Vy+ZsE4WXHGX+umjBqZcsl0KBCq8SVVC3ihr9p4QUxwop/J
iUQSVuTO+nyCMkIDhW6vkSFo1mt5X4LaraU3y4VUMaPKSXNd5T3HxMV7AJtSuzngZFM4oS/+Rp/l
qFke8V/D8uLrU4UyleTvVWS444UMB/SJhs0HEddv8gR6G8A5Ls22UMZOMVIfxuzKLq9L/xzEW0NE
h6qMZCoKOY3dxEgyjua0VmDrzXZgGafK0k+eOAIR0ptnZiC0py8m/F5hixkNJS/T7VxkomseUnDh
dCM7JGBxYVL8XIA7ABiqzrVbW2RkPVWSZQyRznP5olgb2wBExGCeygOJUHgsZy5MS06dxsPm++4Z
sADhUrPOPJ+PzHnI9AK1Kpf+cSjVRyeGgAQwiYClTRBC6kz7T4INyxn8AEMfzO/MgG8TQrCs1BM8
j5vmWc8PKHebgKusszXUjcZO/3S08df+U6dzn1ofNzsutVPnRSqXkZZx3k+9XLI3mfb6BaXQR2he
dhlXLkVh1Q5OdOMlKvVL9JdbPn7vQDTmTKsa+BeePS/rCQ1B+DC9WhsnGYHnCvATYoAh2PrqaKSM
hEuecPy/nL59NSqSLYD4eB6PEf6nH6zbewzU0NJVmNfSHaKY19R2A1d2OSVp4WJ/ByNkdB93aC7z
6KiBmCLExJjdZ1TSp+cn/iXLlBxambQn8dPb0KOenMB+HGbN1LObX2RcTVeg9iBC6b1fBY5824BY
BoGfFaDt1nEmh391l7C1TY2s3SsFhxXD/C1zNnEMSOf7miKXK9NAKBiJApCSg6WNGsRdrQs9pP6q
ZikrIPPYs7CfCxJ916f71heSLSYzjK9CgU7ytGNnsdo4+6BIx6s5P30rwIlGlg5R/ocSMZgDBEIP
vRYLDBhcx7Qe08ud7iN2PM6np7mnOYP0+cmytuzQUpERbMPgkXOxuGayKIJkXWzway/eGLmyJ3yY
kokudsU7D9TROwaZerrBOUuBq7OsawIXWS+H5c25pr+SDdbxhxikLqYrSGv+W0fR368asio/gZr8
IMSTfmrFB7QlAzRgvv0Xv6B8U/t+UJkmtcqrHgB6+rWHrLseXrc5pFgd/+isIxrlOkb6ESxVFVhJ
UJXZC5htMFCwgwtJI/7/bXlWXN38crAW0BsDNWJFqWygTWJ2tElWfyXMJKzFBoN3VFGpQfMEGHP3
bHmEGkllK7wct424PRArdrkYxf6dJYnDtpYRFLad2UnJyOwoaFyNUariOgrle7IDBqETyzQoetEI
BZKfRw6SlZv7cO3Qu6aISlYoE+JuYSelSgou3ju3VGBEMSNAGHODk6/yP7NcG8hsIhcR9nZtVZfJ
G7Xrc+6ZVhpOXRtVGt40x2o0cPzysA1vfa/AqlbJa1/LYVTbRRtB61lkUgm0yvSVKy4D1tzTiklO
phI98ZFFEeDiPjiJb5TXRJdh7Om14jw2qZS+aM45VTnmkcLy6+8KKOWgCJDBxC03aK1pvZ8og6HX
pa09BroiHlV89ZtA75SNL9wMo4fbGyi3qO6a76/UPlK3p7U3XEadY3zF75r9tI/IUdLRmqZalchd
b+dlJg8VOKZOwEwM9GCQLnq+4/YHcH+WlZjuuii+zUvkzXGHcrfxdD/aKf2K5JABusymgTkk8jqO
n3SmbSOyKO2xLL5Twj+zwUAG2iEkQSO9rWAZJlcGfzKsMWXNFKsKklbOwp4YIhLytFWQcULdW8Em
tP4g2f9tfIkozr/neugbdVL5Ni9Zev4hLj5PlVJutgIOhgIfl86PMVqXs/gfqkeiEawQgG1z3VIp
Wwi1gblT9hX+pHrPffHrfVfRqgcW5XKo7cdUYHaxPZ+2kaf9HLwFWkYINqSph5YEhUM81fzCb04V
yvGdMk09naN2DNJe0lAM7QRGLg1HxpGiFcC7yx+AO5IQvoqJthdSdnE8uP5ZK06DGB47DkOJ6rGM
v04Q+Vr7CSMGPxnlmXnOuHWwMxup+3YXmYjCXQ4h4ameTxcktkCZRFY3DvXjV6/f80GBZ2zATU0M
p8SCGI/muz5JFKjk+jHUmOA9NO8E8m+CsCp8aNABOhj56Ysm1GOYxcXOj5rXsRStnDLOUs4eAcKu
E1qJBEwnQRQnBcehJ6IZ0KjRE0+KvK7KK7ml9Sb59e5L/ik1cVBASbqved+o2vPLauDe96oUhPqm
vxOijX8+804HnkBsBYLm48MV99to/eZYxYL6nauwDsEbENtpx5pyzU3UooIUTzPxoycbxHGMhfnq
sChJLsVM7iXt9/HsntBgMcCMaCHnmaWZ2nT7tTuWr0CQENqyCQXmRjynV5gmBVoXOCVEz8NyPSvK
4mYtMTsWDcHE6KtyAuYU5MDEsVLyQo/mVj/L+aY11W+jsbN4wU6yf1YbIeQC8r++Ber6YS7zJavx
jnz9zSe9x28SlW5NQRW49hBtfwMqE08Jx7H+orIuQ72Zyl4nD4gwuIeLT8ClJom8jHYQUFd6LVtZ
zlV+WMKhIdpxaNSWkk22jnWoUkHtzEjZJyrODaSIXBRYyZtXrSCRpAE8zwEEK0EdXxfZe+84r+KE
Y0YWVs1ROX8MNMaVq4JqCqHYzd3IzSJAzHIdVlwBB1uSF2Aldd9/9Rx3GEs/dK1z2INAX0jLbFBc
pRR+9iRUynh4MGMFSq9yUFdnLi0tnWPn8yxpCFjg/N/xTtjXLBUSKauAKT9WJ+uaz5h3h9h/MPjp
f6ZMSQx96lF3B5BOAKtU2ycztuTvIKQj0+SXEL7Y5Dw0p8GvR9WOfDrBOeVKdl2ZAN+2VpGBsyzt
pOJVJmUdIyjJC6eBgS4Ks7rMWjnxhrp3l+iaLgpE4EzogaS2w5twBK1z/1Ko5LFxEWBM/lq/kNmD
ZT4Kw6qQSh16FvukIMtiBRzI92CJEqSjmNWG0ZxD48vltn+k1dxaHvcGk6gjZmBBngXz8hA7ZfA0
JLVqGb29Toh3fjYQSn0lhRzncY7c+bxgxzHL+soJx9JUcryDfCQQXRSM8TWZR3j+IsjlltUfQDzC
II3ll35mmzBUh4iNZVc2d+XhW480SVpA4BwzSXNDAAqxZ5GKMOiSAa4y41UeBJj/mHxjnWeBQIUm
CrTBScbJBA93W3z3VtbqsKg8Fk3sRVcEoXx3Q8N/6KQVd2hJQFF3bDGMY/JDLI8lJgODOQsU7iMI
zs+edvR9b1pc4sruY98Vy+2oWoaRuR3KxuFmsDb2a7Qw1Y4BfePU35BphxyjFzT1Oa4W+AA/VNkn
OB541pXjHcuPFXsOVVj4l3iVFfOrF0udjgYUArxaBCgse179YvNbeo9b6QvS2KKNlDiEv3wOQpkd
nd5a4LCnUqsLYjfviKRSa1Br9yOM6JWSJkpwRLZARnlJ7DBcICPAPPBWt5oU9k18KB5cgVIz2hsx
a/ixDS3wc8by1xxtxwMvq2BdPkZHhtaIbSLg7vc0B5nZVXTeoZpqJl+hJnq16zFO1rSBqOgDdIRU
73oeZO83X3bPZVUGAAHCUzNw41ZzrLuqTh2NuC4y4WItqiR1IxQMCPwG0iZMzX0U4E27L4Webqpz
R4CsjD6TsU10aBOQ2CO/sNECLWl7k7sXUbf70Es3/VJ8nJnNl5ywcpOqdEcbMBb8RImouGJEtBue
Hwj40TtjxQRbFgAhpCCBB0jubSigxBSGb4b0vv9ql07R6YilDBEF7z2XmIQTMjcHv8QHKtOxBcPB
/LiFVxzGseYLr+3rCZit8+8Ju3jbkoVprT6T+o40ZM4CIlJ/ch9WdUIIRnTYFXtJG5jIvjStuHja
L+txZoVRVTKXkZzvWHxLipxnb7qih+jAelSkudt1PDzAy0Jak1jSknlhLDNSpPJ2MLYLkERvHQpT
VyIHuxMk+n7SF1EYgnJDr9fw6dlrybZBblMGfNaIh7hob6+6wcZqy091HdlZ9qBJA9Tre0z70zje
du3nADrEsfV2mrgsssfpr9SaUGSMA7FYtoj5vZrjrNmytJFhiXx2VO0NdXjC3H43sMXPeEekWuIq
lLBpFxMHEWX39ZFHGtV4shhAGLZnCVLFbqIq33oR/YpIp9Ygt5y9JHIP12toO4SBg5STix9f4m+R
MW65tkW4cLpv1HAfRU+v+eCyfB5XXLiex5Ud25Xh71ma+VzoaRubff5CLN5fzR8B1q/aGUX9UOtm
NpA6CegLuB6Lr5CcgFaKc+XsX+77eVvfXSqe/nQ23ZQVGd1x5g/0cHVEh6pPp/OC9YsELQ5h69lz
TWMOFDezghiljN5ExPPJpwZAaYrr7Z7RaLJr0p6MqkeUFzrt+EEH5o/D0ymn0ksCxFJk5UJLYPlp
4TsRplyq3rBdkzrdHMZGa8UtkMMv5VtG7sSeeVTpsncJGF+WThrf0DWcxl02f8yNCAKtf/5hwULc
Aolmr8TlEaytm/1TIMhvC5Ue5FqiPunnoSzvPNtHKoQq6+oUYIZYv4lQZV+bX0b+tSkeRcYcndZN
NR8f2QKcQ6cZSMRuRFQwGydRizByHMsSmGs7Btl7WVB8VfEFOQXRJJXlLQqk+7Mn9zcfaaOKUNQs
5EvstN3lEw02LUZMKhGkTt04pHJW0JvooTM4Z5r+07BvZaZNN5+/2hZKnDomgGayURA1DIfYKvWL
F5LLlKUKmBDOS+pLI+M+OzqUa1Ms1pGfhmqU+mhDHtk8q+C+JGbEhj5ElcG0iVVuO3wvUDXplzkM
jP8s+kA9Da1cSvfeuSTjMFZddOU1uOiHVCVX9S2TAKSL30glb08T7AN/dZJjfNjG9aGtigZkzKQO
WzeXLKmhNAJhe0cXa/+gFGgiKrFDAnt9uSBmniGm821XDtQ7KQqAlNrHvrAgAGU3qIxJNKT07/FU
TN2wfdjX0bbdvRygKX4JcdPzVJXe037Duw9NMU/2xAh7dLA4nh1VgI7U87S9QOOCdM8lr3HkxxNj
eJSYK7AplYb6ZHAgQ91jGQijasmOGlDWgLlFtqw+lfQBAtjmiadv0bg8mV+rBK7lrSe/H1xR4ZCk
seXf5mXY8seCectzPjXHYF7zlVn7GFjJkDA+nHZLJnrdsGCJVcCtzJ+RzpExu4GWOlQT+TQtGKuv
DARrNcf91iTeswzcK6cLtM5H1ZHcUN1YxjKi5U/QcJvzRrMioYtM0IR2NqEMgPjuozgBbgxvqTJl
7LZMSXbHcGg4YLvVVxjkM8Os6tuNSNuc3BqeT0NTGGEkwaA+/rYiC4EsCB1KNLAYlRyP6qlQJ2yY
wmw5TnWMSaUCwz6hMcLc5G7OKEWtnofUEMT8BFbkENwiRnfZ0MBMINZTjFr2feiFhqv0H4lr2XCI
oLDFqkbmblw6HtbVzxGXU4fhs02QbDZRxgatbbjhwzNAnYYE7Eq3STRAOt/yE179dqyXedJOUA3I
pXuePmX7HrsracydGFJPysyjccR/kj/AuzaXWZk5WoWJxkDbBWvHg8BPX5Va0yusWf7muEvI//8J
LydskcgNTraufJOMMzxlvFVqTS3vfhViBFV2LfDo7jvt8uwdYvp2PPDgKGWI7VfW2/zJcamne059
mYnLPie0jkgqlItMRzxk19syyDL6nMmlAH/OswdYJmQa6KkbWvabQAgmWMKbb8jywlR06ixd3QBK
KD3Db1HiOxw5rttITDTJBlFX05be+XbX8jHq6Hdjp+u947FEc4y+GdIjEDNJiaxx91UKQMQ7D/FL
vwvzRkOlKVYmKSyU3XzEJK/KUyxwn880h5KlwJJ0h2pCXXWqidVCA5FqxSdYmvAkoKPFdvADSJyJ
fRpYqjtnUNucL+5Tf/77dE/ybSzKxNtJANAmHWzdz+yH0cxPfegaskiwsxvInQDmwjIEiqZi0uZC
BHgk9QulFfeIUI02gdafZJlIBKbtTVAl6LPS95WJXtDwO4N2CG2sfG/W5nr4BmS9UNPClP6inqur
5g7LYZs4t7cZnlupwL91Cn1J0BpQ1SWQwrNuPTuFsTJpYk9u4drUkY0EjHgv8ARD2Gq0m4dAEOcZ
aCef9ZiDJEOD+FhzzDh7VZ81L63id4BrvKLRQOQFGD5byAlUfbAJtQqSr3PZj4MbomdyB/JB9f/K
JT0uRKgdrJp+T0SCNxF4Ah10D+q2NwDvQ1NuAPtE/1vhFCeRKyUdkDhSIPgNXikSC8wsOMLdZPw6
Ds/XkaTNqo8dzVnfKmAvv3NxG7hAnwb/I8IiLeXBkx5RzrPlDLWn0d9/X/5dFadteWh6indAVfcg
SSNmlGtbFG4yIGlWP9RO7cS1QTfXHGfYYpPB6K4ew/toO2Gpy0T4okmP4JieEfYQE6/hauSWQjDc
NPkdbwtWGnJMXO9+8FP0udlwmjBkvBPJE4PADrNc0bKZNKfqOo6zLHBSS40vmH+aDYwrhyMcGGHP
ya4sOs5cD1tBnzoeOH7Gg86KK4vZR5ZhmjQEPjANnlKmAf+/+0qTYZ4KuU7e5+cDUJX8i4DvlXOz
5nfCywdC9ySXUSEg8l1ykKuqw3X6VYSzSiPXpVfbsZJN6UBH4Bj5idiPQtKPgASRC+In4pS0k26P
mjr+HFqeCRUfkP3uREAizMxpTwIn2ygqqw5SHsEyK93A+f7x+f7A3pfswx/+f8PBImVG5NlTiXiH
mj9hWMqtR70jWXuZsqWdwk5C7eYy8Bg7Ldsu0/510+5COFcUfDoLK1IoLPbg6fSqIPr2+k3A8gLB
ajEt6yIWoh4qQtF89UvmOTuS/2r0/AtQd3aDSVeOgrmAtEjhWN+JR1rA5zWCG3BUhISPJhFim14L
X6Dvg6UgJ37hFrJM5piD2NifgBSJNHdEhsJVBVPGSkqmuwxdUjR/RPqHPNeUZoWALxx8u/Ay7QaI
+/vAwVMEKiE9iIPMn9aSL+UGx6wbnZjDfkHM9Dsa+6onV7XNpe4rxLQk+VECJgWHkAKcHEnWEtBo
zqHAlRBZljfbIA7eVQuCdNKDK2HuR6u0Ke5gNU0FiXQmxPUdGowwb6789s5nlOTOHspqq4ayuhDa
Buh61javEkw0aZ/I1UzamcCGAzdDLh6zDVIQmahkiepLxh/t0gKuemyRmQ3mY9Dtm31sOVyu+p+J
wolNVVRLCnvlIRXpcmD9FqoibdrmHF8g3NWIAb3XzFO/x0wykNfwaIxlvAeCKm8hGwA27FtjugZI
C5vnuNqglS44Q+PFLYUfZbgTYQpPwH6mYS17M16DftI0wnw7mPIoDBgmqeVezvGw8gD81fO8o1BN
wemd7n7ya8/UNEfY+ZAxZgHZUmxbgKlmR4ssK3oOSBE7syqVf3ihsGOQWMr4ZbaCtLWG5618AcvL
DrV5OPvMTvy6l+ZisQ88wsctLW0I+GBU+OahmUQ86+fXALKQvOWvmkIKUVduUAany75NQwiXLzox
z1sx57lztHue0sq5+J5cJUcBqWwgt/IHF0Ja30i0wyEY59BKEtcUumWagugO7rAq3vsM7qQZr5Ar
V/PaVX0Z+HaCK4H3pHjq1bXSic79LMgD7b+2iglMa7OXJpyHLmsb1IiTjJ0YbQUjwwB5QHPDKGLu
oFI+D9A2CTLb9nuM5EJKaZhzznrh7zEC0TWImTGS/wjQN73RiubywdIJsWEkWBy6qhzpZr3W8mTV
Uegm2NI3V1x1MkvedFbKogVBO6yyer4g9umkuDr8h8FAVXYfHk+gY703gJw1/LT0uDfb5NHQVN1g
SXTHzjunk9uIbnwjRZrfFmkagy/OPgYBtF/PVRAfhQRjztj4TBRpJ16luvV8GWs+yNEGVhJ97xS5
mM4F7bMzXrpMxEzOalF/Pg2aBzl8FfVdx1VLSJAEu7+G2hEKpOyOM1M1X2SvRetN9F34JSipfxqS
eP0OVfDmRvPrre2O5KVKkDrAJ1TtYUaYQq6XSCfxlU5am4wrDMwrM3FVuYbaZivCcSwQ9b4w27tf
2QDghcz6fW+QEQq1OPr2fN1g1xWhtEkbg3vYfuWdFg+cTkPp8Je6tuLJ8mxwN/9vFV3Ob2fBXSV4
6MTZiQugnmYN83aWncb1TaFzmDP4nv/D71a5srKJ/kyjfLMj9hnVWUA6PbiA33cifYTRys/OJ8xM
EM+54RZvmnMK1NfRjLX+JjMPXZTyMLCkdnF6cKG1JjsNTpO2d7qR4kgszqjLcq5XEcJb7F5b42MS
SyQjAomCvJ9gEtoOyPGpMoE+k2rLIo2vBlx4ItTk4gi5tc9O+CwKIMoz2DI9Honbl7J4KuwUXkdo
t+vyf1q1FDsDP+gv0s/Tvc/2deuqaya3llDud8QwEP2ISXGrMydc3r6IwQ4/Nw4RWPTW3QbsOZck
F+xRu8lUQIq322DRmQ5D/C2VjnjThQaWOT4Wb6sxEqbA2+P1djbxiZQUHGiSUazPWGwXyk7ZIe8B
ZCdyY4pSQaouzCaj02CnhEnSTSq/lg==
`protect end_protected
